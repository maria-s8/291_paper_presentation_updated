module \$paramod$1e0019554db24e403a85d4260c10a25441229a90\plusarg_reader (out);
  output [31:0] out;
  wire [31:0] out;
  assign out = 32'd0;
endmodule
module ALU(io_fn, io_in2, io_in1, io_out, io_adder_out, io_cmp_out);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire _1340_;
  wire _1341_;
  wire _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  wire _1351_;
  wire _1352_;
  wire _1353_;
  wire _1354_;
  wire _1355_;
  wire _1356_;
  wire _1357_;
  wire _1358_;
  wire _1359_;
  wire _1360_;
  wire _1361_;
  wire _1362_;
  wire _1363_;
  wire _1364_;
  wire _1365_;
  wire _1366_;
  wire _1367_;
  wire _1368_;
  wire _1369_;
  wire _1370_;
  wire _1371_;
  wire _1372_;
  wire _1373_;
  wire _1374_;
  wire _1375_;
  wire _1376_;
  wire _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire _1382_;
  wire _1383_;
  wire _1384_;
  wire _1385_;
  wire _1386_;
  wire _1387_;
  wire _1388_;
  wire _1389_;
  wire _1390_;
  wire _1391_;
  wire _1392_;
  wire _1393_;
  wire _1394_;
  wire _1395_;
  wire _1396_;
  wire _1397_;
  wire _1398_;
  wire _1399_;
  wire _1400_;
  wire _1401_;
  wire _1402_;
  wire _1403_;
  wire _1404_;
  wire _1405_;
  wire _1406_;
  wire _1407_;
  wire _1408_;
  wire _1409_;
  wire _1410_;
  wire _1411_;
  wire _1412_;
  wire _1413_;
  wire _1414_;
  wire _1415_;
  wire _1416_;
  wire _1417_;
  wire _1418_;
  wire _1419_;
  wire _1420_;
  wire _1421_;
  wire _1422_;
  wire _1423_;
  wire _1424_;
  wire _1425_;
  wire _1426_;
  wire _1427_;
  wire _1428_;
  wire _1429_;
  wire _1430_;
  wire _1431_;
  wire _1432_;
  wire _1433_;
  wire _1434_;
  wire _1435_;
  wire _1436_;
  wire _1437_;
  wire _1438_;
  wire _1439_;
  wire _1440_;
  wire _1441_;
  wire _1442_;
  wire _1443_;
  wire _1444_;
  wire _1445_;
  wire _1446_;
  wire _1447_;
  wire _1448_;
  wire _1449_;
  wire _1450_;
  wire _1451_;
  wire _1452_;
  wire _1453_;
  wire _1454_;
  wire _1455_;
  wire _1456_;
  wire _1457_;
  wire _1458_;
  wire _1459_;
  wire _1460_;
  wire _1461_;
  wire _1462_;
  wire _1463_;
  wire _1464_;
  wire _1465_;
  wire _1466_;
  wire _1467_;
  wire _1468_;
  wire _1469_;
  wire _1470_;
  wire _1471_;
  wire _1472_;
  wire _1473_;
  wire _1474_;
  wire _1475_;
  wire _1476_;
  wire _1477_;
  wire _1478_;
  wire _1479_;
  wire _1480_;
  wire _1481_;
  wire _1482_;
  wire _1483_;
  wire _1484_;
  wire _1485_;
  wire _1486_;
  wire _1487_;
  wire _1488_;
  wire _1489_;
  wire _1490_;
  wire _1491_;
  wire _1492_;
  wire _1493_;
  wire _1494_;
  wire _1495_;
  wire _1496_;
  wire _1497_;
  wire _1498_;
  wire _1499_;
  wire _1500_;
  wire _1501_;
  wire _1502_;
  wire _1503_;
  wire _1504_;
  wire _1505_;
  wire _1506_;
  wire _1507_;
  wire _1508_;
  wire _1509_;
  wire _1510_;
  wire _1511_;
  wire _1512_;
  wire _1513_;
  wire _1514_;
  wire _1515_;
  wire _1516_;
  wire _1517_;
  wire _1518_;
  wire _1519_;
  wire _1520_;
  wire _1521_;
  wire _1522_;
  wire _1523_;
  wire _1524_;
  wire _1525_;
  wire _1526_;
  wire _1527_;
  wire _1528_;
  wire _1529_;
  wire _1530_;
  wire _1531_;
  wire _1532_;
  wire _1533_;
  wire _1534_;
  wire _1535_;
  wire _1536_;
  wire _1537_;
  wire _1538_;
  wire _1539_;
  wire _1540_;
  wire _1541_;
  wire _1542_;
  wire _1543_;
  wire _1544_;
  wire _1545_;
  wire _1546_;
  wire _1547_;
  wire _1548_;
  wire _1549_;
  wire _1550_;
  wire _1551_;
  wire _1552_;
  wire _1553_;
  wire _1554_;
  wire _1555_;
  wire _1556_;
  wire _1557_;
  wire _1558_;
  wire _1559_;
  wire _1560_;
  wire _1561_;
  wire _1562_;
  wire _1563_;
  wire _1564_;
  wire _1565_;
  wire _1566_;
  wire _1567_;
  wire _1568_;
  wire _1569_;
  wire _1570_;
  wire _1571_;
  wire _1572_;
  wire _1573_;
  wire _1574_;
  wire _1575_;
  wire _1576_;
  wire _1577_;
  wire _1578_;
  wire _1579_;
  wire _1580_;
  wire _1581_;
  wire _1582_;
  wire _1583_;
  wire _1584_;
  wire _1585_;
  wire _1586_;
  wire _1587_;
  wire _1588_;
  wire _1589_;
  wire _1590_;
  wire _1591_;
  wire _1592_;
  wire _1593_;
  wire _1594_;
  wire _1595_;
  wire _1596_;
  wire _1597_;
  wire _1598_;
  wire _1599_;
  wire _1600_;
  wire _1601_;
  wire _1602_;
  wire _1603_;
  wire _1604_;
  wire _1605_;
  wire _1606_;
  wire _1607_;
  wire _1608_;
  wire _1609_;
  wire _1610_;
  wire _1611_;
  wire _1612_;
  wire _1613_;
  wire _1614_;
  wire _1615_;
  wire _1616_;
  wire _1617_;
  wire _1618_;
  wire _1619_;
  wire _1620_;
  wire _1621_;
  wire _1622_;
  wire _1623_;
  wire _1624_;
  wire _1625_;
  wire _1626_;
  wire _1627_;
  wire _1628_;
  wire _1629_;
  wire _1630_;
  wire _1631_;
  wire _1632_;
  wire _1633_;
  wire _1634_;
  wire _1635_;
  wire _1636_;
  wire _1637_;
  wire _1638_;
  wire _1639_;
  wire _1640_;
  wire _1641_;
  wire _1642_;
  wire _1643_;
  wire _1644_;
  wire _1645_;
  wire _1646_;
  wire _1647_;
  wire _1648_;
  wire _1649_;
  wire _1650_;
  wire _1651_;
  wire _1652_;
  wire _1653_;
  wire _1654_;
  wire _1655_;
  wire _1656_;
  wire _1657_;
  wire _1658_;
  wire _1659_;
  wire _1660_;
  wire _1661_;
  wire _1662_;
  wire _1663_;
  wire _1664_;
  wire _1665_;
  wire _1666_;
  wire _1667_;
  wire _1668_;
  wire _1669_;
  wire _1670_;
  wire _1671_;
  wire _1672_;
  wire _1673_;
  wire _1674_;
  wire _1675_;
  wire _1676_;
  wire _1677_;
  wire _1678_;
  wire _1679_;
  wire _1680_;
  wire _1681_;
  wire _1682_;
  wire _1683_;
  wire _1684_;
  wire _1685_;
  wire _1686_;
  wire _1687_;
  wire _1688_;
  wire _1689_;
  wire _1690_;
  wire _1691_;
  wire _1692_;
  wire _1693_;
  wire _1694_;
  wire _1695_;
  wire _1696_;
  wire _1697_;
  wire _1698_;
  wire _1699_;
  wire _1700_;
  wire _1701_;
  wire _1702_;
  wire _1703_;
  wire _1704_;
  wire _1705_;
  wire _1706_;
  wire _1707_;
  wire _1708_;
  wire _1709_;
  wire _1710_;
  wire _1711_;
  wire _1712_;
  wire _1713_;
  wire _1714_;
  wire _1715_;
  wire _1716_;
  wire _1717_;
  wire _1718_;
  wire _1719_;
  wire _1720_;
  wire _1721_;
  wire _1722_;
  wire _1723_;
  wire _1724_;
  wire _1725_;
  wire _1726_;
  wire _1727_;
  wire _1728_;
  wire _1729_;
  wire _1730_;
  wire _1731_;
  wire _1732_;
  wire _1733_;
  wire _1734_;
  wire _1735_;
  wire _1736_;
  wire _1737_;
  wire _1738_;
  wire _1739_;
  wire [31:0] _GEN_0;
  wire [31:0] _GEN_1;
  wire [31:0] _GEN_10;
  wire [31:0] _GEN_11;
  wire [31:0] _GEN_2;
  wire [31:0] _GEN_3;
  wire [31:0] _GEN_4;
  wire [31:0] _GEN_5;
  wire [31:0] _GEN_6;
  wire [31:0] _GEN_7;
  wire [31:0] _GEN_8;
  wire [31:0] _GEN_9;
  wire _shift_logic_T_1;
  wire [31:0] _shin_T_10;
  wire [31:0] _shin_T_11;
  wire [31:0] _shin_T_16;
  wire [31:0] _shin_T_18;
  wire [31:0] _shin_T_20;
  wire [31:0] _shin_T_21;
  wire [31:0] _shin_T_26;
  wire [31:0] _shin_T_28;
  wire [31:0] _shin_T_30;
  wire [31:0] _shin_T_31;
  wire [31:0] _shin_T_36;
  wire [31:0] _shin_T_38;
  wire [31:0] _shin_T_40;
  wire [31:0] _shin_T_41;
  wire [31:0] _shin_T_46;
  wire [31:0] _shin_T_48;
  wire [31:0] _shin_T_50;
  wire [31:0] _shin_T_51;
  wire [31:0] _shin_T_6;
  wire [31:0] _shin_T_8;
  wire [31:0] _shout_l_T_13;
  wire [31:0] _shout_l_T_15;
  wire [31:0] _shout_l_T_17;
  wire [31:0] _shout_l_T_18;
  wire [31:0] _shout_l_T_23;
  wire [31:0] _shout_l_T_25;
  wire [31:0] _shout_l_T_27;
  wire [31:0] _shout_l_T_28;
  wire [31:0] _shout_l_T_3;
  wire [31:0] _shout_l_T_33;
  wire [31:0] _shout_l_T_35;
  wire [31:0] _shout_l_T_37;
  wire [31:0] _shout_l_T_38;
  wire [31:0] _shout_l_T_43;
  wire [31:0] _shout_l_T_45;
  wire [31:0] _shout_l_T_47;
  wire [31:0] _shout_l_T_5;
  wire [31:0] _shout_l_T_7;
  wire [31:0] _shout_l_T_8;
  wire [32:0] _shout_r_T_5;
  output [31:0] io_adder_out;
  wire [31:0] io_adder_out;
  output io_cmp_out;
  wire io_cmp_out;
  input [3:0] io_fn;
  wire [3:0] io_fn;
  input [31:0] io_in1;
  wire [31:0] io_in1;
  input [31:0] io_in2;
  wire [31:0] io_in2;
  output [31:0] io_out;
  wire [31:0] io_out;
  wire [4:0] shamt;
  wire [31:0] shout_l;
  wire [31:0] shout_r;
  INV_X1 _1740_ (
    .A(io_fn[2]),
    .ZN(_0330_)
  );
  INV_X1 _1741_ (
    .A(io_fn[0]),
    .ZN(_0339_)
  );
  INV_X1 _1742_ (
    .A(io_fn[3]),
    .ZN(_0350_)
  );
  INV_X1 _1743_ (
    .A(io_fn[1]),
    .ZN(_0360_)
  );
  INV_X1 _1744_ (
    .A(io_in2[0]),
    .ZN(_0370_)
  );
  INV_X1 _1745_ (
    .A(io_in2[1]),
    .ZN(_0381_)
  );
  INV_X1 _1746_ (
    .A(io_in2[2]),
    .ZN(_0390_)
  );
  INV_X1 _1747_ (
    .A(io_in2[3]),
    .ZN(_0401_)
  );
  INV_X1 _1748_ (
    .A(io_in2[4]),
    .ZN(_0412_)
  );
  INV_X1 _1749_ (
    .A(io_in2[5]),
    .ZN(_0421_)
  );
  INV_X1 _1750_ (
    .A(io_in2[6]),
    .ZN(_0432_)
  );
  INV_X1 _1751_ (
    .A(io_in2[7]),
    .ZN(_0441_)
  );
  INV_X1 _1752_ (
    .A(io_in2[8]),
    .ZN(_0452_)
  );
  INV_X1 _1753_ (
    .A(io_in2[9]),
    .ZN(_0461_)
  );
  INV_X1 _1754_ (
    .A(io_in2[10]),
    .ZN(_0472_)
  );
  INV_X1 _1755_ (
    .A(io_in2[11]),
    .ZN(_0482_)
  );
  INV_X1 _1756_ (
    .A(io_in2[12]),
    .ZN(_0492_)
  );
  INV_X1 _1757_ (
    .A(io_in2[13]),
    .ZN(_0503_)
  );
  INV_X1 _1758_ (
    .A(io_in2[14]),
    .ZN(_0512_)
  );
  INV_X1 _1759_ (
    .A(io_in2[15]),
    .ZN(_0523_)
  );
  INV_X1 _1760_ (
    .A(io_in2[16]),
    .ZN(_0532_)
  );
  INV_X1 _1761_ (
    .A(io_in2[17]),
    .ZN(_0543_)
  );
  INV_X1 _1762_ (
    .A(io_in2[18]),
    .ZN(_0552_)
  );
  INV_X1 _1763_ (
    .A(io_in2[19]),
    .ZN(_0563_)
  );
  INV_X1 _1764_ (
    .A(io_in2[20]),
    .ZN(_0572_)
  );
  INV_X1 _1765_ (
    .A(io_in2[21]),
    .ZN(_0583_)
  );
  INV_X1 _1766_ (
    .A(io_in2[22]),
    .ZN(_0593_)
  );
  INV_X1 _1767_ (
    .A(io_in2[23]),
    .ZN(_0603_)
  );
  INV_X1 _1768_ (
    .A(io_in2[24]),
    .ZN(_0613_)
  );
  INV_X1 _1769_ (
    .A(io_in2[25]),
    .ZN(_0623_)
  );
  INV_X1 _1770_ (
    .A(io_in2[26]),
    .ZN(_0632_)
  );
  INV_X1 _1771_ (
    .A(io_in2[27]),
    .ZN(_0643_)
  );
  INV_X1 _1772_ (
    .A(io_in2[28]),
    .ZN(_0652_)
  );
  INV_X1 _1773_ (
    .A(io_in2[29]),
    .ZN(_0663_)
  );
  INV_X1 _1774_ (
    .A(io_in2[30]),
    .ZN(_0672_)
  );
  INV_X1 _1775_ (
    .A(io_in2[31]),
    .ZN(_0683_)
  );
  INV_X1 _1776_ (
    .A(io_in1[31]),
    .ZN(_0692_)
  );
  INV_X1 _1777_ (
    .A(io_in1[0]),
    .ZN(_0703_)
  );
  INV_X1 _1778_ (
    .A(io_in1[30]),
    .ZN(_0712_)
  );
  INV_X1 _1779_ (
    .A(io_in1[1]),
    .ZN(_0723_)
  );
  INV_X1 _1780_ (
    .A(io_in1[29]),
    .ZN(_0732_)
  );
  INV_X1 _1781_ (
    .A(io_in1[2]),
    .ZN(_0743_)
  );
  INV_X1 _1782_ (
    .A(io_in1[28]),
    .ZN(_0752_)
  );
  INV_X1 _1783_ (
    .A(io_in1[3]),
    .ZN(_0762_)
  );
  INV_X1 _1784_ (
    .A(io_in1[27]),
    .ZN(_0772_)
  );
  INV_X1 _1785_ (
    .A(io_in1[4]),
    .ZN(_0782_)
  );
  INV_X1 _1786_ (
    .A(io_in1[26]),
    .ZN(_0792_)
  );
  INV_X1 _1787_ (
    .A(io_in1[5]),
    .ZN(_0802_)
  );
  INV_X1 _1788_ (
    .A(io_in1[25]),
    .ZN(_0812_)
  );
  INV_X1 _1789_ (
    .A(io_in1[6]),
    .ZN(_0821_)
  );
  INV_X1 _1790_ (
    .A(io_in1[24]),
    .ZN(_0832_)
  );
  INV_X1 _1791_ (
    .A(io_in1[7]),
    .ZN(_0841_)
  );
  INV_X1 _1792_ (
    .A(io_in1[23]),
    .ZN(_0852_)
  );
  INV_X1 _1793_ (
    .A(io_in1[8]),
    .ZN(_0861_)
  );
  INV_X1 _1794_ (
    .A(io_in1[22]),
    .ZN(_0872_)
  );
  INV_X1 _1795_ (
    .A(io_in1[9]),
    .ZN(_0882_)
  );
  INV_X1 _1796_ (
    .A(io_in1[21]),
    .ZN(_0892_)
  );
  INV_X1 _1797_ (
    .A(io_in1[10]),
    .ZN(_0903_)
  );
  INV_X1 _1798_ (
    .A(io_in1[20]),
    .ZN(_0914_)
  );
  INV_X1 _1799_ (
    .A(io_in1[11]),
    .ZN(_0925_)
  );
  INV_X1 _1800_ (
    .A(io_in1[19]),
    .ZN(_0934_)
  );
  INV_X1 _1801_ (
    .A(io_in1[12]),
    .ZN(_0935_)
  );
  INV_X1 _1802_ (
    .A(io_in1[18]),
    .ZN(_0936_)
  );
  INV_X1 _1803_ (
    .A(io_in1[13]),
    .ZN(_0937_)
  );
  INV_X1 _1804_ (
    .A(io_in1[17]),
    .ZN(_0938_)
  );
  INV_X1 _1805_ (
    .A(io_in1[14]),
    .ZN(_0939_)
  );
  INV_X1 _1806_ (
    .A(io_in1[16]),
    .ZN(_0940_)
  );
  INV_X1 _1807_ (
    .A(io_in1[15]),
    .ZN(_0941_)
  );
  AND2_X1 _1808_ (
    .A1(io_fn[3]),
    .A2(_0593_),
    .ZN(_0942_)
  );
  INV_X1 _1809_ (
    .A(_0942_),
    .ZN(_0943_)
  );
  AND2_X1 _1810_ (
    .A1(_0350_),
    .A2(io_in2[22]),
    .ZN(_0944_)
  );
  INV_X1 _1811_ (
    .A(_0944_),
    .ZN(_0945_)
  );
  AND2_X1 _1812_ (
    .A1(_0350_),
    .A2(_0593_),
    .ZN(_0946_)
  );
  INV_X1 _1813_ (
    .A(_0946_),
    .ZN(_0947_)
  );
  AND2_X1 _1814_ (
    .A1(io_fn[3]),
    .A2(io_in2[22]),
    .ZN(_0948_)
  );
  INV_X1 _1815_ (
    .A(_0948_),
    .ZN(_0949_)
  );
  AND2_X1 _1816_ (
    .A1(_0943_),
    .A2(_0945_),
    .ZN(_0950_)
  );
  AND2_X1 _1817_ (
    .A1(_0947_),
    .A2(_0949_),
    .ZN(_0951_)
  );
  AND2_X1 _1818_ (
    .A1(io_in1[22]),
    .A2(_0951_),
    .ZN(_0952_)
  );
  INV_X1 _1819_ (
    .A(_0952_),
    .ZN(_0953_)
  );
  AND2_X1 _1820_ (
    .A1(_0872_),
    .A2(_0950_),
    .ZN(_0954_)
  );
  INV_X1 _1821_ (
    .A(_0954_),
    .ZN(_0955_)
  );
  AND2_X1 _1822_ (
    .A1(_0953_),
    .A2(_0955_),
    .ZN(_0956_)
  );
  INV_X1 _1823_ (
    .A(_0956_),
    .ZN(_0957_)
  );
  AND2_X1 _1824_ (
    .A1(io_fn[3]),
    .A2(_0583_),
    .ZN(_0958_)
  );
  INV_X1 _1825_ (
    .A(_0958_),
    .ZN(_0959_)
  );
  AND2_X1 _1826_ (
    .A1(_0350_),
    .A2(io_in2[21]),
    .ZN(_0960_)
  );
  INV_X1 _1827_ (
    .A(_0960_),
    .ZN(_0961_)
  );
  AND2_X1 _1828_ (
    .A1(_0350_),
    .A2(_0583_),
    .ZN(_0962_)
  );
  INV_X1 _1829_ (
    .A(_0962_),
    .ZN(_0963_)
  );
  AND2_X1 _1830_ (
    .A1(io_fn[3]),
    .A2(io_in2[21]),
    .ZN(_0964_)
  );
  INV_X1 _1831_ (
    .A(_0964_),
    .ZN(_0965_)
  );
  AND2_X1 _1832_ (
    .A1(_0959_),
    .A2(_0961_),
    .ZN(_0966_)
  );
  AND2_X1 _1833_ (
    .A1(_0963_),
    .A2(_0965_),
    .ZN(_0967_)
  );
  AND2_X1 _1834_ (
    .A1(io_in1[21]),
    .A2(_0967_),
    .ZN(_0968_)
  );
  INV_X1 _1835_ (
    .A(_0968_),
    .ZN(_0969_)
  );
  AND2_X1 _1836_ (
    .A1(_0892_),
    .A2(_0966_),
    .ZN(_0970_)
  );
  INV_X1 _1837_ (
    .A(_0970_),
    .ZN(_0971_)
  );
  AND2_X1 _1838_ (
    .A1(io_fn[3]),
    .A2(_0572_),
    .ZN(_0972_)
  );
  INV_X1 _1839_ (
    .A(_0972_),
    .ZN(_0973_)
  );
  AND2_X1 _1840_ (
    .A1(_0350_),
    .A2(io_in2[20]),
    .ZN(_0974_)
  );
  INV_X1 _1841_ (
    .A(_0974_),
    .ZN(_0975_)
  );
  AND2_X1 _1842_ (
    .A1(_0350_),
    .A2(_0572_),
    .ZN(_0976_)
  );
  INV_X1 _1843_ (
    .A(_0976_),
    .ZN(_0977_)
  );
  AND2_X1 _1844_ (
    .A1(io_fn[3]),
    .A2(io_in2[20]),
    .ZN(_0978_)
  );
  INV_X1 _1845_ (
    .A(_0978_),
    .ZN(_0979_)
  );
  AND2_X1 _1846_ (
    .A1(_0973_),
    .A2(_0975_),
    .ZN(_0980_)
  );
  AND2_X1 _1847_ (
    .A1(_0977_),
    .A2(_0979_),
    .ZN(_0981_)
  );
  AND2_X1 _1848_ (
    .A1(io_in1[20]),
    .A2(_0981_),
    .ZN(_0982_)
  );
  INV_X1 _1849_ (
    .A(_0982_),
    .ZN(_0983_)
  );
  AND2_X1 _1850_ (
    .A1(_0914_),
    .A2(_0980_),
    .ZN(_0984_)
  );
  INV_X1 _1851_ (
    .A(_0984_),
    .ZN(_0985_)
  );
  AND2_X1 _1852_ (
    .A1(_0983_),
    .A2(_0985_),
    .ZN(_0986_)
  );
  INV_X1 _1853_ (
    .A(_0986_),
    .ZN(_0987_)
  );
  AND2_X1 _1854_ (
    .A1(io_fn[3]),
    .A2(_0563_),
    .ZN(_0988_)
  );
  INV_X1 _1855_ (
    .A(_0988_),
    .ZN(_0989_)
  );
  AND2_X1 _1856_ (
    .A1(_0350_),
    .A2(io_in2[19]),
    .ZN(_0990_)
  );
  INV_X1 _1857_ (
    .A(_0990_),
    .ZN(_0991_)
  );
  AND2_X1 _1858_ (
    .A1(_0350_),
    .A2(_0563_),
    .ZN(_0992_)
  );
  INV_X1 _1859_ (
    .A(_0992_),
    .ZN(_0993_)
  );
  AND2_X1 _1860_ (
    .A1(io_fn[3]),
    .A2(io_in2[19]),
    .ZN(_0994_)
  );
  INV_X1 _1861_ (
    .A(_0994_),
    .ZN(_0995_)
  );
  AND2_X1 _1862_ (
    .A1(_0989_),
    .A2(_0991_),
    .ZN(_0996_)
  );
  AND2_X1 _1863_ (
    .A1(_0993_),
    .A2(_0995_),
    .ZN(_0997_)
  );
  AND2_X1 _1864_ (
    .A1(io_in1[19]),
    .A2(_0997_),
    .ZN(_0998_)
  );
  INV_X1 _1865_ (
    .A(_0998_),
    .ZN(_0999_)
  );
  AND2_X1 _1866_ (
    .A1(_0934_),
    .A2(_0996_),
    .ZN(_1000_)
  );
  INV_X1 _1867_ (
    .A(_1000_),
    .ZN(_1001_)
  );
  AND2_X1 _1868_ (
    .A1(_0999_),
    .A2(_1001_),
    .ZN(_1002_)
  );
  INV_X1 _1869_ (
    .A(_1002_),
    .ZN(_1003_)
  );
  AND2_X1 _1870_ (
    .A1(io_fn[3]),
    .A2(_0552_),
    .ZN(_1004_)
  );
  INV_X1 _1871_ (
    .A(_1004_),
    .ZN(_1005_)
  );
  AND2_X1 _1872_ (
    .A1(_0350_),
    .A2(io_in2[18]),
    .ZN(_1006_)
  );
  INV_X1 _1873_ (
    .A(_1006_),
    .ZN(_1007_)
  );
  AND2_X1 _1874_ (
    .A1(_0350_),
    .A2(_0552_),
    .ZN(_1008_)
  );
  INV_X1 _1875_ (
    .A(_1008_),
    .ZN(_1009_)
  );
  AND2_X1 _1876_ (
    .A1(io_fn[3]),
    .A2(io_in2[18]),
    .ZN(_1010_)
  );
  INV_X1 _1877_ (
    .A(_1010_),
    .ZN(_1011_)
  );
  AND2_X1 _1878_ (
    .A1(_1005_),
    .A2(_1007_),
    .ZN(_1012_)
  );
  AND2_X1 _1879_ (
    .A1(_1009_),
    .A2(_1011_),
    .ZN(_1013_)
  );
  AND2_X1 _1880_ (
    .A1(io_in1[18]),
    .A2(_1013_),
    .ZN(_1014_)
  );
  INV_X1 _1881_ (
    .A(_1014_),
    .ZN(_1015_)
  );
  AND2_X1 _1882_ (
    .A1(_0936_),
    .A2(_1012_),
    .ZN(_1016_)
  );
  INV_X1 _1883_ (
    .A(_1016_),
    .ZN(_1017_)
  );
  AND2_X1 _1884_ (
    .A1(_1015_),
    .A2(_1017_),
    .ZN(_1018_)
  );
  INV_X1 _1885_ (
    .A(_1018_),
    .ZN(_1019_)
  );
  AND2_X1 _1886_ (
    .A1(io_fn[3]),
    .A2(_0543_),
    .ZN(_1020_)
  );
  INV_X1 _1887_ (
    .A(_1020_),
    .ZN(_1021_)
  );
  AND2_X1 _1888_ (
    .A1(_0350_),
    .A2(io_in2[17]),
    .ZN(_1022_)
  );
  INV_X1 _1889_ (
    .A(_1022_),
    .ZN(_1023_)
  );
  AND2_X1 _1890_ (
    .A1(_0350_),
    .A2(_0543_),
    .ZN(_1024_)
  );
  INV_X1 _1891_ (
    .A(_1024_),
    .ZN(_1025_)
  );
  AND2_X1 _1892_ (
    .A1(io_fn[3]),
    .A2(io_in2[17]),
    .ZN(_1026_)
  );
  INV_X1 _1893_ (
    .A(_1026_),
    .ZN(_1027_)
  );
  AND2_X1 _1894_ (
    .A1(_1021_),
    .A2(_1023_),
    .ZN(_1028_)
  );
  AND2_X1 _1895_ (
    .A1(_1025_),
    .A2(_1027_),
    .ZN(_1029_)
  );
  AND2_X1 _1896_ (
    .A1(io_in1[17]),
    .A2(_1029_),
    .ZN(_1030_)
  );
  INV_X1 _1897_ (
    .A(_1030_),
    .ZN(_1031_)
  );
  AND2_X1 _1898_ (
    .A1(io_fn[3]),
    .A2(_0532_),
    .ZN(_1032_)
  );
  INV_X1 _1899_ (
    .A(_1032_),
    .ZN(_1033_)
  );
  AND2_X1 _1900_ (
    .A1(_0350_),
    .A2(io_in2[16]),
    .ZN(_1034_)
  );
  INV_X1 _1901_ (
    .A(_1034_),
    .ZN(_1035_)
  );
  AND2_X1 _1902_ (
    .A1(_0350_),
    .A2(_0532_),
    .ZN(_1036_)
  );
  INV_X1 _1903_ (
    .A(_1036_),
    .ZN(_1037_)
  );
  AND2_X1 _1904_ (
    .A1(io_fn[3]),
    .A2(io_in2[16]),
    .ZN(_1038_)
  );
  INV_X1 _1905_ (
    .A(_1038_),
    .ZN(_1039_)
  );
  AND2_X1 _1906_ (
    .A1(_1033_),
    .A2(_1035_),
    .ZN(_1040_)
  );
  AND2_X1 _1907_ (
    .A1(_1037_),
    .A2(_1039_),
    .ZN(_1041_)
  );
  AND2_X1 _1908_ (
    .A1(io_in1[16]),
    .A2(_1041_),
    .ZN(_1042_)
  );
  INV_X1 _1909_ (
    .A(_1042_),
    .ZN(_1043_)
  );
  AND2_X1 _1910_ (
    .A1(io_fn[3]),
    .A2(_0523_),
    .ZN(_1044_)
  );
  INV_X1 _1911_ (
    .A(_1044_),
    .ZN(_1045_)
  );
  AND2_X1 _1912_ (
    .A1(_0350_),
    .A2(io_in2[15]),
    .ZN(_1046_)
  );
  INV_X1 _1913_ (
    .A(_1046_),
    .ZN(_1047_)
  );
  AND2_X1 _1914_ (
    .A1(_0350_),
    .A2(_0523_),
    .ZN(_1048_)
  );
  INV_X1 _1915_ (
    .A(_1048_),
    .ZN(_1049_)
  );
  AND2_X1 _1916_ (
    .A1(io_fn[3]),
    .A2(io_in2[15]),
    .ZN(_1050_)
  );
  INV_X1 _1917_ (
    .A(_1050_),
    .ZN(_1051_)
  );
  AND2_X1 _1918_ (
    .A1(_1045_),
    .A2(_1047_),
    .ZN(_1052_)
  );
  AND2_X1 _1919_ (
    .A1(_1049_),
    .A2(_1051_),
    .ZN(_1053_)
  );
  AND2_X1 _1920_ (
    .A1(_0941_),
    .A2(_1052_),
    .ZN(_1054_)
  );
  INV_X1 _1921_ (
    .A(_1054_),
    .ZN(_1055_)
  );
  AND2_X1 _1922_ (
    .A1(io_in1[15]),
    .A2(_1053_),
    .ZN(_1056_)
  );
  INV_X1 _1923_ (
    .A(_1056_),
    .ZN(_1057_)
  );
  AND2_X1 _1924_ (
    .A1(_1055_),
    .A2(_1057_),
    .ZN(_1058_)
  );
  INV_X1 _1925_ (
    .A(_1058_),
    .ZN(_1059_)
  );
  AND2_X1 _1926_ (
    .A1(io_fn[3]),
    .A2(_0512_),
    .ZN(_1060_)
  );
  INV_X1 _1927_ (
    .A(_1060_),
    .ZN(_1061_)
  );
  AND2_X1 _1928_ (
    .A1(_0350_),
    .A2(io_in2[14]),
    .ZN(_1062_)
  );
  INV_X1 _1929_ (
    .A(_1062_),
    .ZN(_1063_)
  );
  AND2_X1 _1930_ (
    .A1(_0350_),
    .A2(_0512_),
    .ZN(_1064_)
  );
  INV_X1 _1931_ (
    .A(_1064_),
    .ZN(_1065_)
  );
  AND2_X1 _1932_ (
    .A1(io_fn[3]),
    .A2(io_in2[14]),
    .ZN(_1066_)
  );
  INV_X1 _1933_ (
    .A(_1066_),
    .ZN(_1067_)
  );
  AND2_X1 _1934_ (
    .A1(_1061_),
    .A2(_1063_),
    .ZN(_1068_)
  );
  AND2_X1 _1935_ (
    .A1(_1065_),
    .A2(_1067_),
    .ZN(_1069_)
  );
  AND2_X1 _1936_ (
    .A1(io_in1[14]),
    .A2(_1069_),
    .ZN(_1070_)
  );
  INV_X1 _1937_ (
    .A(_1070_),
    .ZN(_1071_)
  );
  AND2_X1 _1938_ (
    .A1(_0939_),
    .A2(_1068_),
    .ZN(_1072_)
  );
  INV_X1 _1939_ (
    .A(_1072_),
    .ZN(_1073_)
  );
  AND2_X1 _1940_ (
    .A1(_1071_),
    .A2(_1073_),
    .ZN(_1074_)
  );
  INV_X1 _1941_ (
    .A(_1074_),
    .ZN(_1075_)
  );
  AND2_X1 _1942_ (
    .A1(io_fn[3]),
    .A2(_0503_),
    .ZN(_1076_)
  );
  INV_X1 _1943_ (
    .A(_1076_),
    .ZN(_1077_)
  );
  AND2_X1 _1944_ (
    .A1(_0350_),
    .A2(io_in2[13]),
    .ZN(_1078_)
  );
  INV_X1 _1945_ (
    .A(_1078_),
    .ZN(_1079_)
  );
  AND2_X1 _1946_ (
    .A1(_0350_),
    .A2(_0503_),
    .ZN(_1080_)
  );
  INV_X1 _1947_ (
    .A(_1080_),
    .ZN(_1081_)
  );
  AND2_X1 _1948_ (
    .A1(io_fn[3]),
    .A2(io_in2[13]),
    .ZN(_1082_)
  );
  INV_X1 _1949_ (
    .A(_1082_),
    .ZN(_1083_)
  );
  AND2_X1 _1950_ (
    .A1(_1077_),
    .A2(_1079_),
    .ZN(_1084_)
  );
  AND2_X1 _1951_ (
    .A1(_1081_),
    .A2(_1083_),
    .ZN(_1085_)
  );
  AND2_X1 _1952_ (
    .A1(io_in1[13]),
    .A2(_1085_),
    .ZN(_1086_)
  );
  INV_X1 _1953_ (
    .A(_1086_),
    .ZN(_1087_)
  );
  AND2_X1 _1954_ (
    .A1(_0937_),
    .A2(_1084_),
    .ZN(_1088_)
  );
  INV_X1 _1955_ (
    .A(_1088_),
    .ZN(_1089_)
  );
  AND2_X1 _1956_ (
    .A1(_1087_),
    .A2(_1089_),
    .ZN(_1090_)
  );
  INV_X1 _1957_ (
    .A(_1090_),
    .ZN(_1091_)
  );
  AND2_X1 _1958_ (
    .A1(io_fn[3]),
    .A2(_0492_),
    .ZN(_1092_)
  );
  INV_X1 _1959_ (
    .A(_1092_),
    .ZN(_1093_)
  );
  AND2_X1 _1960_ (
    .A1(_0350_),
    .A2(io_in2[12]),
    .ZN(_1094_)
  );
  INV_X1 _1961_ (
    .A(_1094_),
    .ZN(_1095_)
  );
  AND2_X1 _1962_ (
    .A1(_0350_),
    .A2(_0492_),
    .ZN(_1096_)
  );
  INV_X1 _1963_ (
    .A(_1096_),
    .ZN(_1097_)
  );
  AND2_X1 _1964_ (
    .A1(io_fn[3]),
    .A2(io_in2[12]),
    .ZN(_1098_)
  );
  INV_X1 _1965_ (
    .A(_1098_),
    .ZN(_1099_)
  );
  AND2_X1 _1966_ (
    .A1(_1093_),
    .A2(_1095_),
    .ZN(_1100_)
  );
  AND2_X1 _1967_ (
    .A1(_1097_),
    .A2(_1099_),
    .ZN(_1101_)
  );
  AND2_X1 _1968_ (
    .A1(io_in1[12]),
    .A2(_1101_),
    .ZN(_1102_)
  );
  INV_X1 _1969_ (
    .A(_1102_),
    .ZN(_1103_)
  );
  AND2_X1 _1970_ (
    .A1(_0935_),
    .A2(_1100_),
    .ZN(_1104_)
  );
  INV_X1 _1971_ (
    .A(_1104_),
    .ZN(_1105_)
  );
  AND2_X1 _1972_ (
    .A1(_1103_),
    .A2(_1105_),
    .ZN(_1106_)
  );
  INV_X1 _1973_ (
    .A(_1106_),
    .ZN(_1107_)
  );
  AND2_X1 _1974_ (
    .A1(io_fn[3]),
    .A2(_0482_),
    .ZN(_1108_)
  );
  INV_X1 _1975_ (
    .A(_1108_),
    .ZN(_1109_)
  );
  AND2_X1 _1976_ (
    .A1(_0350_),
    .A2(io_in2[11]),
    .ZN(_1110_)
  );
  INV_X1 _1977_ (
    .A(_1110_),
    .ZN(_1111_)
  );
  AND2_X1 _1978_ (
    .A1(_0350_),
    .A2(_0482_),
    .ZN(_1112_)
  );
  INV_X1 _1979_ (
    .A(_1112_),
    .ZN(_1113_)
  );
  AND2_X1 _1980_ (
    .A1(io_fn[3]),
    .A2(io_in2[11]),
    .ZN(_1114_)
  );
  INV_X1 _1981_ (
    .A(_1114_),
    .ZN(_1115_)
  );
  AND2_X1 _1982_ (
    .A1(_1109_),
    .A2(_1111_),
    .ZN(_1116_)
  );
  AND2_X1 _1983_ (
    .A1(_1113_),
    .A2(_1115_),
    .ZN(_1117_)
  );
  AND2_X1 _1984_ (
    .A1(io_in1[11]),
    .A2(_1117_),
    .ZN(_1118_)
  );
  INV_X1 _1985_ (
    .A(_1118_),
    .ZN(_1119_)
  );
  AND2_X1 _1986_ (
    .A1(_0925_),
    .A2(_1116_),
    .ZN(_1120_)
  );
  INV_X1 _1987_ (
    .A(_1120_),
    .ZN(_1121_)
  );
  AND2_X1 _1988_ (
    .A1(_1119_),
    .A2(_1121_),
    .ZN(_1122_)
  );
  INV_X1 _1989_ (
    .A(_1122_),
    .ZN(_1123_)
  );
  AND2_X1 _1990_ (
    .A1(io_fn[3]),
    .A2(_0472_),
    .ZN(_1124_)
  );
  INV_X1 _1991_ (
    .A(_1124_),
    .ZN(_1125_)
  );
  AND2_X1 _1992_ (
    .A1(_0350_),
    .A2(io_in2[10]),
    .ZN(_1126_)
  );
  INV_X1 _1993_ (
    .A(_1126_),
    .ZN(_1127_)
  );
  AND2_X1 _1994_ (
    .A1(_0350_),
    .A2(_0472_),
    .ZN(_1128_)
  );
  INV_X1 _1995_ (
    .A(_1128_),
    .ZN(_1129_)
  );
  AND2_X1 _1996_ (
    .A1(io_fn[3]),
    .A2(io_in2[10]),
    .ZN(_1130_)
  );
  INV_X1 _1997_ (
    .A(_1130_),
    .ZN(_1131_)
  );
  AND2_X1 _1998_ (
    .A1(_1125_),
    .A2(_1127_),
    .ZN(_1132_)
  );
  AND2_X1 _1999_ (
    .A1(_1129_),
    .A2(_1131_),
    .ZN(_1133_)
  );
  AND2_X1 _2000_ (
    .A1(io_in1[10]),
    .A2(_1133_),
    .ZN(_1134_)
  );
  INV_X1 _2001_ (
    .A(_1134_),
    .ZN(_1135_)
  );
  AND2_X1 _2002_ (
    .A1(_0903_),
    .A2(_1132_),
    .ZN(_1136_)
  );
  INV_X1 _2003_ (
    .A(_1136_),
    .ZN(_1137_)
  );
  AND2_X1 _2004_ (
    .A1(_1135_),
    .A2(_1137_),
    .ZN(_1138_)
  );
  INV_X1 _2005_ (
    .A(_1138_),
    .ZN(_1139_)
  );
  AND2_X1 _2006_ (
    .A1(io_fn[3]),
    .A2(_0461_),
    .ZN(_1140_)
  );
  INV_X1 _2007_ (
    .A(_1140_),
    .ZN(_1141_)
  );
  AND2_X1 _2008_ (
    .A1(_0350_),
    .A2(io_in2[9]),
    .ZN(_1142_)
  );
  INV_X1 _2009_ (
    .A(_1142_),
    .ZN(_1143_)
  );
  AND2_X1 _2010_ (
    .A1(_0350_),
    .A2(_0461_),
    .ZN(_1144_)
  );
  INV_X1 _2011_ (
    .A(_1144_),
    .ZN(_1145_)
  );
  AND2_X1 _2012_ (
    .A1(io_fn[3]),
    .A2(io_in2[9]),
    .ZN(_1146_)
  );
  INV_X1 _2013_ (
    .A(_1146_),
    .ZN(_1147_)
  );
  AND2_X1 _2014_ (
    .A1(_1141_),
    .A2(_1143_),
    .ZN(_1148_)
  );
  AND2_X1 _2015_ (
    .A1(_1145_),
    .A2(_1147_),
    .ZN(_1149_)
  );
  AND2_X1 _2016_ (
    .A1(io_in1[9]),
    .A2(_1149_),
    .ZN(_1150_)
  );
  INV_X1 _2017_ (
    .A(_1150_),
    .ZN(_1151_)
  );
  AND2_X1 _2018_ (
    .A1(_0882_),
    .A2(_1148_),
    .ZN(_1152_)
  );
  INV_X1 _2019_ (
    .A(_1152_),
    .ZN(_1153_)
  );
  AND2_X1 _2020_ (
    .A1(_1151_),
    .A2(_1153_),
    .ZN(_1154_)
  );
  INV_X1 _2021_ (
    .A(_1154_),
    .ZN(_1155_)
  );
  AND2_X1 _2022_ (
    .A1(io_fn[3]),
    .A2(_0452_),
    .ZN(_1156_)
  );
  INV_X1 _2023_ (
    .A(_1156_),
    .ZN(_1157_)
  );
  AND2_X1 _2024_ (
    .A1(_0350_),
    .A2(io_in2[8]),
    .ZN(_1158_)
  );
  INV_X1 _2025_ (
    .A(_1158_),
    .ZN(_1159_)
  );
  AND2_X1 _2026_ (
    .A1(_0350_),
    .A2(_0452_),
    .ZN(_1160_)
  );
  INV_X1 _2027_ (
    .A(_1160_),
    .ZN(_1161_)
  );
  AND2_X1 _2028_ (
    .A1(io_fn[3]),
    .A2(io_in2[8]),
    .ZN(_1162_)
  );
  INV_X1 _2029_ (
    .A(_1162_),
    .ZN(_1163_)
  );
  AND2_X1 _2030_ (
    .A1(_1157_),
    .A2(_1159_),
    .ZN(_1164_)
  );
  AND2_X1 _2031_ (
    .A1(_1161_),
    .A2(_1163_),
    .ZN(_1165_)
  );
  AND2_X1 _2032_ (
    .A1(io_in1[8]),
    .A2(_1165_),
    .ZN(_1166_)
  );
  INV_X1 _2033_ (
    .A(_1166_),
    .ZN(_1167_)
  );
  AND2_X1 _2034_ (
    .A1(io_fn[3]),
    .A2(_0441_),
    .ZN(_1168_)
  );
  INV_X1 _2035_ (
    .A(_1168_),
    .ZN(_1169_)
  );
  AND2_X1 _2036_ (
    .A1(_0350_),
    .A2(io_in2[7]),
    .ZN(_1170_)
  );
  INV_X1 _2037_ (
    .A(_1170_),
    .ZN(_1171_)
  );
  AND2_X1 _2038_ (
    .A1(_0350_),
    .A2(_0441_),
    .ZN(_1172_)
  );
  INV_X1 _2039_ (
    .A(_1172_),
    .ZN(_1173_)
  );
  AND2_X1 _2040_ (
    .A1(io_fn[3]),
    .A2(io_in2[7]),
    .ZN(_1174_)
  );
  INV_X1 _2041_ (
    .A(_1174_),
    .ZN(_1175_)
  );
  AND2_X1 _2042_ (
    .A1(_1169_),
    .A2(_1171_),
    .ZN(_1176_)
  );
  AND2_X1 _2043_ (
    .A1(_1173_),
    .A2(_1175_),
    .ZN(_1177_)
  );
  AND2_X1 _2044_ (
    .A1(io_in1[7]),
    .A2(_1177_),
    .ZN(_1178_)
  );
  INV_X1 _2045_ (
    .A(_1178_),
    .ZN(_1179_)
  );
  AND2_X1 _2046_ (
    .A1(_0841_),
    .A2(_1176_),
    .ZN(_1180_)
  );
  INV_X1 _2047_ (
    .A(_1180_),
    .ZN(_1181_)
  );
  AND2_X1 _2048_ (
    .A1(_1179_),
    .A2(_1181_),
    .ZN(_1182_)
  );
  INV_X1 _2049_ (
    .A(_1182_),
    .ZN(_1183_)
  );
  AND2_X1 _2050_ (
    .A1(io_fn[3]),
    .A2(_0432_),
    .ZN(_1184_)
  );
  INV_X1 _2051_ (
    .A(_1184_),
    .ZN(_1185_)
  );
  AND2_X1 _2052_ (
    .A1(_0350_),
    .A2(io_in2[6]),
    .ZN(_1186_)
  );
  INV_X1 _2053_ (
    .A(_1186_),
    .ZN(_1187_)
  );
  AND2_X1 _2054_ (
    .A1(_0350_),
    .A2(_0432_),
    .ZN(_1188_)
  );
  INV_X1 _2055_ (
    .A(_1188_),
    .ZN(_1189_)
  );
  AND2_X1 _2056_ (
    .A1(io_fn[3]),
    .A2(io_in2[6]),
    .ZN(_1190_)
  );
  INV_X1 _2057_ (
    .A(_1190_),
    .ZN(_1191_)
  );
  AND2_X1 _2058_ (
    .A1(_1185_),
    .A2(_1187_),
    .ZN(_1192_)
  );
  AND2_X1 _2059_ (
    .A1(_1189_),
    .A2(_1191_),
    .ZN(_1193_)
  );
  AND2_X1 _2060_ (
    .A1(io_in1[6]),
    .A2(_1193_),
    .ZN(_1194_)
  );
  INV_X1 _2061_ (
    .A(_1194_),
    .ZN(_1195_)
  );
  AND2_X1 _2062_ (
    .A1(_0821_),
    .A2(_1192_),
    .ZN(_1196_)
  );
  INV_X1 _2063_ (
    .A(_1196_),
    .ZN(_1197_)
  );
  AND2_X1 _2064_ (
    .A1(_1195_),
    .A2(_1197_),
    .ZN(_1198_)
  );
  INV_X1 _2065_ (
    .A(_1198_),
    .ZN(_1199_)
  );
  AND2_X1 _2066_ (
    .A1(io_fn[3]),
    .A2(_0421_),
    .ZN(_1200_)
  );
  INV_X1 _2067_ (
    .A(_1200_),
    .ZN(_1201_)
  );
  AND2_X1 _2068_ (
    .A1(_0350_),
    .A2(io_in2[5]),
    .ZN(_1202_)
  );
  INV_X1 _2069_ (
    .A(_1202_),
    .ZN(_1203_)
  );
  AND2_X1 _2070_ (
    .A1(_0350_),
    .A2(_0421_),
    .ZN(_1204_)
  );
  INV_X1 _2071_ (
    .A(_1204_),
    .ZN(_1205_)
  );
  AND2_X1 _2072_ (
    .A1(io_fn[3]),
    .A2(io_in2[5]),
    .ZN(_1206_)
  );
  INV_X1 _2073_ (
    .A(_1206_),
    .ZN(_1207_)
  );
  AND2_X1 _2074_ (
    .A1(_1201_),
    .A2(_1203_),
    .ZN(_1208_)
  );
  AND2_X1 _2075_ (
    .A1(_1205_),
    .A2(_1207_),
    .ZN(_1209_)
  );
  AND2_X1 _2076_ (
    .A1(io_in1[5]),
    .A2(_1209_),
    .ZN(_1210_)
  );
  INV_X1 _2077_ (
    .A(_1210_),
    .ZN(_1211_)
  );
  AND2_X1 _2078_ (
    .A1(io_fn[3]),
    .A2(_0412_),
    .ZN(_1212_)
  );
  INV_X1 _2079_ (
    .A(_1212_),
    .ZN(_1213_)
  );
  AND2_X1 _2080_ (
    .A1(_0350_),
    .A2(io_in2[4]),
    .ZN(_1214_)
  );
  INV_X1 _2081_ (
    .A(_1214_),
    .ZN(_1215_)
  );
  AND2_X1 _2082_ (
    .A1(_0350_),
    .A2(_0412_),
    .ZN(_1216_)
  );
  INV_X1 _2083_ (
    .A(_1216_),
    .ZN(_1217_)
  );
  AND2_X1 _2084_ (
    .A1(io_fn[3]),
    .A2(io_in2[4]),
    .ZN(_1218_)
  );
  INV_X1 _2085_ (
    .A(_1218_),
    .ZN(_1219_)
  );
  AND2_X1 _2086_ (
    .A1(_1213_),
    .A2(_1215_),
    .ZN(_1220_)
  );
  AND2_X1 _2087_ (
    .A1(_1217_),
    .A2(_1219_),
    .ZN(_1221_)
  );
  AND2_X1 _2088_ (
    .A1(io_in1[4]),
    .A2(_1221_),
    .ZN(_1222_)
  );
  INV_X1 _2089_ (
    .A(_1222_),
    .ZN(_1223_)
  );
  AND2_X1 _2090_ (
    .A1(io_fn[3]),
    .A2(_0401_),
    .ZN(_1224_)
  );
  INV_X1 _2091_ (
    .A(_1224_),
    .ZN(_1225_)
  );
  AND2_X1 _2092_ (
    .A1(_0350_),
    .A2(io_in2[3]),
    .ZN(_1226_)
  );
  INV_X1 _2093_ (
    .A(_1226_),
    .ZN(_1227_)
  );
  AND2_X1 _2094_ (
    .A1(_0350_),
    .A2(_0401_),
    .ZN(_1228_)
  );
  INV_X1 _2095_ (
    .A(_1228_),
    .ZN(_1229_)
  );
  AND2_X1 _2096_ (
    .A1(io_fn[3]),
    .A2(io_in2[3]),
    .ZN(_1230_)
  );
  INV_X1 _2097_ (
    .A(_1230_),
    .ZN(_1231_)
  );
  AND2_X1 _2098_ (
    .A1(_1225_),
    .A2(_1227_),
    .ZN(_1232_)
  );
  AND2_X1 _2099_ (
    .A1(_1229_),
    .A2(_1231_),
    .ZN(_1233_)
  );
  AND2_X1 _2100_ (
    .A1(io_in1[3]),
    .A2(_1233_),
    .ZN(_1234_)
  );
  INV_X1 _2101_ (
    .A(_1234_),
    .ZN(_1235_)
  );
  AND2_X1 _2102_ (
    .A1(io_fn[3]),
    .A2(_0390_),
    .ZN(_1236_)
  );
  INV_X1 _2103_ (
    .A(_1236_),
    .ZN(_1237_)
  );
  AND2_X1 _2104_ (
    .A1(_0350_),
    .A2(io_in2[2]),
    .ZN(_1238_)
  );
  INV_X1 _2105_ (
    .A(_1238_),
    .ZN(_1239_)
  );
  AND2_X1 _2106_ (
    .A1(_0350_),
    .A2(_0390_),
    .ZN(_1240_)
  );
  INV_X1 _2107_ (
    .A(_1240_),
    .ZN(_1241_)
  );
  AND2_X1 _2108_ (
    .A1(io_fn[3]),
    .A2(io_in2[2]),
    .ZN(_1242_)
  );
  INV_X1 _2109_ (
    .A(_1242_),
    .ZN(_1243_)
  );
  AND2_X1 _2110_ (
    .A1(_1237_),
    .A2(_1239_),
    .ZN(_1244_)
  );
  AND2_X1 _2111_ (
    .A1(_1241_),
    .A2(_1243_),
    .ZN(_1245_)
  );
  AND2_X1 _2112_ (
    .A1(io_in1[2]),
    .A2(_1245_),
    .ZN(_1246_)
  );
  INV_X1 _2113_ (
    .A(_1246_),
    .ZN(_1247_)
  );
  AND2_X1 _2114_ (
    .A1(_0350_),
    .A2(io_in2[1]),
    .ZN(_1248_)
  );
  INV_X1 _2115_ (
    .A(_1248_),
    .ZN(_1249_)
  );
  AND2_X1 _2116_ (
    .A1(io_fn[3]),
    .A2(_0381_),
    .ZN(_1250_)
  );
  INV_X1 _2117_ (
    .A(_1250_),
    .ZN(_1251_)
  );
  AND2_X1 _2118_ (
    .A1(_1249_),
    .A2(_1251_),
    .ZN(_1252_)
  );
  INV_X1 _2119_ (
    .A(_1252_),
    .ZN(_1253_)
  );
  AND2_X1 _2120_ (
    .A1(io_in1[1]),
    .A2(_1253_),
    .ZN(_1254_)
  );
  INV_X1 _2121_ (
    .A(_1254_),
    .ZN(_1255_)
  );
  AND2_X1 _2122_ (
    .A1(_0350_),
    .A2(io_in2[0]),
    .ZN(_1256_)
  );
  INV_X1 _2123_ (
    .A(_1256_),
    .ZN(_1257_)
  );
  AND2_X1 _2124_ (
    .A1(io_fn[3]),
    .A2(_0370_),
    .ZN(_1258_)
  );
  INV_X1 _2125_ (
    .A(_1258_),
    .ZN(_1259_)
  );
  AND2_X1 _2126_ (
    .A1(_1257_),
    .A2(_1259_),
    .ZN(_1260_)
  );
  INV_X1 _2127_ (
    .A(_1260_),
    .ZN(_1261_)
  );
  AND2_X1 _2128_ (
    .A1(io_in1[0]),
    .A2(_1261_),
    .ZN(_1262_)
  );
  INV_X1 _2129_ (
    .A(_1262_),
    .ZN(_1263_)
  );
  AND2_X1 _2130_ (
    .A1(_0723_),
    .A2(_1252_),
    .ZN(_1264_)
  );
  INV_X1 _2131_ (
    .A(_1264_),
    .ZN(_1265_)
  );
  AND2_X1 _2132_ (
    .A1(_1255_),
    .A2(_1265_),
    .ZN(_1266_)
  );
  INV_X1 _2133_ (
    .A(_1266_),
    .ZN(_1267_)
  );
  AND2_X1 _2134_ (
    .A1(_1262_),
    .A2(_1266_),
    .ZN(_1268_)
  );
  INV_X1 _2135_ (
    .A(_1268_),
    .ZN(_1269_)
  );
  AND2_X1 _2136_ (
    .A1(_1255_),
    .A2(_1269_),
    .ZN(_1270_)
  );
  INV_X1 _2137_ (
    .A(_1270_),
    .ZN(_1271_)
  );
  AND2_X1 _2138_ (
    .A1(_0743_),
    .A2(_1244_),
    .ZN(_1272_)
  );
  INV_X1 _2139_ (
    .A(_1272_),
    .ZN(_1273_)
  );
  AND2_X1 _2140_ (
    .A1(_1247_),
    .A2(_1273_),
    .ZN(_1274_)
  );
  INV_X1 _2141_ (
    .A(_1274_),
    .ZN(_1275_)
  );
  AND2_X1 _2142_ (
    .A1(_1271_),
    .A2(_1274_),
    .ZN(_1276_)
  );
  INV_X1 _2143_ (
    .A(_1276_),
    .ZN(_1277_)
  );
  AND2_X1 _2144_ (
    .A1(_1247_),
    .A2(_1277_),
    .ZN(_1278_)
  );
  INV_X1 _2145_ (
    .A(_1278_),
    .ZN(_1279_)
  );
  AND2_X1 _2146_ (
    .A1(_0762_),
    .A2(_1232_),
    .ZN(_1280_)
  );
  INV_X1 _2147_ (
    .A(_1280_),
    .ZN(_1281_)
  );
  AND2_X1 _2148_ (
    .A1(_1235_),
    .A2(_1281_),
    .ZN(_1282_)
  );
  INV_X1 _2149_ (
    .A(_1282_),
    .ZN(_1283_)
  );
  AND2_X1 _2150_ (
    .A1(_1279_),
    .A2(_1282_),
    .ZN(_1284_)
  );
  INV_X1 _2151_ (
    .A(_1284_),
    .ZN(_1285_)
  );
  AND2_X1 _2152_ (
    .A1(_1235_),
    .A2(_1285_),
    .ZN(_1286_)
  );
  INV_X1 _2153_ (
    .A(_1286_),
    .ZN(_1287_)
  );
  AND2_X1 _2154_ (
    .A1(_0782_),
    .A2(_1220_),
    .ZN(_1288_)
  );
  INV_X1 _2155_ (
    .A(_1288_),
    .ZN(_1289_)
  );
  AND2_X1 _2156_ (
    .A1(_1223_),
    .A2(_1289_),
    .ZN(_1290_)
  );
  INV_X1 _2157_ (
    .A(_1290_),
    .ZN(_1291_)
  );
  AND2_X1 _2158_ (
    .A1(_1287_),
    .A2(_1290_),
    .ZN(_1292_)
  );
  INV_X1 _2159_ (
    .A(_1292_),
    .ZN(_1293_)
  );
  AND2_X1 _2160_ (
    .A1(_1223_),
    .A2(_1293_),
    .ZN(_1294_)
  );
  INV_X1 _2161_ (
    .A(_1294_),
    .ZN(_1295_)
  );
  AND2_X1 _2162_ (
    .A1(_0802_),
    .A2(_1208_),
    .ZN(_1296_)
  );
  INV_X1 _2163_ (
    .A(_1296_),
    .ZN(_1297_)
  );
  AND2_X1 _2164_ (
    .A1(_1211_),
    .A2(_1297_),
    .ZN(_1298_)
  );
  INV_X1 _2165_ (
    .A(_1298_),
    .ZN(_1299_)
  );
  AND2_X1 _2166_ (
    .A1(_1295_),
    .A2(_1298_),
    .ZN(_1300_)
  );
  INV_X1 _2167_ (
    .A(_1300_),
    .ZN(_1301_)
  );
  AND2_X1 _2168_ (
    .A1(_1211_),
    .A2(_1301_),
    .ZN(_1302_)
  );
  INV_X1 _2169_ (
    .A(_1302_),
    .ZN(_1303_)
  );
  AND2_X1 _2170_ (
    .A1(_1198_),
    .A2(_1303_),
    .ZN(_1304_)
  );
  INV_X1 _2171_ (
    .A(_1304_),
    .ZN(_1305_)
  );
  AND2_X1 _2172_ (
    .A1(_1195_),
    .A2(_1305_),
    .ZN(_1306_)
  );
  INV_X1 _2173_ (
    .A(_1306_),
    .ZN(_1307_)
  );
  AND2_X1 _2174_ (
    .A1(_1182_),
    .A2(_1307_),
    .ZN(_1308_)
  );
  INV_X1 _2175_ (
    .A(_1308_),
    .ZN(_1309_)
  );
  AND2_X1 _2176_ (
    .A1(_1179_),
    .A2(_1309_),
    .ZN(_1310_)
  );
  INV_X1 _2177_ (
    .A(_1310_),
    .ZN(_1311_)
  );
  AND2_X1 _2178_ (
    .A1(_0861_),
    .A2(_1164_),
    .ZN(_1312_)
  );
  INV_X1 _2179_ (
    .A(_1312_),
    .ZN(_1313_)
  );
  AND2_X1 _2180_ (
    .A1(_1167_),
    .A2(_1313_),
    .ZN(_1314_)
  );
  INV_X1 _2181_ (
    .A(_1314_),
    .ZN(_1315_)
  );
  AND2_X1 _2182_ (
    .A1(_1311_),
    .A2(_1314_),
    .ZN(_1316_)
  );
  INV_X1 _2183_ (
    .A(_1316_),
    .ZN(_1317_)
  );
  AND2_X1 _2184_ (
    .A1(_1167_),
    .A2(_1317_),
    .ZN(_1318_)
  );
  INV_X1 _2185_ (
    .A(_1318_),
    .ZN(_1319_)
  );
  AND2_X1 _2186_ (
    .A1(_1154_),
    .A2(_1319_),
    .ZN(_1320_)
  );
  INV_X1 _2187_ (
    .A(_1320_),
    .ZN(_1321_)
  );
  AND2_X1 _2188_ (
    .A1(_1151_),
    .A2(_1321_),
    .ZN(_1322_)
  );
  INV_X1 _2189_ (
    .A(_1322_),
    .ZN(_1323_)
  );
  AND2_X1 _2190_ (
    .A1(_1138_),
    .A2(_1323_),
    .ZN(_1324_)
  );
  INV_X1 _2191_ (
    .A(_1324_),
    .ZN(_1325_)
  );
  AND2_X1 _2192_ (
    .A1(_1122_),
    .A2(_1324_),
    .ZN(_1326_)
  );
  INV_X1 _2193_ (
    .A(_1326_),
    .ZN(_1327_)
  );
  AND2_X1 _2194_ (
    .A1(_1121_),
    .A2(_1134_),
    .ZN(_1328_)
  );
  INV_X1 _2195_ (
    .A(_1328_),
    .ZN(_1329_)
  );
  AND2_X1 _2196_ (
    .A1(_1119_),
    .A2(_1329_),
    .ZN(_1330_)
  );
  AND2_X1 _2197_ (
    .A1(_1327_),
    .A2(_1330_),
    .ZN(_1331_)
  );
  INV_X1 _2198_ (
    .A(_1331_),
    .ZN(_1332_)
  );
  AND2_X1 _2199_ (
    .A1(_1106_),
    .A2(_1332_),
    .ZN(_1333_)
  );
  INV_X1 _2200_ (
    .A(_1333_),
    .ZN(_1334_)
  );
  AND2_X1 _2201_ (
    .A1(_1090_),
    .A2(_1333_),
    .ZN(_1335_)
  );
  INV_X1 _2202_ (
    .A(_1335_),
    .ZN(_1336_)
  );
  AND2_X1 _2203_ (
    .A1(_1087_),
    .A2(_1103_),
    .ZN(_1337_)
  );
  INV_X1 _2204_ (
    .A(_1337_),
    .ZN(_1338_)
  );
  AND2_X1 _2205_ (
    .A1(_1089_),
    .A2(_1338_),
    .ZN(_1339_)
  );
  INV_X1 _2206_ (
    .A(_1339_),
    .ZN(_1340_)
  );
  AND2_X1 _2207_ (
    .A1(_1336_),
    .A2(_1340_),
    .ZN(_1341_)
  );
  INV_X1 _2208_ (
    .A(_1341_),
    .ZN(_1342_)
  );
  AND2_X1 _2209_ (
    .A1(_1074_),
    .A2(_1342_),
    .ZN(_1343_)
  );
  INV_X1 _2210_ (
    .A(_1343_),
    .ZN(_1344_)
  );
  AND2_X1 _2211_ (
    .A1(_1058_),
    .A2(_1343_),
    .ZN(_1345_)
  );
  INV_X1 _2212_ (
    .A(_1345_),
    .ZN(_1346_)
  );
  AND2_X1 _2213_ (
    .A1(_1057_),
    .A2(_1071_),
    .ZN(_1347_)
  );
  INV_X1 _2214_ (
    .A(_1347_),
    .ZN(_1348_)
  );
  AND2_X1 _2215_ (
    .A1(_1055_),
    .A2(_1348_),
    .ZN(_1349_)
  );
  INV_X1 _2216_ (
    .A(_1349_),
    .ZN(_1350_)
  );
  AND2_X1 _2217_ (
    .A1(_1346_),
    .A2(_1350_),
    .ZN(_1351_)
  );
  INV_X1 _2218_ (
    .A(_1351_),
    .ZN(_1352_)
  );
  AND2_X1 _2219_ (
    .A1(_0940_),
    .A2(_1040_),
    .ZN(_1353_)
  );
  INV_X1 _2220_ (
    .A(_1353_),
    .ZN(_1354_)
  );
  AND2_X1 _2221_ (
    .A1(_1043_),
    .A2(_1354_),
    .ZN(_1355_)
  );
  INV_X1 _2222_ (
    .A(_1355_),
    .ZN(_1356_)
  );
  AND2_X1 _2223_ (
    .A1(_1352_),
    .A2(_1355_),
    .ZN(_1357_)
  );
  INV_X1 _2224_ (
    .A(_1357_),
    .ZN(_1358_)
  );
  AND2_X1 _2225_ (
    .A1(_1043_),
    .A2(_1358_),
    .ZN(_1359_)
  );
  INV_X1 _2226_ (
    .A(_1359_),
    .ZN(_1360_)
  );
  AND2_X1 _2227_ (
    .A1(_0938_),
    .A2(_1028_),
    .ZN(_1361_)
  );
  INV_X1 _2228_ (
    .A(_1361_),
    .ZN(_1362_)
  );
  AND2_X1 _2229_ (
    .A1(_1031_),
    .A2(_1362_),
    .ZN(_1363_)
  );
  INV_X1 _2230_ (
    .A(_1363_),
    .ZN(_1364_)
  );
  AND2_X1 _2231_ (
    .A1(_1360_),
    .A2(_1363_),
    .ZN(_1365_)
  );
  INV_X1 _2232_ (
    .A(_1365_),
    .ZN(_1366_)
  );
  AND2_X1 _2233_ (
    .A1(_1031_),
    .A2(_1366_),
    .ZN(_1367_)
  );
  INV_X1 _2234_ (
    .A(_1367_),
    .ZN(_1368_)
  );
  AND2_X1 _2235_ (
    .A1(_1018_),
    .A2(_1368_),
    .ZN(_1369_)
  );
  INV_X1 _2236_ (
    .A(_1369_),
    .ZN(_1370_)
  );
  AND2_X1 _2237_ (
    .A1(_1015_),
    .A2(_1370_),
    .ZN(_1371_)
  );
  INV_X1 _2238_ (
    .A(_1371_),
    .ZN(_1372_)
  );
  AND2_X1 _2239_ (
    .A1(_1002_),
    .A2(_1372_),
    .ZN(_1373_)
  );
  INV_X1 _2240_ (
    .A(_1373_),
    .ZN(_1374_)
  );
  AND2_X1 _2241_ (
    .A1(_0999_),
    .A2(_1374_),
    .ZN(_1375_)
  );
  INV_X1 _2242_ (
    .A(_1375_),
    .ZN(_1376_)
  );
  AND2_X1 _2243_ (
    .A1(_0986_),
    .A2(_1376_),
    .ZN(_1377_)
  );
  INV_X1 _2244_ (
    .A(_1377_),
    .ZN(_1378_)
  );
  AND2_X1 _2245_ (
    .A1(_0983_),
    .A2(_1378_),
    .ZN(_1379_)
  );
  INV_X1 _2246_ (
    .A(_1379_),
    .ZN(_1380_)
  );
  AND2_X1 _2247_ (
    .A1(_0971_),
    .A2(_1380_),
    .ZN(_1381_)
  );
  INV_X1 _2248_ (
    .A(_1381_),
    .ZN(_1382_)
  );
  AND2_X1 _2249_ (
    .A1(_0969_),
    .A2(_1379_),
    .ZN(_1383_)
  );
  INV_X1 _2250_ (
    .A(_1383_),
    .ZN(_1384_)
  );
  AND2_X1 _2251_ (
    .A1(_0969_),
    .A2(_1382_),
    .ZN(_1385_)
  );
  AND2_X1 _2252_ (
    .A1(_0971_),
    .A2(_1384_),
    .ZN(_1386_)
  );
  AND2_X1 _2253_ (
    .A1(_0956_),
    .A2(_1386_),
    .ZN(_1387_)
  );
  INV_X1 _2254_ (
    .A(_1387_),
    .ZN(_1388_)
  );
  AND2_X1 _2255_ (
    .A1(_0957_),
    .A2(_1385_),
    .ZN(_1389_)
  );
  INV_X1 _2256_ (
    .A(_1389_),
    .ZN(_1390_)
  );
  AND2_X1 _2257_ (
    .A1(_1388_),
    .A2(_1390_),
    .ZN(_1391_)
  );
  INV_X1 _2258_ (
    .A(_1391_),
    .ZN(_1392_)
  );
  AND2_X1 _2259_ (
    .A1(_0987_),
    .A2(_1375_),
    .ZN(_1393_)
  );
  INV_X1 _2260_ (
    .A(_1393_),
    .ZN(_1394_)
  );
  AND2_X1 _2261_ (
    .A1(_1378_),
    .A2(_1394_),
    .ZN(_1395_)
  );
  INV_X1 _2262_ (
    .A(_1395_),
    .ZN(_1396_)
  );
  AND2_X1 _2263_ (
    .A1(_1359_),
    .A2(_1364_),
    .ZN(_1397_)
  );
  INV_X1 _2264_ (
    .A(_1397_),
    .ZN(_1398_)
  );
  AND2_X1 _2265_ (
    .A1(_1366_),
    .A2(_1398_),
    .ZN(_1399_)
  );
  INV_X1 _2266_ (
    .A(_1399_),
    .ZN(_1400_)
  );
  AND2_X1 _2267_ (
    .A1(_1351_),
    .A2(_1356_),
    .ZN(_1401_)
  );
  INV_X1 _2268_ (
    .A(_1401_),
    .ZN(_1402_)
  );
  AND2_X1 _2269_ (
    .A1(_1358_),
    .A2(_1402_),
    .ZN(_1403_)
  );
  INV_X1 _2270_ (
    .A(_1403_),
    .ZN(_1404_)
  );
  AND2_X1 _2271_ (
    .A1(_1075_),
    .A2(_1341_),
    .ZN(_1405_)
  );
  INV_X1 _2272_ (
    .A(_1405_),
    .ZN(_1406_)
  );
  AND2_X1 _2273_ (
    .A1(_1344_),
    .A2(_1406_),
    .ZN(_1407_)
  );
  INV_X1 _2274_ (
    .A(_1407_),
    .ZN(_1408_)
  );
  AND2_X1 _2275_ (
    .A1(_1310_),
    .A2(_1315_),
    .ZN(_1409_)
  );
  INV_X1 _2276_ (
    .A(_1409_),
    .ZN(_1410_)
  );
  AND2_X1 _2277_ (
    .A1(_1317_),
    .A2(_1410_),
    .ZN(_1411_)
  );
  INV_X1 _2278_ (
    .A(_1411_),
    .ZN(_1412_)
  );
  AND2_X1 _2279_ (
    .A1(_0703_),
    .A2(_1260_),
    .ZN(_1413_)
  );
  INV_X1 _2280_ (
    .A(_1413_),
    .ZN(_1414_)
  );
  AND2_X1 _2281_ (
    .A1(_1263_),
    .A2(_1414_),
    .ZN(_1415_)
  );
  INV_X1 _2282_ (
    .A(_1415_),
    .ZN(_1416_)
  );
  AND2_X1 _2283_ (
    .A1(io_fn[3]),
    .A2(_1415_),
    .ZN(_1417_)
  );
  INV_X1 _2284_ (
    .A(_1417_),
    .ZN(_1418_)
  );
  AND2_X1 _2285_ (
    .A1(_1266_),
    .A2(_1417_),
    .ZN(_1419_)
  );
  INV_X1 _2286_ (
    .A(_1419_),
    .ZN(_1420_)
  );
  AND2_X1 _2287_ (
    .A1(_1270_),
    .A2(_1275_),
    .ZN(_1421_)
  );
  INV_X1 _2288_ (
    .A(_1421_),
    .ZN(_1422_)
  );
  AND2_X1 _2289_ (
    .A1(_1277_),
    .A2(_1422_),
    .ZN(_1423_)
  );
  INV_X1 _2290_ (
    .A(_1423_),
    .ZN(_1424_)
  );
  AND2_X1 _2291_ (
    .A1(_1419_),
    .A2(_1423_),
    .ZN(_1425_)
  );
  INV_X1 _2292_ (
    .A(_1425_),
    .ZN(_1426_)
  );
  AND2_X1 _2293_ (
    .A1(_1278_),
    .A2(_1283_),
    .ZN(_1427_)
  );
  INV_X1 _2294_ (
    .A(_1427_),
    .ZN(_1428_)
  );
  AND2_X1 _2295_ (
    .A1(_1285_),
    .A2(_1428_),
    .ZN(_1429_)
  );
  INV_X1 _2296_ (
    .A(_1429_),
    .ZN(_1430_)
  );
  AND2_X1 _2297_ (
    .A1(_1425_),
    .A2(_1429_),
    .ZN(_1431_)
  );
  INV_X1 _2298_ (
    .A(_1431_),
    .ZN(_1432_)
  );
  AND2_X1 _2299_ (
    .A1(_1286_),
    .A2(_1291_),
    .ZN(_1433_)
  );
  INV_X1 _2300_ (
    .A(_1433_),
    .ZN(_1434_)
  );
  AND2_X1 _2301_ (
    .A1(_1293_),
    .A2(_1434_),
    .ZN(_1435_)
  );
  INV_X1 _2302_ (
    .A(_1435_),
    .ZN(_1436_)
  );
  AND2_X1 _2303_ (
    .A1(_1431_),
    .A2(_1435_),
    .ZN(_1437_)
  );
  INV_X1 _2304_ (
    .A(_1437_),
    .ZN(_1438_)
  );
  AND2_X1 _2305_ (
    .A1(_1294_),
    .A2(_1299_),
    .ZN(_1439_)
  );
  INV_X1 _2306_ (
    .A(_1439_),
    .ZN(_1440_)
  );
  AND2_X1 _2307_ (
    .A1(_1301_),
    .A2(_1440_),
    .ZN(_1441_)
  );
  INV_X1 _2308_ (
    .A(_1441_),
    .ZN(_1442_)
  );
  AND2_X1 _2309_ (
    .A1(_1437_),
    .A2(_1441_),
    .ZN(_1443_)
  );
  INV_X1 _2310_ (
    .A(_1443_),
    .ZN(_1444_)
  );
  AND2_X1 _2311_ (
    .A1(_1199_),
    .A2(_1302_),
    .ZN(_1445_)
  );
  INV_X1 _2312_ (
    .A(_1445_),
    .ZN(_1446_)
  );
  AND2_X1 _2313_ (
    .A1(_1305_),
    .A2(_1446_),
    .ZN(_1447_)
  );
  INV_X1 _2314_ (
    .A(_1447_),
    .ZN(_1448_)
  );
  AND2_X1 _2315_ (
    .A1(_1443_),
    .A2(_1447_),
    .ZN(_1449_)
  );
  INV_X1 _2316_ (
    .A(_1449_),
    .ZN(_1450_)
  );
  AND2_X1 _2317_ (
    .A1(_1183_),
    .A2(_1306_),
    .ZN(_1451_)
  );
  INV_X1 _2318_ (
    .A(_1451_),
    .ZN(_1452_)
  );
  AND2_X1 _2319_ (
    .A1(_1309_),
    .A2(_1452_),
    .ZN(_1453_)
  );
  INV_X1 _2320_ (
    .A(_1453_),
    .ZN(_1454_)
  );
  AND2_X1 _2321_ (
    .A1(_1449_),
    .A2(_1453_),
    .ZN(_1455_)
  );
  INV_X1 _2322_ (
    .A(_1455_),
    .ZN(_1456_)
  );
  AND2_X1 _2323_ (
    .A1(_1411_),
    .A2(_1455_),
    .ZN(_1457_)
  );
  INV_X1 _2324_ (
    .A(_1457_),
    .ZN(_1458_)
  );
  AND2_X1 _2325_ (
    .A1(_1155_),
    .A2(_1318_),
    .ZN(_1459_)
  );
  INV_X1 _2326_ (
    .A(_1459_),
    .ZN(_1460_)
  );
  AND2_X1 _2327_ (
    .A1(_1321_),
    .A2(_1460_),
    .ZN(_1461_)
  );
  INV_X1 _2328_ (
    .A(_1461_),
    .ZN(_1462_)
  );
  AND2_X1 _2329_ (
    .A1(_1457_),
    .A2(_1461_),
    .ZN(_1463_)
  );
  INV_X1 _2330_ (
    .A(_1463_),
    .ZN(_1464_)
  );
  AND2_X1 _2331_ (
    .A1(_1139_),
    .A2(_1322_),
    .ZN(_1465_)
  );
  INV_X1 _2332_ (
    .A(_1465_),
    .ZN(_1466_)
  );
  AND2_X1 _2333_ (
    .A1(_1325_),
    .A2(_1466_),
    .ZN(_1467_)
  );
  INV_X1 _2334_ (
    .A(_1467_),
    .ZN(_1468_)
  );
  AND2_X1 _2335_ (
    .A1(_1463_),
    .A2(_1467_),
    .ZN(_1469_)
  );
  INV_X1 _2336_ (
    .A(_1469_),
    .ZN(_1470_)
  );
  AND2_X1 _2337_ (
    .A1(_1135_),
    .A2(_1325_),
    .ZN(_1471_)
  );
  INV_X1 _2338_ (
    .A(_1471_),
    .ZN(_1472_)
  );
  AND2_X1 _2339_ (
    .A1(_1122_),
    .A2(_1471_),
    .ZN(_1473_)
  );
  INV_X1 _2340_ (
    .A(_1473_),
    .ZN(_1474_)
  );
  AND2_X1 _2341_ (
    .A1(_1123_),
    .A2(_1472_),
    .ZN(_1475_)
  );
  INV_X1 _2342_ (
    .A(_1475_),
    .ZN(_1476_)
  );
  AND2_X1 _2343_ (
    .A1(_1123_),
    .A2(_1471_),
    .ZN(_1477_)
  );
  INV_X1 _2344_ (
    .A(_1477_),
    .ZN(_1478_)
  );
  AND2_X1 _2345_ (
    .A1(_1122_),
    .A2(_1472_),
    .ZN(_1479_)
  );
  INV_X1 _2346_ (
    .A(_1479_),
    .ZN(_1480_)
  );
  AND2_X1 _2347_ (
    .A1(_1474_),
    .A2(_1476_),
    .ZN(_1481_)
  );
  AND2_X1 _2348_ (
    .A1(_1478_),
    .A2(_1480_),
    .ZN(_1482_)
  );
  AND2_X1 _2349_ (
    .A1(_1469_),
    .A2(_1482_),
    .ZN(_1483_)
  );
  INV_X1 _2350_ (
    .A(_1483_),
    .ZN(_1484_)
  );
  AND2_X1 _2351_ (
    .A1(_1107_),
    .A2(_1331_),
    .ZN(_1485_)
  );
  INV_X1 _2352_ (
    .A(_1485_),
    .ZN(_1486_)
  );
  AND2_X1 _2353_ (
    .A1(_1334_),
    .A2(_1486_),
    .ZN(_1487_)
  );
  INV_X1 _2354_ (
    .A(_1487_),
    .ZN(_1488_)
  );
  AND2_X1 _2355_ (
    .A1(_1483_),
    .A2(_1487_),
    .ZN(_1489_)
  );
  INV_X1 _2356_ (
    .A(_1489_),
    .ZN(_1490_)
  );
  AND2_X1 _2357_ (
    .A1(_1103_),
    .A2(_1334_),
    .ZN(_1491_)
  );
  INV_X1 _2358_ (
    .A(_1491_),
    .ZN(_1492_)
  );
  AND2_X1 _2359_ (
    .A1(_1090_),
    .A2(_1491_),
    .ZN(_1493_)
  );
  INV_X1 _2360_ (
    .A(_1493_),
    .ZN(_1494_)
  );
  AND2_X1 _2361_ (
    .A1(_1091_),
    .A2(_1492_),
    .ZN(_1495_)
  );
  INV_X1 _2362_ (
    .A(_1495_),
    .ZN(_1496_)
  );
  AND2_X1 _2363_ (
    .A1(_1091_),
    .A2(_1491_),
    .ZN(_1497_)
  );
  INV_X1 _2364_ (
    .A(_1497_),
    .ZN(_1498_)
  );
  AND2_X1 _2365_ (
    .A1(_1090_),
    .A2(_1492_),
    .ZN(_1499_)
  );
  INV_X1 _2366_ (
    .A(_1499_),
    .ZN(_1500_)
  );
  AND2_X1 _2367_ (
    .A1(_1494_),
    .A2(_1496_),
    .ZN(_1501_)
  );
  AND2_X1 _2368_ (
    .A1(_1498_),
    .A2(_1500_),
    .ZN(_1502_)
  );
  AND2_X1 _2369_ (
    .A1(_1489_),
    .A2(_1502_),
    .ZN(_1503_)
  );
  INV_X1 _2370_ (
    .A(_1503_),
    .ZN(_1504_)
  );
  AND2_X1 _2371_ (
    .A1(_1407_),
    .A2(_1503_),
    .ZN(_1505_)
  );
  INV_X1 _2372_ (
    .A(_1505_),
    .ZN(_1506_)
  );
  AND2_X1 _2373_ (
    .A1(_1071_),
    .A2(_1344_),
    .ZN(_1507_)
  );
  INV_X1 _2374_ (
    .A(_1507_),
    .ZN(_1508_)
  );
  AND2_X1 _2375_ (
    .A1(_1058_),
    .A2(_1507_),
    .ZN(_1509_)
  );
  INV_X1 _2376_ (
    .A(_1509_),
    .ZN(_1510_)
  );
  AND2_X1 _2377_ (
    .A1(_1059_),
    .A2(_1508_),
    .ZN(_1511_)
  );
  INV_X1 _2378_ (
    .A(_1511_),
    .ZN(_1512_)
  );
  AND2_X1 _2379_ (
    .A1(_1059_),
    .A2(_1507_),
    .ZN(_1513_)
  );
  INV_X1 _2380_ (
    .A(_1513_),
    .ZN(_1514_)
  );
  AND2_X1 _2381_ (
    .A1(_1058_),
    .A2(_1508_),
    .ZN(_1515_)
  );
  INV_X1 _2382_ (
    .A(_1515_),
    .ZN(_1516_)
  );
  AND2_X1 _2383_ (
    .A1(_1510_),
    .A2(_1512_),
    .ZN(_1517_)
  );
  AND2_X1 _2384_ (
    .A1(_1514_),
    .A2(_1516_),
    .ZN(_1518_)
  );
  AND2_X1 _2385_ (
    .A1(_1505_),
    .A2(_1518_),
    .ZN(_1519_)
  );
  INV_X1 _2386_ (
    .A(_1519_),
    .ZN(_1520_)
  );
  AND2_X1 _2387_ (
    .A1(_1403_),
    .A2(_1519_),
    .ZN(_1521_)
  );
  INV_X1 _2388_ (
    .A(_1521_),
    .ZN(_1522_)
  );
  AND2_X1 _2389_ (
    .A1(_1399_),
    .A2(_1521_),
    .ZN(_1523_)
  );
  INV_X1 _2390_ (
    .A(_1523_),
    .ZN(_1524_)
  );
  AND2_X1 _2391_ (
    .A1(_1019_),
    .A2(_1367_),
    .ZN(_1525_)
  );
  INV_X1 _2392_ (
    .A(_1525_),
    .ZN(_1526_)
  );
  AND2_X1 _2393_ (
    .A1(_1370_),
    .A2(_1526_),
    .ZN(_1527_)
  );
  INV_X1 _2394_ (
    .A(_1527_),
    .ZN(_1528_)
  );
  AND2_X1 _2395_ (
    .A1(_1523_),
    .A2(_1527_),
    .ZN(_1529_)
  );
  INV_X1 _2396_ (
    .A(_1529_),
    .ZN(_1530_)
  );
  AND2_X1 _2397_ (
    .A1(_1003_),
    .A2(_1371_),
    .ZN(_1531_)
  );
  INV_X1 _2398_ (
    .A(_1531_),
    .ZN(_1532_)
  );
  AND2_X1 _2399_ (
    .A1(_1374_),
    .A2(_1532_),
    .ZN(_1533_)
  );
  INV_X1 _2400_ (
    .A(_1533_),
    .ZN(_1534_)
  );
  AND2_X1 _2401_ (
    .A1(_1529_),
    .A2(_1533_),
    .ZN(_1535_)
  );
  INV_X1 _2402_ (
    .A(_1535_),
    .ZN(_1536_)
  );
  AND2_X1 _2403_ (
    .A1(_1395_),
    .A2(_1535_),
    .ZN(_1537_)
  );
  INV_X1 _2404_ (
    .A(_1537_),
    .ZN(_1538_)
  );
  AND2_X1 _2405_ (
    .A1(_0969_),
    .A2(_0971_),
    .ZN(_1539_)
  );
  INV_X1 _2406_ (
    .A(_1539_),
    .ZN(_1540_)
  );
  AND2_X1 _2407_ (
    .A1(_1380_),
    .A2(_1540_),
    .ZN(_1541_)
  );
  INV_X1 _2408_ (
    .A(_1541_),
    .ZN(_1542_)
  );
  AND2_X1 _2409_ (
    .A1(_1379_),
    .A2(_1539_),
    .ZN(_1543_)
  );
  INV_X1 _2410_ (
    .A(_1543_),
    .ZN(_1544_)
  );
  AND2_X1 _2411_ (
    .A1(_1379_),
    .A2(_1540_),
    .ZN(_1545_)
  );
  INV_X1 _2412_ (
    .A(_1545_),
    .ZN(_1546_)
  );
  AND2_X1 _2413_ (
    .A1(_1380_),
    .A2(_1539_),
    .ZN(_1547_)
  );
  INV_X1 _2414_ (
    .A(_1547_),
    .ZN(_1548_)
  );
  AND2_X1 _2415_ (
    .A1(_1542_),
    .A2(_1544_),
    .ZN(_1549_)
  );
  AND2_X1 _2416_ (
    .A1(_1546_),
    .A2(_1548_),
    .ZN(_1550_)
  );
  AND2_X1 _2417_ (
    .A1(_1537_),
    .A2(_1550_),
    .ZN(_1551_)
  );
  INV_X1 _2418_ (
    .A(_1551_),
    .ZN(_1552_)
  );
  AND2_X1 _2419_ (
    .A1(_1391_),
    .A2(_1551_),
    .ZN(_1553_)
  );
  INV_X1 _2420_ (
    .A(_1553_),
    .ZN(_1554_)
  );
  AND2_X1 _2421_ (
    .A1(io_fn[3]),
    .A2(_0603_),
    .ZN(_1555_)
  );
  INV_X1 _2422_ (
    .A(_1555_),
    .ZN(_1556_)
  );
  AND2_X1 _2423_ (
    .A1(_0350_),
    .A2(io_in2[23]),
    .ZN(_1557_)
  );
  INV_X1 _2424_ (
    .A(_1557_),
    .ZN(_1558_)
  );
  AND2_X1 _2425_ (
    .A1(_0350_),
    .A2(_0603_),
    .ZN(_1559_)
  );
  INV_X1 _2426_ (
    .A(_1559_),
    .ZN(_1560_)
  );
  AND2_X1 _2427_ (
    .A1(io_fn[3]),
    .A2(io_in2[23]),
    .ZN(_1561_)
  );
  INV_X1 _2428_ (
    .A(_1561_),
    .ZN(_1562_)
  );
  AND2_X1 _2429_ (
    .A1(_1556_),
    .A2(_1558_),
    .ZN(_1563_)
  );
  AND2_X1 _2430_ (
    .A1(_1560_),
    .A2(_1562_),
    .ZN(_1564_)
  );
  AND2_X1 _2431_ (
    .A1(io_in1[23]),
    .A2(_1564_),
    .ZN(_1565_)
  );
  INV_X1 _2432_ (
    .A(_1565_),
    .ZN(_1566_)
  );
  AND2_X1 _2433_ (
    .A1(_0852_),
    .A2(_1563_),
    .ZN(_1567_)
  );
  INV_X1 _2434_ (
    .A(_1567_),
    .ZN(_1568_)
  );
  AND2_X1 _2435_ (
    .A1(_1566_),
    .A2(_1568_),
    .ZN(_1569_)
  );
  INV_X1 _2436_ (
    .A(_1569_),
    .ZN(_1570_)
  );
  AND2_X1 _2437_ (
    .A1(_0953_),
    .A2(_1388_),
    .ZN(_1571_)
  );
  INV_X1 _2438_ (
    .A(_1571_),
    .ZN(_1572_)
  );
  AND2_X1 _2439_ (
    .A1(_1569_),
    .A2(_1572_),
    .ZN(_1573_)
  );
  INV_X1 _2440_ (
    .A(_1573_),
    .ZN(_1574_)
  );
  AND2_X1 _2441_ (
    .A1(_1570_),
    .A2(_1571_),
    .ZN(_1575_)
  );
  INV_X1 _2442_ (
    .A(_1575_),
    .ZN(_1576_)
  );
  AND2_X1 _2443_ (
    .A1(_1569_),
    .A2(_1571_),
    .ZN(_1577_)
  );
  INV_X1 _2444_ (
    .A(_1577_),
    .ZN(_1578_)
  );
  AND2_X1 _2445_ (
    .A1(_1570_),
    .A2(_1572_),
    .ZN(_1579_)
  );
  INV_X1 _2446_ (
    .A(_1579_),
    .ZN(_1580_)
  );
  AND2_X1 _2447_ (
    .A1(_1574_),
    .A2(_1576_),
    .ZN(_1581_)
  );
  AND2_X1 _2448_ (
    .A1(_1578_),
    .A2(_1580_),
    .ZN(_1582_)
  );
  AND2_X1 _2449_ (
    .A1(_1553_),
    .A2(_1581_),
    .ZN(_1583_)
  );
  INV_X1 _2450_ (
    .A(_1583_),
    .ZN(_1584_)
  );
  AND2_X1 _2451_ (
    .A1(io_fn[3]),
    .A2(_0613_),
    .ZN(_1585_)
  );
  INV_X1 _2452_ (
    .A(_1585_),
    .ZN(_1586_)
  );
  AND2_X1 _2453_ (
    .A1(_0350_),
    .A2(io_in2[24]),
    .ZN(_1587_)
  );
  INV_X1 _2454_ (
    .A(_1587_),
    .ZN(_1588_)
  );
  AND2_X1 _2455_ (
    .A1(_0350_),
    .A2(_0613_),
    .ZN(_1589_)
  );
  INV_X1 _2456_ (
    .A(_1589_),
    .ZN(_1590_)
  );
  AND2_X1 _2457_ (
    .A1(io_fn[3]),
    .A2(io_in2[24]),
    .ZN(_1591_)
  );
  INV_X1 _2458_ (
    .A(_1591_),
    .ZN(_1592_)
  );
  AND2_X1 _2459_ (
    .A1(_1586_),
    .A2(_1588_),
    .ZN(_1593_)
  );
  AND2_X1 _2460_ (
    .A1(_1590_),
    .A2(_1592_),
    .ZN(_1594_)
  );
  AND2_X1 _2461_ (
    .A1(io_in1[24]),
    .A2(_1594_),
    .ZN(_1595_)
  );
  INV_X1 _2462_ (
    .A(_1595_),
    .ZN(_1596_)
  );
  AND2_X1 _2463_ (
    .A1(_0832_),
    .A2(_1593_),
    .ZN(_1597_)
  );
  INV_X1 _2464_ (
    .A(_1597_),
    .ZN(_1598_)
  );
  AND2_X1 _2465_ (
    .A1(_1596_),
    .A2(_1598_),
    .ZN(_1599_)
  );
  INV_X1 _2466_ (
    .A(_1599_),
    .ZN(_1600_)
  );
  AND2_X1 _2467_ (
    .A1(_1568_),
    .A2(_1572_),
    .ZN(_1601_)
  );
  INV_X1 _2468_ (
    .A(_1601_),
    .ZN(_1602_)
  );
  AND2_X1 _2469_ (
    .A1(_1566_),
    .A2(_1571_),
    .ZN(_1603_)
  );
  INV_X1 _2470_ (
    .A(_1603_),
    .ZN(_1604_)
  );
  AND2_X1 _2471_ (
    .A1(_1566_),
    .A2(_1602_),
    .ZN(_1605_)
  );
  AND2_X1 _2472_ (
    .A1(_1568_),
    .A2(_1604_),
    .ZN(_1606_)
  );
  AND2_X1 _2473_ (
    .A1(_1599_),
    .A2(_1606_),
    .ZN(_1607_)
  );
  INV_X1 _2474_ (
    .A(_1607_),
    .ZN(_1608_)
  );
  AND2_X1 _2475_ (
    .A1(_1600_),
    .A2(_1605_),
    .ZN(_1609_)
  );
  INV_X1 _2476_ (
    .A(_1609_),
    .ZN(_1610_)
  );
  AND2_X1 _2477_ (
    .A1(_1608_),
    .A2(_1610_),
    .ZN(_1611_)
  );
  INV_X1 _2478_ (
    .A(_1611_),
    .ZN(_1612_)
  );
  AND2_X1 _2479_ (
    .A1(_1583_),
    .A2(_1611_),
    .ZN(_1613_)
  );
  INV_X1 _2480_ (
    .A(_1613_),
    .ZN(_1614_)
  );
  AND2_X1 _2481_ (
    .A1(io_fn[3]),
    .A2(_0623_),
    .ZN(_1615_)
  );
  INV_X1 _2482_ (
    .A(_1615_),
    .ZN(_1616_)
  );
  AND2_X1 _2483_ (
    .A1(_0350_),
    .A2(io_in2[25]),
    .ZN(_1617_)
  );
  INV_X1 _2484_ (
    .A(_1617_),
    .ZN(_1618_)
  );
  AND2_X1 _2485_ (
    .A1(_0350_),
    .A2(_0623_),
    .ZN(_1619_)
  );
  INV_X1 _2486_ (
    .A(_1619_),
    .ZN(_1620_)
  );
  AND2_X1 _2487_ (
    .A1(io_fn[3]),
    .A2(io_in2[25]),
    .ZN(_1621_)
  );
  INV_X1 _2488_ (
    .A(_1621_),
    .ZN(_1622_)
  );
  AND2_X1 _2489_ (
    .A1(_1616_),
    .A2(_1618_),
    .ZN(_1623_)
  );
  AND2_X1 _2490_ (
    .A1(_1620_),
    .A2(_1622_),
    .ZN(_1624_)
  );
  AND2_X1 _2491_ (
    .A1(io_in1[25]),
    .A2(_1624_),
    .ZN(_1625_)
  );
  INV_X1 _2492_ (
    .A(_1625_),
    .ZN(_1626_)
  );
  AND2_X1 _2493_ (
    .A1(_0812_),
    .A2(_1623_),
    .ZN(_1627_)
  );
  INV_X1 _2494_ (
    .A(_1627_),
    .ZN(_1628_)
  );
  AND2_X1 _2495_ (
    .A1(_1626_),
    .A2(_1628_),
    .ZN(_1629_)
  );
  INV_X1 _2496_ (
    .A(_1629_),
    .ZN(_1630_)
  );
  AND2_X1 _2497_ (
    .A1(_1596_),
    .A2(_1608_),
    .ZN(_1631_)
  );
  INV_X1 _2498_ (
    .A(_1631_),
    .ZN(_1632_)
  );
  AND2_X1 _2499_ (
    .A1(_1629_),
    .A2(_1632_),
    .ZN(_1633_)
  );
  INV_X1 _2500_ (
    .A(_1633_),
    .ZN(_1634_)
  );
  AND2_X1 _2501_ (
    .A1(_1630_),
    .A2(_1631_),
    .ZN(_1635_)
  );
  INV_X1 _2502_ (
    .A(_1635_),
    .ZN(_1636_)
  );
  AND2_X1 _2503_ (
    .A1(_1634_),
    .A2(_1636_),
    .ZN(_1637_)
  );
  INV_X1 _2504_ (
    .A(_1637_),
    .ZN(_1638_)
  );
  AND2_X1 _2505_ (
    .A1(_1613_),
    .A2(_1637_),
    .ZN(_1639_)
  );
  INV_X1 _2506_ (
    .A(_1639_),
    .ZN(_1640_)
  );
  AND2_X1 _2507_ (
    .A1(io_fn[3]),
    .A2(_0632_),
    .ZN(_1641_)
  );
  INV_X1 _2508_ (
    .A(_1641_),
    .ZN(_1642_)
  );
  AND2_X1 _2509_ (
    .A1(_0350_),
    .A2(io_in2[26]),
    .ZN(_1643_)
  );
  INV_X1 _2510_ (
    .A(_1643_),
    .ZN(_1644_)
  );
  AND2_X1 _2511_ (
    .A1(_0350_),
    .A2(_0632_),
    .ZN(_1645_)
  );
  INV_X1 _2512_ (
    .A(_1645_),
    .ZN(_1646_)
  );
  AND2_X1 _2513_ (
    .A1(io_fn[3]),
    .A2(io_in2[26]),
    .ZN(_1647_)
  );
  INV_X1 _2514_ (
    .A(_1647_),
    .ZN(_1648_)
  );
  AND2_X1 _2515_ (
    .A1(_1642_),
    .A2(_1644_),
    .ZN(_1649_)
  );
  AND2_X1 _2516_ (
    .A1(_1646_),
    .A2(_1648_),
    .ZN(_1650_)
  );
  AND2_X1 _2517_ (
    .A1(io_in1[26]),
    .A2(_1650_),
    .ZN(_1651_)
  );
  INV_X1 _2518_ (
    .A(_1651_),
    .ZN(_1652_)
  );
  AND2_X1 _2519_ (
    .A1(_0792_),
    .A2(_1649_),
    .ZN(_1653_)
  );
  INV_X1 _2520_ (
    .A(_1653_),
    .ZN(_1654_)
  );
  AND2_X1 _2521_ (
    .A1(_1652_),
    .A2(_1654_),
    .ZN(_1655_)
  );
  INV_X1 _2522_ (
    .A(_1655_),
    .ZN(_1656_)
  );
  AND2_X1 _2523_ (
    .A1(_1626_),
    .A2(_1634_),
    .ZN(_1657_)
  );
  INV_X1 _2524_ (
    .A(_1657_),
    .ZN(_1658_)
  );
  AND2_X1 _2525_ (
    .A1(_1655_),
    .A2(_1658_),
    .ZN(_1659_)
  );
  INV_X1 _2526_ (
    .A(_1659_),
    .ZN(_1660_)
  );
  AND2_X1 _2527_ (
    .A1(_1656_),
    .A2(_1657_),
    .ZN(_1661_)
  );
  INV_X1 _2528_ (
    .A(_1661_),
    .ZN(_1662_)
  );
  AND2_X1 _2529_ (
    .A1(_1660_),
    .A2(_1662_),
    .ZN(_1663_)
  );
  INV_X1 _2530_ (
    .A(_1663_),
    .ZN(_1664_)
  );
  AND2_X1 _2531_ (
    .A1(_1639_),
    .A2(_1663_),
    .ZN(_1665_)
  );
  INV_X1 _2532_ (
    .A(_1665_),
    .ZN(_1666_)
  );
  AND2_X1 _2533_ (
    .A1(io_fn[3]),
    .A2(_0643_),
    .ZN(_1667_)
  );
  INV_X1 _2534_ (
    .A(_1667_),
    .ZN(_1668_)
  );
  AND2_X1 _2535_ (
    .A1(_0350_),
    .A2(io_in2[27]),
    .ZN(_1669_)
  );
  INV_X1 _2536_ (
    .A(_1669_),
    .ZN(_1670_)
  );
  AND2_X1 _2537_ (
    .A1(_0350_),
    .A2(_0643_),
    .ZN(_1671_)
  );
  INV_X1 _2538_ (
    .A(_1671_),
    .ZN(_1672_)
  );
  AND2_X1 _2539_ (
    .A1(io_fn[3]),
    .A2(io_in2[27]),
    .ZN(_1673_)
  );
  INV_X1 _2540_ (
    .A(_1673_),
    .ZN(_1674_)
  );
  AND2_X1 _2541_ (
    .A1(_1668_),
    .A2(_1670_),
    .ZN(_1675_)
  );
  AND2_X1 _2542_ (
    .A1(_1672_),
    .A2(_1674_),
    .ZN(_1676_)
  );
  AND2_X1 _2543_ (
    .A1(io_in1[27]),
    .A2(_1676_),
    .ZN(_1677_)
  );
  INV_X1 _2544_ (
    .A(_1677_),
    .ZN(_1678_)
  );
  AND2_X1 _2545_ (
    .A1(_0772_),
    .A2(_1675_),
    .ZN(_1679_)
  );
  INV_X1 _2546_ (
    .A(_1679_),
    .ZN(_1680_)
  );
  AND2_X1 _2547_ (
    .A1(_1678_),
    .A2(_1680_),
    .ZN(_1681_)
  );
  INV_X1 _2548_ (
    .A(_1681_),
    .ZN(_1682_)
  );
  AND2_X1 _2549_ (
    .A1(_1652_),
    .A2(_1660_),
    .ZN(_1683_)
  );
  INV_X1 _2550_ (
    .A(_1683_),
    .ZN(_1684_)
  );
  AND2_X1 _2551_ (
    .A1(_1681_),
    .A2(_1684_),
    .ZN(_1685_)
  );
  INV_X1 _2552_ (
    .A(_1685_),
    .ZN(_1686_)
  );
  AND2_X1 _2553_ (
    .A1(_1682_),
    .A2(_1683_),
    .ZN(_1687_)
  );
  INV_X1 _2554_ (
    .A(_1687_),
    .ZN(_1688_)
  );
  AND2_X1 _2555_ (
    .A1(_1686_),
    .A2(_1688_),
    .ZN(_1689_)
  );
  INV_X1 _2556_ (
    .A(_1689_),
    .ZN(_1690_)
  );
  AND2_X1 _2557_ (
    .A1(_1665_),
    .A2(_1689_),
    .ZN(_1691_)
  );
  INV_X1 _2558_ (
    .A(_1691_),
    .ZN(_1692_)
  );
  AND2_X1 _2559_ (
    .A1(_1678_),
    .A2(_1686_),
    .ZN(_1693_)
  );
  INV_X1 _2560_ (
    .A(_1693_),
    .ZN(_1694_)
  );
  AND2_X1 _2561_ (
    .A1(io_fn[3]),
    .A2(_0652_),
    .ZN(_1695_)
  );
  INV_X1 _2562_ (
    .A(_1695_),
    .ZN(_1696_)
  );
  AND2_X1 _2563_ (
    .A1(_0350_),
    .A2(io_in2[28]),
    .ZN(_1697_)
  );
  INV_X1 _2564_ (
    .A(_1697_),
    .ZN(_1698_)
  );
  AND2_X1 _2565_ (
    .A1(_0350_),
    .A2(_0652_),
    .ZN(_1699_)
  );
  INV_X1 _2566_ (
    .A(_1699_),
    .ZN(_1700_)
  );
  AND2_X1 _2567_ (
    .A1(io_fn[3]),
    .A2(io_in2[28]),
    .ZN(_1701_)
  );
  INV_X1 _2568_ (
    .A(_1701_),
    .ZN(_1702_)
  );
  AND2_X1 _2569_ (
    .A1(_1696_),
    .A2(_1698_),
    .ZN(_1703_)
  );
  AND2_X1 _2570_ (
    .A1(_1700_),
    .A2(_1702_),
    .ZN(_1704_)
  );
  AND2_X1 _2571_ (
    .A1(io_in1[28]),
    .A2(_1704_),
    .ZN(_1705_)
  );
  INV_X1 _2572_ (
    .A(_1705_),
    .ZN(_1706_)
  );
  AND2_X1 _2573_ (
    .A1(_0752_),
    .A2(_1703_),
    .ZN(_1707_)
  );
  INV_X1 _2574_ (
    .A(_1707_),
    .ZN(_1708_)
  );
  AND2_X1 _2575_ (
    .A1(_1706_),
    .A2(_1708_),
    .ZN(_1709_)
  );
  INV_X1 _2576_ (
    .A(_1709_),
    .ZN(_1710_)
  );
  AND2_X1 _2577_ (
    .A1(_1694_),
    .A2(_1709_),
    .ZN(_1711_)
  );
  INV_X1 _2578_ (
    .A(_1711_),
    .ZN(_1712_)
  );
  AND2_X1 _2579_ (
    .A1(_1693_),
    .A2(_1710_),
    .ZN(_1713_)
  );
  INV_X1 _2580_ (
    .A(_1713_),
    .ZN(_1714_)
  );
  AND2_X1 _2581_ (
    .A1(_1712_),
    .A2(_1714_),
    .ZN(_1715_)
  );
  INV_X1 _2582_ (
    .A(_1715_),
    .ZN(_1716_)
  );
  AND2_X1 _2583_ (
    .A1(_1691_),
    .A2(_1715_),
    .ZN(_1717_)
  );
  INV_X1 _2584_ (
    .A(_1717_),
    .ZN(_1718_)
  );
  AND2_X1 _2585_ (
    .A1(io_fn[3]),
    .A2(_0663_),
    .ZN(_1719_)
  );
  INV_X1 _2586_ (
    .A(_1719_),
    .ZN(_1720_)
  );
  AND2_X1 _2587_ (
    .A1(_0350_),
    .A2(io_in2[29]),
    .ZN(_1721_)
  );
  INV_X1 _2588_ (
    .A(_1721_),
    .ZN(_1722_)
  );
  AND2_X1 _2589_ (
    .A1(_0350_),
    .A2(_0663_),
    .ZN(_1723_)
  );
  INV_X1 _2590_ (
    .A(_1723_),
    .ZN(_1724_)
  );
  AND2_X1 _2591_ (
    .A1(io_fn[3]),
    .A2(io_in2[29]),
    .ZN(_1725_)
  );
  INV_X1 _2592_ (
    .A(_1725_),
    .ZN(_1726_)
  );
  AND2_X1 _2593_ (
    .A1(_1720_),
    .A2(_1722_),
    .ZN(_1727_)
  );
  AND2_X1 _2594_ (
    .A1(_1724_),
    .A2(_1726_),
    .ZN(_1728_)
  );
  AND2_X1 _2595_ (
    .A1(io_in1[29]),
    .A2(_1728_),
    .ZN(_1729_)
  );
  INV_X1 _2596_ (
    .A(_1729_),
    .ZN(_1730_)
  );
  AND2_X1 _2597_ (
    .A1(_0732_),
    .A2(_1727_),
    .ZN(_1731_)
  );
  INV_X1 _2598_ (
    .A(_1731_),
    .ZN(_1732_)
  );
  AND2_X1 _2599_ (
    .A1(_1730_),
    .A2(_1732_),
    .ZN(_1733_)
  );
  INV_X1 _2600_ (
    .A(_1733_),
    .ZN(_1734_)
  );
  AND2_X1 _2601_ (
    .A1(_1706_),
    .A2(_1712_),
    .ZN(_1735_)
  );
  INV_X1 _2602_ (
    .A(_1735_),
    .ZN(_1736_)
  );
  AND2_X1 _2603_ (
    .A1(_1733_),
    .A2(_1736_),
    .ZN(_1737_)
  );
  INV_X1 _2604_ (
    .A(_1737_),
    .ZN(_1738_)
  );
  AND2_X1 _2605_ (
    .A1(_1734_),
    .A2(_1735_),
    .ZN(_1739_)
  );
  INV_X1 _2606_ (
    .A(_1739_),
    .ZN(_0000_)
  );
  AND2_X1 _2607_ (
    .A1(_1738_),
    .A2(_0000_),
    .ZN(_0001_)
  );
  INV_X1 _2608_ (
    .A(_0001_),
    .ZN(_0002_)
  );
  AND2_X1 _2609_ (
    .A1(_1717_),
    .A2(_0001_),
    .ZN(_0003_)
  );
  INV_X1 _2610_ (
    .A(_0003_),
    .ZN(_0004_)
  );
  AND2_X1 _2611_ (
    .A1(_1730_),
    .A2(_1738_),
    .ZN(_0005_)
  );
  INV_X1 _2612_ (
    .A(_0005_),
    .ZN(_0006_)
  );
  AND2_X1 _2613_ (
    .A1(io_fn[3]),
    .A2(_0672_),
    .ZN(_0007_)
  );
  INV_X1 _2614_ (
    .A(_0007_),
    .ZN(_0008_)
  );
  AND2_X1 _2615_ (
    .A1(_0350_),
    .A2(io_in2[30]),
    .ZN(_0009_)
  );
  INV_X1 _2616_ (
    .A(_0009_),
    .ZN(_0010_)
  );
  AND2_X1 _2617_ (
    .A1(_0350_),
    .A2(_0672_),
    .ZN(_0011_)
  );
  INV_X1 _2618_ (
    .A(_0011_),
    .ZN(_0012_)
  );
  AND2_X1 _2619_ (
    .A1(io_fn[3]),
    .A2(io_in2[30]),
    .ZN(_0013_)
  );
  INV_X1 _2620_ (
    .A(_0013_),
    .ZN(_0014_)
  );
  AND2_X1 _2621_ (
    .A1(_0008_),
    .A2(_0010_),
    .ZN(_0015_)
  );
  AND2_X1 _2622_ (
    .A1(_0012_),
    .A2(_0014_),
    .ZN(_0016_)
  );
  AND2_X1 _2623_ (
    .A1(io_in1[30]),
    .A2(_0016_),
    .ZN(_0017_)
  );
  INV_X1 _2624_ (
    .A(_0017_),
    .ZN(_0018_)
  );
  AND2_X1 _2625_ (
    .A1(_0712_),
    .A2(_0015_),
    .ZN(_0019_)
  );
  INV_X1 _2626_ (
    .A(_0019_),
    .ZN(_0020_)
  );
  AND2_X1 _2627_ (
    .A1(_0018_),
    .A2(_0020_),
    .ZN(_0021_)
  );
  INV_X1 _2628_ (
    .A(_0021_),
    .ZN(_0022_)
  );
  AND2_X1 _2629_ (
    .A1(_0006_),
    .A2(_0021_),
    .ZN(_0023_)
  );
  INV_X1 _2630_ (
    .A(_0023_),
    .ZN(_0024_)
  );
  AND2_X1 _2631_ (
    .A1(_0005_),
    .A2(_0022_),
    .ZN(_0025_)
  );
  INV_X1 _2632_ (
    .A(_0025_),
    .ZN(_0026_)
  );
  AND2_X1 _2633_ (
    .A1(_0024_),
    .A2(_0026_),
    .ZN(_0027_)
  );
  INV_X1 _2634_ (
    .A(_0027_),
    .ZN(_0028_)
  );
  AND2_X1 _2635_ (
    .A1(_0003_),
    .A2(_0027_),
    .ZN(_0029_)
  );
  INV_X1 _2636_ (
    .A(_0029_),
    .ZN(_0030_)
  );
  AND2_X1 _2637_ (
    .A1(_0018_),
    .A2(_0024_),
    .ZN(_0031_)
  );
  INV_X1 _2638_ (
    .A(_0031_),
    .ZN(_0032_)
  );
  AND2_X1 _2639_ (
    .A1(io_in2[31]),
    .A2(_0692_),
    .ZN(_0033_)
  );
  INV_X1 _2640_ (
    .A(_0033_),
    .ZN(_0034_)
  );
  AND2_X1 _2641_ (
    .A1(_0683_),
    .A2(io_in1[31]),
    .ZN(_0035_)
  );
  INV_X1 _2642_ (
    .A(_0035_),
    .ZN(_0036_)
  );
  AND2_X1 _2643_ (
    .A1(_0034_),
    .A2(_0036_),
    .ZN(_0037_)
  );
  INV_X1 _2644_ (
    .A(_0037_),
    .ZN(_0038_)
  );
  AND2_X1 _2645_ (
    .A1(_0350_),
    .A2(_0038_),
    .ZN(_0039_)
  );
  INV_X1 _2646_ (
    .A(_0039_),
    .ZN(_0040_)
  );
  AND2_X1 _2647_ (
    .A1(io_fn[3]),
    .A2(_0037_),
    .ZN(_0041_)
  );
  INV_X1 _2648_ (
    .A(_0041_),
    .ZN(_0042_)
  );
  AND2_X1 _2649_ (
    .A1(_0040_),
    .A2(_0042_),
    .ZN(_0043_)
  );
  INV_X1 _2650_ (
    .A(_0043_),
    .ZN(_0044_)
  );
  AND2_X1 _2651_ (
    .A1(_0031_),
    .A2(_0044_),
    .ZN(_0045_)
  );
  INV_X1 _2652_ (
    .A(_0045_),
    .ZN(_0046_)
  );
  AND2_X1 _2653_ (
    .A1(_0032_),
    .A2(_0043_),
    .ZN(_0047_)
  );
  INV_X1 _2654_ (
    .A(_0047_),
    .ZN(_0048_)
  );
  AND2_X1 _2655_ (
    .A1(_0032_),
    .A2(_0044_),
    .ZN(_0049_)
  );
  INV_X1 _2656_ (
    .A(_0049_),
    .ZN(_0050_)
  );
  AND2_X1 _2657_ (
    .A1(_0031_),
    .A2(_0043_),
    .ZN(_0051_)
  );
  INV_X1 _2658_ (
    .A(_0051_),
    .ZN(_0052_)
  );
  AND2_X1 _2659_ (
    .A1(_0046_),
    .A2(_0048_),
    .ZN(_0053_)
  );
  AND2_X1 _2660_ (
    .A1(_0050_),
    .A2(_0052_),
    .ZN(_0054_)
  );
  AND2_X1 _2661_ (
    .A1(_0029_),
    .A2(_0054_),
    .ZN(_0055_)
  );
  INV_X1 _2662_ (
    .A(_0055_),
    .ZN(_0056_)
  );
  AND2_X1 _2663_ (
    .A1(_0030_),
    .A2(_0053_),
    .ZN(_0057_)
  );
  INV_X1 _2664_ (
    .A(_0057_),
    .ZN(_0058_)
  );
  AND2_X1 _2665_ (
    .A1(_0056_),
    .A2(_0058_),
    .ZN(io_adder_out[31])
  );
  AND2_X1 _2666_ (
    .A1(_0350_),
    .A2(_1416_),
    .ZN(_0059_)
  );
  INV_X1 _2667_ (
    .A(_0059_),
    .ZN(_0060_)
  );
  AND2_X1 _2668_ (
    .A1(_1418_),
    .A2(_0060_),
    .ZN(io_adder_out[0])
  );
  AND2_X1 _2669_ (
    .A1(_0041_),
    .A2(io_adder_out[31]),
    .ZN(_0061_)
  );
  INV_X1 _2670_ (
    .A(_0061_),
    .ZN(_0062_)
  );
  AND2_X1 _2671_ (
    .A1(io_fn[3]),
    .A2(io_fn[1]),
    .ZN(_0063_)
  );
  AND2_X1 _2672_ (
    .A1(_0033_),
    .A2(_0063_),
    .ZN(_0064_)
  );
  INV_X1 _2673_ (
    .A(_0064_),
    .ZN(_0065_)
  );
  AND2_X1 _2674_ (
    .A1(io_fn[3]),
    .A2(_0360_),
    .ZN(_0066_)
  );
  AND2_X1 _2675_ (
    .A1(_0035_),
    .A2(_0066_),
    .ZN(_0067_)
  );
  INV_X1 _2676_ (
    .A(_0067_),
    .ZN(_0068_)
  );
  AND2_X1 _2677_ (
    .A1(_0065_),
    .A2(_0068_),
    .ZN(_0069_)
  );
  AND2_X1 _2678_ (
    .A1(_0062_),
    .A2(_0069_),
    .ZN(_0070_)
  );
  INV_X1 _2679_ (
    .A(_0070_),
    .ZN(_0071_)
  );
  AND2_X1 _2680_ (
    .A1(io_fn[2]),
    .A2(_0071_),
    .ZN(_0072_)
  );
  INV_X1 _2681_ (
    .A(_0072_),
    .ZN(_0073_)
  );
  AND2_X1 _2682_ (
    .A1(_0330_),
    .A2(_0063_),
    .ZN(_0074_)
  );
  INV_X1 _2683_ (
    .A(_0074_),
    .ZN(_0075_)
  );
  AND2_X1 _2684_ (
    .A1(io_fn[2]),
    .A2(_0350_),
    .ZN(_0076_)
  );
  AND2_X1 _2685_ (
    .A1(_0360_),
    .A2(_0076_),
    .ZN(_0077_)
  );
  INV_X1 _2686_ (
    .A(_0077_),
    .ZN(_0078_)
  );
  AND2_X1 _2687_ (
    .A1(_0075_),
    .A2(_0078_),
    .ZN(_0079_)
  );
  INV_X1 _2688_ (
    .A(_0079_),
    .ZN(_0080_)
  );
  AND2_X1 _2689_ (
    .A1(io_fn[0]),
    .A2(_0080_),
    .ZN(_0081_)
  );
  INV_X1 _2690_ (
    .A(_0081_),
    .ZN(_0082_)
  );
  MUX2_X1 _2691_ (
    .A(io_in1[30]),
    .B(io_in1[1]),
    .S(_0081_),
    .Z(_0083_)
  );
  INV_X1 _2692_ (
    .A(_0083_),
    .ZN(_0084_)
  );
  AND2_X1 _2693_ (
    .A1(io_in2[0]),
    .A2(_0084_),
    .ZN(_0085_)
  );
  INV_X1 _2694_ (
    .A(_0085_),
    .ZN(_0086_)
  );
  AND2_X1 _2695_ (
    .A1(io_in1[31]),
    .A2(_0082_),
    .ZN(_0087_)
  );
  INV_X1 _2696_ (
    .A(_0087_),
    .ZN(_0088_)
  );
  AND2_X1 _2697_ (
    .A1(io_in1[0]),
    .A2(_0081_),
    .ZN(_0089_)
  );
  INV_X1 _2698_ (
    .A(_0089_),
    .ZN(_0090_)
  );
  AND2_X1 _2699_ (
    .A1(_0370_),
    .A2(_0090_),
    .ZN(_0091_)
  );
  AND2_X1 _2700_ (
    .A1(_0088_),
    .A2(_0091_),
    .ZN(_0092_)
  );
  INV_X1 _2701_ (
    .A(_0092_),
    .ZN(_0093_)
  );
  AND2_X1 _2702_ (
    .A1(_0086_),
    .A2(_0093_),
    .ZN(_0094_)
  );
  MUX2_X1 _2703_ (
    .A(io_in1[29]),
    .B(io_in1[2]),
    .S(_0081_),
    .Z(_0095_)
  );
  MUX2_X1 _2704_ (
    .A(io_in1[28]),
    .B(io_in1[3]),
    .S(_0081_),
    .Z(_0096_)
  );
  MUX2_X1 _2705_ (
    .A(_0095_),
    .B(_0096_),
    .S(io_in2[0]),
    .Z(_0097_)
  );
  MUX2_X1 _2706_ (
    .A(_0094_),
    .B(_0097_),
    .S(io_in2[1]),
    .Z(_0098_)
  );
  MUX2_X1 _2707_ (
    .A(io_in1[27]),
    .B(io_in1[4]),
    .S(_0081_),
    .Z(_0099_)
  );
  MUX2_X1 _2708_ (
    .A(io_in1[26]),
    .B(io_in1[5]),
    .S(_0081_),
    .Z(_0100_)
  );
  MUX2_X1 _2709_ (
    .A(_0099_),
    .B(_0100_),
    .S(io_in2[0]),
    .Z(_0101_)
  );
  MUX2_X1 _2710_ (
    .A(io_in1[25]),
    .B(io_in1[6]),
    .S(_0081_),
    .Z(_0102_)
  );
  MUX2_X1 _2711_ (
    .A(io_in1[24]),
    .B(io_in1[7]),
    .S(_0081_),
    .Z(_0103_)
  );
  MUX2_X1 _2712_ (
    .A(_0102_),
    .B(_0103_),
    .S(io_in2[0]),
    .Z(_0104_)
  );
  MUX2_X1 _2713_ (
    .A(_0101_),
    .B(_0104_),
    .S(io_in2[1]),
    .Z(_0105_)
  );
  MUX2_X1 _2714_ (
    .A(_0098_),
    .B(_0105_),
    .S(io_in2[2]),
    .Z(_0106_)
  );
  MUX2_X1 _2715_ (
    .A(io_in1[23]),
    .B(io_in1[8]),
    .S(_0081_),
    .Z(_0107_)
  );
  MUX2_X1 _2716_ (
    .A(io_in1[22]),
    .B(io_in1[9]),
    .S(_0081_),
    .Z(_0108_)
  );
  MUX2_X1 _2717_ (
    .A(_0107_),
    .B(_0108_),
    .S(io_in2[0]),
    .Z(_0109_)
  );
  MUX2_X1 _2718_ (
    .A(io_in1[21]),
    .B(io_in1[10]),
    .S(_0081_),
    .Z(_0110_)
  );
  MUX2_X1 _2719_ (
    .A(io_in1[20]),
    .B(io_in1[11]),
    .S(_0081_),
    .Z(_0111_)
  );
  MUX2_X1 _2720_ (
    .A(_0110_),
    .B(_0111_),
    .S(io_in2[0]),
    .Z(_0112_)
  );
  MUX2_X1 _2721_ (
    .A(_0109_),
    .B(_0112_),
    .S(io_in2[1]),
    .Z(_0113_)
  );
  MUX2_X1 _2722_ (
    .A(io_in1[19]),
    .B(io_in1[12]),
    .S(_0081_),
    .Z(_0114_)
  );
  MUX2_X1 _2723_ (
    .A(io_in1[18]),
    .B(io_in1[13]),
    .S(_0081_),
    .Z(_0115_)
  );
  MUX2_X1 _2724_ (
    .A(_0114_),
    .B(_0115_),
    .S(io_in2[0]),
    .Z(_0116_)
  );
  MUX2_X1 _2725_ (
    .A(io_in1[17]),
    .B(io_in1[14]),
    .S(_0081_),
    .Z(_0117_)
  );
  MUX2_X1 _2726_ (
    .A(io_in1[16]),
    .B(io_in1[15]),
    .S(_0081_),
    .Z(_0118_)
  );
  MUX2_X1 _2727_ (
    .A(_0117_),
    .B(_0118_),
    .S(io_in2[0]),
    .Z(_0119_)
  );
  MUX2_X1 _2728_ (
    .A(_0116_),
    .B(_0119_),
    .S(io_in2[1]),
    .Z(_0120_)
  );
  MUX2_X1 _2729_ (
    .A(_0113_),
    .B(_0120_),
    .S(io_in2[2]),
    .Z(_0121_)
  );
  MUX2_X1 _2730_ (
    .A(_0106_),
    .B(_0121_),
    .S(io_in2[3]),
    .Z(_0122_)
  );
  MUX2_X1 _2731_ (
    .A(io_in1[15]),
    .B(io_in1[16]),
    .S(_0081_),
    .Z(_0123_)
  );
  MUX2_X1 _2732_ (
    .A(io_in1[14]),
    .B(io_in1[17]),
    .S(_0081_),
    .Z(_0124_)
  );
  MUX2_X1 _2733_ (
    .A(_0123_),
    .B(_0124_),
    .S(io_in2[0]),
    .Z(_0125_)
  );
  MUX2_X1 _2734_ (
    .A(io_in1[13]),
    .B(io_in1[18]),
    .S(_0081_),
    .Z(_0126_)
  );
  MUX2_X1 _2735_ (
    .A(io_in1[12]),
    .B(io_in1[19]),
    .S(_0081_),
    .Z(_0127_)
  );
  MUX2_X1 _2736_ (
    .A(_0126_),
    .B(_0127_),
    .S(io_in2[0]),
    .Z(_0128_)
  );
  MUX2_X1 _2737_ (
    .A(_0125_),
    .B(_0128_),
    .S(io_in2[1]),
    .Z(_0129_)
  );
  MUX2_X1 _2738_ (
    .A(io_in1[11]),
    .B(io_in1[20]),
    .S(_0081_),
    .Z(_0130_)
  );
  MUX2_X1 _2739_ (
    .A(io_in1[10]),
    .B(io_in1[21]),
    .S(_0081_),
    .Z(_0131_)
  );
  MUX2_X1 _2740_ (
    .A(_0130_),
    .B(_0131_),
    .S(io_in2[0]),
    .Z(_0132_)
  );
  MUX2_X1 _2741_ (
    .A(io_in1[9]),
    .B(io_in1[22]),
    .S(_0081_),
    .Z(_0133_)
  );
  MUX2_X1 _2742_ (
    .A(io_in1[8]),
    .B(io_in1[23]),
    .S(_0081_),
    .Z(_0134_)
  );
  MUX2_X1 _2743_ (
    .A(_0133_),
    .B(_0134_),
    .S(io_in2[0]),
    .Z(_0135_)
  );
  MUX2_X1 _2744_ (
    .A(_0132_),
    .B(_0135_),
    .S(io_in2[1]),
    .Z(_0136_)
  );
  MUX2_X1 _2745_ (
    .A(_0129_),
    .B(_0136_),
    .S(io_in2[2]),
    .Z(_0137_)
  );
  MUX2_X1 _2746_ (
    .A(io_in1[7]),
    .B(io_in1[24]),
    .S(_0081_),
    .Z(_0138_)
  );
  MUX2_X1 _2747_ (
    .A(io_in1[6]),
    .B(io_in1[25]),
    .S(_0081_),
    .Z(_0139_)
  );
  MUX2_X1 _2748_ (
    .A(_0138_),
    .B(_0139_),
    .S(io_in2[0]),
    .Z(_0140_)
  );
  MUX2_X1 _2749_ (
    .A(io_in1[5]),
    .B(io_in1[26]),
    .S(_0081_),
    .Z(_0141_)
  );
  MUX2_X1 _2750_ (
    .A(io_in1[4]),
    .B(io_in1[27]),
    .S(_0081_),
    .Z(_0142_)
  );
  MUX2_X1 _2751_ (
    .A(_0141_),
    .B(_0142_),
    .S(io_in2[0]),
    .Z(_0143_)
  );
  MUX2_X1 _2752_ (
    .A(_0140_),
    .B(_0143_),
    .S(io_in2[1]),
    .Z(_0144_)
  );
  MUX2_X1 _2753_ (
    .A(io_in1[3]),
    .B(io_in1[28]),
    .S(_0081_),
    .Z(_0145_)
  );
  MUX2_X1 _2754_ (
    .A(io_in1[2]),
    .B(io_in1[29]),
    .S(_0081_),
    .Z(_0146_)
  );
  MUX2_X1 _2755_ (
    .A(_0145_),
    .B(_0146_),
    .S(io_in2[0]),
    .Z(_0147_)
  );
  MUX2_X1 _2756_ (
    .A(io_in1[1]),
    .B(io_in1[30]),
    .S(_0081_),
    .Z(_0148_)
  );
  MUX2_X1 _2757_ (
    .A(io_in1[0]),
    .B(io_in1[31]),
    .S(_0081_),
    .Z(_0149_)
  );
  MUX2_X1 _2758_ (
    .A(_0148_),
    .B(_0149_),
    .S(io_in2[0]),
    .Z(_0150_)
  );
  MUX2_X1 _2759_ (
    .A(_0147_),
    .B(_0150_),
    .S(io_in2[1]),
    .Z(_0151_)
  );
  MUX2_X1 _2760_ (
    .A(_0144_),
    .B(_0151_),
    .S(io_in2[2]),
    .Z(_0152_)
  );
  MUX2_X1 _2761_ (
    .A(_0137_),
    .B(_0152_),
    .S(io_in2[3]),
    .Z(_0153_)
  );
  MUX2_X1 _2762_ (
    .A(_0122_),
    .B(_0153_),
    .S(io_in2[4]),
    .Z(_0154_)
  );
  AND2_X1 _2763_ (
    .A1(_0081_),
    .A2(_0154_),
    .ZN(_0155_)
  );
  INV_X1 _2764_ (
    .A(_0155_),
    .ZN(_0156_)
  );
  AND2_X1 _2765_ (
    .A1(_1257_),
    .A2(_0149_),
    .ZN(_0157_)
  );
  AND2_X1 _2766_ (
    .A1(_1249_),
    .A2(_0157_),
    .ZN(_0158_)
  );
  AND2_X1 _2767_ (
    .A1(io_fn[3]),
    .A2(_0149_),
    .ZN(_0159_)
  );
  MUX2_X1 _2768_ (
    .A(_0158_),
    .B(_0159_),
    .S(io_in2[2]),
    .Z(_0160_)
  );
  MUX2_X1 _2769_ (
    .A(_0159_),
    .B(_0160_),
    .S(_0401_),
    .Z(_0161_)
  );
  MUX2_X1 _2770_ (
    .A(_0159_),
    .B(_0161_),
    .S(_0412_),
    .Z(_0162_)
  );
  AND2_X1 _2771_ (
    .A1(_0330_),
    .A2(_0350_),
    .ZN(_0163_)
  );
  AND2_X1 _2772_ (
    .A1(_0360_),
    .A2(_0163_),
    .ZN(_0164_)
  );
  INV_X1 _2773_ (
    .A(_0164_),
    .ZN(_0165_)
  );
  AND2_X1 _2774_ (
    .A1(io_fn[0]),
    .A2(_0164_),
    .ZN(_0166_)
  );
  AND2_X1 _2775_ (
    .A1(_0162_),
    .A2(_0166_),
    .ZN(_0167_)
  );
  INV_X1 _2776_ (
    .A(_0167_),
    .ZN(_0168_)
  );
  AND2_X1 _2777_ (
    .A1(_0075_),
    .A2(_0165_),
    .ZN(_0169_)
  );
  INV_X1 _2778_ (
    .A(_0169_),
    .ZN(_0170_)
  );
  AND2_X1 _2779_ (
    .A1(_0339_),
    .A2(_0170_),
    .ZN(_0171_)
  );
  AND2_X1 _2780_ (
    .A1(io_adder_out[0]),
    .A2(_0171_),
    .ZN(_0172_)
  );
  INV_X1 _2781_ (
    .A(_0172_),
    .ZN(_0173_)
  );
  AND2_X1 _2782_ (
    .A1(io_fn[1]),
    .A2(_0076_),
    .ZN(_0174_)
  );
  AND2_X1 _2783_ (
    .A1(io_in2[0]),
    .A2(io_in1[0]),
    .ZN(_0175_)
  );
  AND2_X1 _2784_ (
    .A1(_0174_),
    .A2(_0175_),
    .ZN(_0176_)
  );
  INV_X1 _2785_ (
    .A(_0176_),
    .ZN(_0177_)
  );
  AND2_X1 _2786_ (
    .A1(_0339_),
    .A2(_0076_),
    .ZN(_0178_)
  );
  AND2_X1 _2787_ (
    .A1(_1415_),
    .A2(_0178_),
    .ZN(_0179_)
  );
  INV_X1 _2788_ (
    .A(_0179_),
    .ZN(_0180_)
  );
  AND2_X1 _2789_ (
    .A1(_0177_),
    .A2(_0180_),
    .ZN(_0181_)
  );
  AND2_X1 _2790_ (
    .A1(_0173_),
    .A2(_0181_),
    .ZN(_0182_)
  );
  AND2_X1 _2791_ (
    .A1(_0168_),
    .A2(_0182_),
    .ZN(_0183_)
  );
  AND2_X1 _2792_ (
    .A1(_0156_),
    .A2(_0183_),
    .ZN(_0184_)
  );
  AND2_X1 _2793_ (
    .A1(_0073_),
    .A2(_0184_),
    .ZN(_0185_)
  );
  INV_X1 _2794_ (
    .A(_0185_),
    .ZN(io_out[0])
  );
  AND2_X1 _2795_ (
    .A1(_1263_),
    .A2(_1267_),
    .ZN(_0186_)
  );
  INV_X1 _2796_ (
    .A(_0186_),
    .ZN(_0187_)
  );
  AND2_X1 _2797_ (
    .A1(_1269_),
    .A2(_0187_),
    .ZN(_0188_)
  );
  MUX2_X1 _2798_ (
    .A(_1267_),
    .B(_0188_),
    .S(_1418_),
    .Z(io_adder_out[1])
  );
  MUX2_X1 _2799_ (
    .A(_0150_),
    .B(_0159_),
    .S(io_in2[1]),
    .Z(_0189_)
  );
  MUX2_X1 _2800_ (
    .A(_0159_),
    .B(_0189_),
    .S(_0390_),
    .Z(_0190_)
  );
  MUX2_X1 _2801_ (
    .A(_0159_),
    .B(_0190_),
    .S(_0401_),
    .Z(_0191_)
  );
  MUX2_X1 _2802_ (
    .A(_0159_),
    .B(_0191_),
    .S(_0412_),
    .Z(_0192_)
  );
  AND2_X1 _2803_ (
    .A1(_0166_),
    .A2(_0192_),
    .ZN(_0193_)
  );
  INV_X1 _2804_ (
    .A(_0193_),
    .ZN(_0194_)
  );
  MUX2_X1 _2805_ (
    .A(_0083_),
    .B(_0095_),
    .S(io_in2[0]),
    .Z(_0195_)
  );
  MUX2_X1 _2806_ (
    .A(_0096_),
    .B(_0099_),
    .S(io_in2[0]),
    .Z(_0196_)
  );
  MUX2_X1 _2807_ (
    .A(_0195_),
    .B(_0196_),
    .S(io_in2[1]),
    .Z(_0197_)
  );
  MUX2_X1 _2808_ (
    .A(_0100_),
    .B(_0102_),
    .S(io_in2[0]),
    .Z(_0198_)
  );
  MUX2_X1 _2809_ (
    .A(_0103_),
    .B(_0107_),
    .S(io_in2[0]),
    .Z(_0199_)
  );
  MUX2_X1 _2810_ (
    .A(_0198_),
    .B(_0199_),
    .S(io_in2[1]),
    .Z(_0200_)
  );
  MUX2_X1 _2811_ (
    .A(_0197_),
    .B(_0200_),
    .S(io_in2[2]),
    .Z(_0201_)
  );
  MUX2_X1 _2812_ (
    .A(_0108_),
    .B(_0110_),
    .S(io_in2[0]),
    .Z(_0202_)
  );
  MUX2_X1 _2813_ (
    .A(_0111_),
    .B(_0114_),
    .S(io_in2[0]),
    .Z(_0203_)
  );
  MUX2_X1 _2814_ (
    .A(_0202_),
    .B(_0203_),
    .S(io_in2[1]),
    .Z(_0204_)
  );
  MUX2_X1 _2815_ (
    .A(_0115_),
    .B(_0117_),
    .S(io_in2[0]),
    .Z(_0205_)
  );
  MUX2_X1 _2816_ (
    .A(_0118_),
    .B(_0123_),
    .S(io_in2[0]),
    .Z(_0206_)
  );
  MUX2_X1 _2817_ (
    .A(_0205_),
    .B(_0206_),
    .S(io_in2[1]),
    .Z(_0207_)
  );
  MUX2_X1 _2818_ (
    .A(_0204_),
    .B(_0207_),
    .S(io_in2[2]),
    .Z(_0208_)
  );
  MUX2_X1 _2819_ (
    .A(_0201_),
    .B(_0208_),
    .S(io_in2[3]),
    .Z(_0209_)
  );
  MUX2_X1 _2820_ (
    .A(_0124_),
    .B(_0126_),
    .S(io_in2[0]),
    .Z(_0210_)
  );
  MUX2_X1 _2821_ (
    .A(_0127_),
    .B(_0130_),
    .S(io_in2[0]),
    .Z(_0211_)
  );
  MUX2_X1 _2822_ (
    .A(_0210_),
    .B(_0211_),
    .S(io_in2[1]),
    .Z(_0212_)
  );
  MUX2_X1 _2823_ (
    .A(_0131_),
    .B(_0133_),
    .S(io_in2[0]),
    .Z(_0213_)
  );
  MUX2_X1 _2824_ (
    .A(_0134_),
    .B(_0138_),
    .S(io_in2[0]),
    .Z(_0214_)
  );
  MUX2_X1 _2825_ (
    .A(_0213_),
    .B(_0214_),
    .S(io_in2[1]),
    .Z(_0215_)
  );
  MUX2_X1 _2826_ (
    .A(_0212_),
    .B(_0215_),
    .S(io_in2[2]),
    .Z(_0216_)
  );
  MUX2_X1 _2827_ (
    .A(_0139_),
    .B(_0141_),
    .S(io_in2[0]),
    .Z(_0217_)
  );
  MUX2_X1 _2828_ (
    .A(_0142_),
    .B(_0145_),
    .S(io_in2[0]),
    .Z(_0218_)
  );
  MUX2_X1 _2829_ (
    .A(_0217_),
    .B(_0218_),
    .S(io_in2[1]),
    .Z(_0219_)
  );
  MUX2_X1 _2830_ (
    .A(_0146_),
    .B(_0148_),
    .S(io_in2[0]),
    .Z(_0220_)
  );
  MUX2_X1 _2831_ (
    .A(_0157_),
    .B(_0220_),
    .S(_0381_),
    .Z(_0221_)
  );
  MUX2_X1 _2832_ (
    .A(_0219_),
    .B(_0221_),
    .S(io_in2[2]),
    .Z(_0222_)
  );
  MUX2_X1 _2833_ (
    .A(_0216_),
    .B(_0222_),
    .S(io_in2[3]),
    .Z(_0223_)
  );
  MUX2_X1 _2834_ (
    .A(_0209_),
    .B(_0223_),
    .S(io_in2[4]),
    .Z(_0224_)
  );
  AND2_X1 _2835_ (
    .A1(_0081_),
    .A2(_0224_),
    .ZN(_0225_)
  );
  INV_X1 _2836_ (
    .A(_0225_),
    .ZN(_0226_)
  );
  AND2_X1 _2837_ (
    .A1(_0171_),
    .A2(io_adder_out[1]),
    .ZN(_0227_)
  );
  INV_X1 _2838_ (
    .A(_0227_),
    .ZN(_0228_)
  );
  AND2_X1 _2839_ (
    .A1(_1266_),
    .A2(_0178_),
    .ZN(_0229_)
  );
  INV_X1 _2840_ (
    .A(_0229_),
    .ZN(_0230_)
  );
  AND2_X1 _2841_ (
    .A1(io_in2[1]),
    .A2(io_in1[1]),
    .ZN(_0231_)
  );
  AND2_X1 _2842_ (
    .A1(_0174_),
    .A2(_0231_),
    .ZN(_0232_)
  );
  INV_X1 _2843_ (
    .A(_0232_),
    .ZN(_0233_)
  );
  AND2_X1 _2844_ (
    .A1(_0230_),
    .A2(_0233_),
    .ZN(_0234_)
  );
  AND2_X1 _2845_ (
    .A1(_0228_),
    .A2(_0234_),
    .ZN(_0235_)
  );
  AND2_X1 _2846_ (
    .A1(_0226_),
    .A2(_0235_),
    .ZN(_0236_)
  );
  AND2_X1 _2847_ (
    .A1(_0194_),
    .A2(_0236_),
    .ZN(_0237_)
  );
  INV_X1 _2848_ (
    .A(_0237_),
    .ZN(io_out[1])
  );
  AND2_X1 _2849_ (
    .A1(_1420_),
    .A2(_1424_),
    .ZN(_0238_)
  );
  INV_X1 _2850_ (
    .A(_0238_),
    .ZN(_0239_)
  );
  AND2_X1 _2851_ (
    .A1(_1426_),
    .A2(_0239_),
    .ZN(io_adder_out[2])
  );
  MUX2_X1 _2852_ (
    .A(_0159_),
    .B(_0221_),
    .S(_0390_),
    .Z(_0240_)
  );
  MUX2_X1 _2853_ (
    .A(_0159_),
    .B(_0240_),
    .S(_0401_),
    .Z(_0241_)
  );
  MUX2_X1 _2854_ (
    .A(_0159_),
    .B(_0241_),
    .S(_0412_),
    .Z(_0242_)
  );
  AND2_X1 _2855_ (
    .A1(_0166_),
    .A2(_0242_),
    .ZN(_0243_)
  );
  INV_X1 _2856_ (
    .A(_0243_),
    .ZN(_0244_)
  );
  MUX2_X1 _2857_ (
    .A(_0097_),
    .B(_0101_),
    .S(io_in2[1]),
    .Z(_0245_)
  );
  MUX2_X1 _2858_ (
    .A(_0104_),
    .B(_0109_),
    .S(io_in2[1]),
    .Z(_0246_)
  );
  MUX2_X1 _2859_ (
    .A(_0245_),
    .B(_0246_),
    .S(io_in2[2]),
    .Z(_0247_)
  );
  MUX2_X1 _2860_ (
    .A(_0112_),
    .B(_0116_),
    .S(io_in2[1]),
    .Z(_0248_)
  );
  MUX2_X1 _2861_ (
    .A(_0119_),
    .B(_0125_),
    .S(io_in2[1]),
    .Z(_0249_)
  );
  MUX2_X1 _2862_ (
    .A(_0248_),
    .B(_0249_),
    .S(io_in2[2]),
    .Z(_0250_)
  );
  MUX2_X1 _2863_ (
    .A(_0247_),
    .B(_0250_),
    .S(io_in2[3]),
    .Z(_0251_)
  );
  MUX2_X1 _2864_ (
    .A(_0128_),
    .B(_0132_),
    .S(io_in2[1]),
    .Z(_0252_)
  );
  MUX2_X1 _2865_ (
    .A(_0135_),
    .B(_0140_),
    .S(io_in2[1]),
    .Z(_0253_)
  );
  MUX2_X1 _2866_ (
    .A(_0252_),
    .B(_0253_),
    .S(io_in2[2]),
    .Z(_0254_)
  );
  MUX2_X1 _2867_ (
    .A(_0143_),
    .B(_0147_),
    .S(io_in2[1]),
    .Z(_0255_)
  );
  MUX2_X1 _2868_ (
    .A(_0189_),
    .B(_0255_),
    .S(_0390_),
    .Z(_0256_)
  );
  MUX2_X1 _2869_ (
    .A(_0254_),
    .B(_0256_),
    .S(io_in2[3]),
    .Z(_0257_)
  );
  MUX2_X1 _2870_ (
    .A(_0251_),
    .B(_0257_),
    .S(io_in2[4]),
    .Z(_0258_)
  );
  AND2_X1 _2871_ (
    .A1(_0081_),
    .A2(_0258_),
    .ZN(_0259_)
  );
  INV_X1 _2872_ (
    .A(_0259_),
    .ZN(_0260_)
  );
  AND2_X1 _2873_ (
    .A1(_0171_),
    .A2(io_adder_out[2]),
    .ZN(_0261_)
  );
  INV_X1 _2874_ (
    .A(_0261_),
    .ZN(_0262_)
  );
  AND2_X1 _2875_ (
    .A1(_1274_),
    .A2(_0178_),
    .ZN(_0263_)
  );
  INV_X1 _2876_ (
    .A(_0263_),
    .ZN(_0264_)
  );
  AND2_X1 _2877_ (
    .A1(io_in2[2]),
    .A2(io_in1[2]),
    .ZN(_0265_)
  );
  AND2_X1 _2878_ (
    .A1(_0174_),
    .A2(_0265_),
    .ZN(_0266_)
  );
  INV_X1 _2879_ (
    .A(_0266_),
    .ZN(_0267_)
  );
  AND2_X1 _2880_ (
    .A1(_0262_),
    .A2(_0264_),
    .ZN(_0268_)
  );
  AND2_X1 _2881_ (
    .A1(_0244_),
    .A2(_0267_),
    .ZN(_0269_)
  );
  AND2_X1 _2882_ (
    .A1(_0260_),
    .A2(_0269_),
    .ZN(_0270_)
  );
  AND2_X1 _2883_ (
    .A1(_0268_),
    .A2(_0270_),
    .ZN(_0271_)
  );
  INV_X1 _2884_ (
    .A(_0271_),
    .ZN(io_out[2])
  );
  AND2_X1 _2885_ (
    .A1(_1426_),
    .A2(_1430_),
    .ZN(_0272_)
  );
  INV_X1 _2886_ (
    .A(_0272_),
    .ZN(_0273_)
  );
  AND2_X1 _2887_ (
    .A1(_1432_),
    .A2(_0273_),
    .ZN(io_adder_out[3])
  );
  MUX2_X1 _2888_ (
    .A(_0151_),
    .B(_0159_),
    .S(io_in2[2]),
    .Z(_0274_)
  );
  MUX2_X1 _2889_ (
    .A(_0159_),
    .B(_0274_),
    .S(_0401_),
    .Z(_0275_)
  );
  MUX2_X1 _2890_ (
    .A(_0159_),
    .B(_0275_),
    .S(_0412_),
    .Z(_0276_)
  );
  AND2_X1 _2891_ (
    .A1(_0166_),
    .A2(_0276_),
    .ZN(_0277_)
  );
  INV_X1 _2892_ (
    .A(_0277_),
    .ZN(_0278_)
  );
  MUX2_X1 _2893_ (
    .A(_0196_),
    .B(_0198_),
    .S(io_in2[1]),
    .Z(_0279_)
  );
  MUX2_X1 _2894_ (
    .A(_0199_),
    .B(_0202_),
    .S(io_in2[1]),
    .Z(_0280_)
  );
  MUX2_X1 _2895_ (
    .A(_0279_),
    .B(_0280_),
    .S(io_in2[2]),
    .Z(_0281_)
  );
  MUX2_X1 _2896_ (
    .A(_0203_),
    .B(_0205_),
    .S(io_in2[1]),
    .Z(_0282_)
  );
  MUX2_X1 _2897_ (
    .A(_0206_),
    .B(_0210_),
    .S(io_in2[1]),
    .Z(_0283_)
  );
  MUX2_X1 _2898_ (
    .A(_0282_),
    .B(_0283_),
    .S(io_in2[2]),
    .Z(_0284_)
  );
  MUX2_X1 _2899_ (
    .A(_0281_),
    .B(_0284_),
    .S(io_in2[3]),
    .Z(_0285_)
  );
  MUX2_X1 _2900_ (
    .A(_0211_),
    .B(_0213_),
    .S(io_in2[1]),
    .Z(_0286_)
  );
  MUX2_X1 _2901_ (
    .A(_0214_),
    .B(_0217_),
    .S(io_in2[1]),
    .Z(_0287_)
  );
  MUX2_X1 _2902_ (
    .A(_0286_),
    .B(_0287_),
    .S(io_in2[2]),
    .Z(_0288_)
  );
  MUX2_X1 _2903_ (
    .A(_0218_),
    .B(_0220_),
    .S(io_in2[1]),
    .Z(_0289_)
  );
  MUX2_X1 _2904_ (
    .A(_0158_),
    .B(_0289_),
    .S(_0390_),
    .Z(_0290_)
  );
  MUX2_X1 _2905_ (
    .A(_0288_),
    .B(_0290_),
    .S(io_in2[3]),
    .Z(_0291_)
  );
  MUX2_X1 _2906_ (
    .A(_0285_),
    .B(_0291_),
    .S(io_in2[4]),
    .Z(_0292_)
  );
  AND2_X1 _2907_ (
    .A1(_0081_),
    .A2(_0292_),
    .ZN(_0293_)
  );
  INV_X1 _2908_ (
    .A(_0293_),
    .ZN(_0294_)
  );
  AND2_X1 _2909_ (
    .A1(_0171_),
    .A2(io_adder_out[3]),
    .ZN(_0295_)
  );
  INV_X1 _2910_ (
    .A(_0295_),
    .ZN(_0296_)
  );
  AND2_X1 _2911_ (
    .A1(_1282_),
    .A2(_0178_),
    .ZN(_0297_)
  );
  INV_X1 _2912_ (
    .A(_0297_),
    .ZN(_0298_)
  );
  AND2_X1 _2913_ (
    .A1(io_in2[3]),
    .A2(io_in1[3]),
    .ZN(_0299_)
  );
  AND2_X1 _2914_ (
    .A1(_0174_),
    .A2(_0299_),
    .ZN(_0300_)
  );
  INV_X1 _2915_ (
    .A(_0300_),
    .ZN(_0301_)
  );
  AND2_X1 _2916_ (
    .A1(_0296_),
    .A2(_0298_),
    .ZN(_0302_)
  );
  AND2_X1 _2917_ (
    .A1(_0278_),
    .A2(_0301_),
    .ZN(_0303_)
  );
  AND2_X1 _2918_ (
    .A1(_0294_),
    .A2(_0303_),
    .ZN(_0304_)
  );
  AND2_X1 _2919_ (
    .A1(_0302_),
    .A2(_0304_),
    .ZN(_0305_)
  );
  INV_X1 _2920_ (
    .A(_0305_),
    .ZN(io_out[3])
  );
  AND2_X1 _2921_ (
    .A1(_1432_),
    .A2(_1436_),
    .ZN(_0306_)
  );
  INV_X1 _2922_ (
    .A(_0306_),
    .ZN(_0307_)
  );
  AND2_X1 _2923_ (
    .A1(_1438_),
    .A2(_0307_),
    .ZN(io_adder_out[4])
  );
  MUX2_X1 _2924_ (
    .A(_0159_),
    .B(_0290_),
    .S(_0401_),
    .Z(_0308_)
  );
  MUX2_X1 _2925_ (
    .A(_0159_),
    .B(_0308_),
    .S(_0412_),
    .Z(_0309_)
  );
  AND2_X1 _2926_ (
    .A1(_0166_),
    .A2(_0309_),
    .ZN(_0310_)
  );
  INV_X1 _2927_ (
    .A(_0310_),
    .ZN(_0311_)
  );
  MUX2_X1 _2928_ (
    .A(_0105_),
    .B(_0113_),
    .S(io_in2[2]),
    .Z(_0312_)
  );
  MUX2_X1 _2929_ (
    .A(_0120_),
    .B(_0129_),
    .S(io_in2[2]),
    .Z(_0313_)
  );
  MUX2_X1 _2930_ (
    .A(_0312_),
    .B(_0313_),
    .S(io_in2[3]),
    .Z(_0314_)
  );
  MUX2_X1 _2931_ (
    .A(_0136_),
    .B(_0144_),
    .S(io_in2[2]),
    .Z(_0315_)
  );
  MUX2_X1 _2932_ (
    .A(_0274_),
    .B(_0315_),
    .S(_0401_),
    .Z(_0316_)
  );
  MUX2_X1 _2933_ (
    .A(_0314_),
    .B(_0316_),
    .S(io_in2[4]),
    .Z(_0317_)
  );
  AND2_X1 _2934_ (
    .A1(_0081_),
    .A2(_0317_),
    .ZN(_0318_)
  );
  INV_X1 _2935_ (
    .A(_0318_),
    .ZN(_0319_)
  );
  AND2_X1 _2936_ (
    .A1(_0171_),
    .A2(io_adder_out[4]),
    .ZN(_0320_)
  );
  INV_X1 _2937_ (
    .A(_0320_),
    .ZN(_0321_)
  );
  AND2_X1 _2938_ (
    .A1(_1290_),
    .A2(_0178_),
    .ZN(_0322_)
  );
  INV_X1 _2939_ (
    .A(_0322_),
    .ZN(_0323_)
  );
  AND2_X1 _2940_ (
    .A1(io_in2[4]),
    .A2(io_in1[4]),
    .ZN(_0324_)
  );
  AND2_X1 _2941_ (
    .A1(_0174_),
    .A2(_0324_),
    .ZN(_0325_)
  );
  INV_X1 _2942_ (
    .A(_0325_),
    .ZN(_0326_)
  );
  AND2_X1 _2943_ (
    .A1(_0321_),
    .A2(_0323_),
    .ZN(_0327_)
  );
  AND2_X1 _2944_ (
    .A1(_0311_),
    .A2(_0326_),
    .ZN(_0328_)
  );
  AND2_X1 _2945_ (
    .A1(_0319_),
    .A2(_0328_),
    .ZN(_0329_)
  );
  AND2_X1 _2946_ (
    .A1(_0327_),
    .A2(_0329_),
    .ZN(_0331_)
  );
  INV_X1 _2947_ (
    .A(_0331_),
    .ZN(io_out[4])
  );
  AND2_X1 _2948_ (
    .A1(_1438_),
    .A2(_1442_),
    .ZN(_0332_)
  );
  INV_X1 _2949_ (
    .A(_0332_),
    .ZN(_0333_)
  );
  AND2_X1 _2950_ (
    .A1(_1444_),
    .A2(_0333_),
    .ZN(io_adder_out[5])
  );
  MUX2_X1 _2951_ (
    .A(_0159_),
    .B(_0256_),
    .S(_0401_),
    .Z(_0334_)
  );
  MUX2_X1 _2952_ (
    .A(_0159_),
    .B(_0334_),
    .S(_0412_),
    .Z(_0335_)
  );
  AND2_X1 _2953_ (
    .A1(_0166_),
    .A2(_0335_),
    .ZN(_0336_)
  );
  INV_X1 _2954_ (
    .A(_0336_),
    .ZN(_0337_)
  );
  AND2_X1 _2955_ (
    .A1(io_in2[5]),
    .A2(io_in1[5]),
    .ZN(_0338_)
  );
  AND2_X1 _2956_ (
    .A1(_0174_),
    .A2(_0338_),
    .ZN(_0340_)
  );
  INV_X1 _2957_ (
    .A(_0340_),
    .ZN(_0341_)
  );
  AND2_X1 _2958_ (
    .A1(_1298_),
    .A2(_0178_),
    .ZN(_0342_)
  );
  INV_X1 _2959_ (
    .A(_0342_),
    .ZN(_0343_)
  );
  AND2_X1 _2960_ (
    .A1(_0341_),
    .A2(_0343_),
    .ZN(_0344_)
  );
  AND2_X1 _2961_ (
    .A1(_0337_),
    .A2(_0344_),
    .ZN(_0345_)
  );
  AND2_X1 _2962_ (
    .A1(_0171_),
    .A2(io_adder_out[5]),
    .ZN(_0346_)
  );
  INV_X1 _2963_ (
    .A(_0346_),
    .ZN(_0347_)
  );
  MUX2_X1 _2964_ (
    .A(_0200_),
    .B(_0204_),
    .S(io_in2[2]),
    .Z(_0348_)
  );
  MUX2_X1 _2965_ (
    .A(_0207_),
    .B(_0212_),
    .S(io_in2[2]),
    .Z(_0349_)
  );
  MUX2_X1 _2966_ (
    .A(_0348_),
    .B(_0349_),
    .S(io_in2[3]),
    .Z(_0351_)
  );
  MUX2_X1 _2967_ (
    .A(_0215_),
    .B(_0219_),
    .S(io_in2[2]),
    .Z(_0352_)
  );
  MUX2_X1 _2968_ (
    .A(_0240_),
    .B(_0352_),
    .S(_0401_),
    .Z(_0353_)
  );
  MUX2_X1 _2969_ (
    .A(_0351_),
    .B(_0353_),
    .S(io_in2[4]),
    .Z(_0354_)
  );
  AND2_X1 _2970_ (
    .A1(_0081_),
    .A2(_0354_),
    .ZN(_0355_)
  );
  INV_X1 _2971_ (
    .A(_0355_),
    .ZN(_0356_)
  );
  AND2_X1 _2972_ (
    .A1(_0347_),
    .A2(_0356_),
    .ZN(_0357_)
  );
  AND2_X1 _2973_ (
    .A1(_0345_),
    .A2(_0357_),
    .ZN(_0358_)
  );
  INV_X1 _2974_ (
    .A(_0358_),
    .ZN(io_out[5])
  );
  AND2_X1 _2975_ (
    .A1(_1444_),
    .A2(_1448_),
    .ZN(_0359_)
  );
  INV_X1 _2976_ (
    .A(_0359_),
    .ZN(_0361_)
  );
  AND2_X1 _2977_ (
    .A1(_1450_),
    .A2(_0361_),
    .ZN(io_adder_out[6])
  );
  AND2_X1 _2978_ (
    .A1(_0171_),
    .A2(io_adder_out[6]),
    .ZN(_0362_)
  );
  INV_X1 _2979_ (
    .A(_0362_),
    .ZN(_0363_)
  );
  MUX2_X1 _2980_ (
    .A(_0246_),
    .B(_0248_),
    .S(io_in2[2]),
    .Z(_0364_)
  );
  MUX2_X1 _2981_ (
    .A(_0249_),
    .B(_0252_),
    .S(io_in2[2]),
    .Z(_0365_)
  );
  MUX2_X1 _2982_ (
    .A(_0364_),
    .B(_0365_),
    .S(io_in2[3]),
    .Z(_0366_)
  );
  MUX2_X1 _2983_ (
    .A(_0253_),
    .B(_0255_),
    .S(io_in2[2]),
    .Z(_0367_)
  );
  MUX2_X1 _2984_ (
    .A(_0190_),
    .B(_0367_),
    .S(_0401_),
    .Z(_0368_)
  );
  MUX2_X1 _2985_ (
    .A(_0366_),
    .B(_0368_),
    .S(io_in2[4]),
    .Z(_0369_)
  );
  AND2_X1 _2986_ (
    .A1(_0081_),
    .A2(_0369_),
    .ZN(_0371_)
  );
  INV_X1 _2987_ (
    .A(_0371_),
    .ZN(_0372_)
  );
  MUX2_X1 _2988_ (
    .A(_0159_),
    .B(_0222_),
    .S(_0401_),
    .Z(_0373_)
  );
  MUX2_X1 _2989_ (
    .A(_0159_),
    .B(_0373_),
    .S(_0412_),
    .Z(_0374_)
  );
  AND2_X1 _2990_ (
    .A1(_0166_),
    .A2(_0374_),
    .ZN(_0375_)
  );
  INV_X1 _2991_ (
    .A(_0375_),
    .ZN(_0376_)
  );
  AND2_X1 _2992_ (
    .A1(io_in2[6]),
    .A2(io_in1[6]),
    .ZN(_0377_)
  );
  AND2_X1 _2993_ (
    .A1(_0174_),
    .A2(_0377_),
    .ZN(_0378_)
  );
  INV_X1 _2994_ (
    .A(_0378_),
    .ZN(_0379_)
  );
  AND2_X1 _2995_ (
    .A1(_1198_),
    .A2(_0178_),
    .ZN(_0380_)
  );
  INV_X1 _2996_ (
    .A(_0380_),
    .ZN(_0382_)
  );
  AND2_X1 _2997_ (
    .A1(_0379_),
    .A2(_0382_),
    .ZN(_0383_)
  );
  AND2_X1 _2998_ (
    .A1(_0376_),
    .A2(_0383_),
    .ZN(_0384_)
  );
  AND2_X1 _2999_ (
    .A1(_0372_),
    .A2(_0384_),
    .ZN(_0385_)
  );
  AND2_X1 _3000_ (
    .A1(_0363_),
    .A2(_0385_),
    .ZN(_0386_)
  );
  INV_X1 _3001_ (
    .A(_0386_),
    .ZN(io_out[6])
  );
  AND2_X1 _3002_ (
    .A1(_1450_),
    .A2(_1454_),
    .ZN(_0387_)
  );
  INV_X1 _3003_ (
    .A(_0387_),
    .ZN(_0388_)
  );
  AND2_X1 _3004_ (
    .A1(_1456_),
    .A2(_0388_),
    .ZN(io_adder_out[7])
  );
  AND2_X1 _3005_ (
    .A1(_0171_),
    .A2(io_adder_out[7]),
    .ZN(_0389_)
  );
  INV_X1 _3006_ (
    .A(_0389_),
    .ZN(_0391_)
  );
  MUX2_X1 _3007_ (
    .A(_0280_),
    .B(_0282_),
    .S(io_in2[2]),
    .Z(_0392_)
  );
  MUX2_X1 _3008_ (
    .A(_0283_),
    .B(_0286_),
    .S(io_in2[2]),
    .Z(_0393_)
  );
  MUX2_X1 _3009_ (
    .A(_0392_),
    .B(_0393_),
    .S(io_in2[3]),
    .Z(_0394_)
  );
  MUX2_X1 _3010_ (
    .A(_0287_),
    .B(_0289_),
    .S(io_in2[2]),
    .Z(_0395_)
  );
  MUX2_X1 _3011_ (
    .A(_0160_),
    .B(_0395_),
    .S(_0401_),
    .Z(_0396_)
  );
  MUX2_X1 _3012_ (
    .A(_0394_),
    .B(_0396_),
    .S(io_in2[4]),
    .Z(_0397_)
  );
  AND2_X1 _3013_ (
    .A1(_0081_),
    .A2(_0397_),
    .ZN(_0398_)
  );
  INV_X1 _3014_ (
    .A(_0398_),
    .ZN(_0399_)
  );
  MUX2_X1 _3015_ (
    .A(_0152_),
    .B(_0159_),
    .S(io_in2[3]),
    .Z(_0400_)
  );
  MUX2_X1 _3016_ (
    .A(_0159_),
    .B(_0400_),
    .S(_0412_),
    .Z(_0402_)
  );
  AND2_X1 _3017_ (
    .A1(_0166_),
    .A2(_0402_),
    .ZN(_0403_)
  );
  INV_X1 _3018_ (
    .A(_0403_),
    .ZN(_0404_)
  );
  AND2_X1 _3019_ (
    .A1(_1182_),
    .A2(_0178_),
    .ZN(_0405_)
  );
  INV_X1 _3020_ (
    .A(_0405_),
    .ZN(_0406_)
  );
  AND2_X1 _3021_ (
    .A1(io_in2[7]),
    .A2(io_in1[7]),
    .ZN(_0407_)
  );
  AND2_X1 _3022_ (
    .A1(_0174_),
    .A2(_0407_),
    .ZN(_0408_)
  );
  INV_X1 _3023_ (
    .A(_0408_),
    .ZN(_0409_)
  );
  AND2_X1 _3024_ (
    .A1(_0406_),
    .A2(_0409_),
    .ZN(_0410_)
  );
  AND2_X1 _3025_ (
    .A1(_0404_),
    .A2(_0410_),
    .ZN(_0411_)
  );
  AND2_X1 _3026_ (
    .A1(_0399_),
    .A2(_0411_),
    .ZN(_0413_)
  );
  AND2_X1 _3027_ (
    .A1(_0391_),
    .A2(_0413_),
    .ZN(_0414_)
  );
  INV_X1 _3028_ (
    .A(_0414_),
    .ZN(io_out[7])
  );
  AND2_X1 _3029_ (
    .A1(_1412_),
    .A2(_1456_),
    .ZN(_0415_)
  );
  INV_X1 _3030_ (
    .A(_0415_),
    .ZN(_0416_)
  );
  AND2_X1 _3031_ (
    .A1(_1458_),
    .A2(_0416_),
    .ZN(io_adder_out[8])
  );
  AND2_X1 _3032_ (
    .A1(_0171_),
    .A2(io_adder_out[8]),
    .ZN(_0417_)
  );
  INV_X1 _3033_ (
    .A(_0417_),
    .ZN(_0418_)
  );
  MUX2_X1 _3034_ (
    .A(_0159_),
    .B(_0396_),
    .S(_0412_),
    .Z(_0419_)
  );
  AND2_X1 _3035_ (
    .A1(_0166_),
    .A2(_0419_),
    .ZN(_0420_)
  );
  INV_X1 _3036_ (
    .A(_0420_),
    .ZN(_0422_)
  );
  MUX2_X1 _3037_ (
    .A(_0121_),
    .B(_0137_),
    .S(io_in2[3]),
    .Z(_0423_)
  );
  MUX2_X1 _3038_ (
    .A(_0400_),
    .B(_0423_),
    .S(_0412_),
    .Z(_0424_)
  );
  AND2_X1 _3039_ (
    .A1(_0081_),
    .A2(_0424_),
    .ZN(_0425_)
  );
  INV_X1 _3040_ (
    .A(_0425_),
    .ZN(_0426_)
  );
  AND2_X1 _3041_ (
    .A1(_1314_),
    .A2(_0178_),
    .ZN(_0427_)
  );
  INV_X1 _3042_ (
    .A(_0427_),
    .ZN(_0428_)
  );
  AND2_X1 _3043_ (
    .A1(io_in2[8]),
    .A2(io_in1[8]),
    .ZN(_0429_)
  );
  AND2_X1 _3044_ (
    .A1(_0174_),
    .A2(_0429_),
    .ZN(_0430_)
  );
  INV_X1 _3045_ (
    .A(_0430_),
    .ZN(_0431_)
  );
  AND2_X1 _3046_ (
    .A1(_0422_),
    .A2(_0428_),
    .ZN(_0433_)
  );
  AND2_X1 _3047_ (
    .A1(_0426_),
    .A2(_0431_),
    .ZN(_0434_)
  );
  AND2_X1 _3048_ (
    .A1(_0433_),
    .A2(_0434_),
    .ZN(_0435_)
  );
  AND2_X1 _3049_ (
    .A1(_0418_),
    .A2(_0435_),
    .ZN(_0436_)
  );
  INV_X1 _3050_ (
    .A(_0436_),
    .ZN(io_out[8])
  );
  AND2_X1 _3051_ (
    .A1(_1458_),
    .A2(_1462_),
    .ZN(_0437_)
  );
  INV_X1 _3052_ (
    .A(_0437_),
    .ZN(_0438_)
  );
  AND2_X1 _3053_ (
    .A1(_1464_),
    .A2(_0438_),
    .ZN(io_adder_out[9])
  );
  AND2_X1 _3054_ (
    .A1(_0171_),
    .A2(io_adder_out[9]),
    .ZN(_0439_)
  );
  INV_X1 _3055_ (
    .A(_0439_),
    .ZN(_0440_)
  );
  MUX2_X1 _3056_ (
    .A(_0159_),
    .B(_0368_),
    .S(_0412_),
    .Z(_0442_)
  );
  AND2_X1 _3057_ (
    .A1(_0166_),
    .A2(_0442_),
    .ZN(_0443_)
  );
  INV_X1 _3058_ (
    .A(_0443_),
    .ZN(_0444_)
  );
  MUX2_X1 _3059_ (
    .A(_0208_),
    .B(_0216_),
    .S(io_in2[3]),
    .Z(_0445_)
  );
  MUX2_X1 _3060_ (
    .A(_0373_),
    .B(_0445_),
    .S(_0412_),
    .Z(_0446_)
  );
  AND2_X1 _3061_ (
    .A1(_0081_),
    .A2(_0446_),
    .ZN(_0447_)
  );
  INV_X1 _3062_ (
    .A(_0447_),
    .ZN(_0448_)
  );
  AND2_X1 _3063_ (
    .A1(_1154_),
    .A2(_0178_),
    .ZN(_0449_)
  );
  INV_X1 _3064_ (
    .A(_0449_),
    .ZN(_0450_)
  );
  AND2_X1 _3065_ (
    .A1(io_in2[9]),
    .A2(io_in1[9]),
    .ZN(_0451_)
  );
  AND2_X1 _3066_ (
    .A1(_0174_),
    .A2(_0451_),
    .ZN(_0453_)
  );
  INV_X1 _3067_ (
    .A(_0453_),
    .ZN(_0454_)
  );
  AND2_X1 _3068_ (
    .A1(_0450_),
    .A2(_0454_),
    .ZN(_0455_)
  );
  AND2_X1 _3069_ (
    .A1(_0448_),
    .A2(_0455_),
    .ZN(_0456_)
  );
  AND2_X1 _3070_ (
    .A1(_0444_),
    .A2(_0456_),
    .ZN(_0457_)
  );
  AND2_X1 _3071_ (
    .A1(_0440_),
    .A2(_0457_),
    .ZN(_0458_)
  );
  INV_X1 _3072_ (
    .A(_0458_),
    .ZN(io_out[9])
  );
  AND2_X1 _3073_ (
    .A1(_1464_),
    .A2(_1468_),
    .ZN(_0459_)
  );
  INV_X1 _3074_ (
    .A(_0459_),
    .ZN(_0460_)
  );
  AND2_X1 _3075_ (
    .A1(_1470_),
    .A2(_0460_),
    .ZN(io_adder_out[10])
  );
  AND2_X1 _3076_ (
    .A1(_0171_),
    .A2(io_adder_out[10]),
    .ZN(_0462_)
  );
  INV_X1 _3077_ (
    .A(_0462_),
    .ZN(_0463_)
  );
  MUX2_X1 _3078_ (
    .A(_0250_),
    .B(_0254_),
    .S(io_in2[3]),
    .Z(_0464_)
  );
  MUX2_X1 _3079_ (
    .A(_0334_),
    .B(_0464_),
    .S(_0412_),
    .Z(_0465_)
  );
  AND2_X1 _3080_ (
    .A1(_0081_),
    .A2(_0465_),
    .ZN(_0466_)
  );
  INV_X1 _3081_ (
    .A(_0466_),
    .ZN(_0467_)
  );
  MUX2_X1 _3082_ (
    .A(_0159_),
    .B(_0353_),
    .S(_0412_),
    .Z(_0468_)
  );
  AND2_X1 _3083_ (
    .A1(_0166_),
    .A2(_0468_),
    .ZN(_0469_)
  );
  INV_X1 _3084_ (
    .A(_0469_),
    .ZN(_0470_)
  );
  AND2_X1 _3085_ (
    .A1(io_in2[10]),
    .A2(io_in1[10]),
    .ZN(_0471_)
  );
  AND2_X1 _3086_ (
    .A1(_0174_),
    .A2(_0471_),
    .ZN(_0473_)
  );
  INV_X1 _3087_ (
    .A(_0473_),
    .ZN(_0474_)
  );
  AND2_X1 _3088_ (
    .A1(_1138_),
    .A2(_0178_),
    .ZN(_0475_)
  );
  INV_X1 _3089_ (
    .A(_0475_),
    .ZN(_0476_)
  );
  AND2_X1 _3090_ (
    .A1(_0474_),
    .A2(_0476_),
    .ZN(_0477_)
  );
  AND2_X1 _3091_ (
    .A1(_0470_),
    .A2(_0477_),
    .ZN(_0478_)
  );
  AND2_X1 _3092_ (
    .A1(_0467_),
    .A2(_0478_),
    .ZN(_0479_)
  );
  AND2_X1 _3093_ (
    .A1(_0463_),
    .A2(_0479_),
    .ZN(_0480_)
  );
  INV_X1 _3094_ (
    .A(_0480_),
    .ZN(io_out[10])
  );
  AND2_X1 _3095_ (
    .A1(_1470_),
    .A2(_1481_),
    .ZN(_0481_)
  );
  INV_X1 _3096_ (
    .A(_0481_),
    .ZN(_0483_)
  );
  AND2_X1 _3097_ (
    .A1(_1484_),
    .A2(_0483_),
    .ZN(io_adder_out[11])
  );
  AND2_X1 _3098_ (
    .A1(_0171_),
    .A2(io_adder_out[11]),
    .ZN(_0484_)
  );
  INV_X1 _3099_ (
    .A(_0484_),
    .ZN(_0485_)
  );
  MUX2_X1 _3100_ (
    .A(_0284_),
    .B(_0288_),
    .S(io_in2[3]),
    .Z(_0486_)
  );
  MUX2_X1 _3101_ (
    .A(_0308_),
    .B(_0486_),
    .S(_0412_),
    .Z(_0487_)
  );
  AND2_X1 _3102_ (
    .A1(_0081_),
    .A2(_0487_),
    .ZN(_0488_)
  );
  INV_X1 _3103_ (
    .A(_0488_),
    .ZN(_0489_)
  );
  AND2_X1 _3104_ (
    .A1(_1122_),
    .A2(_0178_),
    .ZN(_0490_)
  );
  INV_X1 _3105_ (
    .A(_0490_),
    .ZN(_0491_)
  );
  AND2_X1 _3106_ (
    .A1(io_in2[11]),
    .A2(io_in1[11]),
    .ZN(_0493_)
  );
  AND2_X1 _3107_ (
    .A1(_0174_),
    .A2(_0493_),
    .ZN(_0494_)
  );
  INV_X1 _3108_ (
    .A(_0494_),
    .ZN(_0495_)
  );
  AND2_X1 _3109_ (
    .A1(_0491_),
    .A2(_0495_),
    .ZN(_0496_)
  );
  AND2_X1 _3110_ (
    .A1(_0489_),
    .A2(_0496_),
    .ZN(_0497_)
  );
  MUX2_X1 _3111_ (
    .A(_0159_),
    .B(_0316_),
    .S(_0412_),
    .Z(_0498_)
  );
  AND2_X1 _3112_ (
    .A1(_0166_),
    .A2(_0498_),
    .ZN(_0499_)
  );
  INV_X1 _3113_ (
    .A(_0499_),
    .ZN(_0500_)
  );
  AND2_X1 _3114_ (
    .A1(_0497_),
    .A2(_0500_),
    .ZN(_0501_)
  );
  AND2_X1 _3115_ (
    .A1(_0485_),
    .A2(_0501_),
    .ZN(_0502_)
  );
  INV_X1 _3116_ (
    .A(_0502_),
    .ZN(io_out[11])
  );
  AND2_X1 _3117_ (
    .A1(_1484_),
    .A2(_1488_),
    .ZN(_0504_)
  );
  INV_X1 _3118_ (
    .A(_0504_),
    .ZN(_0505_)
  );
  AND2_X1 _3119_ (
    .A1(_1490_),
    .A2(_0505_),
    .ZN(io_adder_out[12])
  );
  AND2_X1 _3120_ (
    .A1(_0171_),
    .A2(io_adder_out[12]),
    .ZN(_0506_)
  );
  INV_X1 _3121_ (
    .A(_0506_),
    .ZN(_0507_)
  );
  MUX2_X1 _3122_ (
    .A(_0313_),
    .B(_0315_),
    .S(io_in2[3]),
    .Z(_0508_)
  );
  MUX2_X1 _3123_ (
    .A(_0275_),
    .B(_0508_),
    .S(_0412_),
    .Z(_0509_)
  );
  AND2_X1 _3124_ (
    .A1(_0081_),
    .A2(_0509_),
    .ZN(_0510_)
  );
  INV_X1 _3125_ (
    .A(_0510_),
    .ZN(_0511_)
  );
  MUX2_X1 _3126_ (
    .A(_0159_),
    .B(_0291_),
    .S(_0412_),
    .Z(_0513_)
  );
  AND2_X1 _3127_ (
    .A1(_0166_),
    .A2(_0513_),
    .ZN(_0514_)
  );
  INV_X1 _3128_ (
    .A(_0514_),
    .ZN(_0515_)
  );
  AND2_X1 _3129_ (
    .A1(io_in2[12]),
    .A2(io_in1[12]),
    .ZN(_0516_)
  );
  AND2_X1 _3130_ (
    .A1(_0174_),
    .A2(_0516_),
    .ZN(_0517_)
  );
  INV_X1 _3131_ (
    .A(_0517_),
    .ZN(_0518_)
  );
  AND2_X1 _3132_ (
    .A1(_1106_),
    .A2(_0178_),
    .ZN(_0519_)
  );
  INV_X1 _3133_ (
    .A(_0519_),
    .ZN(_0520_)
  );
  AND2_X1 _3134_ (
    .A1(_0518_),
    .A2(_0520_),
    .ZN(_0521_)
  );
  AND2_X1 _3135_ (
    .A1(_0515_),
    .A2(_0521_),
    .ZN(_0522_)
  );
  AND2_X1 _3136_ (
    .A1(_0511_),
    .A2(_0522_),
    .ZN(_0524_)
  );
  AND2_X1 _3137_ (
    .A1(_0507_),
    .A2(_0524_),
    .ZN(_0525_)
  );
  INV_X1 _3138_ (
    .A(_0525_),
    .ZN(io_out[12])
  );
  AND2_X1 _3139_ (
    .A1(_1490_),
    .A2(_1501_),
    .ZN(_0526_)
  );
  INV_X1 _3140_ (
    .A(_0526_),
    .ZN(_0527_)
  );
  AND2_X1 _3141_ (
    .A1(_1504_),
    .A2(_0527_),
    .ZN(io_adder_out[13])
  );
  AND2_X1 _3142_ (
    .A1(_0171_),
    .A2(io_adder_out[13]),
    .ZN(_0528_)
  );
  INV_X1 _3143_ (
    .A(_0528_),
    .ZN(_0529_)
  );
  MUX2_X1 _3144_ (
    .A(_0349_),
    .B(_0352_),
    .S(io_in2[3]),
    .Z(_0530_)
  );
  MUX2_X1 _3145_ (
    .A(_0241_),
    .B(_0530_),
    .S(_0412_),
    .Z(_0531_)
  );
  AND2_X1 _3146_ (
    .A1(_0081_),
    .A2(_0531_),
    .ZN(_0533_)
  );
  INV_X1 _3147_ (
    .A(_0533_),
    .ZN(_0534_)
  );
  AND2_X1 _3148_ (
    .A1(_1090_),
    .A2(_0178_),
    .ZN(_0535_)
  );
  INV_X1 _3149_ (
    .A(_0535_),
    .ZN(_0536_)
  );
  AND2_X1 _3150_ (
    .A1(io_in2[13]),
    .A2(io_in1[13]),
    .ZN(_0537_)
  );
  AND2_X1 _3151_ (
    .A1(_0174_),
    .A2(_0537_),
    .ZN(_0538_)
  );
  INV_X1 _3152_ (
    .A(_0538_),
    .ZN(_0539_)
  );
  AND2_X1 _3153_ (
    .A1(_0536_),
    .A2(_0539_),
    .ZN(_0540_)
  );
  AND2_X1 _3154_ (
    .A1(_0534_),
    .A2(_0540_),
    .ZN(_0541_)
  );
  MUX2_X1 _3155_ (
    .A(_0159_),
    .B(_0257_),
    .S(_0412_),
    .Z(_0542_)
  );
  AND2_X1 _3156_ (
    .A1(_0166_),
    .A2(_0542_),
    .ZN(_0544_)
  );
  INV_X1 _3157_ (
    .A(_0544_),
    .ZN(_0545_)
  );
  AND2_X1 _3158_ (
    .A1(_0541_),
    .A2(_0545_),
    .ZN(_0546_)
  );
  AND2_X1 _3159_ (
    .A1(_0529_),
    .A2(_0546_),
    .ZN(_0547_)
  );
  INV_X1 _3160_ (
    .A(_0547_),
    .ZN(io_out[13])
  );
  AND2_X1 _3161_ (
    .A1(_1408_),
    .A2(_1504_),
    .ZN(_0548_)
  );
  INV_X1 _3162_ (
    .A(_0548_),
    .ZN(_0549_)
  );
  AND2_X1 _3163_ (
    .A1(_1506_),
    .A2(_0549_),
    .ZN(io_adder_out[14])
  );
  AND2_X1 _3164_ (
    .A1(_0171_),
    .A2(io_adder_out[14]),
    .ZN(_0550_)
  );
  INV_X1 _3165_ (
    .A(_0550_),
    .ZN(_0551_)
  );
  MUX2_X1 _3166_ (
    .A(_0365_),
    .B(_0367_),
    .S(io_in2[3]),
    .Z(_0553_)
  );
  MUX2_X1 _3167_ (
    .A(_0191_),
    .B(_0553_),
    .S(_0412_),
    .Z(_0554_)
  );
  AND2_X1 _3168_ (
    .A1(_0081_),
    .A2(_0554_),
    .ZN(_0555_)
  );
  INV_X1 _3169_ (
    .A(_0555_),
    .ZN(_0556_)
  );
  AND2_X1 _3170_ (
    .A1(_1074_),
    .A2(_0178_),
    .ZN(_0557_)
  );
  INV_X1 _3171_ (
    .A(_0557_),
    .ZN(_0558_)
  );
  AND2_X1 _3172_ (
    .A1(io_in2[14]),
    .A2(io_in1[14]),
    .ZN(_0559_)
  );
  AND2_X1 _3173_ (
    .A1(_0174_),
    .A2(_0559_),
    .ZN(_0560_)
  );
  INV_X1 _3174_ (
    .A(_0560_),
    .ZN(_0561_)
  );
  AND2_X1 _3175_ (
    .A1(_0558_),
    .A2(_0561_),
    .ZN(_0562_)
  );
  AND2_X1 _3176_ (
    .A1(_0556_),
    .A2(_0562_),
    .ZN(_0564_)
  );
  MUX2_X1 _3177_ (
    .A(_0159_),
    .B(_0223_),
    .S(_0412_),
    .Z(_0565_)
  );
  AND2_X1 _3178_ (
    .A1(_0166_),
    .A2(_0565_),
    .ZN(_0566_)
  );
  INV_X1 _3179_ (
    .A(_0566_),
    .ZN(_0567_)
  );
  AND2_X1 _3180_ (
    .A1(_0564_),
    .A2(_0567_),
    .ZN(_0568_)
  );
  AND2_X1 _3181_ (
    .A1(_0551_),
    .A2(_0568_),
    .ZN(_0569_)
  );
  INV_X1 _3182_ (
    .A(_0569_),
    .ZN(io_out[14])
  );
  AND2_X1 _3183_ (
    .A1(_1506_),
    .A2(_1517_),
    .ZN(_0570_)
  );
  INV_X1 _3184_ (
    .A(_0570_),
    .ZN(_0571_)
  );
  AND2_X1 _3185_ (
    .A1(_1520_),
    .A2(_0571_),
    .ZN(io_adder_out[15])
  );
  AND2_X1 _3186_ (
    .A1(_0171_),
    .A2(io_adder_out[15]),
    .ZN(_0573_)
  );
  INV_X1 _3187_ (
    .A(_0573_),
    .ZN(_0574_)
  );
  MUX2_X1 _3188_ (
    .A(_0393_),
    .B(_0395_),
    .S(io_in2[3]),
    .Z(_0575_)
  );
  MUX2_X1 _3189_ (
    .A(_0161_),
    .B(_0575_),
    .S(_0412_),
    .Z(_0576_)
  );
  AND2_X1 _3190_ (
    .A1(_0081_),
    .A2(_0576_),
    .ZN(_0577_)
  );
  INV_X1 _3191_ (
    .A(_0577_),
    .ZN(_0578_)
  );
  MUX2_X1 _3192_ (
    .A(_0153_),
    .B(_0159_),
    .S(io_in2[4]),
    .Z(_0579_)
  );
  AND2_X1 _3193_ (
    .A1(_0166_),
    .A2(_0579_),
    .ZN(_0580_)
  );
  INV_X1 _3194_ (
    .A(_0580_),
    .ZN(_0581_)
  );
  AND2_X1 _3195_ (
    .A1(_1058_),
    .A2(_0178_),
    .ZN(_0582_)
  );
  INV_X1 _3196_ (
    .A(_0582_),
    .ZN(_0584_)
  );
  AND2_X1 _3197_ (
    .A1(io_in2[15]),
    .A2(io_in1[15]),
    .ZN(_0585_)
  );
  AND2_X1 _3198_ (
    .A1(_0174_),
    .A2(_0585_),
    .ZN(_0586_)
  );
  INV_X1 _3199_ (
    .A(_0586_),
    .ZN(_0587_)
  );
  AND2_X1 _3200_ (
    .A1(_0581_),
    .A2(_0584_),
    .ZN(_0588_)
  );
  AND2_X1 _3201_ (
    .A1(_0578_),
    .A2(_0587_),
    .ZN(_0589_)
  );
  AND2_X1 _3202_ (
    .A1(_0588_),
    .A2(_0589_),
    .ZN(_0590_)
  );
  AND2_X1 _3203_ (
    .A1(_0574_),
    .A2(_0590_),
    .ZN(_0591_)
  );
  INV_X1 _3204_ (
    .A(_0591_),
    .ZN(io_out[15])
  );
  AND2_X1 _3205_ (
    .A1(_1404_),
    .A2(_1520_),
    .ZN(_0592_)
  );
  INV_X1 _3206_ (
    .A(_0592_),
    .ZN(_0594_)
  );
  AND2_X1 _3207_ (
    .A1(_1522_),
    .A2(_0594_),
    .ZN(io_adder_out[16])
  );
  AND2_X1 _3208_ (
    .A1(_0171_),
    .A2(io_adder_out[16]),
    .ZN(_0595_)
  );
  INV_X1 _3209_ (
    .A(_0595_),
    .ZN(_0596_)
  );
  AND2_X1 _3210_ (
    .A1(_0081_),
    .A2(_0579_),
    .ZN(_0597_)
  );
  INV_X1 _3211_ (
    .A(_0597_),
    .ZN(_0598_)
  );
  AND2_X1 _3212_ (
    .A1(_1355_),
    .A2(_0178_),
    .ZN(_0599_)
  );
  INV_X1 _3213_ (
    .A(_0599_),
    .ZN(_0600_)
  );
  AND2_X1 _3214_ (
    .A1(io_in2[16]),
    .A2(io_in1[16]),
    .ZN(_0601_)
  );
  AND2_X1 _3215_ (
    .A1(_0174_),
    .A2(_0601_),
    .ZN(_0602_)
  );
  INV_X1 _3216_ (
    .A(_0602_),
    .ZN(_0604_)
  );
  AND2_X1 _3217_ (
    .A1(_0600_),
    .A2(_0604_),
    .ZN(_0605_)
  );
  AND2_X1 _3218_ (
    .A1(_0598_),
    .A2(_0605_),
    .ZN(_0606_)
  );
  AND2_X1 _3219_ (
    .A1(_0166_),
    .A2(_0576_),
    .ZN(_0607_)
  );
  INV_X1 _3220_ (
    .A(_0607_),
    .ZN(_0608_)
  );
  AND2_X1 _3221_ (
    .A1(_0606_),
    .A2(_0608_),
    .ZN(_0609_)
  );
  AND2_X1 _3222_ (
    .A1(_0596_),
    .A2(_0609_),
    .ZN(_0610_)
  );
  INV_X1 _3223_ (
    .A(_0610_),
    .ZN(io_out[16])
  );
  AND2_X1 _3224_ (
    .A1(_1400_),
    .A2(_1522_),
    .ZN(_0611_)
  );
  INV_X1 _3225_ (
    .A(_0611_),
    .ZN(_0612_)
  );
  AND2_X1 _3226_ (
    .A1(_1524_),
    .A2(_0612_),
    .ZN(io_adder_out[17])
  );
  AND2_X1 _3227_ (
    .A1(_0171_),
    .A2(io_adder_out[17]),
    .ZN(_0614_)
  );
  INV_X1 _3228_ (
    .A(_0614_),
    .ZN(_0615_)
  );
  AND2_X1 _3229_ (
    .A1(_0166_),
    .A2(_0554_),
    .ZN(_0616_)
  );
  INV_X1 _3230_ (
    .A(_0616_),
    .ZN(_0617_)
  );
  AND2_X1 _3231_ (
    .A1(_0081_),
    .A2(_0565_),
    .ZN(_0618_)
  );
  INV_X1 _3232_ (
    .A(_0618_),
    .ZN(_0619_)
  );
  AND2_X1 _3233_ (
    .A1(io_in2[17]),
    .A2(io_in1[17]),
    .ZN(_0620_)
  );
  AND2_X1 _3234_ (
    .A1(_0174_),
    .A2(_0620_),
    .ZN(_0621_)
  );
  INV_X1 _3235_ (
    .A(_0621_),
    .ZN(_0622_)
  );
  AND2_X1 _3236_ (
    .A1(_1363_),
    .A2(_0178_),
    .ZN(_0624_)
  );
  INV_X1 _3237_ (
    .A(_0624_),
    .ZN(_0625_)
  );
  AND2_X1 _3238_ (
    .A1(_0622_),
    .A2(_0625_),
    .ZN(_0626_)
  );
  AND2_X1 _3239_ (
    .A1(_0619_),
    .A2(_0626_),
    .ZN(_0627_)
  );
  AND2_X1 _3240_ (
    .A1(_0617_),
    .A2(_0627_),
    .ZN(_0628_)
  );
  AND2_X1 _3241_ (
    .A1(_0615_),
    .A2(_0628_),
    .ZN(_0629_)
  );
  INV_X1 _3242_ (
    .A(_0629_),
    .ZN(io_out[17])
  );
  AND2_X1 _3243_ (
    .A1(_1524_),
    .A2(_1528_),
    .ZN(_0630_)
  );
  INV_X1 _3244_ (
    .A(_0630_),
    .ZN(_0631_)
  );
  AND2_X1 _3245_ (
    .A1(_1530_),
    .A2(_0631_),
    .ZN(io_adder_out[18])
  );
  AND2_X1 _3246_ (
    .A1(_0171_),
    .A2(io_adder_out[18]),
    .ZN(_0633_)
  );
  INV_X1 _3247_ (
    .A(_0633_),
    .ZN(_0634_)
  );
  AND2_X1 _3248_ (
    .A1(_0081_),
    .A2(_0542_),
    .ZN(_0635_)
  );
  INV_X1 _3249_ (
    .A(_0635_),
    .ZN(_0636_)
  );
  AND2_X1 _3250_ (
    .A1(_1018_),
    .A2(_0178_),
    .ZN(_0637_)
  );
  INV_X1 _3251_ (
    .A(_0637_),
    .ZN(_0638_)
  );
  AND2_X1 _3252_ (
    .A1(io_in2[18]),
    .A2(io_in1[18]),
    .ZN(_0639_)
  );
  AND2_X1 _3253_ (
    .A1(_0174_),
    .A2(_0639_),
    .ZN(_0640_)
  );
  INV_X1 _3254_ (
    .A(_0640_),
    .ZN(_0641_)
  );
  AND2_X1 _3255_ (
    .A1(_0638_),
    .A2(_0641_),
    .ZN(_0642_)
  );
  AND2_X1 _3256_ (
    .A1(_0636_),
    .A2(_0642_),
    .ZN(_0644_)
  );
  AND2_X1 _3257_ (
    .A1(_0166_),
    .A2(_0531_),
    .ZN(_0645_)
  );
  INV_X1 _3258_ (
    .A(_0645_),
    .ZN(_0646_)
  );
  AND2_X1 _3259_ (
    .A1(_0644_),
    .A2(_0646_),
    .ZN(_0647_)
  );
  AND2_X1 _3260_ (
    .A1(_0634_),
    .A2(_0647_),
    .ZN(_0648_)
  );
  INV_X1 _3261_ (
    .A(_0648_),
    .ZN(io_out[18])
  );
  AND2_X1 _3262_ (
    .A1(_1530_),
    .A2(_1534_),
    .ZN(_0649_)
  );
  INV_X1 _3263_ (
    .A(_0649_),
    .ZN(_0650_)
  );
  AND2_X1 _3264_ (
    .A1(_1536_),
    .A2(_0650_),
    .ZN(io_adder_out[19])
  );
  AND2_X1 _3265_ (
    .A1(_0171_),
    .A2(io_adder_out[19]),
    .ZN(_0651_)
  );
  INV_X1 _3266_ (
    .A(_0651_),
    .ZN(_0653_)
  );
  AND2_X1 _3267_ (
    .A1(_0081_),
    .A2(_0513_),
    .ZN(_0654_)
  );
  INV_X1 _3268_ (
    .A(_0654_),
    .ZN(_0655_)
  );
  AND2_X1 _3269_ (
    .A1(_1002_),
    .A2(_0178_),
    .ZN(_0656_)
  );
  INV_X1 _3270_ (
    .A(_0656_),
    .ZN(_0657_)
  );
  AND2_X1 _3271_ (
    .A1(io_in2[19]),
    .A2(io_in1[19]),
    .ZN(_0658_)
  );
  AND2_X1 _3272_ (
    .A1(_0174_),
    .A2(_0658_),
    .ZN(_0659_)
  );
  INV_X1 _3273_ (
    .A(_0659_),
    .ZN(_0660_)
  );
  AND2_X1 _3274_ (
    .A1(_0657_),
    .A2(_0660_),
    .ZN(_0661_)
  );
  AND2_X1 _3275_ (
    .A1(_0655_),
    .A2(_0661_),
    .ZN(_0662_)
  );
  AND2_X1 _3276_ (
    .A1(_0166_),
    .A2(_0509_),
    .ZN(_0664_)
  );
  INV_X1 _3277_ (
    .A(_0664_),
    .ZN(_0665_)
  );
  AND2_X1 _3278_ (
    .A1(_0662_),
    .A2(_0665_),
    .ZN(_0666_)
  );
  AND2_X1 _3279_ (
    .A1(_0653_),
    .A2(_0666_),
    .ZN(_0667_)
  );
  INV_X1 _3280_ (
    .A(_0667_),
    .ZN(io_out[19])
  );
  AND2_X1 _3281_ (
    .A1(_1396_),
    .A2(_1536_),
    .ZN(_0668_)
  );
  INV_X1 _3282_ (
    .A(_0668_),
    .ZN(_0669_)
  );
  AND2_X1 _3283_ (
    .A1(_1538_),
    .A2(_0669_),
    .ZN(io_adder_out[20])
  );
  AND2_X1 _3284_ (
    .A1(_0171_),
    .A2(io_adder_out[20]),
    .ZN(_0670_)
  );
  INV_X1 _3285_ (
    .A(_0670_),
    .ZN(_0671_)
  );
  AND2_X1 _3286_ (
    .A1(_0081_),
    .A2(_0498_),
    .ZN(_0673_)
  );
  INV_X1 _3287_ (
    .A(_0673_),
    .ZN(_0674_)
  );
  AND2_X1 _3288_ (
    .A1(_0986_),
    .A2(_0178_),
    .ZN(_0675_)
  );
  INV_X1 _3289_ (
    .A(_0675_),
    .ZN(_0676_)
  );
  AND2_X1 _3290_ (
    .A1(io_in2[20]),
    .A2(io_in1[20]),
    .ZN(_0677_)
  );
  AND2_X1 _3291_ (
    .A1(_0174_),
    .A2(_0677_),
    .ZN(_0678_)
  );
  INV_X1 _3292_ (
    .A(_0678_),
    .ZN(_0679_)
  );
  AND2_X1 _3293_ (
    .A1(_0676_),
    .A2(_0679_),
    .ZN(_0680_)
  );
  AND2_X1 _3294_ (
    .A1(_0674_),
    .A2(_0680_),
    .ZN(_0681_)
  );
  AND2_X1 _3295_ (
    .A1(_0166_),
    .A2(_0487_),
    .ZN(_0682_)
  );
  INV_X1 _3296_ (
    .A(_0682_),
    .ZN(_0684_)
  );
  AND2_X1 _3297_ (
    .A1(_0681_),
    .A2(_0684_),
    .ZN(_0685_)
  );
  AND2_X1 _3298_ (
    .A1(_0671_),
    .A2(_0685_),
    .ZN(_0686_)
  );
  INV_X1 _3299_ (
    .A(_0686_),
    .ZN(io_out[20])
  );
  AND2_X1 _3300_ (
    .A1(_1538_),
    .A2(_1549_),
    .ZN(_0687_)
  );
  INV_X1 _3301_ (
    .A(_0687_),
    .ZN(_0688_)
  );
  AND2_X1 _3302_ (
    .A1(_1552_),
    .A2(_0688_),
    .ZN(io_adder_out[21])
  );
  AND2_X1 _3303_ (
    .A1(_0171_),
    .A2(io_adder_out[21]),
    .ZN(_0689_)
  );
  INV_X1 _3304_ (
    .A(_0689_),
    .ZN(_0690_)
  );
  AND2_X1 _3305_ (
    .A1(_0081_),
    .A2(_0468_),
    .ZN(_0691_)
  );
  INV_X1 _3306_ (
    .A(_0691_),
    .ZN(_0693_)
  );
  AND2_X1 _3307_ (
    .A1(_1539_),
    .A2(_0178_),
    .ZN(_0694_)
  );
  INV_X1 _3308_ (
    .A(_0694_),
    .ZN(_0695_)
  );
  AND2_X1 _3309_ (
    .A1(io_in2[21]),
    .A2(io_in1[21]),
    .ZN(_0696_)
  );
  AND2_X1 _3310_ (
    .A1(_0174_),
    .A2(_0696_),
    .ZN(_0697_)
  );
  INV_X1 _3311_ (
    .A(_0697_),
    .ZN(_0698_)
  );
  AND2_X1 _3312_ (
    .A1(_0695_),
    .A2(_0698_),
    .ZN(_0699_)
  );
  AND2_X1 _3313_ (
    .A1(_0693_),
    .A2(_0699_),
    .ZN(_0700_)
  );
  AND2_X1 _3314_ (
    .A1(_0166_),
    .A2(_0465_),
    .ZN(_0701_)
  );
  INV_X1 _3315_ (
    .A(_0701_),
    .ZN(_0702_)
  );
  AND2_X1 _3316_ (
    .A1(_0700_),
    .A2(_0702_),
    .ZN(_0704_)
  );
  AND2_X1 _3317_ (
    .A1(_0690_),
    .A2(_0704_),
    .ZN(_0705_)
  );
  INV_X1 _3318_ (
    .A(_0705_),
    .ZN(io_out[21])
  );
  AND2_X1 _3319_ (
    .A1(_1392_),
    .A2(_1552_),
    .ZN(_0706_)
  );
  INV_X1 _3320_ (
    .A(_0706_),
    .ZN(_0707_)
  );
  AND2_X1 _3321_ (
    .A1(_1554_),
    .A2(_0707_),
    .ZN(io_adder_out[22])
  );
  AND2_X1 _3322_ (
    .A1(_0171_),
    .A2(io_adder_out[22]),
    .ZN(_0708_)
  );
  INV_X1 _3323_ (
    .A(_0708_),
    .ZN(_0709_)
  );
  AND2_X1 _3324_ (
    .A1(_0081_),
    .A2(_0442_),
    .ZN(_0710_)
  );
  INV_X1 _3325_ (
    .A(_0710_),
    .ZN(_0711_)
  );
  AND2_X1 _3326_ (
    .A1(_0166_),
    .A2(_0446_),
    .ZN(_0713_)
  );
  INV_X1 _3327_ (
    .A(_0713_),
    .ZN(_0714_)
  );
  AND2_X1 _3328_ (
    .A1(io_in2[22]),
    .A2(io_in1[22]),
    .ZN(_0715_)
  );
  AND2_X1 _3329_ (
    .A1(_0174_),
    .A2(_0715_),
    .ZN(_0716_)
  );
  INV_X1 _3330_ (
    .A(_0716_),
    .ZN(_0717_)
  );
  AND2_X1 _3331_ (
    .A1(_0956_),
    .A2(_0178_),
    .ZN(_0718_)
  );
  INV_X1 _3332_ (
    .A(_0718_),
    .ZN(_0719_)
  );
  AND2_X1 _3333_ (
    .A1(_0717_),
    .A2(_0719_),
    .ZN(_0720_)
  );
  AND2_X1 _3334_ (
    .A1(_0714_),
    .A2(_0720_),
    .ZN(_0721_)
  );
  AND2_X1 _3335_ (
    .A1(_0711_),
    .A2(_0721_),
    .ZN(_0722_)
  );
  AND2_X1 _3336_ (
    .A1(_0709_),
    .A2(_0722_),
    .ZN(_0724_)
  );
  INV_X1 _3337_ (
    .A(_0724_),
    .ZN(io_out[22])
  );
  AND2_X1 _3338_ (
    .A1(_1554_),
    .A2(_1582_),
    .ZN(_0725_)
  );
  INV_X1 _3339_ (
    .A(_0725_),
    .ZN(_0726_)
  );
  AND2_X1 _3340_ (
    .A1(_1584_),
    .A2(_0726_),
    .ZN(io_adder_out[23])
  );
  AND2_X1 _3341_ (
    .A1(_0171_),
    .A2(io_adder_out[23]),
    .ZN(_0727_)
  );
  INV_X1 _3342_ (
    .A(_0727_),
    .ZN(_0728_)
  );
  AND2_X1 _3343_ (
    .A1(_0081_),
    .A2(_0419_),
    .ZN(_0729_)
  );
  INV_X1 _3344_ (
    .A(_0729_),
    .ZN(_0730_)
  );
  AND2_X1 _3345_ (
    .A1(_0166_),
    .A2(_0424_),
    .ZN(_0731_)
  );
  INV_X1 _3346_ (
    .A(_0731_),
    .ZN(_0733_)
  );
  AND2_X1 _3347_ (
    .A1(_1569_),
    .A2(_0178_),
    .ZN(_0734_)
  );
  INV_X1 _3348_ (
    .A(_0734_),
    .ZN(_0735_)
  );
  AND2_X1 _3349_ (
    .A1(io_in2[23]),
    .A2(io_in1[23]),
    .ZN(_0736_)
  );
  AND2_X1 _3350_ (
    .A1(_0174_),
    .A2(_0736_),
    .ZN(_0737_)
  );
  INV_X1 _3351_ (
    .A(_0737_),
    .ZN(_0738_)
  );
  AND2_X1 _3352_ (
    .A1(_0735_),
    .A2(_0738_),
    .ZN(_0739_)
  );
  AND2_X1 _3353_ (
    .A1(_0733_),
    .A2(_0739_),
    .ZN(_0740_)
  );
  AND2_X1 _3354_ (
    .A1(_0730_),
    .A2(_0740_),
    .ZN(_0741_)
  );
  AND2_X1 _3355_ (
    .A1(_0728_),
    .A2(_0741_),
    .ZN(_0742_)
  );
  INV_X1 _3356_ (
    .A(_0742_),
    .ZN(io_out[23])
  );
  AND2_X1 _3357_ (
    .A1(_1584_),
    .A2(_1612_),
    .ZN(_0744_)
  );
  INV_X1 _3358_ (
    .A(_0744_),
    .ZN(_0745_)
  );
  AND2_X1 _3359_ (
    .A1(_1614_),
    .A2(_0745_),
    .ZN(io_adder_out[24])
  );
  AND2_X1 _3360_ (
    .A1(_0171_),
    .A2(io_adder_out[24]),
    .ZN(_0746_)
  );
  INV_X1 _3361_ (
    .A(_0746_),
    .ZN(_0747_)
  );
  AND2_X1 _3362_ (
    .A1(_0081_),
    .A2(_0402_),
    .ZN(_0748_)
  );
  INV_X1 _3363_ (
    .A(_0748_),
    .ZN(_0749_)
  );
  AND2_X1 _3364_ (
    .A1(_1599_),
    .A2(_0178_),
    .ZN(_0750_)
  );
  INV_X1 _3365_ (
    .A(_0750_),
    .ZN(_0751_)
  );
  AND2_X1 _3366_ (
    .A1(io_in2[24]),
    .A2(io_in1[24]),
    .ZN(_0753_)
  );
  AND2_X1 _3367_ (
    .A1(_0174_),
    .A2(_0753_),
    .ZN(_0754_)
  );
  INV_X1 _3368_ (
    .A(_0754_),
    .ZN(_0755_)
  );
  AND2_X1 _3369_ (
    .A1(_0751_),
    .A2(_0755_),
    .ZN(_0756_)
  );
  AND2_X1 _3370_ (
    .A1(_0749_),
    .A2(_0756_),
    .ZN(_0757_)
  );
  AND2_X1 _3371_ (
    .A1(_0166_),
    .A2(_0397_),
    .ZN(_0758_)
  );
  INV_X1 _3372_ (
    .A(_0758_),
    .ZN(_0759_)
  );
  AND2_X1 _3373_ (
    .A1(_0757_),
    .A2(_0759_),
    .ZN(_0760_)
  );
  AND2_X1 _3374_ (
    .A1(_0747_),
    .A2(_0760_),
    .ZN(_0761_)
  );
  INV_X1 _3375_ (
    .A(_0761_),
    .ZN(io_out[24])
  );
  AND2_X1 _3376_ (
    .A1(_1614_),
    .A2(_1638_),
    .ZN(_0763_)
  );
  INV_X1 _3377_ (
    .A(_0763_),
    .ZN(_0764_)
  );
  AND2_X1 _3378_ (
    .A1(_1640_),
    .A2(_0764_),
    .ZN(io_adder_out[25])
  );
  AND2_X1 _3379_ (
    .A1(_0171_),
    .A2(io_adder_out[25]),
    .ZN(_0765_)
  );
  INV_X1 _3380_ (
    .A(_0765_),
    .ZN(_0766_)
  );
  AND2_X1 _3381_ (
    .A1(_0081_),
    .A2(_0374_),
    .ZN(_0767_)
  );
  INV_X1 _3382_ (
    .A(_0767_),
    .ZN(_0768_)
  );
  AND2_X1 _3383_ (
    .A1(_1629_),
    .A2(_0178_),
    .ZN(_0769_)
  );
  INV_X1 _3384_ (
    .A(_0769_),
    .ZN(_0770_)
  );
  AND2_X1 _3385_ (
    .A1(io_in2[25]),
    .A2(io_in1[25]),
    .ZN(_0771_)
  );
  AND2_X1 _3386_ (
    .A1(_0174_),
    .A2(_0771_),
    .ZN(_0773_)
  );
  INV_X1 _3387_ (
    .A(_0773_),
    .ZN(_0774_)
  );
  AND2_X1 _3388_ (
    .A1(_0770_),
    .A2(_0774_),
    .ZN(_0775_)
  );
  AND2_X1 _3389_ (
    .A1(_0768_),
    .A2(_0775_),
    .ZN(_0776_)
  );
  AND2_X1 _3390_ (
    .A1(_0166_),
    .A2(_0369_),
    .ZN(_0777_)
  );
  INV_X1 _3391_ (
    .A(_0777_),
    .ZN(_0778_)
  );
  AND2_X1 _3392_ (
    .A1(_0776_),
    .A2(_0778_),
    .ZN(_0779_)
  );
  AND2_X1 _3393_ (
    .A1(_0766_),
    .A2(_0779_),
    .ZN(_0780_)
  );
  INV_X1 _3394_ (
    .A(_0780_),
    .ZN(io_out[25])
  );
  AND2_X1 _3395_ (
    .A1(_1640_),
    .A2(_1664_),
    .ZN(_0781_)
  );
  INV_X1 _3396_ (
    .A(_0781_),
    .ZN(_0783_)
  );
  AND2_X1 _3397_ (
    .A1(_1666_),
    .A2(_0783_),
    .ZN(io_adder_out[26])
  );
  AND2_X1 _3398_ (
    .A1(_0171_),
    .A2(io_adder_out[26]),
    .ZN(_0784_)
  );
  INV_X1 _3399_ (
    .A(_0784_),
    .ZN(_0785_)
  );
  AND2_X1 _3400_ (
    .A1(_0081_),
    .A2(_0335_),
    .ZN(_0786_)
  );
  INV_X1 _3401_ (
    .A(_0786_),
    .ZN(_0787_)
  );
  AND2_X1 _3402_ (
    .A1(_0166_),
    .A2(_0354_),
    .ZN(_0788_)
  );
  INV_X1 _3403_ (
    .A(_0788_),
    .ZN(_0789_)
  );
  AND2_X1 _3404_ (
    .A1(_1655_),
    .A2(_0178_),
    .ZN(_0790_)
  );
  INV_X1 _3405_ (
    .A(_0790_),
    .ZN(_0791_)
  );
  AND2_X1 _3406_ (
    .A1(io_in2[26]),
    .A2(io_in1[26]),
    .ZN(_0793_)
  );
  AND2_X1 _3407_ (
    .A1(_0174_),
    .A2(_0793_),
    .ZN(_0794_)
  );
  INV_X1 _3408_ (
    .A(_0794_),
    .ZN(_0795_)
  );
  AND2_X1 _3409_ (
    .A1(_0791_),
    .A2(_0795_),
    .ZN(_0796_)
  );
  AND2_X1 _3410_ (
    .A1(_0789_),
    .A2(_0796_),
    .ZN(_0797_)
  );
  AND2_X1 _3411_ (
    .A1(_0787_),
    .A2(_0797_),
    .ZN(_0798_)
  );
  AND2_X1 _3412_ (
    .A1(_0785_),
    .A2(_0798_),
    .ZN(_0799_)
  );
  INV_X1 _3413_ (
    .A(_0799_),
    .ZN(io_out[26])
  );
  AND2_X1 _3414_ (
    .A1(_1666_),
    .A2(_1690_),
    .ZN(_0800_)
  );
  INV_X1 _3415_ (
    .A(_0800_),
    .ZN(_0801_)
  );
  AND2_X1 _3416_ (
    .A1(_1692_),
    .A2(_0801_),
    .ZN(io_adder_out[27])
  );
  AND2_X1 _3417_ (
    .A1(_0171_),
    .A2(io_adder_out[27]),
    .ZN(_0803_)
  );
  INV_X1 _3418_ (
    .A(_0803_),
    .ZN(_0804_)
  );
  AND2_X1 _3419_ (
    .A1(_0081_),
    .A2(_0309_),
    .ZN(_0805_)
  );
  INV_X1 _3420_ (
    .A(_0805_),
    .ZN(_0806_)
  );
  AND2_X1 _3421_ (
    .A1(_1681_),
    .A2(_0178_),
    .ZN(_0807_)
  );
  INV_X1 _3422_ (
    .A(_0807_),
    .ZN(_0808_)
  );
  AND2_X1 _3423_ (
    .A1(io_in2[27]),
    .A2(io_in1[27]),
    .ZN(_0809_)
  );
  AND2_X1 _3424_ (
    .A1(_0174_),
    .A2(_0809_),
    .ZN(_0810_)
  );
  INV_X1 _3425_ (
    .A(_0810_),
    .ZN(_0811_)
  );
  AND2_X1 _3426_ (
    .A1(_0808_),
    .A2(_0811_),
    .ZN(_0813_)
  );
  AND2_X1 _3427_ (
    .A1(_0806_),
    .A2(_0813_),
    .ZN(_0814_)
  );
  AND2_X1 _3428_ (
    .A1(_0166_),
    .A2(_0317_),
    .ZN(_0815_)
  );
  INV_X1 _3429_ (
    .A(_0815_),
    .ZN(_0816_)
  );
  AND2_X1 _3430_ (
    .A1(_0814_),
    .A2(_0816_),
    .ZN(_0817_)
  );
  AND2_X1 _3431_ (
    .A1(_0804_),
    .A2(_0817_),
    .ZN(_0818_)
  );
  INV_X1 _3432_ (
    .A(_0818_),
    .ZN(io_out[27])
  );
  AND2_X1 _3433_ (
    .A1(_1692_),
    .A2(_1716_),
    .ZN(_0819_)
  );
  INV_X1 _3434_ (
    .A(_0819_),
    .ZN(_0820_)
  );
  AND2_X1 _3435_ (
    .A1(_1718_),
    .A2(_0820_),
    .ZN(io_adder_out[28])
  );
  AND2_X1 _3436_ (
    .A1(_0171_),
    .A2(io_adder_out[28]),
    .ZN(_0822_)
  );
  INV_X1 _3437_ (
    .A(_0822_),
    .ZN(_0823_)
  );
  AND2_X1 _3438_ (
    .A1(_0081_),
    .A2(_0276_),
    .ZN(_0824_)
  );
  INV_X1 _3439_ (
    .A(_0824_),
    .ZN(_0825_)
  );
  AND2_X1 _3440_ (
    .A1(_1709_),
    .A2(_0178_),
    .ZN(_0826_)
  );
  INV_X1 _3441_ (
    .A(_0826_),
    .ZN(_0827_)
  );
  AND2_X1 _3442_ (
    .A1(io_in2[28]),
    .A2(io_in1[28]),
    .ZN(_0828_)
  );
  AND2_X1 _3443_ (
    .A1(_0174_),
    .A2(_0828_),
    .ZN(_0829_)
  );
  INV_X1 _3444_ (
    .A(_0829_),
    .ZN(_0830_)
  );
  AND2_X1 _3445_ (
    .A1(_0827_),
    .A2(_0830_),
    .ZN(_0831_)
  );
  AND2_X1 _3446_ (
    .A1(_0825_),
    .A2(_0831_),
    .ZN(_0833_)
  );
  AND2_X1 _3447_ (
    .A1(_0166_),
    .A2(_0292_),
    .ZN(_0834_)
  );
  INV_X1 _3448_ (
    .A(_0834_),
    .ZN(_0835_)
  );
  AND2_X1 _3449_ (
    .A1(_0833_),
    .A2(_0835_),
    .ZN(_0836_)
  );
  AND2_X1 _3450_ (
    .A1(_0823_),
    .A2(_0836_),
    .ZN(_0837_)
  );
  INV_X1 _3451_ (
    .A(_0837_),
    .ZN(io_out[28])
  );
  AND2_X1 _3452_ (
    .A1(_1718_),
    .A2(_0002_),
    .ZN(_0838_)
  );
  INV_X1 _3453_ (
    .A(_0838_),
    .ZN(_0839_)
  );
  AND2_X1 _3454_ (
    .A1(_0004_),
    .A2(_0839_),
    .ZN(io_adder_out[29])
  );
  AND2_X1 _3455_ (
    .A1(_0171_),
    .A2(io_adder_out[29]),
    .ZN(_0840_)
  );
  INV_X1 _3456_ (
    .A(_0840_),
    .ZN(_0842_)
  );
  AND2_X1 _3457_ (
    .A1(_0166_),
    .A2(_0258_),
    .ZN(_0843_)
  );
  INV_X1 _3458_ (
    .A(_0843_),
    .ZN(_0844_)
  );
  AND2_X1 _3459_ (
    .A1(_0081_),
    .A2(_0242_),
    .ZN(_0845_)
  );
  INV_X1 _3460_ (
    .A(_0845_),
    .ZN(_0846_)
  );
  AND2_X1 _3461_ (
    .A1(_1733_),
    .A2(_0178_),
    .ZN(_0847_)
  );
  INV_X1 _3462_ (
    .A(_0847_),
    .ZN(_0848_)
  );
  AND2_X1 _3463_ (
    .A1(io_in2[29]),
    .A2(io_in1[29]),
    .ZN(_0849_)
  );
  AND2_X1 _3464_ (
    .A1(_0174_),
    .A2(_0849_),
    .ZN(_0850_)
  );
  INV_X1 _3465_ (
    .A(_0850_),
    .ZN(_0851_)
  );
  AND2_X1 _3466_ (
    .A1(_0848_),
    .A2(_0851_),
    .ZN(_0853_)
  );
  AND2_X1 _3467_ (
    .A1(_0846_),
    .A2(_0853_),
    .ZN(_0854_)
  );
  AND2_X1 _3468_ (
    .A1(_0844_),
    .A2(_0854_),
    .ZN(_0855_)
  );
  AND2_X1 _3469_ (
    .A1(_0842_),
    .A2(_0855_),
    .ZN(_0856_)
  );
  INV_X1 _3470_ (
    .A(_0856_),
    .ZN(io_out[29])
  );
  AND2_X1 _3471_ (
    .A1(_0004_),
    .A2(_0028_),
    .ZN(_0857_)
  );
  INV_X1 _3472_ (
    .A(_0857_),
    .ZN(_0858_)
  );
  AND2_X1 _3473_ (
    .A1(_0030_),
    .A2(_0858_),
    .ZN(io_adder_out[30])
  );
  AND2_X1 _3474_ (
    .A1(_0171_),
    .A2(io_adder_out[30]),
    .ZN(_0859_)
  );
  INV_X1 _3475_ (
    .A(_0859_),
    .ZN(_0860_)
  );
  AND2_X1 _3476_ (
    .A1(_0166_),
    .A2(_0224_),
    .ZN(_0862_)
  );
  INV_X1 _3477_ (
    .A(_0862_),
    .ZN(_0863_)
  );
  AND2_X1 _3478_ (
    .A1(_0081_),
    .A2(_0192_),
    .ZN(_0864_)
  );
  INV_X1 _3479_ (
    .A(_0864_),
    .ZN(_0865_)
  );
  AND2_X1 _3480_ (
    .A1(_0021_),
    .A2(_0178_),
    .ZN(_0866_)
  );
  INV_X1 _3481_ (
    .A(_0866_),
    .ZN(_0867_)
  );
  AND2_X1 _3482_ (
    .A1(io_in2[30]),
    .A2(io_in1[30]),
    .ZN(_0868_)
  );
  AND2_X1 _3483_ (
    .A1(_0174_),
    .A2(_0868_),
    .ZN(_0869_)
  );
  INV_X1 _3484_ (
    .A(_0869_),
    .ZN(_0870_)
  );
  AND2_X1 _3485_ (
    .A1(_0867_),
    .A2(_0870_),
    .ZN(_0871_)
  );
  AND2_X1 _3486_ (
    .A1(_0865_),
    .A2(_0871_),
    .ZN(_0873_)
  );
  AND2_X1 _3487_ (
    .A1(_0863_),
    .A2(_0873_),
    .ZN(_0874_)
  );
  AND2_X1 _3488_ (
    .A1(_0860_),
    .A2(_0874_),
    .ZN(_0875_)
  );
  INV_X1 _3489_ (
    .A(_0875_),
    .ZN(io_out[30])
  );
  AND2_X1 _3490_ (
    .A1(io_adder_out[31]),
    .A2(_0171_),
    .ZN(_0876_)
  );
  INV_X1 _3491_ (
    .A(_0876_),
    .ZN(_0877_)
  );
  AND2_X1 _3492_ (
    .A1(_0154_),
    .A2(_0166_),
    .ZN(_0878_)
  );
  INV_X1 _3493_ (
    .A(_0878_),
    .ZN(_0879_)
  );
  AND2_X1 _3494_ (
    .A1(_0081_),
    .A2(_0162_),
    .ZN(_0880_)
  );
  INV_X1 _3495_ (
    .A(_0880_),
    .ZN(_0881_)
  );
  AND2_X1 _3496_ (
    .A1(_0038_),
    .A2(_0178_),
    .ZN(_0883_)
  );
  INV_X1 _3497_ (
    .A(_0883_),
    .ZN(_0884_)
  );
  AND2_X1 _3498_ (
    .A1(io_in2[31]),
    .A2(io_in1[31]),
    .ZN(_0885_)
  );
  AND2_X1 _3499_ (
    .A1(_0174_),
    .A2(_0885_),
    .ZN(_0886_)
  );
  INV_X1 _3500_ (
    .A(_0886_),
    .ZN(_0887_)
  );
  AND2_X1 _3501_ (
    .A1(_0884_),
    .A2(_0887_),
    .ZN(_0888_)
  );
  AND2_X1 _3502_ (
    .A1(_0881_),
    .A2(_0888_),
    .ZN(_0889_)
  );
  AND2_X1 _3503_ (
    .A1(_0879_),
    .A2(_0889_),
    .ZN(_0890_)
  );
  AND2_X1 _3504_ (
    .A1(_0877_),
    .A2(_0890_),
    .ZN(_0891_)
  );
  INV_X1 _3505_ (
    .A(_0891_),
    .ZN(io_out[31])
  );
  AND2_X1 _3506_ (
    .A1(_0022_),
    .A2(_0043_),
    .ZN(_0893_)
  );
  AND2_X1 _3507_ (
    .A1(_1734_),
    .A2(_0893_),
    .ZN(_0894_)
  );
  AND2_X1 _3508_ (
    .A1(_1630_),
    .A2(_1656_),
    .ZN(_0895_)
  );
  AND2_X1 _3509_ (
    .A1(_1682_),
    .A2(_1710_),
    .ZN(_0896_)
  );
  AND2_X1 _3510_ (
    .A1(_0895_),
    .A2(_0896_),
    .ZN(_0897_)
  );
  AND2_X1 _3511_ (
    .A1(_1364_),
    .A2(_1540_),
    .ZN(_0898_)
  );
  AND2_X1 _3512_ (
    .A1(_1570_),
    .A2(_1600_),
    .ZN(_0899_)
  );
  AND2_X1 _3513_ (
    .A1(_0898_),
    .A2(_0899_),
    .ZN(_0900_)
  );
  AND2_X1 _3514_ (
    .A1(_0897_),
    .A2(_0900_),
    .ZN(_0901_)
  );
  AND2_X1 _3515_ (
    .A1(_0894_),
    .A2(_0901_),
    .ZN(_0902_)
  );
  AND2_X1 _3516_ (
    .A1(_0957_),
    .A2(_0987_),
    .ZN(_0904_)
  );
  AND2_X1 _3517_ (
    .A1(_1003_),
    .A2(_1019_),
    .ZN(_0905_)
  );
  AND2_X1 _3518_ (
    .A1(_0904_),
    .A2(_0905_),
    .ZN(_0906_)
  );
  AND2_X1 _3519_ (
    .A1(_0059_),
    .A2(_0906_),
    .ZN(_0907_)
  );
  AND2_X1 _3520_ (
    .A1(_1123_),
    .A2(_1139_),
    .ZN(_0908_)
  );
  AND2_X1 _3521_ (
    .A1(_1155_),
    .A2(_1183_),
    .ZN(_0909_)
  );
  AND2_X1 _3522_ (
    .A1(_0908_),
    .A2(_0909_),
    .ZN(_0910_)
  );
  AND2_X1 _3523_ (
    .A1(_1059_),
    .A2(_1075_),
    .ZN(_0911_)
  );
  AND2_X1 _3524_ (
    .A1(_1091_),
    .A2(_1107_),
    .ZN(_0912_)
  );
  AND2_X1 _3525_ (
    .A1(_0911_),
    .A2(_0912_),
    .ZN(_0913_)
  );
  AND2_X1 _3526_ (
    .A1(_0910_),
    .A2(_0913_),
    .ZN(_0915_)
  );
  AND2_X1 _3527_ (
    .A1(_1291_),
    .A2(_1299_),
    .ZN(_0916_)
  );
  AND2_X1 _3528_ (
    .A1(_1315_),
    .A2(_1356_),
    .ZN(_0917_)
  );
  AND2_X1 _3529_ (
    .A1(_0916_),
    .A2(_0917_),
    .ZN(_0918_)
  );
  AND2_X1 _3530_ (
    .A1(_1199_),
    .A2(_1267_),
    .ZN(_0919_)
  );
  AND2_X1 _3531_ (
    .A1(_1275_),
    .A2(_1283_),
    .ZN(_0920_)
  );
  AND2_X1 _3532_ (
    .A1(_0919_),
    .A2(_0920_),
    .ZN(_0921_)
  );
  AND2_X1 _3533_ (
    .A1(_0918_),
    .A2(_0921_),
    .ZN(_0922_)
  );
  AND2_X1 _3534_ (
    .A1(_0915_),
    .A2(_0922_),
    .ZN(_0923_)
  );
  AND2_X1 _3535_ (
    .A1(_0907_),
    .A2(_0923_),
    .ZN(_0924_)
  );
  AND2_X1 _3536_ (
    .A1(_0902_),
    .A2(_0924_),
    .ZN(_0926_)
  );
  INV_X1 _3537_ (
    .A(_0926_),
    .ZN(_0927_)
  );
  AND2_X1 _3538_ (
    .A1(_0070_),
    .A2(_0927_),
    .ZN(_0928_)
  );
  INV_X1 _3539_ (
    .A(_0928_),
    .ZN(_0929_)
  );
  AND2_X1 _3540_ (
    .A1(_0339_),
    .A2(_0928_),
    .ZN(_0930_)
  );
  INV_X1 _3541_ (
    .A(_0930_),
    .ZN(_0931_)
  );
  AND2_X1 _3542_ (
    .A1(io_fn[0]),
    .A2(_0929_),
    .ZN(_0932_)
  );
  INV_X1 _3543_ (
    .A(_0932_),
    .ZN(_0933_)
  );
  AND2_X1 _3544_ (
    .A1(_0931_),
    .A2(_0933_),
    .ZN(io_cmp_out)
  );
  assign _GEN_0 = { 31'h00000000, io_fn[3] };
  assign _GEN_1 = { 16'h0000, io_in1[31:16] };
  assign _GEN_10[31] = 1'h0;
  assign _GEN_11[31:1] = 31'h00000000;
  assign _GEN_2 = { 8'h00, io_in1[15:0], io_in1[31:24] };
  assign _GEN_3 = { 4'h0, io_in1[7:0], io_in1[15:8], io_in1[23:16], io_in1[31:28] };
  assign _GEN_4 = { 2'h0, io_in1[3:0], io_in1[7:4], io_in1[11:8], io_in1[15:12], io_in1[19:16], io_in1[23:20], io_in1[27:24], io_in1[31:30] };
  assign _GEN_5 = { 1'h0, io_in1[1:0], io_in1[3:2], io_in1[5:4], io_in1[7:6], io_in1[9:8], io_in1[11:10], io_in1[13:12], io_in1[15:14], io_in1[17:16], io_in1[19:18], io_in1[21:20], io_in1[23:22], io_in1[25:24], io_in1[27:26], io_in1[29:28], io_in1[31] };
  assign { _GEN_6[31:15], _GEN_6[13:0] } = { 16'h0000, _GEN_10[0], _GEN_10[2:1], _GEN_10[4:3], _GEN_10[6:5], _GEN_10[8:7], _GEN_10[10:9], _GEN_10[12:11], _GEN_10[14:13] };
  assign _GEN_7 = { 8'h00, _GEN_10[16:15], _GEN_10[18:17], _GEN_10[20:19], _GEN_10[22:21], _GEN_10[24:23], _GEN_10[26:25], _GEN_10[28:27], _GEN_10[30:29], _GEN_10[0], _GEN_6[14], _GEN_10[2:1], _GEN_10[4:3], _GEN_10[6:5] };
  assign _GEN_8 = { 4'h0, _GEN_10[24:23], _GEN_10[26:25], _GEN_10[28:27], _GEN_10[30:29], _GEN_10[16:15], _GEN_10[18:17], _GEN_10[20:19], _GEN_10[22:21], _GEN_10[8:7], _GEN_10[10:9], _GEN_10[12:11], _GEN_10[14:13], _GEN_10[0], _GEN_6[14], _GEN_10[2:1] };
  assign _GEN_9 = { 2'h0, _GEN_10[28:27], _GEN_10[30:29], _GEN_10[24:23], _GEN_10[26:25], _GEN_10[20:19], _GEN_10[22:21], _GEN_10[16:15], _GEN_10[18:17], _GEN_10[12:11], _GEN_10[14:13], _GEN_10[8:7], _GEN_10[10:9], _GEN_10[4:3], _GEN_10[6:5], _GEN_10[0], _GEN_6[14] };
  assign _shift_logic_T_1 = _GEN_11[0];
  assign _shin_T_10 = { io_in1[15:0], 16'h0000 };
  assign _shin_T_11 = { io_in1[15:0], io_in1[31:16] };
  assign _shin_T_16 = { 8'h00, io_in1[15:8], 8'h00, io_in1[31:24] };
  assign _shin_T_18 = { io_in1[7:0], io_in1[31:16], 8'h00 };
  assign _shin_T_20 = { io_in1[7:0], 8'h00, io_in1[23:16], 8'h00 };
  assign _shin_T_21 = { io_in1[7:0], io_in1[15:8], io_in1[23:16], io_in1[31:24] };
  assign _shin_T_26 = { 4'h0, io_in1[7:4], 4'h0, io_in1[15:12], 4'h0, io_in1[23:20], 4'h0, io_in1[31:28] };
  assign _shin_T_28 = { io_in1[3:0], io_in1[15:8], io_in1[23:16], io_in1[31:24], 4'h0 };
  assign _shin_T_30 = { io_in1[3:0], 4'h0, io_in1[11:8], 4'h0, io_in1[19:16], 4'h0, io_in1[27:24], 4'h0 };
  assign _shin_T_31 = { io_in1[3:0], io_in1[7:4], io_in1[11:8], io_in1[15:12], io_in1[19:16], io_in1[23:20], io_in1[27:24], io_in1[31:28] };
  assign _shin_T_36 = { 2'h0, io_in1[3:2], 2'h0, io_in1[7:6], 2'h0, io_in1[11:10], 2'h0, io_in1[15:14], 2'h0, io_in1[19:18], 2'h0, io_in1[23:22], 2'h0, io_in1[27:26], 2'h0, io_in1[31:30] };
  assign _shin_T_38 = { io_in1[1:0], io_in1[7:4], io_in1[11:8], io_in1[15:12], io_in1[19:16], io_in1[23:20], io_in1[27:24], io_in1[31:28], 2'h0 };
  assign _shin_T_40 = { io_in1[1:0], 2'h0, io_in1[5:4], 2'h0, io_in1[9:8], 2'h0, io_in1[13:12], 2'h0, io_in1[17:16], 2'h0, io_in1[21:20], 2'h0, io_in1[25:24], 2'h0, io_in1[29:28], 2'h0 };
  assign _shin_T_41 = { io_in1[1:0], io_in1[3:2], io_in1[5:4], io_in1[7:6], io_in1[9:8], io_in1[11:10], io_in1[13:12], io_in1[15:14], io_in1[17:16], io_in1[19:18], io_in1[21:20], io_in1[23:22], io_in1[25:24], io_in1[27:26], io_in1[29:28], io_in1[31:30] };
  assign _shin_T_46 = { 1'h0, io_in1[1], 1'h0, io_in1[3], 1'h0, io_in1[5], 1'h0, io_in1[7], 1'h0, io_in1[9], 1'h0, io_in1[11], 1'h0, io_in1[13], 1'h0, io_in1[15], 1'h0, io_in1[17], 1'h0, io_in1[19], 1'h0, io_in1[21], 1'h0, io_in1[23], 1'h0, io_in1[25], 1'h0, io_in1[27], 1'h0, io_in1[29], 1'h0, io_in1[31] };
  assign _shin_T_48 = { io_in1[0], io_in1[3:2], io_in1[5:4], io_in1[7:6], io_in1[9:8], io_in1[11:10], io_in1[13:12], io_in1[15:14], io_in1[17:16], io_in1[19:18], io_in1[21:20], io_in1[23:22], io_in1[25:24], io_in1[27:26], io_in1[29:28], io_in1[31:30], 1'h0 };
  assign _shin_T_50 = { io_in1[0], 1'h0, io_in1[2], 1'h0, io_in1[4], 1'h0, io_in1[6], 1'h0, io_in1[8], 1'h0, io_in1[10], 1'h0, io_in1[12], 1'h0, io_in1[14], 1'h0, io_in1[16], 1'h0, io_in1[18], 1'h0, io_in1[20], 1'h0, io_in1[22], 1'h0, io_in1[24], 1'h0, io_in1[26], 1'h0, io_in1[28], 1'h0, io_in1[30], 1'h0 };
  assign _shin_T_51 = { io_in1[0], io_in1[1], io_in1[2], io_in1[3], io_in1[4], io_in1[5], io_in1[6], io_in1[7], io_in1[8], io_in1[9], io_in1[10], io_in1[11], io_in1[12], io_in1[13], io_in1[14], io_in1[15], io_in1[16], io_in1[17], io_in1[18], io_in1[19], io_in1[20], io_in1[21], io_in1[22], io_in1[23], io_in1[24], io_in1[25], io_in1[26], io_in1[27], io_in1[28], io_in1[29], io_in1[30], io_in1[31] };
  assign _shin_T_6 = { 16'h0000, io_in1[31:16] };
  assign _shin_T_8 = { io_in1[15:0], 16'h0000 };
  assign _shout_l_T_13 = { 8'h00, _GEN_10[16:15], _GEN_10[18:17], _GEN_10[20:19], _GEN_10[22:21], 8'h00, _GEN_10[0], _GEN_6[14], _GEN_10[2:1], _GEN_10[4:3], _GEN_10[6:5] };
  assign _shout_l_T_15 = { _GEN_10[24:23], _GEN_10[26:25], _GEN_10[28:27], _GEN_10[30:29], _GEN_10[0], _GEN_6[14], _GEN_10[2:1], _GEN_10[4:3], _GEN_10[6:5], _GEN_10[8:7], _GEN_10[10:9], _GEN_10[12:11], _GEN_10[14:13], 8'h00 };
  assign _shout_l_T_17 = { _GEN_10[24:23], _GEN_10[26:25], _GEN_10[28:27], _GEN_10[30:29], 8'h00, _GEN_10[8:7], _GEN_10[10:9], _GEN_10[12:11], _GEN_10[14:13], 8'h00 };
  assign _shout_l_T_18 = { _GEN_10[24:23], _GEN_10[26:25], _GEN_10[28:27], _GEN_10[30:29], _GEN_10[16:15], _GEN_10[18:17], _GEN_10[20:19], _GEN_10[22:21], _GEN_10[8:7], _GEN_10[10:9], _GEN_10[12:11], _GEN_10[14:13], _GEN_10[0], _GEN_6[14], _GEN_10[2:1], _GEN_10[4:3], _GEN_10[6:5] };
  assign _shout_l_T_23 = { 4'h0, _GEN_10[24:23], _GEN_10[26:25], 4'h0, _GEN_10[16:15], _GEN_10[18:17], 4'h0, _GEN_10[8:7], _GEN_10[10:9], 4'h0, _GEN_10[0], _GEN_6[14], _GEN_10[2:1] };
  assign _shout_l_T_25 = { _GEN_10[28:27], _GEN_10[30:29], _GEN_10[16:15], _GEN_10[18:17], _GEN_10[20:19], _GEN_10[22:21], _GEN_10[8:7], _GEN_10[10:9], _GEN_10[12:11], _GEN_10[14:13], _GEN_10[0], _GEN_6[14], _GEN_10[2:1], _GEN_10[4:3], _GEN_10[6:5], 4'h0 };
  assign _shout_l_T_27 = { _GEN_10[28:27], _GEN_10[30:29], 4'h0, _GEN_10[20:19], _GEN_10[22:21], 4'h0, _GEN_10[12:11], _GEN_10[14:13], 4'h0, _GEN_10[4:3], _GEN_10[6:5], 4'h0 };
  assign _shout_l_T_28 = { _GEN_10[28:27], _GEN_10[30:29], _GEN_10[24:23], _GEN_10[26:25], _GEN_10[20:19], _GEN_10[22:21], _GEN_10[16:15], _GEN_10[18:17], _GEN_10[12:11], _GEN_10[14:13], _GEN_10[8:7], _GEN_10[10:9], _GEN_10[4:3], _GEN_10[6:5], _GEN_10[0], _GEN_6[14], _GEN_10[2:1] };
  assign _shout_l_T_3 = { 16'h0000, _GEN_10[0], _GEN_6[14], _GEN_10[2:1], _GEN_10[4:3], _GEN_10[6:5], _GEN_10[8:7], _GEN_10[10:9], _GEN_10[12:11], _GEN_10[14:13] };
  assign _shout_l_T_33 = { 2'h0, _GEN_10[28:27], 2'h0, _GEN_10[24:23], 2'h0, _GEN_10[20:19], 2'h0, _GEN_10[16:15], 2'h0, _GEN_10[12:11], 2'h0, _GEN_10[8:7], 2'h0, _GEN_10[4:3], 2'h0, _GEN_10[0], _GEN_6[14] };
  assign _shout_l_T_35 = { _GEN_10[30:29], _GEN_10[24:23], _GEN_10[26:25], _GEN_10[20:19], _GEN_10[22:21], _GEN_10[16:15], _GEN_10[18:17], _GEN_10[12:11], _GEN_10[14:13], _GEN_10[8:7], _GEN_10[10:9], _GEN_10[4:3], _GEN_10[6:5], _GEN_10[0], _GEN_6[14], _GEN_10[2:1], 2'h0 };
  assign _shout_l_T_37 = { _GEN_10[30:29], 2'h0, _GEN_10[26:25], 2'h0, _GEN_10[22:21], 2'h0, _GEN_10[18:17], 2'h0, _GEN_10[14:13], 2'h0, _GEN_10[10:9], 2'h0, _GEN_10[6:5], 2'h0, _GEN_10[2:1], 2'h0 };
  assign _shout_l_T_38 = { _GEN_10[30:0], _GEN_6[14] };
  assign _shout_l_T_43 = { 1'h0, _GEN_10[30], 1'h0, _GEN_10[28], 1'h0, _GEN_10[26], 1'h0, _GEN_10[24], 1'h0, _GEN_10[22], 1'h0, _GEN_10[20], 1'h0, _GEN_10[18], 1'h0, _GEN_10[16], 1'h0, _GEN_10[14], 1'h0, _GEN_10[12], 1'h0, _GEN_10[10], 1'h0, _GEN_10[8], 1'h0, _GEN_10[6], 1'h0, _GEN_10[4], 1'h0, _GEN_10[2], 1'h0, _GEN_10[0] };
  assign _shout_l_T_45 = { _GEN_10[29:0], _GEN_6[14], 1'h0 };
  assign _shout_l_T_47 = { _GEN_10[29], 1'h0, _GEN_10[27], 1'h0, _GEN_10[25], 1'h0, _GEN_10[23], 1'h0, _GEN_10[21], 1'h0, _GEN_10[19], 1'h0, _GEN_10[17], 1'h0, _GEN_10[15], 1'h0, _GEN_10[13], 1'h0, _GEN_10[11], 1'h0, _GEN_10[9], 1'h0, _GEN_10[7], 1'h0, _GEN_10[5], 1'h0, _GEN_10[3], 1'h0, _GEN_10[1], 1'h0, _GEN_6[14], 1'h0 };
  assign _shout_l_T_5 = { _GEN_10[16:15], _GEN_10[18:17], _GEN_10[20:19], _GEN_10[22:21], _GEN_10[24:23], _GEN_10[26:25], _GEN_10[28:27], _GEN_10[30:29], 16'h0000 };
  assign _shout_l_T_7 = { _GEN_10[16:15], _GEN_10[18:17], _GEN_10[20:19], _GEN_10[22:21], _GEN_10[24:23], _GEN_10[26:25], _GEN_10[28:27], _GEN_10[30:29], 16'h0000 };
  assign _shout_l_T_8 = { _GEN_10[16:15], _GEN_10[18:17], _GEN_10[20:19], _GEN_10[22:21], _GEN_10[24:23], _GEN_10[26:25], _GEN_10[28:27], _GEN_10[30:29], _GEN_10[0], _GEN_6[14], _GEN_10[2:1], _GEN_10[4:3], _GEN_10[6:5], _GEN_10[8:7], _GEN_10[10:9], _GEN_10[12:11], _GEN_10[14:13] };
  assign _shout_r_T_5[31:0] = { _GEN_10[0], _GEN_6[14], _GEN_10[2:1], _GEN_10[4:3], _GEN_10[6:5], _GEN_10[8:7], _GEN_10[10:9], _GEN_10[12:11], _GEN_10[14:13], _GEN_10[16:15], _GEN_10[18:17], _GEN_10[20:19], _GEN_10[22:21], _GEN_10[24:23], _GEN_10[26:25], _GEN_10[28:27], _GEN_10[30:29] };
  assign shamt = io_in2[4:0];
  assign shout_l = { _GEN_10[29], _GEN_10[30], _GEN_10[27], _GEN_10[28], _GEN_10[25], _GEN_10[26], _GEN_10[23], _GEN_10[24], _GEN_10[21], _GEN_10[22], _GEN_10[19], _GEN_10[20], _GEN_10[17], _GEN_10[18], _GEN_10[15], _GEN_10[16], _GEN_10[13], _GEN_10[14], _GEN_10[11], _GEN_10[12], _GEN_10[9], _GEN_10[10], _GEN_10[7], _GEN_10[8], _GEN_10[5], _GEN_10[6], _GEN_10[3], _GEN_10[4], _GEN_10[1], _GEN_10[2], _GEN_6[14], _GEN_10[0] };
  assign shout_r = { _GEN_10[0], _GEN_6[14], _GEN_10[2:1], _GEN_10[4:3], _GEN_10[6:5], _GEN_10[8:7], _GEN_10[10:9], _GEN_10[12:11], _GEN_10[14:13], _GEN_10[16:15], _GEN_10[18:17], _GEN_10[20:19], _GEN_10[22:21], _GEN_10[24:23], _GEN_10[26:25], _GEN_10[28:27], _GEN_10[30:29] };
endmodule
module BreakpointUnit(io_status_debug, io_bp_0_control_action, io_bp_0_control_tmatch, io_bp_0_control_x, io_bp_0_control_w, io_bp_0_control_r, io_bp_0_address, io_pc, io_ea, io_xcpt_if, io_xcpt_ld, io_xcpt_st, io_debug_if, io_debug_ld, io_debug_st);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire [31:0] _GEN_11;
  wire _r_T_10;
  wire _r_T_12;
  wire [3:0] _r_T_13;
  wire _r_T_8;
  input [31:0] io_bp_0_address;
  wire [31:0] io_bp_0_address;
  input io_bp_0_control_action;
  wire io_bp_0_control_action;
  input io_bp_0_control_r;
  wire io_bp_0_control_r;
  input [1:0] io_bp_0_control_tmatch;
  wire [1:0] io_bp_0_control_tmatch;
  input io_bp_0_control_w;
  wire io_bp_0_control_w;
  input io_bp_0_control_x;
  wire io_bp_0_control_x;
  output io_debug_if;
  wire io_debug_if;
  output io_debug_ld;
  wire io_debug_ld;
  output io_debug_st;
  wire io_debug_st;
  input [31:0] io_ea;
  wire [31:0] io_ea;
  input [31:0] io_pc;
  wire [31:0] io_pc;
  input io_status_debug;
  wire io_status_debug;
  output io_xcpt_if;
  wire io_xcpt_if;
  output io_xcpt_ld;
  wire io_xcpt_ld;
  output io_xcpt_st;
  wire io_xcpt_st;
  INV_X1 _0723_ (
    .A(io_bp_0_control_tmatch[1]),
    .ZN(_0000_)
  );
  INV_X1 _0724_ (
    .A(io_status_debug),
    .ZN(_0001_)
  );
  INV_X1 _0725_ (
    .A(io_ea[0]),
    .ZN(_0002_)
  );
  INV_X1 _0726_ (
    .A(io_ea[1]),
    .ZN(_0003_)
  );
  INV_X1 _0727_ (
    .A(io_ea[2]),
    .ZN(_0004_)
  );
  INV_X1 _0728_ (
    .A(io_ea[3]),
    .ZN(_0005_)
  );
  INV_X1 _0729_ (
    .A(io_ea[4]),
    .ZN(_0006_)
  );
  INV_X1 _0730_ (
    .A(io_ea[5]),
    .ZN(_0007_)
  );
  INV_X1 _0731_ (
    .A(io_ea[6]),
    .ZN(_0008_)
  );
  INV_X1 _0732_ (
    .A(io_ea[7]),
    .ZN(_0009_)
  );
  INV_X1 _0733_ (
    .A(io_ea[8]),
    .ZN(_0010_)
  );
  INV_X1 _0734_ (
    .A(io_ea[9]),
    .ZN(_0011_)
  );
  INV_X1 _0735_ (
    .A(io_ea[10]),
    .ZN(_0012_)
  );
  INV_X1 _0736_ (
    .A(io_ea[11]),
    .ZN(_0013_)
  );
  INV_X1 _0737_ (
    .A(io_ea[12]),
    .ZN(_0014_)
  );
  INV_X1 _0738_ (
    .A(io_ea[13]),
    .ZN(_0015_)
  );
  INV_X1 _0739_ (
    .A(io_ea[14]),
    .ZN(_0016_)
  );
  INV_X1 _0740_ (
    .A(io_ea[15]),
    .ZN(_0017_)
  );
  INV_X1 _0741_ (
    .A(io_ea[16]),
    .ZN(_0018_)
  );
  INV_X1 _0742_ (
    .A(io_ea[17]),
    .ZN(_0019_)
  );
  INV_X1 _0743_ (
    .A(io_ea[18]),
    .ZN(_0020_)
  );
  INV_X1 _0744_ (
    .A(io_ea[19]),
    .ZN(_0021_)
  );
  INV_X1 _0745_ (
    .A(io_ea[20]),
    .ZN(_0022_)
  );
  INV_X1 _0746_ (
    .A(io_ea[21]),
    .ZN(_0023_)
  );
  INV_X1 _0747_ (
    .A(io_ea[22]),
    .ZN(_0024_)
  );
  INV_X1 _0748_ (
    .A(io_ea[23]),
    .ZN(_0025_)
  );
  INV_X1 _0749_ (
    .A(io_ea[24]),
    .ZN(_0026_)
  );
  INV_X1 _0750_ (
    .A(io_ea[25]),
    .ZN(_0027_)
  );
  INV_X1 _0751_ (
    .A(io_ea[26]),
    .ZN(_0028_)
  );
  INV_X1 _0752_ (
    .A(io_ea[27]),
    .ZN(_0029_)
  );
  INV_X1 _0753_ (
    .A(io_ea[28]),
    .ZN(_0030_)
  );
  INV_X1 _0754_ (
    .A(io_ea[29]),
    .ZN(_0031_)
  );
  INV_X1 _0755_ (
    .A(io_ea[30]),
    .ZN(_0032_)
  );
  INV_X1 _0756_ (
    .A(io_ea[31]),
    .ZN(_0033_)
  );
  INV_X1 _0757_ (
    .A(io_pc[0]),
    .ZN(_0034_)
  );
  INV_X1 _0758_ (
    .A(io_pc[1]),
    .ZN(_0035_)
  );
  INV_X1 _0759_ (
    .A(io_pc[2]),
    .ZN(_0036_)
  );
  INV_X1 _0760_ (
    .A(io_pc[3]),
    .ZN(_0037_)
  );
  INV_X1 _0761_ (
    .A(io_pc[4]),
    .ZN(_0038_)
  );
  INV_X1 _0762_ (
    .A(io_pc[5]),
    .ZN(_0039_)
  );
  INV_X1 _0763_ (
    .A(io_pc[6]),
    .ZN(_0040_)
  );
  INV_X1 _0764_ (
    .A(io_pc[7]),
    .ZN(_0041_)
  );
  INV_X1 _0765_ (
    .A(io_pc[8]),
    .ZN(_0042_)
  );
  INV_X1 _0766_ (
    .A(io_pc[9]),
    .ZN(_0043_)
  );
  INV_X1 _0767_ (
    .A(io_pc[10]),
    .ZN(_0044_)
  );
  INV_X1 _0768_ (
    .A(io_pc[11]),
    .ZN(_0045_)
  );
  INV_X1 _0769_ (
    .A(io_pc[12]),
    .ZN(_0046_)
  );
  INV_X1 _0770_ (
    .A(io_pc[13]),
    .ZN(_0047_)
  );
  INV_X1 _0771_ (
    .A(io_pc[14]),
    .ZN(_0048_)
  );
  INV_X1 _0772_ (
    .A(io_pc[15]),
    .ZN(_0049_)
  );
  INV_X1 _0773_ (
    .A(io_pc[16]),
    .ZN(_0050_)
  );
  INV_X1 _0774_ (
    .A(io_pc[17]),
    .ZN(_0051_)
  );
  INV_X1 _0775_ (
    .A(io_pc[18]),
    .ZN(_0052_)
  );
  INV_X1 _0776_ (
    .A(io_pc[19]),
    .ZN(_0053_)
  );
  INV_X1 _0777_ (
    .A(io_pc[20]),
    .ZN(_0054_)
  );
  INV_X1 _0778_ (
    .A(io_pc[21]),
    .ZN(_0055_)
  );
  INV_X1 _0779_ (
    .A(io_pc[22]),
    .ZN(_0056_)
  );
  INV_X1 _0780_ (
    .A(io_pc[23]),
    .ZN(_0057_)
  );
  INV_X1 _0781_ (
    .A(io_pc[24]),
    .ZN(_0058_)
  );
  INV_X1 _0782_ (
    .A(io_pc[25]),
    .ZN(_0059_)
  );
  INV_X1 _0783_ (
    .A(io_pc[26]),
    .ZN(_0060_)
  );
  INV_X1 _0784_ (
    .A(io_pc[27]),
    .ZN(_0061_)
  );
  INV_X1 _0785_ (
    .A(io_pc[28]),
    .ZN(_0062_)
  );
  INV_X1 _0786_ (
    .A(io_pc[29]),
    .ZN(_0063_)
  );
  INV_X1 _0787_ (
    .A(io_pc[30]),
    .ZN(_0064_)
  );
  INV_X1 _0788_ (
    .A(io_pc[31]),
    .ZN(_0065_)
  );
  INV_X1 _0789_ (
    .A(io_bp_0_control_action),
    .ZN(_0066_)
  );
  INV_X1 _0790_ (
    .A(io_bp_0_address[0]),
    .ZN(_0067_)
  );
  INV_X1 _0791_ (
    .A(io_bp_0_address[1]),
    .ZN(_0068_)
  );
  INV_X1 _0792_ (
    .A(io_bp_0_address[2]),
    .ZN(_0069_)
  );
  INV_X1 _0793_ (
    .A(io_bp_0_address[3]),
    .ZN(_0070_)
  );
  INV_X1 _0794_ (
    .A(io_bp_0_address[4]),
    .ZN(_0071_)
  );
  INV_X1 _0795_ (
    .A(io_bp_0_address[5]),
    .ZN(_0072_)
  );
  INV_X1 _0796_ (
    .A(io_bp_0_address[6]),
    .ZN(_0073_)
  );
  INV_X1 _0797_ (
    .A(io_bp_0_address[7]),
    .ZN(_0074_)
  );
  INV_X1 _0798_ (
    .A(io_bp_0_address[8]),
    .ZN(_0075_)
  );
  INV_X1 _0799_ (
    .A(io_bp_0_address[9]),
    .ZN(_0076_)
  );
  INV_X1 _0800_ (
    .A(io_bp_0_address[10]),
    .ZN(_0077_)
  );
  INV_X1 _0801_ (
    .A(io_bp_0_address[11]),
    .ZN(_0078_)
  );
  INV_X1 _0802_ (
    .A(io_bp_0_address[12]),
    .ZN(_0079_)
  );
  INV_X1 _0803_ (
    .A(io_bp_0_address[13]),
    .ZN(_0080_)
  );
  INV_X1 _0804_ (
    .A(io_bp_0_address[14]),
    .ZN(_0081_)
  );
  INV_X1 _0805_ (
    .A(io_bp_0_address[15]),
    .ZN(_0082_)
  );
  INV_X1 _0806_ (
    .A(io_bp_0_address[16]),
    .ZN(_0083_)
  );
  INV_X1 _0807_ (
    .A(io_bp_0_address[17]),
    .ZN(_0084_)
  );
  INV_X1 _0808_ (
    .A(io_bp_0_address[18]),
    .ZN(_0085_)
  );
  INV_X1 _0809_ (
    .A(io_bp_0_address[19]),
    .ZN(_0086_)
  );
  INV_X1 _0810_ (
    .A(io_bp_0_address[20]),
    .ZN(_0087_)
  );
  INV_X1 _0811_ (
    .A(io_bp_0_address[21]),
    .ZN(_0088_)
  );
  INV_X1 _0812_ (
    .A(io_bp_0_address[22]),
    .ZN(_0089_)
  );
  INV_X1 _0813_ (
    .A(io_bp_0_address[23]),
    .ZN(_0090_)
  );
  INV_X1 _0814_ (
    .A(io_bp_0_address[24]),
    .ZN(_0091_)
  );
  INV_X1 _0815_ (
    .A(io_bp_0_address[25]),
    .ZN(_0092_)
  );
  INV_X1 _0816_ (
    .A(io_bp_0_address[26]),
    .ZN(_0093_)
  );
  INV_X1 _0817_ (
    .A(io_bp_0_address[27]),
    .ZN(_0094_)
  );
  INV_X1 _0818_ (
    .A(io_bp_0_address[28]),
    .ZN(_0095_)
  );
  INV_X1 _0819_ (
    .A(io_bp_0_address[29]),
    .ZN(_0096_)
  );
  INV_X1 _0820_ (
    .A(io_bp_0_address[30]),
    .ZN(_0097_)
  );
  INV_X1 _0821_ (
    .A(io_bp_0_address[31]),
    .ZN(_0098_)
  );
  INV_X1 _0822_ (
    .A(io_bp_0_control_tmatch[0]),
    .ZN(_0099_)
  );
  AND2_X1 _0823_ (
    .A1(io_pc[31]),
    .A2(_0098_),
    .ZN(_0100_)
  );
  INV_X1 _0824_ (
    .A(_0100_),
    .ZN(_0101_)
  );
  AND2_X1 _0825_ (
    .A1(io_pc[30]),
    .A2(_0097_),
    .ZN(_0102_)
  );
  INV_X1 _0826_ (
    .A(_0102_),
    .ZN(_0103_)
  );
  AND2_X1 _0827_ (
    .A1(_0101_),
    .A2(_0103_),
    .ZN(_0104_)
  );
  INV_X1 _0828_ (
    .A(_0104_),
    .ZN(_0105_)
  );
  AND2_X1 _0829_ (
    .A1(_0064_),
    .A2(io_bp_0_address[30]),
    .ZN(_0106_)
  );
  INV_X1 _0830_ (
    .A(_0106_),
    .ZN(_0107_)
  );
  AND2_X1 _0831_ (
    .A1(_0065_),
    .A2(io_bp_0_address[31]),
    .ZN(_0108_)
  );
  INV_X1 _0832_ (
    .A(_0108_),
    .ZN(_0109_)
  );
  AND2_X1 _0833_ (
    .A1(_0063_),
    .A2(io_bp_0_address[29]),
    .ZN(_0110_)
  );
  INV_X1 _0834_ (
    .A(_0110_),
    .ZN(_0111_)
  );
  AND2_X1 _0835_ (
    .A1(_0062_),
    .A2(io_bp_0_address[28]),
    .ZN(_0112_)
  );
  INV_X1 _0836_ (
    .A(_0112_),
    .ZN(_0113_)
  );
  AND2_X1 _0837_ (
    .A1(io_pc[28]),
    .A2(_0095_),
    .ZN(_0114_)
  );
  INV_X1 _0838_ (
    .A(_0114_),
    .ZN(_0115_)
  );
  AND2_X1 _0839_ (
    .A1(io_pc[29]),
    .A2(_0096_),
    .ZN(_0116_)
  );
  INV_X1 _0840_ (
    .A(_0116_),
    .ZN(_0117_)
  );
  AND2_X1 _0841_ (
    .A1(_0115_),
    .A2(_0117_),
    .ZN(_0118_)
  );
  INV_X1 _0842_ (
    .A(_0118_),
    .ZN(_0119_)
  );
  AND2_X1 _0843_ (
    .A1(_0111_),
    .A2(_0113_),
    .ZN(_0120_)
  );
  AND2_X1 _0844_ (
    .A1(_0107_),
    .A2(_0109_),
    .ZN(_0121_)
  );
  AND2_X1 _0845_ (
    .A1(_0104_),
    .A2(_0121_),
    .ZN(_0122_)
  );
  AND2_X1 _0846_ (
    .A1(_0118_),
    .A2(_0122_),
    .ZN(_0123_)
  );
  AND2_X1 _0847_ (
    .A1(_0120_),
    .A2(_0123_),
    .ZN(_0124_)
  );
  AND2_X1 _0848_ (
    .A1(io_pc[17]),
    .A2(_0084_),
    .ZN(_0125_)
  );
  INV_X1 _0849_ (
    .A(_0125_),
    .ZN(_0126_)
  );
  AND2_X1 _0850_ (
    .A1(_0050_),
    .A2(io_bp_0_address[16]),
    .ZN(_0127_)
  );
  INV_X1 _0851_ (
    .A(_0127_),
    .ZN(_0128_)
  );
  AND2_X1 _0852_ (
    .A1(_0126_),
    .A2(_0128_),
    .ZN(_0129_)
  );
  AND2_X1 _0853_ (
    .A1(io_pc[16]),
    .A2(_0083_),
    .ZN(_0130_)
  );
  INV_X1 _0854_ (
    .A(_0130_),
    .ZN(_0131_)
  );
  AND2_X1 _0855_ (
    .A1(_0054_),
    .A2(io_bp_0_address[20]),
    .ZN(_0132_)
  );
  INV_X1 _0856_ (
    .A(_0132_),
    .ZN(_0133_)
  );
  AND2_X1 _0857_ (
    .A1(_0131_),
    .A2(_0133_),
    .ZN(_0134_)
  );
  AND2_X1 _0858_ (
    .A1(_0129_),
    .A2(_0134_),
    .ZN(_0135_)
  );
  AND2_X1 _0859_ (
    .A1(_0055_),
    .A2(io_bp_0_address[21]),
    .ZN(_0136_)
  );
  INV_X1 _0860_ (
    .A(_0136_),
    .ZN(_0137_)
  );
  AND2_X1 _0861_ (
    .A1(_0056_),
    .A2(io_bp_0_address[22]),
    .ZN(_0138_)
  );
  INV_X1 _0862_ (
    .A(_0138_),
    .ZN(_0139_)
  );
  AND2_X1 _0863_ (
    .A1(_0137_),
    .A2(_0139_),
    .ZN(_0140_)
  );
  AND2_X1 _0864_ (
    .A1(io_pc[23]),
    .A2(_0090_),
    .ZN(_0141_)
  );
  INV_X1 _0865_ (
    .A(_0141_),
    .ZN(_0142_)
  );
  AND2_X1 _0866_ (
    .A1(io_pc[22]),
    .A2(_0089_),
    .ZN(_0143_)
  );
  INV_X1 _0867_ (
    .A(_0143_),
    .ZN(_0144_)
  );
  AND2_X1 _0868_ (
    .A1(_0142_),
    .A2(_0144_),
    .ZN(_0145_)
  );
  AND2_X1 _0869_ (
    .A1(_0140_),
    .A2(_0145_),
    .ZN(_0146_)
  );
  AND2_X1 _0870_ (
    .A1(_0135_),
    .A2(_0146_),
    .ZN(_0147_)
  );
  AND2_X1 _0871_ (
    .A1(io_pc[19]),
    .A2(_0086_),
    .ZN(_0148_)
  );
  INV_X1 _0872_ (
    .A(_0148_),
    .ZN(_0149_)
  );
  AND2_X1 _0873_ (
    .A1(_0053_),
    .A2(io_bp_0_address[19]),
    .ZN(_0150_)
  );
  INV_X1 _0874_ (
    .A(_0150_),
    .ZN(_0151_)
  );
  AND2_X1 _0875_ (
    .A1(_0149_),
    .A2(_0151_),
    .ZN(_0152_)
  );
  AND2_X1 _0876_ (
    .A1(_0052_),
    .A2(io_bp_0_address[18]),
    .ZN(_0153_)
  );
  INV_X1 _0877_ (
    .A(_0153_),
    .ZN(_0154_)
  );
  AND2_X1 _0878_ (
    .A1(io_pc[18]),
    .A2(_0085_),
    .ZN(_0155_)
  );
  INV_X1 _0879_ (
    .A(_0155_),
    .ZN(_0156_)
  );
  AND2_X1 _0880_ (
    .A1(_0154_),
    .A2(_0156_),
    .ZN(_0157_)
  );
  AND2_X1 _0881_ (
    .A1(_0152_),
    .A2(_0157_),
    .ZN(_0158_)
  );
  AND2_X1 _0882_ (
    .A1(_0057_),
    .A2(io_bp_0_address[23]),
    .ZN(_0159_)
  );
  INV_X1 _0883_ (
    .A(_0159_),
    .ZN(_0160_)
  );
  AND2_X1 _0884_ (
    .A1(io_pc[21]),
    .A2(_0088_),
    .ZN(_0161_)
  );
  INV_X1 _0885_ (
    .A(_0161_),
    .ZN(_0162_)
  );
  AND2_X1 _0886_ (
    .A1(_0160_),
    .A2(_0162_),
    .ZN(_0163_)
  );
  AND2_X1 _0887_ (
    .A1(_0051_),
    .A2(io_bp_0_address[17]),
    .ZN(_0164_)
  );
  INV_X1 _0888_ (
    .A(_0164_),
    .ZN(_0165_)
  );
  AND2_X1 _0889_ (
    .A1(io_pc[20]),
    .A2(_0087_),
    .ZN(_0166_)
  );
  INV_X1 _0890_ (
    .A(_0166_),
    .ZN(_0167_)
  );
  AND2_X1 _0891_ (
    .A1(_0165_),
    .A2(_0167_),
    .ZN(_0168_)
  );
  AND2_X1 _0892_ (
    .A1(_0163_),
    .A2(_0168_),
    .ZN(_0169_)
  );
  AND2_X1 _0893_ (
    .A1(_0158_),
    .A2(_0169_),
    .ZN(_0170_)
  );
  AND2_X1 _0894_ (
    .A1(_0147_),
    .A2(_0170_),
    .ZN(_0171_)
  );
  AND2_X1 _0895_ (
    .A1(io_pc[27]),
    .A2(_0094_),
    .ZN(_0172_)
  );
  INV_X1 _0896_ (
    .A(_0172_),
    .ZN(_0173_)
  );
  AND2_X1 _0897_ (
    .A1(_0061_),
    .A2(io_bp_0_address[27]),
    .ZN(_0174_)
  );
  INV_X1 _0898_ (
    .A(_0174_),
    .ZN(_0175_)
  );
  AND2_X1 _0899_ (
    .A1(_0173_),
    .A2(_0175_),
    .ZN(_0176_)
  );
  AND2_X1 _0900_ (
    .A1(_0060_),
    .A2(io_bp_0_address[26]),
    .ZN(_0177_)
  );
  INV_X1 _0901_ (
    .A(_0177_),
    .ZN(_0178_)
  );
  AND2_X1 _0902_ (
    .A1(io_pc[26]),
    .A2(_0093_),
    .ZN(_0179_)
  );
  INV_X1 _0903_ (
    .A(_0179_),
    .ZN(_0180_)
  );
  AND2_X1 _0904_ (
    .A1(_0178_),
    .A2(_0180_),
    .ZN(_0181_)
  );
  AND2_X1 _0905_ (
    .A1(_0176_),
    .A2(_0181_),
    .ZN(_0182_)
  );
  AND2_X1 _0906_ (
    .A1(_0059_),
    .A2(io_bp_0_address[25]),
    .ZN(_0183_)
  );
  INV_X1 _0907_ (
    .A(_0183_),
    .ZN(_0184_)
  );
  AND2_X1 _0908_ (
    .A1(_0058_),
    .A2(io_bp_0_address[24]),
    .ZN(_0185_)
  );
  INV_X1 _0909_ (
    .A(_0185_),
    .ZN(_0186_)
  );
  AND2_X1 _0910_ (
    .A1(_0184_),
    .A2(_0186_),
    .ZN(_0187_)
  );
  AND2_X1 _0911_ (
    .A1(io_pc[25]),
    .A2(_0092_),
    .ZN(_0188_)
  );
  INV_X1 _0912_ (
    .A(_0188_),
    .ZN(_0189_)
  );
  AND2_X1 _0913_ (
    .A1(io_pc[24]),
    .A2(_0091_),
    .ZN(_0190_)
  );
  INV_X1 _0914_ (
    .A(_0190_),
    .ZN(_0191_)
  );
  AND2_X1 _0915_ (
    .A1(_0189_),
    .A2(_0191_),
    .ZN(_0192_)
  );
  INV_X1 _0916_ (
    .A(_0192_),
    .ZN(_0193_)
  );
  AND2_X1 _0917_ (
    .A1(_0187_),
    .A2(_0192_),
    .ZN(_0194_)
  );
  AND2_X1 _0918_ (
    .A1(_0182_),
    .A2(_0194_),
    .ZN(_0195_)
  );
  AND2_X1 _0919_ (
    .A1(_0124_),
    .A2(_0195_),
    .ZN(_0196_)
  );
  AND2_X1 _0920_ (
    .A1(_0171_),
    .A2(_0196_),
    .ZN(_0197_)
  );
  AND2_X1 _0921_ (
    .A1(io_pc[5]),
    .A2(_0072_),
    .ZN(_0198_)
  );
  INV_X1 _0922_ (
    .A(_0198_),
    .ZN(_0199_)
  );
  AND2_X1 _0923_ (
    .A1(io_pc[6]),
    .A2(_0073_),
    .ZN(_0200_)
  );
  INV_X1 _0924_ (
    .A(_0200_),
    .ZN(_0201_)
  );
  AND2_X1 _0925_ (
    .A1(_0199_),
    .A2(_0201_),
    .ZN(_0202_)
  );
  AND2_X1 _0926_ (
    .A1(_0041_),
    .A2(io_bp_0_address[7]),
    .ZN(_0203_)
  );
  INV_X1 _0927_ (
    .A(_0203_),
    .ZN(_0204_)
  );
  AND2_X1 _0928_ (
    .A1(_0040_),
    .A2(io_bp_0_address[6]),
    .ZN(_0205_)
  );
  INV_X1 _0929_ (
    .A(_0205_),
    .ZN(_0206_)
  );
  AND2_X1 _0930_ (
    .A1(_0204_),
    .A2(_0206_),
    .ZN(_0207_)
  );
  AND2_X1 _0931_ (
    .A1(_0039_),
    .A2(io_bp_0_address[5]),
    .ZN(_0208_)
  );
  INV_X1 _0932_ (
    .A(_0208_),
    .ZN(_0209_)
  );
  AND2_X1 _0933_ (
    .A1(_0038_),
    .A2(io_bp_0_address[4]),
    .ZN(_0210_)
  );
  INV_X1 _0934_ (
    .A(_0210_),
    .ZN(_0211_)
  );
  AND2_X1 _0935_ (
    .A1(_0209_),
    .A2(_0211_),
    .ZN(_0212_)
  );
  AND2_X1 _0936_ (
    .A1(_0207_),
    .A2(_0212_),
    .ZN(_0213_)
  );
  AND2_X1 _0937_ (
    .A1(_0202_),
    .A2(_0213_),
    .ZN(_0214_)
  );
  AND2_X1 _0938_ (
    .A1(_0034_),
    .A2(io_bp_0_address[0]),
    .ZN(_0215_)
  );
  INV_X1 _0939_ (
    .A(_0215_),
    .ZN(_0216_)
  );
  AND2_X1 _0940_ (
    .A1(io_pc[0]),
    .A2(_0067_),
    .ZN(_0217_)
  );
  INV_X1 _0941_ (
    .A(_0217_),
    .ZN(_0218_)
  );
  AND2_X1 _0942_ (
    .A1(_0216_),
    .A2(_0218_),
    .ZN(_0219_)
  );
  INV_X1 _0943_ (
    .A(_0219_),
    .ZN(_0220_)
  );
  AND2_X1 _0944_ (
    .A1(_0099_),
    .A2(_0220_),
    .ZN(_0221_)
  );
  INV_X1 _0945_ (
    .A(_0221_),
    .ZN(_0222_)
  );
  AND2_X1 _0946_ (
    .A1(io_pc[4]),
    .A2(_0071_),
    .ZN(_0223_)
  );
  INV_X1 _0947_ (
    .A(_0223_),
    .ZN(_0224_)
  );
  AND2_X1 _0948_ (
    .A1(io_pc[7]),
    .A2(_0074_),
    .ZN(_0225_)
  );
  INV_X1 _0949_ (
    .A(_0225_),
    .ZN(_0226_)
  );
  AND2_X1 _0950_ (
    .A1(_0000_),
    .A2(_0226_),
    .ZN(_0227_)
  );
  AND2_X1 _0951_ (
    .A1(_0224_),
    .A2(_0227_),
    .ZN(_0228_)
  );
  AND2_X1 _0952_ (
    .A1(_0222_),
    .A2(_0228_),
    .ZN(_0229_)
  );
  AND2_X1 _0953_ (
    .A1(_0214_),
    .A2(_0229_),
    .ZN(_0230_)
  );
  AND2_X1 _0954_ (
    .A1(io_pc[11]),
    .A2(_0078_),
    .ZN(_0231_)
  );
  INV_X1 _0955_ (
    .A(_0231_),
    .ZN(_0232_)
  );
  AND2_X1 _0956_ (
    .A1(io_pc[10]),
    .A2(_0077_),
    .ZN(_0233_)
  );
  INV_X1 _0957_ (
    .A(_0233_),
    .ZN(_0234_)
  );
  AND2_X1 _0958_ (
    .A1(_0232_),
    .A2(_0234_),
    .ZN(_0235_)
  );
  INV_X1 _0959_ (
    .A(_0235_),
    .ZN(_0236_)
  );
  AND2_X1 _0960_ (
    .A1(_0045_),
    .A2(io_bp_0_address[11]),
    .ZN(_0237_)
  );
  INV_X1 _0961_ (
    .A(_0237_),
    .ZN(_0238_)
  );
  AND2_X1 _0962_ (
    .A1(_0044_),
    .A2(io_bp_0_address[10]),
    .ZN(_0239_)
  );
  INV_X1 _0963_ (
    .A(_0239_),
    .ZN(_0240_)
  );
  AND2_X1 _0964_ (
    .A1(_0238_),
    .A2(_0240_),
    .ZN(_0241_)
  );
  AND2_X1 _0965_ (
    .A1(_0235_),
    .A2(_0241_),
    .ZN(_0242_)
  );
  AND2_X1 _0966_ (
    .A1(_0043_),
    .A2(io_bp_0_address[9]),
    .ZN(_0243_)
  );
  INV_X1 _0967_ (
    .A(_0243_),
    .ZN(_0244_)
  );
  AND2_X1 _0968_ (
    .A1(_0042_),
    .A2(io_bp_0_address[8]),
    .ZN(_0245_)
  );
  INV_X1 _0969_ (
    .A(_0245_),
    .ZN(_0246_)
  );
  AND2_X1 _0970_ (
    .A1(_0244_),
    .A2(_0246_),
    .ZN(_0247_)
  );
  AND2_X1 _0971_ (
    .A1(io_pc[9]),
    .A2(_0076_),
    .ZN(_0248_)
  );
  INV_X1 _0972_ (
    .A(_0248_),
    .ZN(_0249_)
  );
  AND2_X1 _0973_ (
    .A1(io_pc[8]),
    .A2(_0075_),
    .ZN(_0250_)
  );
  INV_X1 _0974_ (
    .A(_0250_),
    .ZN(_0251_)
  );
  AND2_X1 _0975_ (
    .A1(_0249_),
    .A2(_0251_),
    .ZN(_0252_)
  );
  INV_X1 _0976_ (
    .A(_0252_),
    .ZN(_0253_)
  );
  AND2_X1 _0977_ (
    .A1(_0247_),
    .A2(_0252_),
    .ZN(_0254_)
  );
  AND2_X1 _0978_ (
    .A1(_0242_),
    .A2(_0254_),
    .ZN(_0255_)
  );
  AND2_X1 _0979_ (
    .A1(io_bp_0_address[0]),
    .A2(io_bp_0_control_tmatch[0]),
    .ZN(_0256_)
  );
  INV_X1 _0980_ (
    .A(_0256_),
    .ZN(_0257_)
  );
  AND2_X1 _0981_ (
    .A1(io_bp_0_address[1]),
    .A2(_0256_),
    .ZN(_0258_)
  );
  INV_X1 _0982_ (
    .A(_0258_),
    .ZN(_0259_)
  );
  AND2_X1 _0983_ (
    .A1(io_bp_0_address[2]),
    .A2(_0258_),
    .ZN(_0260_)
  );
  INV_X1 _0984_ (
    .A(_0260_),
    .ZN(_0261_)
  );
  AND2_X1 _0985_ (
    .A1(_0037_),
    .A2(io_bp_0_address[3]),
    .ZN(_0262_)
  );
  INV_X1 _0986_ (
    .A(_0262_),
    .ZN(_0263_)
  );
  AND2_X1 _0987_ (
    .A1(io_pc[3]),
    .A2(_0070_),
    .ZN(_0264_)
  );
  INV_X1 _0988_ (
    .A(_0264_),
    .ZN(_0265_)
  );
  AND2_X1 _0989_ (
    .A1(_0263_),
    .A2(_0265_),
    .ZN(_0266_)
  );
  INV_X1 _0990_ (
    .A(_0266_),
    .ZN(_0267_)
  );
  AND2_X1 _0991_ (
    .A1(_0261_),
    .A2(_0267_),
    .ZN(_0268_)
  );
  INV_X1 _0992_ (
    .A(_0268_),
    .ZN(_0269_)
  );
  AND2_X1 _0993_ (
    .A1(_0048_),
    .A2(io_bp_0_address[14]),
    .ZN(_0270_)
  );
  INV_X1 _0994_ (
    .A(_0270_),
    .ZN(_0271_)
  );
  AND2_X1 _0995_ (
    .A1(_0049_),
    .A2(io_bp_0_address[15]),
    .ZN(_0272_)
  );
  INV_X1 _0996_ (
    .A(_0272_),
    .ZN(_0273_)
  );
  AND2_X1 _0997_ (
    .A1(io_pc[14]),
    .A2(_0081_),
    .ZN(_0274_)
  );
  INV_X1 _0998_ (
    .A(_0274_),
    .ZN(_0275_)
  );
  AND2_X1 _0999_ (
    .A1(_0047_),
    .A2(io_bp_0_address[13]),
    .ZN(_0276_)
  );
  INV_X1 _1000_ (
    .A(_0276_),
    .ZN(_0277_)
  );
  AND2_X1 _1001_ (
    .A1(io_pc[15]),
    .A2(_0082_),
    .ZN(_0278_)
  );
  INV_X1 _1002_ (
    .A(_0278_),
    .ZN(_0279_)
  );
  AND2_X1 _1003_ (
    .A1(_0277_),
    .A2(_0279_),
    .ZN(_0280_)
  );
  AND2_X1 _1004_ (
    .A1(_0271_),
    .A2(_0275_),
    .ZN(_0281_)
  );
  AND2_X1 _1005_ (
    .A1(_0273_),
    .A2(_0281_),
    .ZN(_0282_)
  );
  AND2_X1 _1006_ (
    .A1(_0280_),
    .A2(_0282_),
    .ZN(_0283_)
  );
  AND2_X1 _1007_ (
    .A1(_0046_),
    .A2(io_bp_0_address[12]),
    .ZN(_0284_)
  );
  INV_X1 _1008_ (
    .A(_0284_),
    .ZN(_0285_)
  );
  AND2_X1 _1009_ (
    .A1(io_pc[13]),
    .A2(_0080_),
    .ZN(_0286_)
  );
  INV_X1 _1010_ (
    .A(_0286_),
    .ZN(_0287_)
  );
  AND2_X1 _1011_ (
    .A1(io_pc[12]),
    .A2(_0079_),
    .ZN(_0288_)
  );
  INV_X1 _1012_ (
    .A(_0288_),
    .ZN(_0289_)
  );
  AND2_X1 _1013_ (
    .A1(_0287_),
    .A2(_0289_),
    .ZN(_0290_)
  );
  INV_X1 _1014_ (
    .A(_0290_),
    .ZN(_0291_)
  );
  AND2_X1 _1015_ (
    .A1(_0285_),
    .A2(_0290_),
    .ZN(_0292_)
  );
  AND2_X1 _1016_ (
    .A1(_0283_),
    .A2(_0292_),
    .ZN(_0293_)
  );
  AND2_X1 _1017_ (
    .A1(io_pc[1]),
    .A2(_0068_),
    .ZN(_0294_)
  );
  INV_X1 _1018_ (
    .A(_0294_),
    .ZN(_0295_)
  );
  AND2_X1 _1019_ (
    .A1(_0035_),
    .A2(io_bp_0_address[1]),
    .ZN(_0296_)
  );
  INV_X1 _1020_ (
    .A(_0296_),
    .ZN(_0297_)
  );
  AND2_X1 _1021_ (
    .A1(_0295_),
    .A2(_0297_),
    .ZN(_0298_)
  );
  INV_X1 _1022_ (
    .A(_0298_),
    .ZN(_0299_)
  );
  AND2_X1 _1023_ (
    .A1(_0257_),
    .A2(_0299_),
    .ZN(_0300_)
  );
  INV_X1 _1024_ (
    .A(_0300_),
    .ZN(_0301_)
  );
  AND2_X1 _1025_ (
    .A1(_0036_),
    .A2(io_bp_0_address[2]),
    .ZN(_0302_)
  );
  INV_X1 _1026_ (
    .A(_0302_),
    .ZN(_0303_)
  );
  AND2_X1 _1027_ (
    .A1(io_pc[2]),
    .A2(_0069_),
    .ZN(_0304_)
  );
  INV_X1 _1028_ (
    .A(_0304_),
    .ZN(_0305_)
  );
  AND2_X1 _1029_ (
    .A1(_0303_),
    .A2(_0305_),
    .ZN(_0306_)
  );
  AND2_X1 _1030_ (
    .A1(_0301_),
    .A2(_0306_),
    .ZN(_0307_)
  );
  INV_X1 _1031_ (
    .A(_0307_),
    .ZN(_0308_)
  );
  AND2_X1 _1032_ (
    .A1(_0259_),
    .A2(_0308_),
    .ZN(_0309_)
  );
  INV_X1 _1033_ (
    .A(_0309_),
    .ZN(_0310_)
  );
  AND2_X1 _1034_ (
    .A1(_0269_),
    .A2(_0310_),
    .ZN(_0311_)
  );
  AND2_X1 _1035_ (
    .A1(_0230_),
    .A2(_0255_),
    .ZN(_0312_)
  );
  AND2_X1 _1036_ (
    .A1(_0293_),
    .A2(_0312_),
    .ZN(_0313_)
  );
  AND2_X1 _1037_ (
    .A1(_0311_),
    .A2(_0313_),
    .ZN(_0314_)
  );
  AND2_X1 _1038_ (
    .A1(_0197_),
    .A2(_0314_),
    .ZN(_0315_)
  );
  INV_X1 _1039_ (
    .A(_0315_),
    .ZN(_0316_)
  );
  AND2_X1 _1040_ (
    .A1(_0215_),
    .A2(_0295_),
    .ZN(_0317_)
  );
  INV_X1 _1041_ (
    .A(_0317_),
    .ZN(_0318_)
  );
  AND2_X1 _1042_ (
    .A1(_0297_),
    .A2(_0303_),
    .ZN(_0319_)
  );
  AND2_X1 _1043_ (
    .A1(_0318_),
    .A2(_0319_),
    .ZN(_0320_)
  );
  INV_X1 _1044_ (
    .A(_0320_),
    .ZN(_0321_)
  );
  AND2_X1 _1045_ (
    .A1(_0265_),
    .A2(_0305_),
    .ZN(_0322_)
  );
  AND2_X1 _1046_ (
    .A1(_0321_),
    .A2(_0322_),
    .ZN(_0323_)
  );
  INV_X1 _1047_ (
    .A(_0323_),
    .ZN(_0324_)
  );
  AND2_X1 _1048_ (
    .A1(_0263_),
    .A2(_0324_),
    .ZN(_0325_)
  );
  INV_X1 _1049_ (
    .A(_0325_),
    .ZN(_0326_)
  );
  AND2_X1 _1050_ (
    .A1(_0224_),
    .A2(_0326_),
    .ZN(_0327_)
  );
  INV_X1 _1051_ (
    .A(_0327_),
    .ZN(_0328_)
  );
  AND2_X1 _1052_ (
    .A1(_0212_),
    .A2(_0328_),
    .ZN(_0329_)
  );
  INV_X1 _1053_ (
    .A(_0329_),
    .ZN(_0330_)
  );
  AND2_X1 _1054_ (
    .A1(_0202_),
    .A2(_0330_),
    .ZN(_0331_)
  );
  INV_X1 _1055_ (
    .A(_0331_),
    .ZN(_0332_)
  );
  AND2_X1 _1056_ (
    .A1(_0207_),
    .A2(_0332_),
    .ZN(_0333_)
  );
  INV_X1 _1057_ (
    .A(_0333_),
    .ZN(_0334_)
  );
  AND2_X1 _1058_ (
    .A1(_0226_),
    .A2(_0334_),
    .ZN(_0335_)
  );
  INV_X1 _1059_ (
    .A(_0335_),
    .ZN(_0336_)
  );
  AND2_X1 _1060_ (
    .A1(_0255_),
    .A2(_0336_),
    .ZN(_0337_)
  );
  INV_X1 _1061_ (
    .A(_0337_),
    .ZN(_0338_)
  );
  AND2_X1 _1062_ (
    .A1(_0236_),
    .A2(_0238_),
    .ZN(_0339_)
  );
  INV_X1 _1063_ (
    .A(_0339_),
    .ZN(_0340_)
  );
  AND2_X1 _1064_ (
    .A1(_0244_),
    .A2(_0253_),
    .ZN(_0341_)
  );
  AND2_X1 _1065_ (
    .A1(_0242_),
    .A2(_0341_),
    .ZN(_0342_)
  );
  INV_X1 _1066_ (
    .A(_0342_),
    .ZN(_0343_)
  );
  AND2_X1 _1067_ (
    .A1(_0340_),
    .A2(_0343_),
    .ZN(_0344_)
  );
  AND2_X1 _1068_ (
    .A1(_0338_),
    .A2(_0344_),
    .ZN(_0345_)
  );
  INV_X1 _1069_ (
    .A(_0345_),
    .ZN(_0346_)
  );
  AND2_X1 _1070_ (
    .A1(_0293_),
    .A2(_0346_),
    .ZN(_0347_)
  );
  INV_X1 _1071_ (
    .A(_0347_),
    .ZN(_0348_)
  );
  AND2_X1 _1072_ (
    .A1(_0283_),
    .A2(_0291_),
    .ZN(_0349_)
  );
  INV_X1 _1073_ (
    .A(_0349_),
    .ZN(_0350_)
  );
  AND2_X1 _1074_ (
    .A1(_0273_),
    .A2(_0274_),
    .ZN(_0351_)
  );
  INV_X1 _1075_ (
    .A(_0351_),
    .ZN(_0352_)
  );
  AND2_X1 _1076_ (
    .A1(_0279_),
    .A2(_0352_),
    .ZN(_0353_)
  );
  AND2_X1 _1077_ (
    .A1(_0350_),
    .A2(_0353_),
    .ZN(_0354_)
  );
  AND2_X1 _1078_ (
    .A1(_0348_),
    .A2(_0354_),
    .ZN(_0355_)
  );
  INV_X1 _1079_ (
    .A(_0355_),
    .ZN(_0356_)
  );
  AND2_X1 _1080_ (
    .A1(_0197_),
    .A2(_0356_),
    .ZN(_0357_)
  );
  INV_X1 _1081_ (
    .A(_0357_),
    .ZN(_0358_)
  );
  AND2_X1 _1082_ (
    .A1(_0175_),
    .A2(_0179_),
    .ZN(_0359_)
  );
  INV_X1 _1083_ (
    .A(_0359_),
    .ZN(_0360_)
  );
  AND2_X1 _1084_ (
    .A1(_0173_),
    .A2(_0360_),
    .ZN(_0361_)
  );
  AND2_X1 _1085_ (
    .A1(_0184_),
    .A2(_0193_),
    .ZN(_0362_)
  );
  AND2_X1 _1086_ (
    .A1(_0182_),
    .A2(_0362_),
    .ZN(_0363_)
  );
  INV_X1 _1087_ (
    .A(_0363_),
    .ZN(_0364_)
  );
  AND2_X1 _1088_ (
    .A1(_0361_),
    .A2(_0364_),
    .ZN(_0365_)
  );
  INV_X1 _1089_ (
    .A(_0365_),
    .ZN(_0366_)
  );
  AND2_X1 _1090_ (
    .A1(_0130_),
    .A2(_0165_),
    .ZN(_0367_)
  );
  INV_X1 _1091_ (
    .A(_0367_),
    .ZN(_0368_)
  );
  AND2_X1 _1092_ (
    .A1(_0126_),
    .A2(_0368_),
    .ZN(_0369_)
  );
  INV_X1 _1093_ (
    .A(_0369_),
    .ZN(_0370_)
  );
  AND2_X1 _1094_ (
    .A1(_0158_),
    .A2(_0370_),
    .ZN(_0371_)
  );
  INV_X1 _1095_ (
    .A(_0371_),
    .ZN(_0372_)
  );
  AND2_X1 _1096_ (
    .A1(_0151_),
    .A2(_0155_),
    .ZN(_0373_)
  );
  INV_X1 _1097_ (
    .A(_0373_),
    .ZN(_0374_)
  );
  AND2_X1 _1098_ (
    .A1(_0149_),
    .A2(_0167_),
    .ZN(_0375_)
  );
  AND2_X1 _1099_ (
    .A1(_0374_),
    .A2(_0375_),
    .ZN(_0376_)
  );
  AND2_X1 _1100_ (
    .A1(_0372_),
    .A2(_0376_),
    .ZN(_0377_)
  );
  INV_X1 _1101_ (
    .A(_0377_),
    .ZN(_0378_)
  );
  AND2_X1 _1102_ (
    .A1(_0133_),
    .A2(_0378_),
    .ZN(_0379_)
  );
  INV_X1 _1103_ (
    .A(_0379_),
    .ZN(_0380_)
  );
  AND2_X1 _1104_ (
    .A1(_0162_),
    .A2(_0380_),
    .ZN(_0381_)
  );
  INV_X1 _1105_ (
    .A(_0381_),
    .ZN(_0382_)
  );
  AND2_X1 _1106_ (
    .A1(_0140_),
    .A2(_0382_),
    .ZN(_0383_)
  );
  INV_X1 _1107_ (
    .A(_0383_),
    .ZN(_0384_)
  );
  AND2_X1 _1108_ (
    .A1(_0145_),
    .A2(_0384_),
    .ZN(_0385_)
  );
  INV_X1 _1109_ (
    .A(_0385_),
    .ZN(_0386_)
  );
  AND2_X1 _1110_ (
    .A1(_0119_),
    .A2(_0122_),
    .ZN(_0387_)
  );
  AND2_X1 _1111_ (
    .A1(_0111_),
    .A2(_0387_),
    .ZN(_0388_)
  );
  INV_X1 _1112_ (
    .A(_0388_),
    .ZN(_0389_)
  );
  AND2_X1 _1113_ (
    .A1(_0105_),
    .A2(_0109_),
    .ZN(_0390_)
  );
  INV_X1 _1114_ (
    .A(_0390_),
    .ZN(_0391_)
  );
  AND2_X1 _1115_ (
    .A1(_0124_),
    .A2(_0366_),
    .ZN(_0392_)
  );
  INV_X1 _1116_ (
    .A(_0392_),
    .ZN(_0393_)
  );
  AND2_X1 _1117_ (
    .A1(_0389_),
    .A2(_0393_),
    .ZN(_0394_)
  );
  AND2_X1 _1118_ (
    .A1(_0160_),
    .A2(_0196_),
    .ZN(_0395_)
  );
  AND2_X1 _1119_ (
    .A1(_0386_),
    .A2(_0395_),
    .ZN(_0396_)
  );
  INV_X1 _1120_ (
    .A(_0396_),
    .ZN(_0397_)
  );
  AND2_X1 _1121_ (
    .A1(_0391_),
    .A2(_0397_),
    .ZN(_0398_)
  );
  AND2_X1 _1122_ (
    .A1(_0394_),
    .A2(_0398_),
    .ZN(_0399_)
  );
  AND2_X1 _1123_ (
    .A1(_0358_),
    .A2(_0399_),
    .ZN(_0400_)
  );
  INV_X1 _1124_ (
    .A(_0400_),
    .ZN(_0401_)
  );
  AND2_X1 _1125_ (
    .A1(_0099_),
    .A2(_0400_),
    .ZN(_0402_)
  );
  INV_X1 _1126_ (
    .A(_0402_),
    .ZN(_0403_)
  );
  AND2_X1 _1127_ (
    .A1(io_bp_0_control_tmatch[0]),
    .A2(_0401_),
    .ZN(_0404_)
  );
  INV_X1 _1128_ (
    .A(_0404_),
    .ZN(_0405_)
  );
  AND2_X1 _1129_ (
    .A1(_0403_),
    .A2(_0405_),
    .ZN(_0406_)
  );
  AND2_X1 _1130_ (
    .A1(io_bp_0_control_tmatch[1]),
    .A2(_0406_),
    .ZN(_0407_)
  );
  INV_X1 _1131_ (
    .A(_0407_),
    .ZN(_0408_)
  );
  AND2_X1 _1132_ (
    .A1(_0316_),
    .A2(_0408_),
    .ZN(_0409_)
  );
  INV_X1 _1133_ (
    .A(_0409_),
    .ZN(_0410_)
  );
  AND2_X1 _1134_ (
    .A1(_0001_),
    .A2(io_bp_0_control_x),
    .ZN(_0411_)
  );
  AND2_X1 _1135_ (
    .A1(_0410_),
    .A2(_0411_),
    .ZN(_0412_)
  );
  AND2_X1 _1136_ (
    .A1(_0066_),
    .A2(_0412_),
    .ZN(io_xcpt_if)
  );
  AND2_X1 _1137_ (
    .A1(io_ea[31]),
    .A2(_0098_),
    .ZN(_0413_)
  );
  INV_X1 _1138_ (
    .A(_0413_),
    .ZN(_0414_)
  );
  AND2_X1 _1139_ (
    .A1(io_ea[28]),
    .A2(_0095_),
    .ZN(_0415_)
  );
  INV_X1 _1140_ (
    .A(_0415_),
    .ZN(_0416_)
  );
  AND2_X1 _1141_ (
    .A1(_0414_),
    .A2(_0416_),
    .ZN(_0417_)
  );
  AND2_X1 _1142_ (
    .A1(io_ea[30]),
    .A2(_0097_),
    .ZN(_0418_)
  );
  INV_X1 _1143_ (
    .A(_0418_),
    .ZN(_0419_)
  );
  AND2_X1 _1144_ (
    .A1(_0027_),
    .A2(io_bp_0_address[25]),
    .ZN(_0420_)
  );
  INV_X1 _1145_ (
    .A(_0420_),
    .ZN(_0421_)
  );
  AND2_X1 _1146_ (
    .A1(_0419_),
    .A2(_0421_),
    .ZN(_0422_)
  );
  AND2_X1 _1147_ (
    .A1(_0417_),
    .A2(_0422_),
    .ZN(_0423_)
  );
  AND2_X1 _1148_ (
    .A1(_0033_),
    .A2(io_bp_0_address[31]),
    .ZN(_0424_)
  );
  INV_X1 _1149_ (
    .A(_0424_),
    .ZN(_0425_)
  );
  AND2_X1 _1150_ (
    .A1(_0032_),
    .A2(io_bp_0_address[30]),
    .ZN(_0426_)
  );
  INV_X1 _1151_ (
    .A(_0426_),
    .ZN(_0427_)
  );
  AND2_X1 _1152_ (
    .A1(_0425_),
    .A2(_0427_),
    .ZN(_0428_)
  );
  AND2_X1 _1153_ (
    .A1(_0031_),
    .A2(io_bp_0_address[29]),
    .ZN(_0429_)
  );
  INV_X1 _1154_ (
    .A(_0429_),
    .ZN(_0430_)
  );
  AND2_X1 _1155_ (
    .A1(_0030_),
    .A2(io_bp_0_address[28]),
    .ZN(_0431_)
  );
  INV_X1 _1156_ (
    .A(_0431_),
    .ZN(_0432_)
  );
  AND2_X1 _1157_ (
    .A1(_0430_),
    .A2(_0432_),
    .ZN(_0433_)
  );
  AND2_X1 _1158_ (
    .A1(_0428_),
    .A2(_0433_),
    .ZN(_0434_)
  );
  AND2_X1 _1159_ (
    .A1(_0423_),
    .A2(_0434_),
    .ZN(_0435_)
  );
  AND2_X1 _1160_ (
    .A1(io_ea[27]),
    .A2(_0094_),
    .ZN(_0436_)
  );
  INV_X1 _1161_ (
    .A(_0436_),
    .ZN(_0437_)
  );
  AND2_X1 _1162_ (
    .A1(_0029_),
    .A2(io_bp_0_address[27]),
    .ZN(_0438_)
  );
  INV_X1 _1163_ (
    .A(_0438_),
    .ZN(_0439_)
  );
  AND2_X1 _1164_ (
    .A1(_0437_),
    .A2(_0439_),
    .ZN(_0440_)
  );
  AND2_X1 _1165_ (
    .A1(_0028_),
    .A2(io_bp_0_address[26]),
    .ZN(_0441_)
  );
  INV_X1 _1166_ (
    .A(_0441_),
    .ZN(_0442_)
  );
  AND2_X1 _1167_ (
    .A1(io_ea[26]),
    .A2(_0093_),
    .ZN(_0443_)
  );
  INV_X1 _1168_ (
    .A(_0443_),
    .ZN(_0444_)
  );
  AND2_X1 _1169_ (
    .A1(_0442_),
    .A2(_0444_),
    .ZN(_0445_)
  );
  AND2_X1 _1170_ (
    .A1(_0440_),
    .A2(_0445_),
    .ZN(_0446_)
  );
  AND2_X1 _1171_ (
    .A1(_0026_),
    .A2(io_bp_0_address[24]),
    .ZN(_0447_)
  );
  INV_X1 _1172_ (
    .A(_0447_),
    .ZN(_0448_)
  );
  AND2_X1 _1173_ (
    .A1(io_ea[25]),
    .A2(_0092_),
    .ZN(_0449_)
  );
  INV_X1 _1174_ (
    .A(_0449_),
    .ZN(_0450_)
  );
  AND2_X1 _1175_ (
    .A1(_0448_),
    .A2(_0450_),
    .ZN(_0451_)
  );
  AND2_X1 _1176_ (
    .A1(io_ea[29]),
    .A2(_0096_),
    .ZN(_0452_)
  );
  INV_X1 _1177_ (
    .A(_0452_),
    .ZN(_0453_)
  );
  AND2_X1 _1178_ (
    .A1(io_ea[24]),
    .A2(_0091_),
    .ZN(_0454_)
  );
  INV_X1 _1179_ (
    .A(_0454_),
    .ZN(_0455_)
  );
  AND2_X1 _1180_ (
    .A1(_0453_),
    .A2(_0455_),
    .ZN(_0456_)
  );
  AND2_X1 _1181_ (
    .A1(_0451_),
    .A2(_0456_),
    .ZN(_0457_)
  );
  AND2_X1 _1182_ (
    .A1(_0446_),
    .A2(_0457_),
    .ZN(_0458_)
  );
  AND2_X1 _1183_ (
    .A1(_0435_),
    .A2(_0458_),
    .ZN(_0459_)
  );
  AND2_X1 _1184_ (
    .A1(_0024_),
    .A2(io_bp_0_address[22]),
    .ZN(_0460_)
  );
  INV_X1 _1185_ (
    .A(_0460_),
    .ZN(_0461_)
  );
  AND2_X1 _1186_ (
    .A1(_0023_),
    .A2(io_bp_0_address[21]),
    .ZN(_0462_)
  );
  INV_X1 _1187_ (
    .A(_0462_),
    .ZN(_0463_)
  );
  AND2_X1 _1188_ (
    .A1(_0461_),
    .A2(_0463_),
    .ZN(_0464_)
  );
  AND2_X1 _1189_ (
    .A1(io_ea[21]),
    .A2(_0088_),
    .ZN(_0465_)
  );
  INV_X1 _1190_ (
    .A(_0465_),
    .ZN(_0466_)
  );
  AND2_X1 _1191_ (
    .A1(_0018_),
    .A2(io_bp_0_address[16]),
    .ZN(_0467_)
  );
  INV_X1 _1192_ (
    .A(_0467_),
    .ZN(_0468_)
  );
  AND2_X1 _1193_ (
    .A1(_0466_),
    .A2(_0468_),
    .ZN(_0469_)
  );
  AND2_X1 _1194_ (
    .A1(_0464_),
    .A2(_0469_),
    .ZN(_0470_)
  );
  AND2_X1 _1195_ (
    .A1(io_ea[23]),
    .A2(_0090_),
    .ZN(_0471_)
  );
  INV_X1 _1196_ (
    .A(_0471_),
    .ZN(_0472_)
  );
  AND2_X1 _1197_ (
    .A1(io_ea[22]),
    .A2(_0089_),
    .ZN(_0473_)
  );
  INV_X1 _1198_ (
    .A(_0473_),
    .ZN(_0474_)
  );
  AND2_X1 _1199_ (
    .A1(_0472_),
    .A2(_0474_),
    .ZN(_0475_)
  );
  AND2_X1 _1200_ (
    .A1(io_ea[17]),
    .A2(_0084_),
    .ZN(_0476_)
  );
  INV_X1 _1201_ (
    .A(_0476_),
    .ZN(_0477_)
  );
  AND2_X1 _1202_ (
    .A1(io_ea[16]),
    .A2(_0083_),
    .ZN(_0478_)
  );
  INV_X1 _1203_ (
    .A(_0478_),
    .ZN(_0479_)
  );
  AND2_X1 _1204_ (
    .A1(_0477_),
    .A2(_0479_),
    .ZN(_0480_)
  );
  INV_X1 _1205_ (
    .A(_0480_),
    .ZN(_0481_)
  );
  AND2_X1 _1206_ (
    .A1(_0475_),
    .A2(_0480_),
    .ZN(_0482_)
  );
  AND2_X1 _1207_ (
    .A1(_0470_),
    .A2(_0482_),
    .ZN(_0483_)
  );
  AND2_X1 _1208_ (
    .A1(io_ea[19]),
    .A2(_0086_),
    .ZN(_0484_)
  );
  INV_X1 _1209_ (
    .A(_0484_),
    .ZN(_0485_)
  );
  AND2_X1 _1210_ (
    .A1(io_ea[18]),
    .A2(_0085_),
    .ZN(_0486_)
  );
  INV_X1 _1211_ (
    .A(_0486_),
    .ZN(_0487_)
  );
  AND2_X1 _1212_ (
    .A1(_0485_),
    .A2(_0487_),
    .ZN(_0488_)
  );
  INV_X1 _1213_ (
    .A(_0488_),
    .ZN(_0489_)
  );
  AND2_X1 _1214_ (
    .A1(_0021_),
    .A2(io_bp_0_address[19]),
    .ZN(_0490_)
  );
  INV_X1 _1215_ (
    .A(_0490_),
    .ZN(_0491_)
  );
  AND2_X1 _1216_ (
    .A1(_0020_),
    .A2(io_bp_0_address[18]),
    .ZN(_0492_)
  );
  INV_X1 _1217_ (
    .A(_0492_),
    .ZN(_0493_)
  );
  AND2_X1 _1218_ (
    .A1(_0491_),
    .A2(_0493_),
    .ZN(_0494_)
  );
  AND2_X1 _1219_ (
    .A1(_0488_),
    .A2(_0494_),
    .ZN(_0495_)
  );
  AND2_X1 _1220_ (
    .A1(_0025_),
    .A2(io_bp_0_address[23]),
    .ZN(_0496_)
  );
  INV_X1 _1221_ (
    .A(_0496_),
    .ZN(_0497_)
  );
  AND2_X1 _1222_ (
    .A1(io_ea[20]),
    .A2(_0087_),
    .ZN(_0498_)
  );
  INV_X1 _1223_ (
    .A(_0498_),
    .ZN(_0499_)
  );
  AND2_X1 _1224_ (
    .A1(_0497_),
    .A2(_0499_),
    .ZN(_0500_)
  );
  AND2_X1 _1225_ (
    .A1(_0022_),
    .A2(io_bp_0_address[20]),
    .ZN(_0501_)
  );
  INV_X1 _1226_ (
    .A(_0501_),
    .ZN(_0502_)
  );
  AND2_X1 _1227_ (
    .A1(_0019_),
    .A2(io_bp_0_address[17]),
    .ZN(_0503_)
  );
  INV_X1 _1228_ (
    .A(_0503_),
    .ZN(_0504_)
  );
  AND2_X1 _1229_ (
    .A1(_0502_),
    .A2(_0504_),
    .ZN(_0505_)
  );
  AND2_X1 _1230_ (
    .A1(_0500_),
    .A2(_0505_),
    .ZN(_0506_)
  );
  AND2_X1 _1231_ (
    .A1(_0495_),
    .A2(_0506_),
    .ZN(_0507_)
  );
  AND2_X1 _1232_ (
    .A1(_0483_),
    .A2(_0507_),
    .ZN(_0508_)
  );
  AND2_X1 _1233_ (
    .A1(_0459_),
    .A2(_0508_),
    .ZN(_0509_)
  );
  AND2_X1 _1234_ (
    .A1(io_ea[14]),
    .A2(_0081_),
    .ZN(_0510_)
  );
  INV_X1 _1235_ (
    .A(_0510_),
    .ZN(_0511_)
  );
  AND2_X1 _1236_ (
    .A1(_0011_),
    .A2(io_bp_0_address[9]),
    .ZN(_0512_)
  );
  INV_X1 _1237_ (
    .A(_0512_),
    .ZN(_0513_)
  );
  AND2_X1 _1238_ (
    .A1(_0511_),
    .A2(_0513_),
    .ZN(_0514_)
  );
  AND2_X1 _1239_ (
    .A1(_0015_),
    .A2(io_bp_0_address[13]),
    .ZN(_0515_)
  );
  INV_X1 _1240_ (
    .A(_0515_),
    .ZN(_0516_)
  );
  AND2_X1 _1241_ (
    .A1(io_ea[12]),
    .A2(_0079_),
    .ZN(_0517_)
  );
  INV_X1 _1242_ (
    .A(_0517_),
    .ZN(_0518_)
  );
  AND2_X1 _1243_ (
    .A1(_0516_),
    .A2(_0518_),
    .ZN(_0519_)
  );
  AND2_X1 _1244_ (
    .A1(_0514_),
    .A2(_0519_),
    .ZN(_0520_)
  );
  AND2_X1 _1245_ (
    .A1(_0017_),
    .A2(io_bp_0_address[15]),
    .ZN(_0521_)
  );
  INV_X1 _1246_ (
    .A(_0521_),
    .ZN(_0522_)
  );
  AND2_X1 _1247_ (
    .A1(_0016_),
    .A2(io_bp_0_address[14]),
    .ZN(_0523_)
  );
  INV_X1 _1248_ (
    .A(_0523_),
    .ZN(_0524_)
  );
  AND2_X1 _1249_ (
    .A1(_0522_),
    .A2(_0524_),
    .ZN(_0525_)
  );
  AND2_X1 _1250_ (
    .A1(io_ea[15]),
    .A2(_0082_),
    .ZN(_0526_)
  );
  INV_X1 _1251_ (
    .A(_0526_),
    .ZN(_0527_)
  );
  AND2_X1 _1252_ (
    .A1(io_ea[13]),
    .A2(_0080_),
    .ZN(_0528_)
  );
  INV_X1 _1253_ (
    .A(_0528_),
    .ZN(_0529_)
  );
  AND2_X1 _1254_ (
    .A1(_0527_),
    .A2(_0529_),
    .ZN(_0530_)
  );
  AND2_X1 _1255_ (
    .A1(_0525_),
    .A2(_0530_),
    .ZN(_0531_)
  );
  AND2_X1 _1256_ (
    .A1(_0520_),
    .A2(_0531_),
    .ZN(_0532_)
  );
  AND2_X1 _1257_ (
    .A1(io_ea[11]),
    .A2(_0078_),
    .ZN(_0533_)
  );
  INV_X1 _1258_ (
    .A(_0533_),
    .ZN(_0534_)
  );
  AND2_X1 _1259_ (
    .A1(_0013_),
    .A2(io_bp_0_address[11]),
    .ZN(_0535_)
  );
  INV_X1 _1260_ (
    .A(_0535_),
    .ZN(_0536_)
  );
  AND2_X1 _1261_ (
    .A1(_0534_),
    .A2(_0536_),
    .ZN(_0537_)
  );
  AND2_X1 _1262_ (
    .A1(_0012_),
    .A2(io_bp_0_address[10]),
    .ZN(_0538_)
  );
  INV_X1 _1263_ (
    .A(_0538_),
    .ZN(_0539_)
  );
  AND2_X1 _1264_ (
    .A1(io_ea[10]),
    .A2(_0077_),
    .ZN(_0540_)
  );
  INV_X1 _1265_ (
    .A(_0540_),
    .ZN(_0541_)
  );
  AND2_X1 _1266_ (
    .A1(_0539_),
    .A2(_0541_),
    .ZN(_0542_)
  );
  AND2_X1 _1267_ (
    .A1(_0537_),
    .A2(_0542_),
    .ZN(_0543_)
  );
  AND2_X1 _1268_ (
    .A1(_0010_),
    .A2(io_bp_0_address[8]),
    .ZN(_0544_)
  );
  INV_X1 _1269_ (
    .A(_0544_),
    .ZN(_0545_)
  );
  AND2_X1 _1270_ (
    .A1(io_ea[9]),
    .A2(_0076_),
    .ZN(_0546_)
  );
  INV_X1 _1271_ (
    .A(_0546_),
    .ZN(_0547_)
  );
  AND2_X1 _1272_ (
    .A1(_0545_),
    .A2(_0547_),
    .ZN(_0548_)
  );
  AND2_X1 _1273_ (
    .A1(_0014_),
    .A2(io_bp_0_address[12]),
    .ZN(_0549_)
  );
  INV_X1 _1274_ (
    .A(_0549_),
    .ZN(_0550_)
  );
  AND2_X1 _1275_ (
    .A1(io_ea[8]),
    .A2(_0075_),
    .ZN(_0551_)
  );
  INV_X1 _1276_ (
    .A(_0551_),
    .ZN(_0552_)
  );
  AND2_X1 _1277_ (
    .A1(_0550_),
    .A2(_0552_),
    .ZN(_0553_)
  );
  AND2_X1 _1278_ (
    .A1(_0548_),
    .A2(_0553_),
    .ZN(_0554_)
  );
  AND2_X1 _1279_ (
    .A1(_0543_),
    .A2(_0554_),
    .ZN(_0555_)
  );
  AND2_X1 _1280_ (
    .A1(_0532_),
    .A2(_0555_),
    .ZN(_0556_)
  );
  AND2_X1 _1281_ (
    .A1(io_ea[7]),
    .A2(_0074_),
    .ZN(_0557_)
  );
  INV_X1 _1282_ (
    .A(_0557_),
    .ZN(_0558_)
  );
  AND2_X1 _1283_ (
    .A1(_0009_),
    .A2(io_bp_0_address[7]),
    .ZN(_0559_)
  );
  INV_X1 _1284_ (
    .A(_0559_),
    .ZN(_0560_)
  );
  AND2_X1 _1285_ (
    .A1(_0008_),
    .A2(io_bp_0_address[6]),
    .ZN(_0561_)
  );
  INV_X1 _1286_ (
    .A(_0561_),
    .ZN(_0562_)
  );
  AND2_X1 _1287_ (
    .A1(_0560_),
    .A2(_0562_),
    .ZN(_0563_)
  );
  AND2_X1 _1288_ (
    .A1(io_ea[6]),
    .A2(_0073_),
    .ZN(_0564_)
  );
  INV_X1 _1289_ (
    .A(_0564_),
    .ZN(_0565_)
  );
  AND2_X1 _1290_ (
    .A1(io_ea[5]),
    .A2(_0072_),
    .ZN(_0566_)
  );
  INV_X1 _1291_ (
    .A(_0566_),
    .ZN(_0567_)
  );
  AND2_X1 _1292_ (
    .A1(_0565_),
    .A2(_0567_),
    .ZN(_0568_)
  );
  AND2_X1 _1293_ (
    .A1(io_ea[4]),
    .A2(_0071_),
    .ZN(_0569_)
  );
  INV_X1 _1294_ (
    .A(_0569_),
    .ZN(_0570_)
  );
  AND2_X1 _1295_ (
    .A1(_0005_),
    .A2(io_bp_0_address[3]),
    .ZN(_0571_)
  );
  INV_X1 _1296_ (
    .A(_0571_),
    .ZN(_0572_)
  );
  AND2_X1 _1297_ (
    .A1(io_ea[1]),
    .A2(_0068_),
    .ZN(_0573_)
  );
  INV_X1 _1298_ (
    .A(_0573_),
    .ZN(_0574_)
  );
  AND2_X1 _1299_ (
    .A1(_0002_),
    .A2(io_bp_0_address[0]),
    .ZN(_0575_)
  );
  INV_X1 _1300_ (
    .A(_0575_),
    .ZN(_0576_)
  );
  AND2_X1 _1301_ (
    .A1(_0574_),
    .A2(_0575_),
    .ZN(_0577_)
  );
  INV_X1 _1302_ (
    .A(_0577_),
    .ZN(_0578_)
  );
  AND2_X1 _1303_ (
    .A1(_0004_),
    .A2(io_bp_0_address[2]),
    .ZN(_0579_)
  );
  INV_X1 _1304_ (
    .A(_0579_),
    .ZN(_0580_)
  );
  AND2_X1 _1305_ (
    .A1(_0003_),
    .A2(io_bp_0_address[1]),
    .ZN(_0581_)
  );
  INV_X1 _1306_ (
    .A(_0581_),
    .ZN(_0582_)
  );
  AND2_X1 _1307_ (
    .A1(_0580_),
    .A2(_0582_),
    .ZN(_0583_)
  );
  AND2_X1 _1308_ (
    .A1(_0578_),
    .A2(_0583_),
    .ZN(_0584_)
  );
  INV_X1 _1309_ (
    .A(_0584_),
    .ZN(_0585_)
  );
  AND2_X1 _1310_ (
    .A1(io_ea[3]),
    .A2(_0070_),
    .ZN(_0586_)
  );
  INV_X1 _1311_ (
    .A(_0586_),
    .ZN(_0587_)
  );
  AND2_X1 _1312_ (
    .A1(io_ea[2]),
    .A2(_0069_),
    .ZN(_0588_)
  );
  INV_X1 _1313_ (
    .A(_0588_),
    .ZN(_0589_)
  );
  AND2_X1 _1314_ (
    .A1(_0587_),
    .A2(_0589_),
    .ZN(_0590_)
  );
  AND2_X1 _1315_ (
    .A1(_0585_),
    .A2(_0590_),
    .ZN(_0591_)
  );
  INV_X1 _1316_ (
    .A(_0591_),
    .ZN(_0592_)
  );
  AND2_X1 _1317_ (
    .A1(_0572_),
    .A2(_0592_),
    .ZN(_0593_)
  );
  INV_X1 _1318_ (
    .A(_0593_),
    .ZN(_0594_)
  );
  AND2_X1 _1319_ (
    .A1(_0570_),
    .A2(_0594_),
    .ZN(_0595_)
  );
  INV_X1 _1320_ (
    .A(_0595_),
    .ZN(_0596_)
  );
  AND2_X1 _1321_ (
    .A1(_0007_),
    .A2(io_bp_0_address[5]),
    .ZN(_0597_)
  );
  INV_X1 _1322_ (
    .A(_0597_),
    .ZN(_0598_)
  );
  AND2_X1 _1323_ (
    .A1(_0006_),
    .A2(io_bp_0_address[4]),
    .ZN(_0599_)
  );
  INV_X1 _1324_ (
    .A(_0599_),
    .ZN(_0600_)
  );
  AND2_X1 _1325_ (
    .A1(_0598_),
    .A2(_0600_),
    .ZN(_0601_)
  );
  AND2_X1 _1326_ (
    .A1(_0596_),
    .A2(_0601_),
    .ZN(_0602_)
  );
  INV_X1 _1327_ (
    .A(_0602_),
    .ZN(_0603_)
  );
  AND2_X1 _1328_ (
    .A1(_0568_),
    .A2(_0603_),
    .ZN(_0604_)
  );
  INV_X1 _1329_ (
    .A(_0604_),
    .ZN(_0605_)
  );
  AND2_X1 _1330_ (
    .A1(_0563_),
    .A2(_0605_),
    .ZN(_0606_)
  );
  INV_X1 _1331_ (
    .A(_0606_),
    .ZN(_0607_)
  );
  AND2_X1 _1332_ (
    .A1(_0558_),
    .A2(_0607_),
    .ZN(_0608_)
  );
  INV_X1 _1333_ (
    .A(_0608_),
    .ZN(_0609_)
  );
  AND2_X1 _1334_ (
    .A1(_0556_),
    .A2(_0609_),
    .ZN(_0610_)
  );
  INV_X1 _1335_ (
    .A(_0610_),
    .ZN(_0611_)
  );
  AND2_X1 _1336_ (
    .A1(_0513_),
    .A2(_0551_),
    .ZN(_0612_)
  );
  INV_X1 _1337_ (
    .A(_0612_),
    .ZN(_0613_)
  );
  AND2_X1 _1338_ (
    .A1(_0547_),
    .A2(_0613_),
    .ZN(_0614_)
  );
  INV_X1 _1339_ (
    .A(_0614_),
    .ZN(_0615_)
  );
  AND2_X1 _1340_ (
    .A1(_0543_),
    .A2(_0615_),
    .ZN(_0616_)
  );
  INV_X1 _1341_ (
    .A(_0616_),
    .ZN(_0617_)
  );
  AND2_X1 _1342_ (
    .A1(_0536_),
    .A2(_0540_),
    .ZN(_0618_)
  );
  INV_X1 _1343_ (
    .A(_0618_),
    .ZN(_0619_)
  );
  AND2_X1 _1344_ (
    .A1(_0534_),
    .A2(_0619_),
    .ZN(_0620_)
  );
  AND2_X1 _1345_ (
    .A1(_0518_),
    .A2(_0620_),
    .ZN(_0621_)
  );
  AND2_X1 _1346_ (
    .A1(_0617_),
    .A2(_0621_),
    .ZN(_0622_)
  );
  INV_X1 _1347_ (
    .A(_0622_),
    .ZN(_0623_)
  );
  AND2_X1 _1348_ (
    .A1(_0516_),
    .A2(_0550_),
    .ZN(_0624_)
  );
  AND2_X1 _1349_ (
    .A1(_0623_),
    .A2(_0624_),
    .ZN(_0625_)
  );
  INV_X1 _1350_ (
    .A(_0625_),
    .ZN(_0626_)
  );
  AND2_X1 _1351_ (
    .A1(_0511_),
    .A2(_0529_),
    .ZN(_0627_)
  );
  AND2_X1 _1352_ (
    .A1(_0626_),
    .A2(_0627_),
    .ZN(_0628_)
  );
  INV_X1 _1353_ (
    .A(_0628_),
    .ZN(_0629_)
  );
  AND2_X1 _1354_ (
    .A1(_0525_),
    .A2(_0629_),
    .ZN(_0630_)
  );
  INV_X1 _1355_ (
    .A(_0630_),
    .ZN(_0631_)
  );
  AND2_X1 _1356_ (
    .A1(_0527_),
    .A2(_0631_),
    .ZN(_0632_)
  );
  AND2_X1 _1357_ (
    .A1(_0611_),
    .A2(_0632_),
    .ZN(_0633_)
  );
  INV_X1 _1358_ (
    .A(_0633_),
    .ZN(_0634_)
  );
  AND2_X1 _1359_ (
    .A1(_0509_),
    .A2(_0634_),
    .ZN(_0635_)
  );
  INV_X1 _1360_ (
    .A(_0635_),
    .ZN(_0636_)
  );
  AND2_X1 _1361_ (
    .A1(_0481_),
    .A2(_0504_),
    .ZN(_0637_)
  );
  AND2_X1 _1362_ (
    .A1(_0495_),
    .A2(_0637_),
    .ZN(_0638_)
  );
  INV_X1 _1363_ (
    .A(_0638_),
    .ZN(_0639_)
  );
  AND2_X1 _1364_ (
    .A1(_0489_),
    .A2(_0491_),
    .ZN(_0640_)
  );
  INV_X1 _1365_ (
    .A(_0640_),
    .ZN(_0641_)
  );
  AND2_X1 _1366_ (
    .A1(_0499_),
    .A2(_0641_),
    .ZN(_0642_)
  );
  AND2_X1 _1367_ (
    .A1(_0639_),
    .A2(_0642_),
    .ZN(_0643_)
  );
  INV_X1 _1368_ (
    .A(_0643_),
    .ZN(_0644_)
  );
  AND2_X1 _1369_ (
    .A1(_0502_),
    .A2(_0644_),
    .ZN(_0645_)
  );
  INV_X1 _1370_ (
    .A(_0645_),
    .ZN(_0646_)
  );
  AND2_X1 _1371_ (
    .A1(_0466_),
    .A2(_0646_),
    .ZN(_0647_)
  );
  INV_X1 _1372_ (
    .A(_0647_),
    .ZN(_0648_)
  );
  AND2_X1 _1373_ (
    .A1(_0464_),
    .A2(_0648_),
    .ZN(_0649_)
  );
  INV_X1 _1374_ (
    .A(_0649_),
    .ZN(_0650_)
  );
  AND2_X1 _1375_ (
    .A1(_0475_),
    .A2(_0650_),
    .ZN(_0651_)
  );
  INV_X1 _1376_ (
    .A(_0651_),
    .ZN(_0652_)
  );
  AND2_X1 _1377_ (
    .A1(_0459_),
    .A2(_0497_),
    .ZN(_0653_)
  );
  AND2_X1 _1378_ (
    .A1(_0652_),
    .A2(_0653_),
    .ZN(_0654_)
  );
  INV_X1 _1379_ (
    .A(_0654_),
    .ZN(_0655_)
  );
  AND2_X1 _1380_ (
    .A1(_0421_),
    .A2(_0454_),
    .ZN(_0656_)
  );
  INV_X1 _1381_ (
    .A(_0656_),
    .ZN(_0657_)
  );
  AND2_X1 _1382_ (
    .A1(_0450_),
    .A2(_0657_),
    .ZN(_0658_)
  );
  INV_X1 _1383_ (
    .A(_0658_),
    .ZN(_0659_)
  );
  AND2_X1 _1384_ (
    .A1(_0446_),
    .A2(_0659_),
    .ZN(_0660_)
  );
  INV_X1 _1385_ (
    .A(_0660_),
    .ZN(_0661_)
  );
  AND2_X1 _1386_ (
    .A1(_0439_),
    .A2(_0443_),
    .ZN(_0662_)
  );
  INV_X1 _1387_ (
    .A(_0662_),
    .ZN(_0663_)
  );
  AND2_X1 _1388_ (
    .A1(_0416_),
    .A2(_0437_),
    .ZN(_0664_)
  );
  AND2_X1 _1389_ (
    .A1(_0663_),
    .A2(_0664_),
    .ZN(_0665_)
  );
  AND2_X1 _1390_ (
    .A1(_0661_),
    .A2(_0665_),
    .ZN(_0666_)
  );
  INV_X1 _1391_ (
    .A(_0666_),
    .ZN(_0667_)
  );
  AND2_X1 _1392_ (
    .A1(_0433_),
    .A2(_0667_),
    .ZN(_0668_)
  );
  INV_X1 _1393_ (
    .A(_0668_),
    .ZN(_0669_)
  );
  AND2_X1 _1394_ (
    .A1(_0419_),
    .A2(_0453_),
    .ZN(_0670_)
  );
  AND2_X1 _1395_ (
    .A1(_0669_),
    .A2(_0670_),
    .ZN(_0671_)
  );
  INV_X1 _1396_ (
    .A(_0671_),
    .ZN(_0672_)
  );
  AND2_X1 _1397_ (
    .A1(_0428_),
    .A2(_0672_),
    .ZN(_0673_)
  );
  INV_X1 _1398_ (
    .A(_0673_),
    .ZN(_0674_)
  );
  AND2_X1 _1399_ (
    .A1(_0414_),
    .A2(_0674_),
    .ZN(_0675_)
  );
  AND2_X1 _1400_ (
    .A1(_0655_),
    .A2(_0675_),
    .ZN(_0676_)
  );
  AND2_X1 _1401_ (
    .A1(_0636_),
    .A2(_0676_),
    .ZN(_0677_)
  );
  INV_X1 _1402_ (
    .A(_0677_),
    .ZN(_0678_)
  );
  AND2_X1 _1403_ (
    .A1(io_bp_0_control_tmatch[0]),
    .A2(_0678_),
    .ZN(_0679_)
  );
  INV_X1 _1404_ (
    .A(_0679_),
    .ZN(_0680_)
  );
  AND2_X1 _1405_ (
    .A1(_0099_),
    .A2(_0677_),
    .ZN(_0681_)
  );
  INV_X1 _1406_ (
    .A(_0681_),
    .ZN(_0682_)
  );
  AND2_X1 _1407_ (
    .A1(io_bp_0_control_tmatch[1]),
    .A2(_0682_),
    .ZN(_0683_)
  );
  AND2_X1 _1408_ (
    .A1(_0680_),
    .A2(_0683_),
    .ZN(_0684_)
  );
  INV_X1 _1409_ (
    .A(_0684_),
    .ZN(_0685_)
  );
  AND2_X1 _1410_ (
    .A1(_0572_),
    .A2(_0587_),
    .ZN(_0686_)
  );
  INV_X1 _1411_ (
    .A(_0686_),
    .ZN(_0687_)
  );
  AND2_X1 _1412_ (
    .A1(_0261_),
    .A2(_0687_),
    .ZN(_0688_)
  );
  INV_X1 _1413_ (
    .A(_0688_),
    .ZN(_0689_)
  );
  AND2_X1 _1414_ (
    .A1(io_ea[0]),
    .A2(_0067_),
    .ZN(_0690_)
  );
  INV_X1 _1415_ (
    .A(_0690_),
    .ZN(_0691_)
  );
  AND2_X1 _1416_ (
    .A1(_0576_),
    .A2(_0691_),
    .ZN(_0692_)
  );
  INV_X1 _1417_ (
    .A(_0692_),
    .ZN(_0693_)
  );
  AND2_X1 _1418_ (
    .A1(_0099_),
    .A2(_0693_),
    .ZN(_0694_)
  );
  INV_X1 _1419_ (
    .A(_0694_),
    .ZN(_0695_)
  );
  AND2_X1 _1420_ (
    .A1(_0568_),
    .A2(_0600_),
    .ZN(_0696_)
  );
  AND2_X1 _1421_ (
    .A1(_0695_),
    .A2(_0696_),
    .ZN(_0697_)
  );
  AND2_X1 _1422_ (
    .A1(_0558_),
    .A2(_0570_),
    .ZN(_0698_)
  );
  AND2_X1 _1423_ (
    .A1(_0000_),
    .A2(_0598_),
    .ZN(_0699_)
  );
  AND2_X1 _1424_ (
    .A1(_0563_),
    .A2(_0699_),
    .ZN(_0700_)
  );
  AND2_X1 _1425_ (
    .A1(_0698_),
    .A2(_0700_),
    .ZN(_0701_)
  );
  AND2_X1 _1426_ (
    .A1(_0689_),
    .A2(_0701_),
    .ZN(_0702_)
  );
  AND2_X1 _1427_ (
    .A1(_0697_),
    .A2(_0702_),
    .ZN(_0703_)
  );
  AND2_X1 _1428_ (
    .A1(_0574_),
    .A2(_0582_),
    .ZN(_0704_)
  );
  INV_X1 _1429_ (
    .A(_0704_),
    .ZN(_0705_)
  );
  AND2_X1 _1430_ (
    .A1(_0257_),
    .A2(_0705_),
    .ZN(_0706_)
  );
  INV_X1 _1431_ (
    .A(_0706_),
    .ZN(_0707_)
  );
  AND2_X1 _1432_ (
    .A1(_0580_),
    .A2(_0589_),
    .ZN(_0708_)
  );
  AND2_X1 _1433_ (
    .A1(_0707_),
    .A2(_0708_),
    .ZN(_0709_)
  );
  INV_X1 _1434_ (
    .A(_0709_),
    .ZN(_0710_)
  );
  AND2_X1 _1435_ (
    .A1(_0259_),
    .A2(_0710_),
    .ZN(_0711_)
  );
  INV_X1 _1436_ (
    .A(_0711_),
    .ZN(_0712_)
  );
  AND2_X1 _1437_ (
    .A1(_0556_),
    .A2(_0703_),
    .ZN(_0713_)
  );
  AND2_X1 _1438_ (
    .A1(_0509_),
    .A2(_0712_),
    .ZN(_0714_)
  );
  AND2_X1 _1439_ (
    .A1(_0713_),
    .A2(_0714_),
    .ZN(_0715_)
  );
  INV_X1 _1440_ (
    .A(_0715_),
    .ZN(_0716_)
  );
  AND2_X1 _1441_ (
    .A1(_0685_),
    .A2(_0716_),
    .ZN(_0717_)
  );
  INV_X1 _1442_ (
    .A(_0717_),
    .ZN(_0718_)
  );
  AND2_X1 _1443_ (
    .A1(_0001_),
    .A2(io_bp_0_control_r),
    .ZN(_0719_)
  );
  AND2_X1 _1444_ (
    .A1(_0718_),
    .A2(_0719_),
    .ZN(_0720_)
  );
  AND2_X1 _1445_ (
    .A1(_0066_),
    .A2(_0720_),
    .ZN(io_xcpt_ld)
  );
  AND2_X1 _1446_ (
    .A1(_0001_),
    .A2(io_bp_0_control_w),
    .ZN(_0721_)
  );
  AND2_X1 _1447_ (
    .A1(_0718_),
    .A2(_0721_),
    .ZN(_0722_)
  );
  AND2_X1 _1448_ (
    .A1(_0066_),
    .A2(_0722_),
    .ZN(io_xcpt_st)
  );
  AND2_X1 _1449_ (
    .A1(io_bp_0_control_action),
    .A2(_0412_),
    .ZN(io_debug_if)
  );
  AND2_X1 _1450_ (
    .A1(io_bp_0_control_action),
    .A2(_0720_),
    .ZN(io_debug_ld)
  );
  AND2_X1 _1451_ (
    .A1(io_bp_0_control_action),
    .A2(_0722_),
    .ZN(io_debug_st)
  );
  assign { _GEN_11[31:4], _GEN_11[0] } = { 28'h0000000, io_bp_0_control_tmatch[0] };
  assign _r_T_10 = _GEN_11[2];
  assign _r_T_12 = _GEN_11[3];
  assign _r_T_13 = { _GEN_11[3:1], io_bp_0_control_tmatch[0] };
  assign _r_T_8 = _GEN_11[1];
endmodule
module CSRFile(clock, reset, io_ungated_clock, io_interrupts_debug, io_interrupts_mtip, io_interrupts_msip, io_interrupts_meip, io_hartid, io_rw_addr, io_rw_cmd, io_rw_rdata, io_rw_wdata, io_decode_0_inst, io_decode_0_fp_illegal, io_decode_0_fp_csr, io_decode_0_rocc_illegal, io_decode_0_read_illegal, io_decode_0_write_illegal, io_decode_0_write_flush, io_decode_0_system_illegal, io_csr_stall
, io_eret, io_singleStep, io_status_debug, io_status_cease, io_status_wfi, io_status_isa, io_status_dprv, io_status_dv, io_status_prv, io_status_v, io_status_sd, io_status_zero2, io_status_mpv, io_status_gva, io_status_mbe, io_status_sbe, io_status_sxl, io_status_uxl, io_status_sd_rv32, io_status_zero1, io_status_tsr
, io_status_tw, io_status_tvm, io_status_mxr, io_status_sum, io_status_mprv, io_status_xs, io_status_fs, io_status_mpp, io_status_vs, io_status_spp, io_status_mpie, io_status_ube, io_status_spie, io_status_upie, io_status_mie, io_status_hie, io_status_sie, io_status_uie, io_evec, io_exception, io_retire
, io_cause, io_pc, io_tval, io_gva, io_time, io_interrupt, io_interrupt_cause, io_bp_0_control_action, io_bp_0_control_tmatch, io_bp_0_control_x, io_bp_0_control_w, io_bp_0_control_r, io_bp_0_address, io_pmp_0_cfg_l, io_pmp_0_cfg_a, io_pmp_0_cfg_x, io_pmp_0_cfg_w, io_pmp_0_cfg_r, io_pmp_0_addr, io_pmp_0_mask, io_pmp_1_cfg_l
, io_pmp_1_cfg_a, io_pmp_1_cfg_x, io_pmp_1_cfg_w, io_pmp_1_cfg_r, io_pmp_1_addr, io_pmp_1_mask, io_pmp_2_cfg_l, io_pmp_2_cfg_a, io_pmp_2_cfg_x, io_pmp_2_cfg_w, io_pmp_2_cfg_r, io_pmp_2_addr, io_pmp_2_mask, io_pmp_3_cfg_l, io_pmp_3_cfg_a, io_pmp_3_cfg_x, io_pmp_3_cfg_w, io_pmp_3_cfg_r, io_pmp_3_addr, io_pmp_3_mask, io_pmp_4_cfg_l
, io_pmp_4_cfg_a, io_pmp_4_cfg_x, io_pmp_4_cfg_w, io_pmp_4_cfg_r, io_pmp_4_addr, io_pmp_4_mask, io_pmp_5_cfg_l, io_pmp_5_cfg_a, io_pmp_5_cfg_x, io_pmp_5_cfg_w, io_pmp_5_cfg_r, io_pmp_5_addr, io_pmp_5_mask, io_pmp_6_cfg_l, io_pmp_6_cfg_a, io_pmp_6_cfg_x, io_pmp_6_cfg_w, io_pmp_6_cfg_r, io_pmp_6_addr, io_pmp_6_mask, io_pmp_7_cfg_l
, io_pmp_7_cfg_a, io_pmp_7_cfg_x, io_pmp_7_cfg_w, io_pmp_7_cfg_r, io_pmp_7_addr, io_pmp_7_mask, io_inhibit_cycle, io_inst_0, io_trace_0_valid, io_trace_0_iaddr, io_trace_0_insn, io_trace_0_exception, io_customCSRs_0_value);
  wire [31:0] _00000_;
  wire [31:0] _00001_;
  wire [31:0] _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire [1:0] _GEN_170;
  wire [1:0] _GEN_207;
  wire [31:0] _GEN_239;
  wire [5:0] _GEN_34;
  wire [5:0] _GEN_35;
  wire [31:0] _GEN_40;
  wire [31:0] _GEN_41;
  wire _GEN_51;
  wire [31:0] _GEN_586;
  wire [31:0] _GEN_592;
  wire [31:0] _GEN_593;
  wire [31:0] _GEN_594;
  wire [63:0] _GEN_595;
  wire [63:0] _GEN_596;
  wire [63:0] _GEN_597;
  wire [63:0] _GEN_598;
  wire [63:0] _GEN_599;
  wire [63:0] _GEN_600;
  wire [63:0] _GEN_601;
  wire [63:0] _GEN_602;
  wire [63:0] _GEN_603;
  wire [63:0] _GEN_604;
  wire [63:0] _GEN_605;
  wire [63:0] _GEN_606;
  wire [63:0] _GEN_607;
  wire [63:0] _GEN_608;
  wire [63:0] _GEN_609;
  wire [63:0] _GEN_610;
  wire [31:0] _GEN_611;
  wire [1:0] _GEN_73;
  wire _T_14;
  wire _T_15;
  wire [31:0] _T_16;
  wire [31:0] _T_18;
  wire [1:0] _T_20;
  wire [63:0] _T_2000;
  wire [63:0] _T_2003;
  wire [63:0] _T_2005;
  wire [63:0] _T_2008;
  wire [31:0] _T_21;
  wire [31:0] _T_213;
  wire [31:0] _T_22;
  wire [31:0] _T_23;
  wire [31:0] _T_24;
  wire [31:0] _T_27;
  wire [31:0] _T_28;
  wire [7:0] _T_60;
  wire [7:0] _T_62;
  wire [31:0] _T_64;
  wire [7:0] _T_65;
  wire [7:0] _T_67;
  wire [31:0] _T_69;
  wire _any_T_78;
  wire [3:0] _causeIsDebugBreak_T_3;
  wire [3:0] _causeIsDebugBreak_T_4;
  wire [11:0] _debugTVec_T;
  wire [1:0] _decoded_T_10;
  wire [11:0] _decoded_T_14;
  wire [3:0] _decoded_T_16;
  wire [9:0] _decoded_T_18;
  wire [11:0] _decoded_T_2;
  wire [9:0] _decoded_T_20;
  wire [1:0] _decoded_T_22;
  wire [3:0] _decoded_T_4;
  wire [9:0] _decoded_T_6;
  wire [9:0] _decoded_T_8;
  wire [11:0] _decoded_decoded_T;
  wire [10:0] _decoded_decoded_T_10;
  wire [11:0] _decoded_decoded_T_100;
  wire [11:0] _decoded_decoded_T_102;
  wire [11:0] _decoded_decoded_T_104;
  wire [11:0] _decoded_decoded_T_106;
  wire [11:0] _decoded_decoded_T_108;
  wire [11:0] _decoded_decoded_T_110;
  wire [11:0] _decoded_decoded_T_112;
  wire [11:0] _decoded_decoded_T_114;
  wire [11:0] _decoded_decoded_T_116;
  wire [11:0] _decoded_decoded_T_118;
  wire [11:0] _decoded_decoded_T_12;
  wire [11:0] _decoded_decoded_T_120;
  wire [11:0] _decoded_decoded_T_122;
  wire [11:0] _decoded_decoded_T_124;
  wire [11:0] _decoded_decoded_T_126;
  wire [11:0] _decoded_decoded_T_128;
  wire [10:0] _decoded_decoded_T_130;
  wire [5:0] _decoded_decoded_T_132;
  wire [10:0] _decoded_decoded_T_134;
  wire [11:0] _decoded_decoded_T_136;
  wire [11:0] _decoded_decoded_T_138;
  wire [11:0] _decoded_decoded_T_14;
  wire [11:0] _decoded_decoded_T_140;
  wire [11:0] _decoded_decoded_T_142;
  wire [11:0] _decoded_decoded_T_144;
  wire [11:0] _decoded_decoded_T_146;
  wire [11:0] _decoded_decoded_T_148;
  wire [11:0] _decoded_decoded_T_150;
  wire [11:0] _decoded_decoded_T_152;
  wire [11:0] _decoded_decoded_T_154;
  wire [11:0] _decoded_decoded_T_156;
  wire [11:0] _decoded_decoded_T_158;
  wire [11:0] _decoded_decoded_T_16;
  wire [11:0] _decoded_decoded_T_160;
  wire [11:0] _decoded_decoded_T_162;
  wire [11:0] _decoded_decoded_T_164;
  wire [11:0] _decoded_decoded_T_166;
  wire [11:0] _decoded_decoded_T_168;
  wire [11:0] _decoded_decoded_T_170;
  wire [11:0] _decoded_decoded_T_172;
  wire [11:0] _decoded_decoded_T_174;
  wire [11:0] _decoded_decoded_T_176;
  wire [11:0] _decoded_decoded_T_178;
  wire [11:0] _decoded_decoded_T_18;
  wire [11:0] _decoded_decoded_T_180;
  wire [11:0] _decoded_decoded_T_182;
  wire [11:0] _decoded_decoded_T_184;
  wire [11:0] _decoded_decoded_T_186;
  wire [11:0] _decoded_decoded_T_188;
  wire [11:0] _decoded_decoded_T_190;
  wire [11:0] _decoded_decoded_T_192;
  wire [11:0] _decoded_decoded_T_194;
  wire [10:0] _decoded_decoded_T_196;
  wire [11:0] _decoded_decoded_T_198;
  wire [11:0] _decoded_decoded_T_2;
  wire [11:0] _decoded_decoded_T_20;
  wire [11:0] _decoded_decoded_T_200;
  wire [11:0] _decoded_decoded_T_202;
  wire [11:0] _decoded_decoded_T_204;
  wire [11:0] _decoded_decoded_T_206;
  wire [11:0] _decoded_decoded_T_208;
  wire [11:0] _decoded_decoded_T_210;
  wire [11:0] _decoded_decoded_T_212;
  wire [11:0] _decoded_decoded_T_214;
  wire [11:0] _decoded_decoded_T_216;
  wire [11:0] _decoded_decoded_T_218;
  wire [11:0] _decoded_decoded_T_22;
  wire [11:0] _decoded_decoded_T_220;
  wire [11:0] _decoded_decoded_T_222;
  wire [11:0] _decoded_decoded_T_224;
  wire [11:0] _decoded_decoded_T_226;
  wire [11:0] _decoded_decoded_T_228;
  wire [11:0] _decoded_decoded_T_230;
  wire [11:0] _decoded_decoded_T_232;
  wire [11:0] _decoded_decoded_T_234;
  wire [11:0] _decoded_decoded_T_236;
  wire [11:0] _decoded_decoded_T_238;
  wire [11:0] _decoded_decoded_T_24;
  wire [11:0] _decoded_decoded_T_240;
  wire [11:0] _decoded_decoded_T_242;
  wire [11:0] _decoded_decoded_T_244;
  wire [11:0] _decoded_decoded_T_246;
  wire [11:0] _decoded_decoded_T_248;
  wire [11:0] _decoded_decoded_T_250;
  wire [11:0] _decoded_decoded_T_252;
  wire [11:0] _decoded_decoded_T_254;
  wire [11:0] _decoded_decoded_T_256;
  wire [10:0] _decoded_decoded_T_258;
  wire [11:0] _decoded_decoded_T_26;
  wire [11:0] _decoded_decoded_T_260;
  wire _decoded_decoded_T_261;
  wire [11:0] _decoded_decoded_T_262;
  wire _decoded_decoded_T_263;
  wire [9:0] _decoded_decoded_T_264;
  wire [11:0] _decoded_decoded_T_28;
  wire [11:0] _decoded_decoded_T_30;
  wire [11:0] _decoded_decoded_T_32;
  wire [11:0] _decoded_decoded_T_34;
  wire [11:0] _decoded_decoded_T_36;
  wire [11:0] _decoded_decoded_T_38;
  wire [11:0] _decoded_decoded_T_4;
  wire [11:0] _decoded_decoded_T_40;
  wire [11:0] _decoded_decoded_T_42;
  wire [11:0] _decoded_decoded_T_44;
  wire [11:0] _decoded_decoded_T_46;
  wire [11:0] _decoded_decoded_T_48;
  wire [11:0] _decoded_decoded_T_50;
  wire [11:0] _decoded_decoded_T_52;
  wire [11:0] _decoded_decoded_T_54;
  wire [11:0] _decoded_decoded_T_56;
  wire [11:0] _decoded_decoded_T_58;
  wire [11:0] _decoded_decoded_T_6;
  wire [11:0] _decoded_decoded_T_60;
  wire [11:0] _decoded_decoded_T_62;
  wire [11:0] _decoded_decoded_T_64;
  wire [11:0] _decoded_decoded_T_66;
  wire [11:0] _decoded_decoded_T_68;
  wire [11:0] _decoded_decoded_T_70;
  wire [11:0] _decoded_decoded_T_72;
  wire [11:0] _decoded_decoded_T_74;
  wire [9:0] _decoded_decoded_T_76;
  wire [11:0] _decoded_decoded_T_78;
  wire [10:0] _decoded_decoded_T_8;
  wire [11:0] _decoded_decoded_T_80;
  wire [11:0] _decoded_decoded_T_82;
  wire [11:0] _decoded_decoded_T_84;
  wire [11:0] _decoded_decoded_T_86;
  wire [11:0] _decoded_decoded_T_88;
  wire [11:0] _decoded_decoded_T_90;
  wire [11:0] _decoded_decoded_T_92;
  wire [11:0] _decoded_decoded_T_94;
  wire [11:0] _decoded_decoded_T_96;
  wire [11:0] _decoded_decoded_T_98;
  wire _decoded_decoded_orMatrixOutputs_T;
  wire _decoded_decoded_orMatrixOutputs_T_2;
  wire [31:0] _epc_T_1;
  wire [7:0] _io_decode_0_read_illegal_T_12;
  wire _io_decode_0_read_illegal_T_15;
  wire _io_decode_0_read_illegal_T_17;
  wire _io_decode_0_read_illegal_T_21;
  wire [31:0] _io_rw_rdata_T_1;
  wire [31:0] _io_rw_rdata_T_10;
  wire [31:0] _io_rw_rdata_T_107;
  wire [31:0] _io_rw_rdata_T_108;
  wire [31:0] _io_rw_rdata_T_109;
  wire [31:0] _io_rw_rdata_T_110;
  wire [29:0] _io_rw_rdata_T_113;
  wire [29:0] _io_rw_rdata_T_114;
  wire [29:0] _io_rw_rdata_T_115;
  wire [29:0] _io_rw_rdata_T_116;
  wire [29:0] _io_rw_rdata_T_117;
  wire [29:0] _io_rw_rdata_T_118;
  wire [29:0] _io_rw_rdata_T_119;
  wire [29:0] _io_rw_rdata_T_120;
  wire [31:0] _io_rw_rdata_T_129;
  wire _io_rw_rdata_T_13;
  wire [31:0] _io_rw_rdata_T_130;
  wire [31:0] _io_rw_rdata_T_132;
  wire [31:0] _io_rw_rdata_T_14;
  wire [31:0] _io_rw_rdata_T_148;
  wire [31:0] _io_rw_rdata_T_149;
  wire [31:0] _io_rw_rdata_T_15;
  wire [2:0] _io_rw_rdata_T_17;
  wire [63:0] _io_rw_rdata_T_240;
  wire [63:0] _io_rw_rdata_T_241;
  wire [63:0] _io_rw_rdata_T_242;
  wire [63:0] _io_rw_rdata_T_245;
  wire [63:0] _io_rw_rdata_T_246;
  wire [63:0] _io_rw_rdata_T_247;
  wire [63:0] _io_rw_rdata_T_248;
  wire [63:0] _io_rw_rdata_T_249;
  wire [63:0] _io_rw_rdata_T_250;
  wire [63:0] _io_rw_rdata_T_251;
  wire [63:0] _io_rw_rdata_T_252;
  wire [63:0] _io_rw_rdata_T_261;
  wire [63:0] _io_rw_rdata_T_262;
  wire [63:0] _io_rw_rdata_T_264;
  wire [31:0] _io_rw_rdata_T_4;
  wire [31:0] _io_rw_rdata_T_5;
  wire [31:0] _io_rw_rdata_T_6;
  wire [15:0] _io_rw_rdata_T_7;
  wire [31:0] _io_rw_rdata_T_8;
  wire [57:0] _large_r_T_1;
  wire [57:0] _large_r_T_3;
  wire [31:0] _m_interrupts_T_3;
  wire [31:0] _m_interrupts_T_5;
  wire [31:0] _newBPC_T_2;
  wire [31:0] _newBPC_T_3;
  wire [104:0] _new_mstatus_WIRE;
  wire [31:0] _notDebugTVec_T_1;
  wire [30:0] _pmp_mask_T_12;
  wire [30:0] _pmp_mask_T_13;
  wire [32:0] _pmp_mask_T_14;
  wire [30:0] _pmp_mask_T_17;
  wire [30:0] _pmp_mask_T_18;
  wire [32:0] _pmp_mask_T_19;
  wire [30:0] _pmp_mask_T_2;
  wire [30:0] _pmp_mask_T_22;
  wire [30:0] _pmp_mask_T_23;
  wire [32:0] _pmp_mask_T_24;
  wire [30:0] _pmp_mask_T_27;
  wire [30:0] _pmp_mask_T_28;
  wire [32:0] _pmp_mask_T_29;
  wire [30:0] _pmp_mask_T_3;
  wire [30:0] _pmp_mask_T_32;
  wire [30:0] _pmp_mask_T_33;
  wire [32:0] _pmp_mask_T_34;
  wire [30:0] _pmp_mask_T_37;
  wire [30:0] _pmp_mask_T_38;
  wire [32:0] _pmp_mask_T_39;
  wire [32:0] _pmp_mask_T_4;
  wire [30:0] _pmp_mask_T_7;
  wire [30:0] _pmp_mask_T_8;
  wire [32:0] _pmp_mask_T_9;
  wire [15:0] _read_mip_T;
  wire [104:0] _read_mstatus_T;
  wire [6:0] _read_mtvec_T_1;
  wire [31:0] _read_mtvec_T_3;
  wire [31:0] _read_mtvec_T_4;
  wire [31:0] _reg_custom_0_T;
  wire [31:0] _reg_custom_0_T_2;
  wire [31:0] _reg_custom_0_T_3;
  wire [2:0] _reg_dcsr_cause_T_2;
  wire [31:0] _reg_mcause_T;
  wire [31:0] _reg_mcountinhibit_T_1;
  wire [31:0] _reg_mepc_T_1;
  wire [31:0] _reg_mepc_T_2;
  wire [31:0] _reg_mie_T;
  wire [31:0] _reg_misa_T;
  wire _reg_misa_T_1;
  wire [3:0] _reg_misa_T_2;
  wire [31:0] _reg_misa_T_3;
  wire [31:0] _reg_misa_T_4;
  wire [31:0] _reg_misa_T_5;
  wire [31:0] _reg_misa_T_7;
  wire [31:0] _reg_misa_T_8;
  wire [3:0] _which_T_100;
  wire [3:0] _which_T_101;
  wire [3:0] _which_T_102;
  wire [3:0] _which_T_103;
  wire [3:0] _which_T_104;
  wire [3:0] _which_T_105;
  wire [3:0] _which_T_106;
  wire [3:0] _which_T_107;
  wire [3:0] _which_T_108;
  wire [3:0] _which_T_109;
  wire [3:0] _which_T_111;
  wire [3:0] _which_T_112;
  wire [3:0] _which_T_113;
  wire [3:0] _which_T_114;
  wire [3:0] _which_T_115;
  wire [3:0] _which_T_116;
  wire [3:0] _which_T_117;
  wire [3:0] _which_T_118;
  wire [3:0] _which_T_119;
  wire [3:0] _which_T_120;
  wire [3:0] _which_T_121;
  wire [3:0] _which_T_122;
  wire [3:0] _which_T_123;
  wire [3:0] _which_T_124;
  wire [3:0] _which_T_95;
  wire [3:0] _which_T_96;
  wire [3:0] _which_T_97;
  wire [3:0] _which_T_98;
  wire [3:0] _which_T_99;
  wire [12:0] addr;
  wire [11:0] addr_1;
  input clock;
  wire clock;
  wire [14:0] d_interrupts;
  wire [11:0] debugTVec;
  wire decoded_130;
  wire decoded_132;
  wire decoded_andMatrixInput_0_1;
  wire decoded_andMatrixInput_0_10;
  wire decoded_andMatrixInput_0_11;
  wire decoded_andMatrixInput_0_2;
  wire decoded_andMatrixInput_0_4;
  wire decoded_andMatrixInput_0_5;
  wire decoded_andMatrixInput_0_7;
  wire decoded_andMatrixInput_0_8;
  wire decoded_andMatrixInput_7_2;
  wire decoded_andMatrixInput_7_6;
  wire decoded_decoded_andMatrixInput_0_1;
  wire decoded_decoded_andMatrixInput_0_5;
  wire decoded_decoded_andMatrixInput_10_58;
  wire decoded_decoded_andMatrixInput_10_65;
  wire decoded_decoded_andMatrixInput_2_2;
  wire decoded_decoded_andMatrixInput_3_10;
  wire decoded_decoded_andMatrixInput_4_18;
  wire decoded_decoded_andMatrixInput_4_4;
  wire decoded_decoded_andMatrixInput_6_34;
  wire decoded_decoded_andMatrixInput_7_39;
  wire decoded_decoded_andMatrixInput_8;
  wire decoded_decoded_andMatrixInput_9;
  wire [132:0] decoded_decoded_invMatrixOutputs;
  wire [32:0] decoded_decoded_invMatrixOutputs_lo_lo;
  wire [7:0] decoded_decoded_invMatrixOutputs_lo_lo_lo_lo;
  wire [5:0] decoded_decoded_lo;
  wire [4:0] decoded_decoded_lo_129;
  wire [5:0] decoded_decoded_lo_130;
  wire [5:0] decoded_decoded_lo_34;
  wire [5:0] decoded_decoded_lo_39;
  wire [4:0] decoded_decoded_lo_4;
  wire [5:0] decoded_decoded_lo_59;
  wire [4:0] decoded_decoded_lo_65;
  wire [4:0] decoded_decoded_lo_67;
  wire [5:0] decoded_decoded_lo_68;
  wire [4:0] decoded_decoded_lo_98;
  wire [5:0] decoded_decoded_lo_99;
  wire [132:0] decoded_decoded_orMatrixOutputs;
  wire [32:0] decoded_decoded_orMatrixOutputs_lo_lo;
  wire [7:0] decoded_decoded_orMatrixOutputs_lo_lo_lo_lo;
  wire [11:0] decoded_decoded_plaInput;
  wire [31:0] decoded_invInputs;
  wire [8:0] decoded_invMatrixOutputs;
  wire [8:0] decoded_invMatrixOutputs_1;
  wire [8:0] decoded_orMatrixOutputs;
  wire [8:0] decoded_orMatrixOutputs_1;
  wire [31:0] decoded_plaInput;
  wire [31:0] epc;
  wire exception;
  wire f;
  output [31:0] io_bp_0_address;
  wire [31:0] io_bp_0_address;
  output io_bp_0_control_action;
  wire io_bp_0_control_action;
  output io_bp_0_control_r;
  wire io_bp_0_control_r;
  output [1:0] io_bp_0_control_tmatch;
  wire [1:0] io_bp_0_control_tmatch;
  output io_bp_0_control_w;
  wire io_bp_0_control_w;
  output io_bp_0_control_x;
  wire io_bp_0_control_x;
  input [31:0] io_cause;
  wire [31:0] io_cause;
  output io_csr_stall;
  wire io_csr_stall;
  output [31:0] io_customCSRs_0_value;
  wire [31:0] io_customCSRs_0_value;
  output io_decode_0_fp_csr;
  wire io_decode_0_fp_csr;
  output io_decode_0_fp_illegal;
  wire io_decode_0_fp_illegal;
  input [31:0] io_decode_0_inst;
  wire [31:0] io_decode_0_inst;
  output io_decode_0_read_illegal;
  wire io_decode_0_read_illegal;
  wire io_decode_0_read_illegal_andMatrixInput_0;
  wire io_decode_0_read_illegal_andMatrixInput_1;
  wire io_decode_0_read_illegal_andMatrixInput_3;
  wire io_decode_0_read_illegal_andMatrixInput_4;
  wire io_decode_0_read_illegal_andMatrixInput_5;
  wire io_decode_0_read_illegal_andMatrixInput_6;
  output io_decode_0_rocc_illegal;
  wire io_decode_0_rocc_illegal;
  output io_decode_0_system_illegal;
  wire io_decode_0_system_illegal;
  output io_decode_0_write_flush;
  wire io_decode_0_write_flush;
  wire [11:0] io_decode_0_write_flush_addr_m;
  output io_decode_0_write_illegal;
  wire io_decode_0_write_illegal;
  output io_eret;
  wire io_eret;
  output [31:0] io_evec;
  wire [31:0] io_evec;
  input io_exception;
  wire io_exception;
  input io_gva;
  wire io_gva;
  input io_hartid;
  wire io_hartid;
  output io_inhibit_cycle;
  wire io_inhibit_cycle;
  input [31:0] io_inst_0;
  wire [31:0] io_inst_0;
  output io_interrupt;
  wire io_interrupt;
  output [31:0] io_interrupt_cause;
  wire [31:0] io_interrupt_cause;
  input io_interrupts_debug;
  wire io_interrupts_debug;
  input io_interrupts_meip;
  wire io_interrupts_meip;
  input io_interrupts_msip;
  wire io_interrupts_msip;
  input io_interrupts_mtip;
  wire io_interrupts_mtip;
  input [31:0] io_pc;
  wire [31:0] io_pc;
  output [29:0] io_pmp_0_addr;
  wire [29:0] io_pmp_0_addr;
  output [1:0] io_pmp_0_cfg_a;
  wire [1:0] io_pmp_0_cfg_a;
  output io_pmp_0_cfg_l;
  wire io_pmp_0_cfg_l;
  output io_pmp_0_cfg_r;
  wire io_pmp_0_cfg_r;
  output io_pmp_0_cfg_w;
  wire io_pmp_0_cfg_w;
  output io_pmp_0_cfg_x;
  wire io_pmp_0_cfg_x;
  output [31:0] io_pmp_0_mask;
  wire [31:0] io_pmp_0_mask;
  output [29:0] io_pmp_1_addr;
  wire [29:0] io_pmp_1_addr;
  output [1:0] io_pmp_1_cfg_a;
  wire [1:0] io_pmp_1_cfg_a;
  output io_pmp_1_cfg_l;
  wire io_pmp_1_cfg_l;
  output io_pmp_1_cfg_r;
  wire io_pmp_1_cfg_r;
  output io_pmp_1_cfg_w;
  wire io_pmp_1_cfg_w;
  output io_pmp_1_cfg_x;
  wire io_pmp_1_cfg_x;
  output [31:0] io_pmp_1_mask;
  wire [31:0] io_pmp_1_mask;
  output [29:0] io_pmp_2_addr;
  wire [29:0] io_pmp_2_addr;
  output [1:0] io_pmp_2_cfg_a;
  wire [1:0] io_pmp_2_cfg_a;
  output io_pmp_2_cfg_l;
  wire io_pmp_2_cfg_l;
  output io_pmp_2_cfg_r;
  wire io_pmp_2_cfg_r;
  output io_pmp_2_cfg_w;
  wire io_pmp_2_cfg_w;
  output io_pmp_2_cfg_x;
  wire io_pmp_2_cfg_x;
  output [31:0] io_pmp_2_mask;
  wire [31:0] io_pmp_2_mask;
  output [29:0] io_pmp_3_addr;
  wire [29:0] io_pmp_3_addr;
  output [1:0] io_pmp_3_cfg_a;
  wire [1:0] io_pmp_3_cfg_a;
  output io_pmp_3_cfg_l;
  wire io_pmp_3_cfg_l;
  output io_pmp_3_cfg_r;
  wire io_pmp_3_cfg_r;
  output io_pmp_3_cfg_w;
  wire io_pmp_3_cfg_w;
  output io_pmp_3_cfg_x;
  wire io_pmp_3_cfg_x;
  output [31:0] io_pmp_3_mask;
  wire [31:0] io_pmp_3_mask;
  output [29:0] io_pmp_4_addr;
  wire [29:0] io_pmp_4_addr;
  output [1:0] io_pmp_4_cfg_a;
  wire [1:0] io_pmp_4_cfg_a;
  output io_pmp_4_cfg_l;
  wire io_pmp_4_cfg_l;
  output io_pmp_4_cfg_r;
  wire io_pmp_4_cfg_r;
  output io_pmp_4_cfg_w;
  wire io_pmp_4_cfg_w;
  output io_pmp_4_cfg_x;
  wire io_pmp_4_cfg_x;
  output [31:0] io_pmp_4_mask;
  wire [31:0] io_pmp_4_mask;
  output [29:0] io_pmp_5_addr;
  wire [29:0] io_pmp_5_addr;
  output [1:0] io_pmp_5_cfg_a;
  wire [1:0] io_pmp_5_cfg_a;
  output io_pmp_5_cfg_l;
  wire io_pmp_5_cfg_l;
  output io_pmp_5_cfg_r;
  wire io_pmp_5_cfg_r;
  output io_pmp_5_cfg_w;
  wire io_pmp_5_cfg_w;
  output io_pmp_5_cfg_x;
  wire io_pmp_5_cfg_x;
  output [31:0] io_pmp_5_mask;
  wire [31:0] io_pmp_5_mask;
  output [29:0] io_pmp_6_addr;
  wire [29:0] io_pmp_6_addr;
  output [1:0] io_pmp_6_cfg_a;
  wire [1:0] io_pmp_6_cfg_a;
  output io_pmp_6_cfg_l;
  wire io_pmp_6_cfg_l;
  output io_pmp_6_cfg_r;
  wire io_pmp_6_cfg_r;
  output io_pmp_6_cfg_w;
  wire io_pmp_6_cfg_w;
  output io_pmp_6_cfg_x;
  wire io_pmp_6_cfg_x;
  output [31:0] io_pmp_6_mask;
  wire [31:0] io_pmp_6_mask;
  output [29:0] io_pmp_7_addr;
  wire [29:0] io_pmp_7_addr;
  output [1:0] io_pmp_7_cfg_a;
  wire [1:0] io_pmp_7_cfg_a;
  output io_pmp_7_cfg_l;
  wire io_pmp_7_cfg_l;
  output io_pmp_7_cfg_r;
  wire io_pmp_7_cfg_r;
  output io_pmp_7_cfg_w;
  wire io_pmp_7_cfg_w;
  output io_pmp_7_cfg_x;
  wire io_pmp_7_cfg_x;
  output [31:0] io_pmp_7_mask;
  wire [31:0] io_pmp_7_mask;
  input io_retire;
  wire io_retire;
  input [11:0] io_rw_addr;
  wire [11:0] io_rw_addr;
  input [2:0] io_rw_cmd;
  wire [2:0] io_rw_cmd;
  output [31:0] io_rw_rdata;
  wire [31:0] io_rw_rdata;
  input [31:0] io_rw_wdata;
  wire [31:0] io_rw_wdata;
  output io_singleStep;
  wire io_singleStep;
  output io_status_cease;
  wire io_status_cease;
  wire io_status_cease_r;
  output io_status_debug;
  wire io_status_debug;
  output [1:0] io_status_dprv;
  wire [1:0] io_status_dprv;
  output io_status_dv;
  wire io_status_dv;
  output [1:0] io_status_fs;
  wire [1:0] io_status_fs;
  output io_status_gva;
  wire io_status_gva;
  output io_status_hie;
  wire io_status_hie;
  output [31:0] io_status_isa;
  wire [31:0] io_status_isa;
  output io_status_mbe;
  wire io_status_mbe;
  output io_status_mie;
  wire io_status_mie;
  output io_status_mpie;
  wire io_status_mpie;
  output [1:0] io_status_mpp;
  wire [1:0] io_status_mpp;
  output io_status_mprv;
  wire io_status_mprv;
  output io_status_mpv;
  wire io_status_mpv;
  output io_status_mxr;
  wire io_status_mxr;
  output [1:0] io_status_prv;
  wire [1:0] io_status_prv;
  output io_status_sbe;
  wire io_status_sbe;
  output io_status_sd;
  wire io_status_sd;
  output io_status_sd_rv32;
  wire io_status_sd_rv32;
  output io_status_sie;
  wire io_status_sie;
  output io_status_spie;
  wire io_status_spie;
  output io_status_spp;
  wire io_status_spp;
  output io_status_sum;
  wire io_status_sum;
  output [1:0] io_status_sxl;
  wire [1:0] io_status_sxl;
  output io_status_tsr;
  wire io_status_tsr;
  output io_status_tvm;
  wire io_status_tvm;
  output io_status_tw;
  wire io_status_tw;
  output io_status_ube;
  wire io_status_ube;
  output io_status_uie;
  wire io_status_uie;
  output io_status_upie;
  wire io_status_upie;
  output [1:0] io_status_uxl;
  wire [1:0] io_status_uxl;
  output io_status_v;
  wire io_status_v;
  output [1:0] io_status_vs;
  wire [1:0] io_status_vs;
  output io_status_wfi;
  wire io_status_wfi;
  output [1:0] io_status_xs;
  wire [1:0] io_status_xs;
  output [7:0] io_status_zero1;
  wire [7:0] io_status_zero1;
  output [22:0] io_status_zero2;
  wire [22:0] io_status_zero2;
  output [31:0] io_time;
  wire [31:0] io_time;
  output io_trace_0_exception;
  wire io_trace_0_exception;
  output [31:0] io_trace_0_iaddr;
  wire [31:0] io_trace_0_iaddr;
  output [31:0] io_trace_0_insn;
  wire [31:0] io_trace_0_insn;
  output io_trace_0_valid;
  wire io_trace_0_valid;
  input [31:0] io_tval;
  wire [31:0] io_tval;
  input io_ungated_clock;
  wire io_ungated_clock;
  wire [57:0] large_;
  wire [57:0] large_1;
  wire [15:0] lo_11;
  wire [15:0] lo_16;
  wire [6:0] lo_4;
  wire [31:0] m_interrupts;
  wire [1:0] newCfg_1_a;
  wire newCfg_1_l;
  wire newCfg_1_r;
  wire newCfg_1_w;
  wire newCfg_1_x;
  wire [1:0] newCfg_2_a;
  wire newCfg_2_l;
  wire newCfg_2_r;
  wire newCfg_2_w;
  wire newCfg_2_x;
  wire [1:0] newCfg_3_a;
  wire newCfg_3_l;
  wire newCfg_3_r;
  wire newCfg_3_w;
  wire newCfg_3_x;
  wire [1:0] newCfg_a;
  wire newCfg_l;
  wire newCfg_r;
  wire newCfg_w;
  wire newCfg_x;
  wire new_dcsr_ebreakm;
  wire new_mstatus_mie;
  wire new_mstatus_mpie;
  wire [31:0] notDebugTVec;
  wire [6:0] notDebugTVec_interruptOffset;
  wire [31:0] notDebugTVec_interruptVec;
  wire [31:0] pending_interrupts;
  wire [30:0] pmp_mask_base;
  wire [30:0] pmp_mask_base_1;
  wire [30:0] pmp_mask_base_2;
  wire [30:0] pmp_mask_base_3;
  wire [30:0] pmp_mask_base_4;
  wire [30:0] pmp_mask_base_5;
  wire [30:0] pmp_mask_base_6;
  wire [30:0] pmp_mask_base_7;
  wire [15:0] read_mip;
  wire [31:0] read_mstatus;
  wire [82:0] read_mstatus_hi;
  wire [64:0] read_mstatus_hi_hi;
  wire [21:0] read_mstatus_lo;
  wire [8:0] read_mstatus_lo_lo;
  wire [31:0] read_mtvec;
  wire [31:0] reg_bp_0_address;
  wire reg_bp_0_control_action;
  wire reg_bp_0_control_dmode;
  wire reg_bp_0_control_r;
  wire [1:0] reg_bp_0_control_tmatch;
  wire reg_bp_0_control_w;
  wire reg_bp_0_control_x;
  wire [31:0] reg_custom_0;
  wire [2:0] reg_dcsr_cause;
  wire reg_dcsr_ebreakm;
  wire reg_dcsr_step;
  wire reg_debug;
  wire [31:0] reg_dpc;
  wire [31:0] reg_dscratch0;
  wire [31:0] reg_mcause;
  wire [2:0] reg_mcountinhibit;
  wire [31:0] reg_mepc;
  wire [31:0] reg_mie;
  wire [31:0] reg_misa;
  wire [31:0] reg_mscratch;
  wire reg_mstatus_gva;
  wire reg_mstatus_mie;
  wire reg_mstatus_mpie;
  wire reg_mstatus_spp;
  wire [31:0] reg_mtval;
  wire [31:0] reg_mtvec;
  wire [29:0] reg_pmp_0_addr;
  wire [1:0] reg_pmp_0_cfg_a;
  wire reg_pmp_0_cfg_l;
  wire reg_pmp_0_cfg_r;
  wire reg_pmp_0_cfg_w;
  wire reg_pmp_0_cfg_x;
  wire [29:0] reg_pmp_1_addr;
  wire [1:0] reg_pmp_1_cfg_a;
  wire reg_pmp_1_cfg_l;
  wire reg_pmp_1_cfg_r;
  wire reg_pmp_1_cfg_w;
  wire reg_pmp_1_cfg_x;
  wire [29:0] reg_pmp_2_addr;
  wire [1:0] reg_pmp_2_cfg_a;
  wire reg_pmp_2_cfg_l;
  wire reg_pmp_2_cfg_r;
  wire reg_pmp_2_cfg_w;
  wire reg_pmp_2_cfg_x;
  wire [29:0] reg_pmp_3_addr;
  wire [1:0] reg_pmp_3_cfg_a;
  wire reg_pmp_3_cfg_l;
  wire reg_pmp_3_cfg_r;
  wire reg_pmp_3_cfg_w;
  wire reg_pmp_3_cfg_x;
  wire [29:0] reg_pmp_4_addr;
  wire [1:0] reg_pmp_4_cfg_a;
  wire reg_pmp_4_cfg_l;
  wire reg_pmp_4_cfg_r;
  wire reg_pmp_4_cfg_w;
  wire reg_pmp_4_cfg_x;
  wire [29:0] reg_pmp_5_addr;
  wire [1:0] reg_pmp_5_cfg_a;
  wire reg_pmp_5_cfg_l;
  wire reg_pmp_5_cfg_r;
  wire reg_pmp_5_cfg_w;
  wire reg_pmp_5_cfg_x;
  wire [29:0] reg_pmp_6_addr;
  wire [1:0] reg_pmp_6_cfg_a;
  wire reg_pmp_6_cfg_l;
  wire reg_pmp_6_cfg_r;
  wire reg_pmp_6_cfg_w;
  wire reg_pmp_6_cfg_x;
  wire [29:0] reg_pmp_7_addr;
  wire [1:0] reg_pmp_7_cfg_a;
  wire reg_pmp_7_cfg_l;
  wire reg_pmp_7_cfg_r;
  wire reg_pmp_7_cfg_w;
  wire reg_pmp_7_cfg_x;
  wire reg_singleStepped;
  wire reg_wfi;
  input reset;
  wire reset;
  wire [5:0] small_;
  wire [5:0] small_1;
  wire [31:0] tvec;
  wire [63:0] value;
  wire [63:0] value_1;
  wire [31:0] wdata;
  wire [3:0] whichInterrupt;
  wire x79;
  wire x86;
  AND2_X1 _07165_ (
    .A1(_02165_),
    .A2(_02233_),
    .ZN(_02234_)
  );
  INV_X1 _07166_ (
    .A(_02234_),
    .ZN(_02235_)
  );
  MUX2_X1 _07167_ (
    .A(reg_pmp_5_addr[10]),
    .B(_02235_),
    .S(_01525_),
    .Z(_00037_)
  );
  AND2_X1 _07168_ (
    .A1(io_rw_wdata[11]),
    .A2(_00903_),
    .ZN(_02236_)
  );
  INV_X1 _07169_ (
    .A(_02236_),
    .ZN(_02237_)
  );
  AND2_X1 _07170_ (
    .A1(reg_mtval[11]),
    .A2(_00926_),
    .ZN(_02238_)
  );
  INV_X1 _07171_ (
    .A(_02238_),
    .ZN(_02239_)
  );
  AND2_X1 _07172_ (
    .A1(reg_mscratch[11]),
    .A2(_00929_),
    .ZN(_02240_)
  );
  INV_X1 _07173_ (
    .A(_02240_),
    .ZN(_02241_)
  );
  AND2_X1 _07174_ (
    .A1(_02239_),
    .A2(_02241_),
    .ZN(_02242_)
  );
  AND2_X1 _07175_ (
    .A1(reg_mtvec[11]),
    .A2(_00940_),
    .ZN(_02243_)
  );
  INV_X1 _07176_ (
    .A(_02243_),
    .ZN(_02244_)
  );
  AND2_X1 _07177_ (
    .A1(reg_mepc[11]),
    .A2(_00943_),
    .ZN(_02245_)
  );
  INV_X1 _07178_ (
    .A(_02245_),
    .ZN(_02246_)
  );
  AND2_X1 _07179_ (
    .A1(_02244_),
    .A2(_02246_),
    .ZN(_02247_)
  );
  AND2_X1 _07180_ (
    .A1(_02242_),
    .A2(_02247_),
    .ZN(_02248_)
  );
  AND2_X1 _07181_ (
    .A1(reg_pmp_5_addr[11]),
    .A2(_00948_),
    .ZN(_02249_)
  );
  INV_X1 _07182_ (
    .A(_02249_),
    .ZN(_02250_)
  );
  AND2_X1 _07183_ (
    .A1(reg_pmp_4_addr[11]),
    .A2(_00968_),
    .ZN(_02251_)
  );
  INV_X1 _07184_ (
    .A(_02251_),
    .ZN(_02252_)
  );
  AND2_X1 _07185_ (
    .A1(_02250_),
    .A2(_02252_),
    .ZN(_02253_)
  );
  AND2_X1 _07186_ (
    .A1(reg_mcause[11]),
    .A2(_01001_),
    .ZN(_02254_)
  );
  INV_X1 _07187_ (
    .A(_02254_),
    .ZN(_02255_)
  );
  AND2_X1 _07188_ (
    .A1(reg_dscratch0[11]),
    .A2(_00958_),
    .ZN(_02256_)
  );
  INV_X1 _07189_ (
    .A(_02256_),
    .ZN(_02257_)
  );
  AND2_X1 _07190_ (
    .A1(_02255_),
    .A2(_02257_),
    .ZN(_02258_)
  );
  AND2_X1 _07191_ (
    .A1(_02253_),
    .A2(_02258_),
    .ZN(_02259_)
  );
  AND2_X1 _07192_ (
    .A1(_02248_),
    .A2(_02259_),
    .ZN(_02260_)
  );
  AND2_X1 _07193_ (
    .A1(reg_bp_0_address[11]),
    .A2(_00962_),
    .ZN(_02261_)
  );
  INV_X1 _07194_ (
    .A(_02261_),
    .ZN(_02262_)
  );
  AND2_X1 _07195_ (
    .A1(reg_pmp_1_cfg_a[0]),
    .A2(_00916_),
    .ZN(_02263_)
  );
  INV_X1 _07196_ (
    .A(_02263_),
    .ZN(_02264_)
  );
  AND2_X1 _07197_ (
    .A1(reg_pmp_5_cfg_a[0]),
    .A2(_00894_),
    .ZN(_02265_)
  );
  INV_X1 _07198_ (
    .A(_02265_),
    .ZN(_02266_)
  );
  AND2_X1 _07199_ (
    .A1(_02264_),
    .A2(_02266_),
    .ZN(_02267_)
  );
  AND2_X1 _07200_ (
    .A1(_02262_),
    .A2(_02267_),
    .ZN(_02268_)
  );
  AND2_X1 _07201_ (
    .A1(io_interrupts_meip),
    .A2(_01803_),
    .ZN(_02269_)
  );
  INV_X1 _07202_ (
    .A(_02269_),
    .ZN(_02270_)
  );
  AND2_X1 _07203_ (
    .A1(reg_pmp_2_addr[11]),
    .A2(_00953_),
    .ZN(_02271_)
  );
  INV_X1 _07204_ (
    .A(_02271_),
    .ZN(_02272_)
  );
  AND2_X1 _07205_ (
    .A1(_02270_),
    .A2(_02272_),
    .ZN(_02273_)
  );
  AND2_X1 _07206_ (
    .A1(reg_dpc[11]),
    .A2(_00912_),
    .ZN(_02274_)
  );
  INV_X1 _07207_ (
    .A(_02274_),
    .ZN(_02275_)
  );
  AND2_X1 _07208_ (
    .A1(reg_pmp_1_addr[11]),
    .A2(_01008_),
    .ZN(_02276_)
  );
  INV_X1 _07209_ (
    .A(_02276_),
    .ZN(_02277_)
  );
  AND2_X1 _07210_ (
    .A1(_02275_),
    .A2(_02277_),
    .ZN(_02278_)
  );
  AND2_X1 _07211_ (
    .A1(_02273_),
    .A2(_02278_),
    .ZN(_02279_)
  );
  AND2_X1 _07212_ (
    .A1(_02268_),
    .A2(_02279_),
    .ZN(_02280_)
  );
  AND2_X1 _07213_ (
    .A1(_02260_),
    .A2(_02280_),
    .ZN(_02281_)
  );
  AND2_X1 _07214_ (
    .A1(reg_pmp_7_addr[11]),
    .A2(_01016_),
    .ZN(_02282_)
  );
  INV_X1 _07215_ (
    .A(_02282_),
    .ZN(_02283_)
  );
  AND2_X1 _07216_ (
    .A1(large_1[37]),
    .A2(_01019_),
    .ZN(_02284_)
  );
  INV_X1 _07217_ (
    .A(_02284_),
    .ZN(_02285_)
  );
  AND2_X1 _07218_ (
    .A1(_02283_),
    .A2(_02285_),
    .ZN(_02286_)
  );
  AND2_X1 _07219_ (
    .A1(large_[37]),
    .A2(_00991_),
    .ZN(_02287_)
  );
  INV_X1 _07220_ (
    .A(_02287_),
    .ZN(_02288_)
  );
  AND2_X1 _07221_ (
    .A1(large_1[5]),
    .A2(_00995_),
    .ZN(_02289_)
  );
  INV_X1 _07222_ (
    .A(_02289_),
    .ZN(_02290_)
  );
  AND2_X1 _07223_ (
    .A1(_02288_),
    .A2(_02290_),
    .ZN(_02291_)
  );
  AND2_X1 _07224_ (
    .A1(_02286_),
    .A2(_02291_),
    .ZN(_02292_)
  );
  AND2_X1 _07225_ (
    .A1(reg_pmp_0_addr[11]),
    .A2(_01004_),
    .ZN(_02293_)
  );
  INV_X1 _07226_ (
    .A(_02293_),
    .ZN(_02294_)
  );
  AND2_X1 _07227_ (
    .A1(_01814_),
    .A2(_02294_),
    .ZN(_02295_)
  );
  AND2_X1 _07228_ (
    .A1(reg_mie[11]),
    .A2(_01782_),
    .ZN(_02296_)
  );
  INV_X1 _07229_ (
    .A(_02296_),
    .ZN(_02297_)
  );
  AND2_X1 _07230_ (
    .A1(reg_pmp_3_addr[11]),
    .A2(_01011_),
    .ZN(_02298_)
  );
  INV_X1 _07231_ (
    .A(_02298_),
    .ZN(_02299_)
  );
  AND2_X1 _07232_ (
    .A1(_02297_),
    .A2(_02299_),
    .ZN(_02300_)
  );
  AND2_X1 _07233_ (
    .A1(_02295_),
    .A2(_02300_),
    .ZN(_02301_)
  );
  AND2_X1 _07234_ (
    .A1(reg_pmp_6_addr[11]),
    .A2(_00978_),
    .ZN(_02302_)
  );
  INV_X1 _07235_ (
    .A(_02302_),
    .ZN(_02303_)
  );
  AND2_X1 _07236_ (
    .A1(large_[5]),
    .A2(_00985_),
    .ZN(_02304_)
  );
  INV_X1 _07237_ (
    .A(_02304_),
    .ZN(_02305_)
  );
  AND2_X1 _07238_ (
    .A1(_02303_),
    .A2(_02305_),
    .ZN(_02306_)
  );
  AND2_X1 _07239_ (
    .A1(_02301_),
    .A2(_02306_),
    .ZN(_02307_)
  );
  AND2_X1 _07240_ (
    .A1(_02292_),
    .A2(_02307_),
    .ZN(_02308_)
  );
  AND2_X1 _07241_ (
    .A1(_02281_),
    .A2(_02308_),
    .ZN(_02309_)
  );
  INV_X1 _07242_ (
    .A(_02309_),
    .ZN(io_rw_rdata[11])
  );
  AND2_X1 _07243_ (
    .A1(io_rw_cmd[1]),
    .A2(_00847_),
    .ZN(_02310_)
  );
  AND2_X1 _07244_ (
    .A1(io_rw_rdata[11]),
    .A2(_02310_),
    .ZN(_02311_)
  );
  INV_X1 _07245_ (
    .A(_02311_),
    .ZN(_02312_)
  );
  AND2_X1 _07246_ (
    .A1(_02237_),
    .A2(_02312_),
    .ZN(_02313_)
  );
  INV_X1 _07247_ (
    .A(_02313_),
    .ZN(_02314_)
  );
  MUX2_X1 _07248_ (
    .A(reg_pmp_5_addr[11]),
    .B(_02314_),
    .S(_01525_),
    .Z(_00038_)
  );
  AND2_X1 _07249_ (
    .A1(reg_pmp_1_addr[12]),
    .A2(_01008_),
    .ZN(_02315_)
  );
  INV_X1 _07250_ (
    .A(_02315_),
    .ZN(_02316_)
  );
  AND2_X1 _07251_ (
    .A1(reg_mepc[12]),
    .A2(_00943_),
    .ZN(_02317_)
  );
  INV_X1 _07252_ (
    .A(_02317_),
    .ZN(_02318_)
  );
  AND2_X1 _07253_ (
    .A1(_02316_),
    .A2(_02318_),
    .ZN(_02319_)
  );
  AND2_X1 _07254_ (
    .A1(reg_dscratch0[12]),
    .A2(_00958_),
    .ZN(_02320_)
  );
  INV_X1 _07255_ (
    .A(_02320_),
    .ZN(_02321_)
  );
  AND2_X1 _07256_ (
    .A1(reg_dpc[12]),
    .A2(_00912_),
    .ZN(_02322_)
  );
  INV_X1 _07257_ (
    .A(_02322_),
    .ZN(_02323_)
  );
  AND2_X1 _07258_ (
    .A1(_02321_),
    .A2(_02323_),
    .ZN(_02324_)
  );
  AND2_X1 _07259_ (
    .A1(_02319_),
    .A2(_02324_),
    .ZN(_02325_)
  );
  AND2_X1 _07260_ (
    .A1(reg_pmp_2_addr[12]),
    .A2(_00953_),
    .ZN(_02326_)
  );
  INV_X1 _07261_ (
    .A(_02326_),
    .ZN(_02327_)
  );
  AND2_X1 _07262_ (
    .A1(reg_pmp_0_addr[12]),
    .A2(_01004_),
    .ZN(_02328_)
  );
  INV_X1 _07263_ (
    .A(_02328_),
    .ZN(_02329_)
  );
  AND2_X1 _07264_ (
    .A1(_02327_),
    .A2(_02329_),
    .ZN(_02330_)
  );
  AND2_X1 _07265_ (
    .A1(reg_pmp_5_addr[12]),
    .A2(_00948_),
    .ZN(_02331_)
  );
  INV_X1 _07266_ (
    .A(_02331_),
    .ZN(_02332_)
  );
  AND2_X1 _07267_ (
    .A1(reg_pmp_4_addr[12]),
    .A2(_00968_),
    .ZN(_02333_)
  );
  INV_X1 _07268_ (
    .A(_02333_),
    .ZN(_02334_)
  );
  AND2_X1 _07269_ (
    .A1(_02332_),
    .A2(_02334_),
    .ZN(_02335_)
  );
  AND2_X1 _07270_ (
    .A1(_02330_),
    .A2(_02335_),
    .ZN(_02336_)
  );
  AND2_X1 _07271_ (
    .A1(_02325_),
    .A2(_02336_),
    .ZN(_02337_)
  );
  AND2_X1 _07272_ (
    .A1(reg_mtval[12]),
    .A2(_00926_),
    .ZN(_02338_)
  );
  INV_X1 _07273_ (
    .A(_02338_),
    .ZN(_02339_)
  );
  AND2_X1 _07274_ (
    .A1(reg_mcause[12]),
    .A2(_01001_),
    .ZN(_02340_)
  );
  INV_X1 _07275_ (
    .A(_02340_),
    .ZN(_02341_)
  );
  AND2_X1 _07276_ (
    .A1(_02339_),
    .A2(_02341_),
    .ZN(_02342_)
  );
  AND2_X1 _07277_ (
    .A1(reg_mscratch[12]),
    .A2(_00929_),
    .ZN(_02343_)
  );
  INV_X1 _07278_ (
    .A(_02343_),
    .ZN(_02344_)
  );
  AND2_X1 _07279_ (
    .A1(reg_mtvec[12]),
    .A2(_00940_),
    .ZN(_02345_)
  );
  INV_X1 _07280_ (
    .A(_02345_),
    .ZN(_02346_)
  );
  AND2_X1 _07281_ (
    .A1(_02344_),
    .A2(_02346_),
    .ZN(_02347_)
  );
  AND2_X1 _07282_ (
    .A1(_02342_),
    .A2(_02347_),
    .ZN(_02348_)
  );
  AND2_X1 _07283_ (
    .A1(reg_bp_0_control_action),
    .A2(_01341_),
    .ZN(_02349_)
  );
  INV_X1 _07284_ (
    .A(_02349_),
    .ZN(_02350_)
  );
  AND2_X1 _07285_ (
    .A1(reg_pmp_3_addr[12]),
    .A2(_01011_),
    .ZN(_02351_)
  );
  INV_X1 _07286_ (
    .A(_02351_),
    .ZN(_02352_)
  );
  AND2_X1 _07287_ (
    .A1(_02350_),
    .A2(_02352_),
    .ZN(_02353_)
  );
  AND2_X1 _07288_ (
    .A1(reg_misa[12]),
    .A2(_01339_),
    .ZN(_02354_)
  );
  INV_X1 _07289_ (
    .A(_02354_),
    .ZN(_02355_)
  );
  AND2_X1 _07290_ (
    .A1(reg_pmp_5_cfg_a[1]),
    .A2(_00894_),
    .ZN(_02356_)
  );
  INV_X1 _07291_ (
    .A(_02356_),
    .ZN(_02357_)
  );
  AND2_X1 _07292_ (
    .A1(_02355_),
    .A2(_02357_),
    .ZN(_02358_)
  );
  AND2_X1 _07293_ (
    .A1(_02353_),
    .A2(_02358_),
    .ZN(_02359_)
  );
  AND2_X1 _07294_ (
    .A1(_02348_),
    .A2(_02359_),
    .ZN(_02360_)
  );
  AND2_X1 _07295_ (
    .A1(_02337_),
    .A2(_02360_),
    .ZN(_02361_)
  );
  AND2_X1 _07296_ (
    .A1(reg_pmp_7_addr[12]),
    .A2(_01016_),
    .ZN(_02362_)
  );
  INV_X1 _07297_ (
    .A(_02362_),
    .ZN(_02363_)
  );
  AND2_X1 _07298_ (
    .A1(large_[6]),
    .A2(_00985_),
    .ZN(_02364_)
  );
  INV_X1 _07299_ (
    .A(_02364_),
    .ZN(_02365_)
  );
  AND2_X1 _07300_ (
    .A1(_02363_),
    .A2(_02365_),
    .ZN(_02366_)
  );
  AND2_X1 _07301_ (
    .A1(large_1[38]),
    .A2(_01019_),
    .ZN(_02367_)
  );
  INV_X1 _07302_ (
    .A(_02367_),
    .ZN(_02368_)
  );
  AND2_X1 _07303_ (
    .A1(reg_pmp_6_addr[12]),
    .A2(_00978_),
    .ZN(_02369_)
  );
  INV_X1 _07304_ (
    .A(_02369_),
    .ZN(_02370_)
  );
  AND2_X1 _07305_ (
    .A1(_02368_),
    .A2(_02370_),
    .ZN(_02371_)
  );
  AND2_X1 _07306_ (
    .A1(_02366_),
    .A2(_02371_),
    .ZN(_02372_)
  );
  AND2_X1 _07307_ (
    .A1(_01132_),
    .A2(_01814_),
    .ZN(_02373_)
  );
  AND2_X1 _07308_ (
    .A1(reg_bp_0_address[12]),
    .A2(_00962_),
    .ZN(_02374_)
  );
  INV_X1 _07309_ (
    .A(_02374_),
    .ZN(_02375_)
  );
  AND2_X1 _07310_ (
    .A1(reg_pmp_1_cfg_a[1]),
    .A2(_00916_),
    .ZN(_02376_)
  );
  INV_X1 _07311_ (
    .A(_02376_),
    .ZN(_02377_)
  );
  AND2_X1 _07312_ (
    .A1(_02375_),
    .A2(_02377_),
    .ZN(_02378_)
  );
  AND2_X1 _07313_ (
    .A1(_02373_),
    .A2(_02378_),
    .ZN(_02379_)
  );
  AND2_X1 _07314_ (
    .A1(large_[38]),
    .A2(_00991_),
    .ZN(_02380_)
  );
  INV_X1 _07315_ (
    .A(_02380_),
    .ZN(_02381_)
  );
  AND2_X1 _07316_ (
    .A1(large_1[6]),
    .A2(_00995_),
    .ZN(_02382_)
  );
  INV_X1 _07317_ (
    .A(_02382_),
    .ZN(_02383_)
  );
  AND2_X1 _07318_ (
    .A1(_02381_),
    .A2(_02383_),
    .ZN(_02384_)
  );
  AND2_X1 _07319_ (
    .A1(_02379_),
    .A2(_02384_),
    .ZN(_02385_)
  );
  AND2_X1 _07320_ (
    .A1(_02372_),
    .A2(_02385_),
    .ZN(_02386_)
  );
  AND2_X1 _07321_ (
    .A1(_02361_),
    .A2(_02386_),
    .ZN(_02387_)
  );
  INV_X1 _07322_ (
    .A(_02387_),
    .ZN(io_rw_rdata[12])
  );
  AND2_X1 _07323_ (
    .A1(io_rw_cmd[1]),
    .A2(io_rw_rdata[12]),
    .ZN(_02388_)
  );
  MUX2_X1 _07324_ (
    .A(_02388_),
    .B(_00903_),
    .S(io_rw_wdata[12]),
    .Z(_02389_)
  );
  INV_X1 _07325_ (
    .A(_02389_),
    .ZN(_02390_)
  );
  MUX2_X1 _07326_ (
    .A(reg_pmp_5_addr[12]),
    .B(_02389_),
    .S(_01525_),
    .Z(_00039_)
  );
  AND2_X1 _07327_ (
    .A1(io_rw_wdata[13]),
    .A2(_00903_),
    .ZN(_02391_)
  );
  INV_X1 _07328_ (
    .A(_02391_),
    .ZN(_02392_)
  );
  AND2_X1 _07329_ (
    .A1(reg_pmp_3_addr[13]),
    .A2(_01011_),
    .ZN(_02393_)
  );
  INV_X1 _07330_ (
    .A(_02393_),
    .ZN(_02394_)
  );
  AND2_X1 _07331_ (
    .A1(reg_mepc[13]),
    .A2(_00943_),
    .ZN(_02395_)
  );
  INV_X1 _07332_ (
    .A(_02395_),
    .ZN(_02396_)
  );
  AND2_X1 _07333_ (
    .A1(_02394_),
    .A2(_02396_),
    .ZN(_02397_)
  );
  AND2_X1 _07334_ (
    .A1(reg_mtval[13]),
    .A2(_00926_),
    .ZN(_02398_)
  );
  INV_X1 _07335_ (
    .A(_02398_),
    .ZN(_02399_)
  );
  AND2_X1 _07336_ (
    .A1(reg_pmp_4_addr[13]),
    .A2(_00968_),
    .ZN(_02400_)
  );
  INV_X1 _07337_ (
    .A(_02400_),
    .ZN(_02401_)
  );
  AND2_X1 _07338_ (
    .A1(_02399_),
    .A2(_02401_),
    .ZN(_02402_)
  );
  AND2_X1 _07339_ (
    .A1(_02397_),
    .A2(_02402_),
    .ZN(_02403_)
  );
  AND2_X1 _07340_ (
    .A1(reg_dscratch0[13]),
    .A2(_00958_),
    .ZN(_02404_)
  );
  INV_X1 _07341_ (
    .A(_02404_),
    .ZN(_02405_)
  );
  AND2_X1 _07342_ (
    .A1(reg_pmp_1_addr[13]),
    .A2(_01008_),
    .ZN(_02406_)
  );
  INV_X1 _07343_ (
    .A(_02406_),
    .ZN(_02407_)
  );
  AND2_X1 _07344_ (
    .A1(_02405_),
    .A2(_02407_),
    .ZN(_02408_)
  );
  AND2_X1 _07345_ (
    .A1(reg_mscratch[13]),
    .A2(_00929_),
    .ZN(_02409_)
  );
  INV_X1 _07346_ (
    .A(_02409_),
    .ZN(_02410_)
  );
  AND2_X1 _07347_ (
    .A1(reg_mtvec[13]),
    .A2(_00940_),
    .ZN(_02411_)
  );
  INV_X1 _07348_ (
    .A(_02411_),
    .ZN(_02412_)
  );
  AND2_X1 _07349_ (
    .A1(_02410_),
    .A2(_02412_),
    .ZN(_02413_)
  );
  AND2_X1 _07350_ (
    .A1(_02408_),
    .A2(_02413_),
    .ZN(_02414_)
  );
  AND2_X1 _07351_ (
    .A1(reg_bp_0_address[13]),
    .A2(_00962_),
    .ZN(_02415_)
  );
  INV_X1 _07352_ (
    .A(_02415_),
    .ZN(_02416_)
  );
  AND2_X1 _07353_ (
    .A1(reg_pmp_5_addr[13]),
    .A2(_00948_),
    .ZN(_02417_)
  );
  INV_X1 _07354_ (
    .A(_02417_),
    .ZN(_02418_)
  );
  AND2_X1 _07355_ (
    .A1(_02416_),
    .A2(_02418_),
    .ZN(_02419_)
  );
  AND2_X1 _07356_ (
    .A1(reg_pmp_0_addr[13]),
    .A2(_01004_),
    .ZN(_02420_)
  );
  INV_X1 _07357_ (
    .A(_02420_),
    .ZN(_02421_)
  );
  AND2_X1 _07358_ (
    .A1(reg_dpc[13]),
    .A2(_00912_),
    .ZN(_02422_)
  );
  INV_X1 _07359_ (
    .A(_02422_),
    .ZN(_02423_)
  );
  AND2_X1 _07360_ (
    .A1(_02421_),
    .A2(_02423_),
    .ZN(_02424_)
  );
  AND2_X1 _07361_ (
    .A1(_02419_),
    .A2(_02424_),
    .ZN(_02425_)
  );
  AND2_X1 _07362_ (
    .A1(_02414_),
    .A2(_02425_),
    .ZN(_02426_)
  );
  AND2_X1 _07363_ (
    .A1(_02403_),
    .A2(_02426_),
    .ZN(_02427_)
  );
  AND2_X1 _07364_ (
    .A1(reg_pmp_7_addr[13]),
    .A2(_01016_),
    .ZN(_02428_)
  );
  INV_X1 _07365_ (
    .A(_02428_),
    .ZN(_02429_)
  );
  AND2_X1 _07366_ (
    .A1(large_[39]),
    .A2(_00991_),
    .ZN(_02430_)
  );
  INV_X1 _07367_ (
    .A(_02430_),
    .ZN(_02431_)
  );
  AND2_X1 _07368_ (
    .A1(large_1[7]),
    .A2(_00995_),
    .ZN(_02432_)
  );
  INV_X1 _07369_ (
    .A(_02432_),
    .ZN(_02433_)
  );
  AND2_X1 _07370_ (
    .A1(_02431_),
    .A2(_02433_),
    .ZN(_02434_)
  );
  AND2_X1 _07371_ (
    .A1(_02429_),
    .A2(_02434_),
    .ZN(_02435_)
  );
  AND2_X1 _07372_ (
    .A1(large_1[39]),
    .A2(_01019_),
    .ZN(_02436_)
  );
  INV_X1 _07373_ (
    .A(_02436_),
    .ZN(_02437_)
  );
  AND2_X1 _07374_ (
    .A1(reg_pmp_2_addr[13]),
    .A2(_00953_),
    .ZN(_02438_)
  );
  INV_X1 _07375_ (
    .A(_02438_),
    .ZN(_02439_)
  );
  AND2_X1 _07376_ (
    .A1(reg_mcause[13]),
    .A2(_01001_),
    .ZN(_02440_)
  );
  INV_X1 _07377_ (
    .A(_02440_),
    .ZN(_02441_)
  );
  AND2_X1 _07378_ (
    .A1(_02439_),
    .A2(_02441_),
    .ZN(_02442_)
  );
  AND2_X1 _07379_ (
    .A1(_02437_),
    .A2(_02442_),
    .ZN(_02443_)
  );
  AND2_X1 _07380_ (
    .A1(reg_pmp_6_addr[13]),
    .A2(_00978_),
    .ZN(_02444_)
  );
  INV_X1 _07381_ (
    .A(_02444_),
    .ZN(_02445_)
  );
  AND2_X1 _07382_ (
    .A1(large_[7]),
    .A2(_00985_),
    .ZN(_02446_)
  );
  INV_X1 _07383_ (
    .A(_02446_),
    .ZN(_02447_)
  );
  AND2_X1 _07384_ (
    .A1(_02445_),
    .A2(_02447_),
    .ZN(_02448_)
  );
  AND2_X1 _07385_ (
    .A1(_02443_),
    .A2(_02448_),
    .ZN(_02449_)
  );
  AND2_X1 _07386_ (
    .A1(_02435_),
    .A2(_02449_),
    .ZN(_02450_)
  );
  AND2_X1 _07387_ (
    .A1(_02427_),
    .A2(_02450_),
    .ZN(_02451_)
  );
  INV_X1 _07388_ (
    .A(_02451_),
    .ZN(io_rw_rdata[13])
  );
  AND2_X1 _07389_ (
    .A1(io_rw_cmd[1]),
    .A2(_00848_),
    .ZN(_02452_)
  );
  AND2_X1 _07390_ (
    .A1(io_rw_rdata[13]),
    .A2(_02452_),
    .ZN(_02453_)
  );
  INV_X1 _07391_ (
    .A(_02453_),
    .ZN(_02454_)
  );
  AND2_X1 _07392_ (
    .A1(_02392_),
    .A2(_02454_),
    .ZN(_02455_)
  );
  INV_X1 _07393_ (
    .A(_02455_),
    .ZN(_02456_)
  );
  MUX2_X1 _07394_ (
    .A(reg_pmp_5_addr[13]),
    .B(_02456_),
    .S(_01525_),
    .Z(_00040_)
  );
  AND2_X1 _07395_ (
    .A1(io_rw_wdata[14]),
    .A2(_00903_),
    .ZN(_02457_)
  );
  INV_X1 _07396_ (
    .A(_02457_),
    .ZN(_02458_)
  );
  AND2_X1 _07397_ (
    .A1(reg_pmp_0_addr[14]),
    .A2(_01004_),
    .ZN(_02459_)
  );
  INV_X1 _07398_ (
    .A(_02459_),
    .ZN(_02460_)
  );
  AND2_X1 _07399_ (
    .A1(reg_dscratch0[14]),
    .A2(_00958_),
    .ZN(_02461_)
  );
  INV_X1 _07400_ (
    .A(_02461_),
    .ZN(_02462_)
  );
  AND2_X1 _07401_ (
    .A1(_02460_),
    .A2(_02462_),
    .ZN(_02463_)
  );
  AND2_X1 _07402_ (
    .A1(reg_pmp_3_addr[14]),
    .A2(_01011_),
    .ZN(_02464_)
  );
  INV_X1 _07403_ (
    .A(_02464_),
    .ZN(_02465_)
  );
  AND2_X1 _07404_ (
    .A1(reg_mtvec[14]),
    .A2(_00940_),
    .ZN(_02466_)
  );
  INV_X1 _07405_ (
    .A(_02466_),
    .ZN(_02467_)
  );
  AND2_X1 _07406_ (
    .A1(_02465_),
    .A2(_02467_),
    .ZN(_02468_)
  );
  AND2_X1 _07407_ (
    .A1(_02463_),
    .A2(_02468_),
    .ZN(_02469_)
  );
  AND2_X1 _07408_ (
    .A1(reg_dpc[14]),
    .A2(_00912_),
    .ZN(_02470_)
  );
  INV_X1 _07409_ (
    .A(_02470_),
    .ZN(_02471_)
  );
  AND2_X1 _07410_ (
    .A1(reg_bp_0_address[14]),
    .A2(_00962_),
    .ZN(_02472_)
  );
  INV_X1 _07411_ (
    .A(_02472_),
    .ZN(_02473_)
  );
  AND2_X1 _07412_ (
    .A1(_02471_),
    .A2(_02473_),
    .ZN(_02474_)
  );
  AND2_X1 _07413_ (
    .A1(reg_pmp_5_addr[14]),
    .A2(_00948_),
    .ZN(_02475_)
  );
  INV_X1 _07414_ (
    .A(_02475_),
    .ZN(_02476_)
  );
  AND2_X1 _07415_ (
    .A1(reg_pmp_1_addr[14]),
    .A2(_01008_),
    .ZN(_02477_)
  );
  INV_X1 _07416_ (
    .A(_02477_),
    .ZN(_02478_)
  );
  AND2_X1 _07417_ (
    .A1(_02476_),
    .A2(_02478_),
    .ZN(_02479_)
  );
  AND2_X1 _07418_ (
    .A1(_02474_),
    .A2(_02479_),
    .ZN(_02480_)
  );
  AND2_X1 _07419_ (
    .A1(reg_mscratch[14]),
    .A2(_00929_),
    .ZN(_02481_)
  );
  INV_X1 _07420_ (
    .A(_02481_),
    .ZN(_02482_)
  );
  AND2_X1 _07421_ (
    .A1(reg_mcause[14]),
    .A2(_01001_),
    .ZN(_02483_)
  );
  INV_X1 _07422_ (
    .A(_02483_),
    .ZN(_02484_)
  );
  AND2_X1 _07423_ (
    .A1(_02482_),
    .A2(_02484_),
    .ZN(_02485_)
  );
  AND2_X1 _07424_ (
    .A1(reg_mepc[14]),
    .A2(_00943_),
    .ZN(_02486_)
  );
  INV_X1 _07425_ (
    .A(_02486_),
    .ZN(_02487_)
  );
  AND2_X1 _07426_ (
    .A1(reg_mtval[14]),
    .A2(_00926_),
    .ZN(_02488_)
  );
  INV_X1 _07427_ (
    .A(_02488_),
    .ZN(_02489_)
  );
  AND2_X1 _07428_ (
    .A1(_02487_),
    .A2(_02489_),
    .ZN(_02490_)
  );
  AND2_X1 _07429_ (
    .A1(_02485_),
    .A2(_02490_),
    .ZN(_02491_)
  );
  AND2_X1 _07430_ (
    .A1(_02480_),
    .A2(_02491_),
    .ZN(_02492_)
  );
  AND2_X1 _07431_ (
    .A1(_02469_),
    .A2(_02492_),
    .ZN(_02493_)
  );
  AND2_X1 _07432_ (
    .A1(large_1[8]),
    .A2(_00995_),
    .ZN(_02494_)
  );
  INV_X1 _07433_ (
    .A(_02494_),
    .ZN(_02495_)
  );
  AND2_X1 _07434_ (
    .A1(reg_pmp_6_addr[14]),
    .A2(_00978_),
    .ZN(_02496_)
  );
  INV_X1 _07435_ (
    .A(_02496_),
    .ZN(_02497_)
  );
  AND2_X1 _07436_ (
    .A1(reg_pmp_7_addr[14]),
    .A2(_01016_),
    .ZN(_02498_)
  );
  INV_X1 _07437_ (
    .A(_02498_),
    .ZN(_02499_)
  );
  AND2_X1 _07438_ (
    .A1(_02497_),
    .A2(_02499_),
    .ZN(_02500_)
  );
  AND2_X1 _07439_ (
    .A1(_02495_),
    .A2(_02500_),
    .ZN(_02501_)
  );
  AND2_X1 _07440_ (
    .A1(large_[8]),
    .A2(_00985_),
    .ZN(_02502_)
  );
  INV_X1 _07441_ (
    .A(_02502_),
    .ZN(_02503_)
  );
  AND2_X1 _07442_ (
    .A1(reg_pmp_4_addr[14]),
    .A2(_00968_),
    .ZN(_02504_)
  );
  INV_X1 _07443_ (
    .A(_02504_),
    .ZN(_02505_)
  );
  AND2_X1 _07444_ (
    .A1(reg_pmp_2_addr[14]),
    .A2(_00953_),
    .ZN(_02506_)
  );
  INV_X1 _07445_ (
    .A(_02506_),
    .ZN(_02507_)
  );
  AND2_X1 _07446_ (
    .A1(_02505_),
    .A2(_02507_),
    .ZN(_02508_)
  );
  AND2_X1 _07447_ (
    .A1(_02503_),
    .A2(_02508_),
    .ZN(_02509_)
  );
  AND2_X1 _07448_ (
    .A1(large_1[40]),
    .A2(_01019_),
    .ZN(_02510_)
  );
  INV_X1 _07449_ (
    .A(_02510_),
    .ZN(_02511_)
  );
  AND2_X1 _07450_ (
    .A1(large_[40]),
    .A2(_00991_),
    .ZN(_02512_)
  );
  INV_X1 _07451_ (
    .A(_02512_),
    .ZN(_02513_)
  );
  AND2_X1 _07452_ (
    .A1(_02511_),
    .A2(_02513_),
    .ZN(_02514_)
  );
  AND2_X1 _07453_ (
    .A1(_02509_),
    .A2(_02514_),
    .ZN(_02515_)
  );
  AND2_X1 _07454_ (
    .A1(_02501_),
    .A2(_02515_),
    .ZN(_02516_)
  );
  AND2_X1 _07455_ (
    .A1(_02493_),
    .A2(_02516_),
    .ZN(_02517_)
  );
  INV_X1 _07456_ (
    .A(_02517_),
    .ZN(io_rw_rdata[14])
  );
  AND2_X1 _07457_ (
    .A1(io_rw_cmd[1]),
    .A2(_00849_),
    .ZN(_02518_)
  );
  AND2_X1 _07458_ (
    .A1(io_rw_rdata[14]),
    .A2(_02518_),
    .ZN(_02519_)
  );
  INV_X1 _07459_ (
    .A(_02519_),
    .ZN(_02520_)
  );
  AND2_X1 _07460_ (
    .A1(_02458_),
    .A2(_02520_),
    .ZN(_02521_)
  );
  INV_X1 _07461_ (
    .A(_02521_),
    .ZN(_02522_)
  );
  MUX2_X1 _07462_ (
    .A(reg_pmp_5_addr[14]),
    .B(_02522_),
    .S(_01525_),
    .Z(_00041_)
  );
  AND2_X1 _07463_ (
    .A1(io_rw_wdata[15]),
    .A2(_00903_),
    .ZN(_02523_)
  );
  INV_X1 _07464_ (
    .A(_02523_),
    .ZN(_02524_)
  );
  AND2_X1 _07465_ (
    .A1(reg_pmp_5_cfg_l),
    .A2(_00894_),
    .ZN(_02525_)
  );
  INV_X1 _07466_ (
    .A(_02525_),
    .ZN(_02526_)
  );
  AND2_X1 _07467_ (
    .A1(reg_pmp_1_cfg_l),
    .A2(_00916_),
    .ZN(_02527_)
  );
  INV_X1 _07468_ (
    .A(_02527_),
    .ZN(_02528_)
  );
  AND2_X1 _07469_ (
    .A1(_02526_),
    .A2(_02528_),
    .ZN(_02529_)
  );
  AND2_X1 _07470_ (
    .A1(reg_pmp_2_addr[15]),
    .A2(_00953_),
    .ZN(_02530_)
  );
  INV_X1 _07471_ (
    .A(_02530_),
    .ZN(_02531_)
  );
  AND2_X1 _07472_ (
    .A1(reg_bp_0_address[15]),
    .A2(_00962_),
    .ZN(_02532_)
  );
  INV_X1 _07473_ (
    .A(_02532_),
    .ZN(_02533_)
  );
  AND2_X1 _07474_ (
    .A1(_02531_),
    .A2(_02533_),
    .ZN(_02534_)
  );
  AND2_X1 _07475_ (
    .A1(_02529_),
    .A2(_02534_),
    .ZN(_02535_)
  );
  AND2_X1 _07476_ (
    .A1(reg_pmp_1_addr[15]),
    .A2(_01008_),
    .ZN(_02536_)
  );
  INV_X1 _07477_ (
    .A(_02536_),
    .ZN(_02537_)
  );
  AND2_X1 _07478_ (
    .A1(reg_pmp_3_addr[15]),
    .A2(_01011_),
    .ZN(_02538_)
  );
  INV_X1 _07479_ (
    .A(_02538_),
    .ZN(_02539_)
  );
  AND2_X1 _07480_ (
    .A1(_02537_),
    .A2(_02539_),
    .ZN(_02540_)
  );
  AND2_X1 _07481_ (
    .A1(reg_dcsr_ebreakm),
    .A2(_01381_),
    .ZN(_02541_)
  );
  INV_X1 _07482_ (
    .A(_02541_),
    .ZN(_02542_)
  );
  AND2_X1 _07483_ (
    .A1(reg_pmp_5_addr[15]),
    .A2(_00948_),
    .ZN(_02543_)
  );
  INV_X1 _07484_ (
    .A(_02543_),
    .ZN(_02544_)
  );
  AND2_X1 _07485_ (
    .A1(_02542_),
    .A2(_02544_),
    .ZN(_02545_)
  );
  AND2_X1 _07486_ (
    .A1(_02540_),
    .A2(_02545_),
    .ZN(_02546_)
  );
  AND2_X1 _07487_ (
    .A1(_02535_),
    .A2(_02546_),
    .ZN(_02547_)
  );
  AND2_X1 _07488_ (
    .A1(reg_mtvec[15]),
    .A2(_00940_),
    .ZN(_02548_)
  );
  INV_X1 _07489_ (
    .A(_02548_),
    .ZN(_02549_)
  );
  AND2_X1 _07490_ (
    .A1(reg_dscratch0[15]),
    .A2(_00958_),
    .ZN(_02550_)
  );
  INV_X1 _07491_ (
    .A(_02550_),
    .ZN(_02551_)
  );
  AND2_X1 _07492_ (
    .A1(reg_mtval[15]),
    .A2(_00926_),
    .ZN(_02552_)
  );
  INV_X1 _07493_ (
    .A(_02552_),
    .ZN(_02553_)
  );
  AND2_X1 _07494_ (
    .A1(_02551_),
    .A2(_02553_),
    .ZN(_02554_)
  );
  AND2_X1 _07495_ (
    .A1(_02549_),
    .A2(_02554_),
    .ZN(_02555_)
  );
  AND2_X1 _07496_ (
    .A1(reg_dpc[15]),
    .A2(_00912_),
    .ZN(_02556_)
  );
  INV_X1 _07497_ (
    .A(_02556_),
    .ZN(_02557_)
  );
  AND2_X1 _07498_ (
    .A1(reg_mepc[15]),
    .A2(_00943_),
    .ZN(_02558_)
  );
  INV_X1 _07499_ (
    .A(_02558_),
    .ZN(_02559_)
  );
  AND2_X1 _07500_ (
    .A1(_02557_),
    .A2(_02559_),
    .ZN(_02560_)
  );
  AND2_X1 _07501_ (
    .A1(reg_mscratch[15]),
    .A2(_00929_),
    .ZN(_02561_)
  );
  INV_X1 _07502_ (
    .A(_02561_),
    .ZN(_02562_)
  );
  AND2_X1 _07503_ (
    .A1(reg_mcause[15]),
    .A2(_01001_),
    .ZN(_02563_)
  );
  INV_X1 _07504_ (
    .A(_02563_),
    .ZN(_02564_)
  );
  AND2_X1 _07505_ (
    .A1(_02562_),
    .A2(_02564_),
    .ZN(_02565_)
  );
  AND2_X1 _07506_ (
    .A1(_02560_),
    .A2(_02565_),
    .ZN(_02566_)
  );
  AND2_X1 _07507_ (
    .A1(_02555_),
    .A2(_02566_),
    .ZN(_02567_)
  );
  AND2_X1 _07508_ (
    .A1(_02547_),
    .A2(_02567_),
    .ZN(_02568_)
  );
  AND2_X1 _07509_ (
    .A1(large_1[9]),
    .A2(_00995_),
    .ZN(_02569_)
  );
  INV_X1 _07510_ (
    .A(_02569_),
    .ZN(_02570_)
  );
  AND2_X1 _07511_ (
    .A1(large_1[41]),
    .A2(_01019_),
    .ZN(_02571_)
  );
  INV_X1 _07512_ (
    .A(_02571_),
    .ZN(_02572_)
  );
  AND2_X1 _07513_ (
    .A1(large_[9]),
    .A2(_00985_),
    .ZN(_02573_)
  );
  INV_X1 _07514_ (
    .A(_02573_),
    .ZN(_02574_)
  );
  AND2_X1 _07515_ (
    .A1(_02572_),
    .A2(_02574_),
    .ZN(_02575_)
  );
  AND2_X1 _07516_ (
    .A1(_02570_),
    .A2(_02575_),
    .ZN(_02576_)
  );
  AND2_X1 _07517_ (
    .A1(reg_pmp_6_addr[15]),
    .A2(_00978_),
    .ZN(_02577_)
  );
  INV_X1 _07518_ (
    .A(_02577_),
    .ZN(_02578_)
  );
  AND2_X1 _07519_ (
    .A1(reg_pmp_4_addr[15]),
    .A2(_00968_),
    .ZN(_02579_)
  );
  INV_X1 _07520_ (
    .A(_02579_),
    .ZN(_02580_)
  );
  AND2_X1 _07521_ (
    .A1(reg_pmp_0_addr[15]),
    .A2(_01004_),
    .ZN(_02581_)
  );
  INV_X1 _07522_ (
    .A(_02581_),
    .ZN(_02582_)
  );
  AND2_X1 _07523_ (
    .A1(_02580_),
    .A2(_02582_),
    .ZN(_02583_)
  );
  AND2_X1 _07524_ (
    .A1(_02578_),
    .A2(_02583_),
    .ZN(_02584_)
  );
  AND2_X1 _07525_ (
    .A1(reg_pmp_7_addr[15]),
    .A2(_01016_),
    .ZN(_02585_)
  );
  INV_X1 _07526_ (
    .A(_02585_),
    .ZN(_02586_)
  );
  AND2_X1 _07527_ (
    .A1(large_[41]),
    .A2(_00991_),
    .ZN(_02587_)
  );
  INV_X1 _07528_ (
    .A(_02587_),
    .ZN(_02588_)
  );
  AND2_X1 _07529_ (
    .A1(_02586_),
    .A2(_02588_),
    .ZN(_02589_)
  );
  AND2_X1 _07530_ (
    .A1(_02584_),
    .A2(_02589_),
    .ZN(_02590_)
  );
  AND2_X1 _07531_ (
    .A1(_02576_),
    .A2(_02590_),
    .ZN(_02591_)
  );
  AND2_X1 _07532_ (
    .A1(_02568_),
    .A2(_02591_),
    .ZN(_02592_)
  );
  INV_X1 _07533_ (
    .A(_02592_),
    .ZN(io_rw_rdata[15])
  );
  AND2_X1 _07534_ (
    .A1(io_rw_cmd[1]),
    .A2(_00850_),
    .ZN(_02593_)
  );
  AND2_X1 _07535_ (
    .A1(io_rw_rdata[15]),
    .A2(_02593_),
    .ZN(_02594_)
  );
  INV_X1 _07536_ (
    .A(_02594_),
    .ZN(_02595_)
  );
  AND2_X1 _07537_ (
    .A1(_02524_),
    .A2(_02595_),
    .ZN(_02596_)
  );
  INV_X1 _07538_ (
    .A(_02596_),
    .ZN(_02597_)
  );
  MUX2_X1 _07539_ (
    .A(reg_pmp_5_addr[15]),
    .B(_02597_),
    .S(_01525_),
    .Z(_00042_)
  );
  MUX2_X1 _07540_ (
    .A(reg_pmp_5_addr[16]),
    .B(_01035_),
    .S(_01525_),
    .Z(_00043_)
  );
  AND2_X1 _07541_ (
    .A1(io_rw_wdata[17]),
    .A2(_00903_),
    .ZN(_02598_)
  );
  INV_X1 _07542_ (
    .A(_02598_),
    .ZN(_02599_)
  );
  AND2_X1 _07543_ (
    .A1(reg_mcause[17]),
    .A2(_01001_),
    .ZN(_02600_)
  );
  INV_X1 _07544_ (
    .A(_02600_),
    .ZN(_02601_)
  );
  AND2_X1 _07545_ (
    .A1(reg_mscratch[17]),
    .A2(_00929_),
    .ZN(_02602_)
  );
  INV_X1 _07546_ (
    .A(_02602_),
    .ZN(_02603_)
  );
  AND2_X1 _07547_ (
    .A1(_02601_),
    .A2(_02603_),
    .ZN(_02604_)
  );
  AND2_X1 _07548_ (
    .A1(reg_mtvec[17]),
    .A2(_00940_),
    .ZN(_02605_)
  );
  INV_X1 _07549_ (
    .A(_02605_),
    .ZN(_02606_)
  );
  AND2_X1 _07550_ (
    .A1(reg_mepc[17]),
    .A2(_00943_),
    .ZN(_02607_)
  );
  INV_X1 _07551_ (
    .A(_02607_),
    .ZN(_02608_)
  );
  AND2_X1 _07552_ (
    .A1(_02606_),
    .A2(_02608_),
    .ZN(_02609_)
  );
  AND2_X1 _07553_ (
    .A1(_02604_),
    .A2(_02609_),
    .ZN(_02610_)
  );
  AND2_X1 _07554_ (
    .A1(reg_mtval[17]),
    .A2(_00926_),
    .ZN(_02611_)
  );
  INV_X1 _07555_ (
    .A(_02611_),
    .ZN(_02612_)
  );
  AND2_X1 _07556_ (
    .A1(reg_dpc[17]),
    .A2(_00912_),
    .ZN(_02613_)
  );
  INV_X1 _07557_ (
    .A(_02613_),
    .ZN(_02614_)
  );
  AND2_X1 _07558_ (
    .A1(_02612_),
    .A2(_02614_),
    .ZN(_02615_)
  );
  AND2_X1 _07559_ (
    .A1(reg_pmp_4_addr[17]),
    .A2(_00968_),
    .ZN(_02616_)
  );
  INV_X1 _07560_ (
    .A(_02616_),
    .ZN(_02617_)
  );
  AND2_X1 _07561_ (
    .A1(reg_pmp_6_cfg_w),
    .A2(_00894_),
    .ZN(_02618_)
  );
  INV_X1 _07562_ (
    .A(_02618_),
    .ZN(_02619_)
  );
  AND2_X1 _07563_ (
    .A1(_02617_),
    .A2(_02619_),
    .ZN(_02620_)
  );
  AND2_X1 _07564_ (
    .A1(_02615_),
    .A2(_02620_),
    .ZN(_02621_)
  );
  AND2_X1 _07565_ (
    .A1(reg_bp_0_address[17]),
    .A2(_00962_),
    .ZN(_02622_)
  );
  INV_X1 _07566_ (
    .A(_02622_),
    .ZN(_02623_)
  );
  AND2_X1 _07567_ (
    .A1(reg_pmp_5_addr[17]),
    .A2(_00948_),
    .ZN(_02624_)
  );
  INV_X1 _07568_ (
    .A(_02624_),
    .ZN(_02625_)
  );
  AND2_X1 _07569_ (
    .A1(_02623_),
    .A2(_02625_),
    .ZN(_02626_)
  );
  AND2_X1 _07570_ (
    .A1(reg_pmp_2_cfg_w),
    .A2(_00916_),
    .ZN(_02627_)
  );
  INV_X1 _07571_ (
    .A(_02627_),
    .ZN(_02628_)
  );
  AND2_X1 _07572_ (
    .A1(reg_dscratch0[17]),
    .A2(_00958_),
    .ZN(_02629_)
  );
  INV_X1 _07573_ (
    .A(_02629_),
    .ZN(_02630_)
  );
  AND2_X1 _07574_ (
    .A1(_02628_),
    .A2(_02630_),
    .ZN(_02631_)
  );
  AND2_X1 _07575_ (
    .A1(_02626_),
    .A2(_02631_),
    .ZN(_02632_)
  );
  AND2_X1 _07576_ (
    .A1(_02621_),
    .A2(_02632_),
    .ZN(_02633_)
  );
  AND2_X1 _07577_ (
    .A1(_02610_),
    .A2(_02633_),
    .ZN(_02634_)
  );
  AND2_X1 _07578_ (
    .A1(reg_pmp_7_addr[17]),
    .A2(_01016_),
    .ZN(_02635_)
  );
  INV_X1 _07579_ (
    .A(_02635_),
    .ZN(_02636_)
  );
  AND2_X1 _07580_ (
    .A1(large_[11]),
    .A2(_00985_),
    .ZN(_02637_)
  );
  INV_X1 _07581_ (
    .A(_02637_),
    .ZN(_02638_)
  );
  AND2_X1 _07582_ (
    .A1(_02636_),
    .A2(_02638_),
    .ZN(_02639_)
  );
  AND2_X1 _07583_ (
    .A1(reg_pmp_6_addr[17]),
    .A2(_00978_),
    .ZN(_02640_)
  );
  INV_X1 _07584_ (
    .A(_02640_),
    .ZN(_02641_)
  );
  AND2_X1 _07585_ (
    .A1(large_1[11]),
    .A2(_00995_),
    .ZN(_02642_)
  );
  INV_X1 _07586_ (
    .A(_02642_),
    .ZN(_02643_)
  );
  AND2_X1 _07587_ (
    .A1(_02641_),
    .A2(_02643_),
    .ZN(_02644_)
  );
  AND2_X1 _07588_ (
    .A1(_02639_),
    .A2(_02644_),
    .ZN(_02645_)
  );
  AND2_X1 _07589_ (
    .A1(reg_pmp_3_addr[17]),
    .A2(_01011_),
    .ZN(_02646_)
  );
  INV_X1 _07590_ (
    .A(_02646_),
    .ZN(_02647_)
  );
  AND2_X1 _07591_ (
    .A1(reg_pmp_1_addr[17]),
    .A2(_01008_),
    .ZN(_02648_)
  );
  INV_X1 _07592_ (
    .A(_02648_),
    .ZN(_02649_)
  );
  AND2_X1 _07593_ (
    .A1(_02647_),
    .A2(_02649_),
    .ZN(_02650_)
  );
  AND2_X1 _07594_ (
    .A1(reg_pmp_0_addr[17]),
    .A2(_01004_),
    .ZN(_02651_)
  );
  INV_X1 _07595_ (
    .A(_02651_),
    .ZN(_02652_)
  );
  AND2_X1 _07596_ (
    .A1(reg_pmp_2_addr[17]),
    .A2(_00953_),
    .ZN(_02653_)
  );
  INV_X1 _07597_ (
    .A(_02653_),
    .ZN(_02654_)
  );
  AND2_X1 _07598_ (
    .A1(_02652_),
    .A2(_02654_),
    .ZN(_02655_)
  );
  AND2_X1 _07599_ (
    .A1(_02650_),
    .A2(_02655_),
    .ZN(_02656_)
  );
  AND2_X1 _07600_ (
    .A1(large_[43]),
    .A2(_00991_),
    .ZN(_02657_)
  );
  INV_X1 _07601_ (
    .A(_02657_),
    .ZN(_02658_)
  );
  AND2_X1 _07602_ (
    .A1(large_1[43]),
    .A2(_01019_),
    .ZN(_02659_)
  );
  INV_X1 _07603_ (
    .A(_02659_),
    .ZN(_02660_)
  );
  AND2_X1 _07604_ (
    .A1(_02658_),
    .A2(_02660_),
    .ZN(_02661_)
  );
  AND2_X1 _07605_ (
    .A1(_02656_),
    .A2(_02661_),
    .ZN(_02662_)
  );
  AND2_X1 _07606_ (
    .A1(_02645_),
    .A2(_02662_),
    .ZN(_02663_)
  );
  AND2_X1 _07607_ (
    .A1(_02634_),
    .A2(_02663_),
    .ZN(_02664_)
  );
  INV_X1 _07608_ (
    .A(_02664_),
    .ZN(io_rw_rdata[17])
  );
  AND2_X1 _07609_ (
    .A1(io_rw_cmd[1]),
    .A2(_00852_),
    .ZN(_02665_)
  );
  AND2_X1 _07610_ (
    .A1(io_rw_rdata[17]),
    .A2(_02665_),
    .ZN(_02666_)
  );
  INV_X1 _07611_ (
    .A(_02666_),
    .ZN(_02667_)
  );
  AND2_X1 _07612_ (
    .A1(_02599_),
    .A2(_02667_),
    .ZN(_02668_)
  );
  INV_X1 _07613_ (
    .A(_02668_),
    .ZN(_02669_)
  );
  MUX2_X1 _07614_ (
    .A(reg_pmp_5_addr[17]),
    .B(_02669_),
    .S(_01525_),
    .Z(_00044_)
  );
  MUX2_X1 _07615_ (
    .A(reg_pmp_5_addr[18]),
    .B(_01107_),
    .S(_01525_),
    .Z(_00045_)
  );
  MUX2_X1 _07616_ (
    .A(reg_pmp_5_addr[19]),
    .B(_01199_),
    .S(_01525_),
    .Z(_00046_)
  );
  MUX2_X1 _07617_ (
    .A(reg_pmp_5_addr[20]),
    .B(_01277_),
    .S(_01525_),
    .Z(_00047_)
  );
  AND2_X1 _07618_ (
    .A1(io_rw_wdata[21]),
    .A2(_00903_),
    .ZN(_02670_)
  );
  INV_X1 _07619_ (
    .A(_02670_),
    .ZN(_02671_)
  );
  AND2_X1 _07620_ (
    .A1(reg_dpc[21]),
    .A2(_00912_),
    .ZN(_02672_)
  );
  INV_X1 _07621_ (
    .A(_02672_),
    .ZN(_02673_)
  );
  AND2_X1 _07622_ (
    .A1(reg_bp_0_address[21]),
    .A2(_00962_),
    .ZN(_02674_)
  );
  INV_X1 _07623_ (
    .A(_02674_),
    .ZN(_02675_)
  );
  AND2_X1 _07624_ (
    .A1(_02673_),
    .A2(_02675_),
    .ZN(_02676_)
  );
  AND2_X1 _07625_ (
    .A1(reg_pmp_2_addr[21]),
    .A2(_00953_),
    .ZN(_02677_)
  );
  INV_X1 _07626_ (
    .A(_02677_),
    .ZN(_02678_)
  );
  AND2_X1 _07627_ (
    .A1(reg_dscratch0[21]),
    .A2(_00958_),
    .ZN(_02679_)
  );
  INV_X1 _07628_ (
    .A(_02679_),
    .ZN(_02680_)
  );
  AND2_X1 _07629_ (
    .A1(_02678_),
    .A2(_02680_),
    .ZN(_02681_)
  );
  AND2_X1 _07630_ (
    .A1(_02676_),
    .A2(_02681_),
    .ZN(_02682_)
  );
  AND2_X1 _07631_ (
    .A1(reg_pmp_5_addr[21]),
    .A2(_00948_),
    .ZN(_02683_)
  );
  INV_X1 _07632_ (
    .A(_02683_),
    .ZN(_02684_)
  );
  AND2_X1 _07633_ (
    .A1(reg_pmp_1_addr[21]),
    .A2(_01008_),
    .ZN(_02685_)
  );
  INV_X1 _07634_ (
    .A(_02685_),
    .ZN(_02686_)
  );
  AND2_X1 _07635_ (
    .A1(_02684_),
    .A2(_02686_),
    .ZN(_02687_)
  );
  AND2_X1 _07636_ (
    .A1(reg_mepc[21]),
    .A2(_00943_),
    .ZN(_02688_)
  );
  INV_X1 _07637_ (
    .A(_02688_),
    .ZN(_02689_)
  );
  AND2_X1 _07638_ (
    .A1(reg_mtval[21]),
    .A2(_00926_),
    .ZN(_02690_)
  );
  INV_X1 _07639_ (
    .A(_02690_),
    .ZN(_02691_)
  );
  AND2_X1 _07640_ (
    .A1(_02689_),
    .A2(_02691_),
    .ZN(_02692_)
  );
  AND2_X1 _07641_ (
    .A1(_02687_),
    .A2(_02692_),
    .ZN(_02693_)
  );
  AND2_X1 _07642_ (
    .A1(reg_pmp_4_addr[21]),
    .A2(_00968_),
    .ZN(_02694_)
  );
  INV_X1 _07643_ (
    .A(_02694_),
    .ZN(_02695_)
  );
  AND2_X1 _07644_ (
    .A1(reg_mtvec[21]),
    .A2(_00940_),
    .ZN(_02696_)
  );
  INV_X1 _07645_ (
    .A(_02696_),
    .ZN(_02697_)
  );
  AND2_X1 _07646_ (
    .A1(_02695_),
    .A2(_02697_),
    .ZN(_02698_)
  );
  AND2_X1 _07647_ (
    .A1(reg_pmp_0_addr[21]),
    .A2(_01004_),
    .ZN(_02699_)
  );
  INV_X1 _07648_ (
    .A(_02699_),
    .ZN(_02700_)
  );
  AND2_X1 _07649_ (
    .A1(reg_mcause[21]),
    .A2(_01001_),
    .ZN(_02701_)
  );
  INV_X1 _07650_ (
    .A(_02701_),
    .ZN(_02702_)
  );
  AND2_X1 _07651_ (
    .A1(_02700_),
    .A2(_02702_),
    .ZN(_02703_)
  );
  AND2_X1 _07652_ (
    .A1(_02698_),
    .A2(_02703_),
    .ZN(_02704_)
  );
  AND2_X1 _07653_ (
    .A1(_02693_),
    .A2(_02704_),
    .ZN(_02705_)
  );
  AND2_X1 _07654_ (
    .A1(_02682_),
    .A2(_02705_),
    .ZN(_02706_)
  );
  AND2_X1 _07655_ (
    .A1(large_1[47]),
    .A2(_01019_),
    .ZN(_02707_)
  );
  INV_X1 _07656_ (
    .A(_02707_),
    .ZN(_02708_)
  );
  AND2_X1 _07657_ (
    .A1(reg_pmp_7_addr[21]),
    .A2(_01016_),
    .ZN(_02709_)
  );
  INV_X1 _07658_ (
    .A(_02709_),
    .ZN(_02710_)
  );
  AND2_X1 _07659_ (
    .A1(large_[47]),
    .A2(_00991_),
    .ZN(_02711_)
  );
  INV_X1 _07660_ (
    .A(_02711_),
    .ZN(_02712_)
  );
  AND2_X1 _07661_ (
    .A1(_02710_),
    .A2(_02712_),
    .ZN(_02713_)
  );
  AND2_X1 _07662_ (
    .A1(_02708_),
    .A2(_02713_),
    .ZN(_02714_)
  );
  AND2_X1 _07663_ (
    .A1(large_[15]),
    .A2(_00985_),
    .ZN(_02715_)
  );
  INV_X1 _07664_ (
    .A(_02715_),
    .ZN(_02716_)
  );
  AND2_X1 _07665_ (
    .A1(reg_mscratch[21]),
    .A2(_00929_),
    .ZN(_02717_)
  );
  INV_X1 _07666_ (
    .A(_02717_),
    .ZN(_02718_)
  );
  AND2_X1 _07667_ (
    .A1(reg_pmp_3_addr[21]),
    .A2(_01011_),
    .ZN(_02719_)
  );
  INV_X1 _07668_ (
    .A(_02719_),
    .ZN(_02720_)
  );
  AND2_X1 _07669_ (
    .A1(_02718_),
    .A2(_02720_),
    .ZN(_02721_)
  );
  AND2_X1 _07670_ (
    .A1(_02716_),
    .A2(_02721_),
    .ZN(_02722_)
  );
  AND2_X1 _07671_ (
    .A1(reg_pmp_6_addr[21]),
    .A2(_00978_),
    .ZN(_02723_)
  );
  INV_X1 _07672_ (
    .A(_02723_),
    .ZN(_02724_)
  );
  AND2_X1 _07673_ (
    .A1(large_1[15]),
    .A2(_00995_),
    .ZN(_02725_)
  );
  INV_X1 _07674_ (
    .A(_02725_),
    .ZN(_02726_)
  );
  AND2_X1 _07675_ (
    .A1(_02724_),
    .A2(_02726_),
    .ZN(_02727_)
  );
  AND2_X1 _07676_ (
    .A1(_02722_),
    .A2(_02727_),
    .ZN(_02728_)
  );
  AND2_X1 _07677_ (
    .A1(_02714_),
    .A2(_02728_),
    .ZN(_02729_)
  );
  AND2_X1 _07678_ (
    .A1(_02706_),
    .A2(_02729_),
    .ZN(_02730_)
  );
  INV_X1 _07679_ (
    .A(_02730_),
    .ZN(io_rw_rdata[21])
  );
  AND2_X1 _07680_ (
    .A1(io_rw_cmd[1]),
    .A2(_00856_),
    .ZN(_02731_)
  );
  AND2_X1 _07681_ (
    .A1(io_rw_rdata[21]),
    .A2(_02731_),
    .ZN(_02732_)
  );
  INV_X1 _07682_ (
    .A(_02732_),
    .ZN(_02733_)
  );
  AND2_X1 _07683_ (
    .A1(_02671_),
    .A2(_02733_),
    .ZN(_02734_)
  );
  INV_X1 _07684_ (
    .A(_02734_),
    .ZN(_02735_)
  );
  MUX2_X1 _07685_ (
    .A(reg_pmp_5_addr[21]),
    .B(_02735_),
    .S(_01525_),
    .Z(_00048_)
  );
  AND2_X1 _07686_ (
    .A1(io_rw_wdata[22]),
    .A2(_00903_),
    .ZN(_02736_)
  );
  INV_X1 _07687_ (
    .A(_02736_),
    .ZN(_02737_)
  );
  AND2_X1 _07688_ (
    .A1(reg_pmp_1_addr[22]),
    .A2(_01008_),
    .ZN(_02738_)
  );
  INV_X1 _07689_ (
    .A(_02738_),
    .ZN(_02739_)
  );
  AND2_X1 _07690_ (
    .A1(reg_pmp_5_addr[22]),
    .A2(_00948_),
    .ZN(_02740_)
  );
  INV_X1 _07691_ (
    .A(_02740_),
    .ZN(_02741_)
  );
  AND2_X1 _07692_ (
    .A1(reg_pmp_2_addr[22]),
    .A2(_00953_),
    .ZN(_02742_)
  );
  INV_X1 _07693_ (
    .A(_02742_),
    .ZN(_02743_)
  );
  AND2_X1 _07694_ (
    .A1(reg_dscratch0[22]),
    .A2(_00958_),
    .ZN(_02744_)
  );
  INV_X1 _07695_ (
    .A(_02744_),
    .ZN(_02745_)
  );
  AND2_X1 _07696_ (
    .A1(reg_mtvec[22]),
    .A2(_00940_),
    .ZN(_02746_)
  );
  INV_X1 _07697_ (
    .A(_02746_),
    .ZN(_02747_)
  );
  AND2_X1 _07698_ (
    .A1(reg_pmp_4_addr[22]),
    .A2(_00968_),
    .ZN(_02748_)
  );
  INV_X1 _07699_ (
    .A(_02748_),
    .ZN(_02749_)
  );
  AND2_X1 _07700_ (
    .A1(_02747_),
    .A2(_02749_),
    .ZN(_02750_)
  );
  AND2_X1 _07701_ (
    .A1(reg_mscratch[22]),
    .A2(_00929_),
    .ZN(_02751_)
  );
  INV_X1 _07702_ (
    .A(_02751_),
    .ZN(_02752_)
  );
  AND2_X1 _07703_ (
    .A1(reg_bp_0_address[22]),
    .A2(_00962_),
    .ZN(_02753_)
  );
  INV_X1 _07704_ (
    .A(_02753_),
    .ZN(_02754_)
  );
  AND2_X1 _07705_ (
    .A1(reg_pmp_3_addr[22]),
    .A2(_01011_),
    .ZN(_02755_)
  );
  INV_X1 _07706_ (
    .A(_02755_),
    .ZN(_02756_)
  );
  AND2_X1 _07707_ (
    .A1(reg_dpc[22]),
    .A2(_00912_),
    .ZN(_02757_)
  );
  INV_X1 _07708_ (
    .A(_02757_),
    .ZN(_02758_)
  );
  AND2_X1 _07709_ (
    .A1(reg_pmp_0_addr[22]),
    .A2(_01004_),
    .ZN(_02759_)
  );
  INV_X1 _07710_ (
    .A(_02759_),
    .ZN(_02760_)
  );
  AND2_X1 _07711_ (
    .A1(reg_mepc[22]),
    .A2(_00943_),
    .ZN(_02761_)
  );
  INV_X1 _07712_ (
    .A(_02761_),
    .ZN(_02762_)
  );
  AND2_X1 _07713_ (
    .A1(reg_pmp_7_addr[22]),
    .A2(_01016_),
    .ZN(_02763_)
  );
  INV_X1 _07714_ (
    .A(_02763_),
    .ZN(_02764_)
  );
  AND2_X1 _07715_ (
    .A1(reg_pmp_6_addr[22]),
    .A2(_00978_),
    .ZN(_02765_)
  );
  INV_X1 _07716_ (
    .A(_02765_),
    .ZN(_02766_)
  );
  AND2_X1 _07717_ (
    .A1(large_[48]),
    .A2(_00991_),
    .ZN(_02767_)
  );
  INV_X1 _07718_ (
    .A(_02767_),
    .ZN(_02768_)
  );
  AND2_X1 _07719_ (
    .A1(large_1[48]),
    .A2(_01019_),
    .ZN(_02769_)
  );
  INV_X1 _07720_ (
    .A(_02769_),
    .ZN(_02770_)
  );
  AND2_X1 _07721_ (
    .A1(reg_mtval[22]),
    .A2(_00926_),
    .ZN(_02771_)
  );
  INV_X1 _07722_ (
    .A(_02771_),
    .ZN(_02772_)
  );
  AND2_X1 _07723_ (
    .A1(reg_mcause[22]),
    .A2(_01001_),
    .ZN(_02773_)
  );
  INV_X1 _07724_ (
    .A(_02773_),
    .ZN(_02774_)
  );
  AND2_X1 _07725_ (
    .A1(_02752_),
    .A2(_02772_),
    .ZN(_02775_)
  );
  AND2_X1 _07726_ (
    .A1(_02774_),
    .A2(_02775_),
    .ZN(_02776_)
  );
  AND2_X1 _07727_ (
    .A1(_02739_),
    .A2(_02760_),
    .ZN(_02777_)
  );
  AND2_X1 _07728_ (
    .A1(large_[16]),
    .A2(_01027_),
    .ZN(_02778_)
  );
  INV_X1 _07729_ (
    .A(_02778_),
    .ZN(_02779_)
  );
  AND2_X1 _07730_ (
    .A1(large_1[16]),
    .A2(_01029_),
    .ZN(_02780_)
  );
  INV_X1 _07731_ (
    .A(_02780_),
    .ZN(_02781_)
  );
  AND2_X1 _07732_ (
    .A1(_02743_),
    .A2(_02766_),
    .ZN(_02782_)
  );
  AND2_X1 _07733_ (
    .A1(_02776_),
    .A2(_02782_),
    .ZN(_02783_)
  );
  AND2_X1 _07734_ (
    .A1(_02756_),
    .A2(_02777_),
    .ZN(_02784_)
  );
  AND2_X1 _07735_ (
    .A1(_02768_),
    .A2(_02770_),
    .ZN(_02785_)
  );
  AND2_X1 _07736_ (
    .A1(_02784_),
    .A2(_02785_),
    .ZN(_02786_)
  );
  AND2_X1 _07737_ (
    .A1(_02783_),
    .A2(_02786_),
    .ZN(_02787_)
  );
  AND2_X1 _07738_ (
    .A1(_02750_),
    .A2(_02764_),
    .ZN(_02788_)
  );
  AND2_X1 _07739_ (
    .A1(_02754_),
    .A2(_02762_),
    .ZN(_02789_)
  );
  AND2_X1 _07740_ (
    .A1(_02788_),
    .A2(_02789_),
    .ZN(_02790_)
  );
  AND2_X1 _07741_ (
    .A1(_02741_),
    .A2(_02745_),
    .ZN(_02791_)
  );
  AND2_X1 _07742_ (
    .A1(_02758_),
    .A2(_02779_),
    .ZN(_02792_)
  );
  AND2_X1 _07743_ (
    .A1(_02781_),
    .A2(_02792_),
    .ZN(_02793_)
  );
  AND2_X1 _07744_ (
    .A1(_02791_),
    .A2(_02793_),
    .ZN(_02794_)
  );
  AND2_X1 _07745_ (
    .A1(_02790_),
    .A2(_02794_),
    .ZN(_02795_)
  );
  AND2_X1 _07746_ (
    .A1(_02787_),
    .A2(_02795_),
    .ZN(_02796_)
  );
  INV_X1 _07747_ (
    .A(_02796_),
    .ZN(io_rw_rdata[22])
  );
  AND2_X1 _07748_ (
    .A1(io_rw_cmd[1]),
    .A2(_00857_),
    .ZN(_02797_)
  );
  AND2_X1 _07749_ (
    .A1(io_rw_rdata[22]),
    .A2(_02797_),
    .ZN(_02798_)
  );
  INV_X1 _07750_ (
    .A(_02798_),
    .ZN(_02799_)
  );
  AND2_X1 _07751_ (
    .A1(_02737_),
    .A2(_02799_),
    .ZN(_02800_)
  );
  INV_X1 _07752_ (
    .A(_02800_),
    .ZN(_02801_)
  );
  MUX2_X1 _07753_ (
    .A(reg_pmp_5_addr[22]),
    .B(_02801_),
    .S(_01525_),
    .Z(_00049_)
  );
  MUX2_X1 _07754_ (
    .A(reg_pmp_5_addr[23]),
    .B(_01360_),
    .S(_01525_),
    .Z(_00050_)
  );
  AND2_X1 _07755_ (
    .A1(io_rw_wdata[24]),
    .A2(_00903_),
    .ZN(_02802_)
  );
  INV_X1 _07756_ (
    .A(_02802_),
    .ZN(_02803_)
  );
  AND2_X1 _07757_ (
    .A1(reg_mcause[24]),
    .A2(_01001_),
    .ZN(_02804_)
  );
  INV_X1 _07758_ (
    .A(_02804_),
    .ZN(_02805_)
  );
  AND2_X1 _07759_ (
    .A1(reg_pmp_1_addr[24]),
    .A2(_01008_),
    .ZN(_02806_)
  );
  INV_X1 _07760_ (
    .A(_02806_),
    .ZN(_02807_)
  );
  AND2_X1 _07761_ (
    .A1(_02805_),
    .A2(_02807_),
    .ZN(_02808_)
  );
  AND2_X1 _07762_ (
    .A1(reg_mtvec[24]),
    .A2(_00940_),
    .ZN(_02809_)
  );
  INV_X1 _07763_ (
    .A(_02809_),
    .ZN(_02810_)
  );
  AND2_X1 _07764_ (
    .A1(reg_mscratch[24]),
    .A2(_00929_),
    .ZN(_02811_)
  );
  INV_X1 _07765_ (
    .A(_02811_),
    .ZN(_02812_)
  );
  AND2_X1 _07766_ (
    .A1(_02810_),
    .A2(_02812_),
    .ZN(_02813_)
  );
  AND2_X1 _07767_ (
    .A1(_02808_),
    .A2(_02813_),
    .ZN(_02814_)
  );
  AND2_X1 _07768_ (
    .A1(reg_mtval[24]),
    .A2(_00926_),
    .ZN(_02815_)
  );
  INV_X1 _07769_ (
    .A(_02815_),
    .ZN(_02816_)
  );
  AND2_X1 _07770_ (
    .A1(reg_pmp_0_addr[24]),
    .A2(_01004_),
    .ZN(_02817_)
  );
  INV_X1 _07771_ (
    .A(_02817_),
    .ZN(_02818_)
  );
  AND2_X1 _07772_ (
    .A1(_02816_),
    .A2(_02818_),
    .ZN(_02819_)
  );
  AND2_X1 _07773_ (
    .A1(reg_pmp_2_addr[24]),
    .A2(_00953_),
    .ZN(_02820_)
  );
  INV_X1 _07774_ (
    .A(_02820_),
    .ZN(_02821_)
  );
  AND2_X1 _07775_ (
    .A1(reg_dscratch0[24]),
    .A2(_00958_),
    .ZN(_02822_)
  );
  INV_X1 _07776_ (
    .A(_02822_),
    .ZN(_02823_)
  );
  AND2_X1 _07777_ (
    .A1(_02821_),
    .A2(_02823_),
    .ZN(_02824_)
  );
  AND2_X1 _07778_ (
    .A1(_02819_),
    .A2(_02824_),
    .ZN(_02825_)
  );
  AND2_X1 _07779_ (
    .A1(reg_mepc[24]),
    .A2(_00943_),
    .ZN(_02826_)
  );
  INV_X1 _07780_ (
    .A(_02826_),
    .ZN(_02827_)
  );
  AND2_X1 _07781_ (
    .A1(reg_pmp_4_addr[24]),
    .A2(_00968_),
    .ZN(_02828_)
  );
  INV_X1 _07782_ (
    .A(_02828_),
    .ZN(_02829_)
  );
  AND2_X1 _07783_ (
    .A1(_02827_),
    .A2(_02829_),
    .ZN(_02830_)
  );
  AND2_X1 _07784_ (
    .A1(reg_pmp_5_addr[24]),
    .A2(_00948_),
    .ZN(_02831_)
  );
  INV_X1 _07785_ (
    .A(_02831_),
    .ZN(_02832_)
  );
  AND2_X1 _07786_ (
    .A1(reg_dpc[24]),
    .A2(_00912_),
    .ZN(_02833_)
  );
  INV_X1 _07787_ (
    .A(_02833_),
    .ZN(_02834_)
  );
  AND2_X1 _07788_ (
    .A1(_02832_),
    .A2(_02834_),
    .ZN(_02835_)
  );
  AND2_X1 _07789_ (
    .A1(_02830_),
    .A2(_02835_),
    .ZN(_02836_)
  );
  AND2_X1 _07790_ (
    .A1(_02825_),
    .A2(_02836_),
    .ZN(_02837_)
  );
  AND2_X1 _07791_ (
    .A1(_02814_),
    .A2(_02837_),
    .ZN(_02838_)
  );
  AND2_X1 _07792_ (
    .A1(large_[18]),
    .A2(_00985_),
    .ZN(_02839_)
  );
  INV_X1 _07793_ (
    .A(_02839_),
    .ZN(_02840_)
  );
  AND2_X1 _07794_ (
    .A1(large_1[18]),
    .A2(_00995_),
    .ZN(_02841_)
  );
  INV_X1 _07795_ (
    .A(_02841_),
    .ZN(_02842_)
  );
  AND2_X1 _07796_ (
    .A1(_02840_),
    .A2(_02842_),
    .ZN(_02843_)
  );
  AND2_X1 _07797_ (
    .A1(reg_pmp_6_addr[24]),
    .A2(_00978_),
    .ZN(_02844_)
  );
  INV_X1 _07798_ (
    .A(_02844_),
    .ZN(_02845_)
  );
  AND2_X1 _07799_ (
    .A1(reg_pmp_7_addr[24]),
    .A2(_01016_),
    .ZN(_02846_)
  );
  INV_X1 _07800_ (
    .A(_02846_),
    .ZN(_02847_)
  );
  AND2_X1 _07801_ (
    .A1(_02845_),
    .A2(_02847_),
    .ZN(_02848_)
  );
  AND2_X1 _07802_ (
    .A1(_02843_),
    .A2(_02848_),
    .ZN(_02849_)
  );
  AND2_X1 _07803_ (
    .A1(large_1[50]),
    .A2(_01019_),
    .ZN(_02850_)
  );
  INV_X1 _07804_ (
    .A(_02850_),
    .ZN(_02851_)
  );
  AND2_X1 _07805_ (
    .A1(large_[50]),
    .A2(_00991_),
    .ZN(_02852_)
  );
  INV_X1 _07806_ (
    .A(_02852_),
    .ZN(_02853_)
  );
  AND2_X1 _07807_ (
    .A1(_02851_),
    .A2(_02853_),
    .ZN(_02854_)
  );
  AND2_X1 _07808_ (
    .A1(reg_pmp_3_cfg_r),
    .A2(_00916_),
    .ZN(_02855_)
  );
  INV_X1 _07809_ (
    .A(_02855_),
    .ZN(_02856_)
  );
  AND2_X1 _07810_ (
    .A1(reg_bp_0_address[24]),
    .A2(_00962_),
    .ZN(_02857_)
  );
  INV_X1 _07811_ (
    .A(_02857_),
    .ZN(_02858_)
  );
  AND2_X1 _07812_ (
    .A1(_02856_),
    .A2(_02858_),
    .ZN(_02859_)
  );
  AND2_X1 _07813_ (
    .A1(reg_pmp_7_cfg_r),
    .A2(_00894_),
    .ZN(_02860_)
  );
  INV_X1 _07814_ (
    .A(_02860_),
    .ZN(_02861_)
  );
  AND2_X1 _07815_ (
    .A1(reg_pmp_3_addr[24]),
    .A2(_01011_),
    .ZN(_02862_)
  );
  INV_X1 _07816_ (
    .A(_02862_),
    .ZN(_02863_)
  );
  AND2_X1 _07817_ (
    .A1(_02861_),
    .A2(_02863_),
    .ZN(_02864_)
  );
  AND2_X1 _07818_ (
    .A1(_02859_),
    .A2(_02864_),
    .ZN(_02865_)
  );
  AND2_X1 _07819_ (
    .A1(_02854_),
    .A2(_02865_),
    .ZN(_02866_)
  );
  AND2_X1 _07820_ (
    .A1(_02849_),
    .A2(_02866_),
    .ZN(_02867_)
  );
  AND2_X1 _07821_ (
    .A1(_02838_),
    .A2(_02867_),
    .ZN(_02868_)
  );
  INV_X1 _07822_ (
    .A(_02868_),
    .ZN(io_rw_rdata[24])
  );
  AND2_X1 _07823_ (
    .A1(io_rw_cmd[1]),
    .A2(_00859_),
    .ZN(_02869_)
  );
  AND2_X1 _07824_ (
    .A1(io_rw_rdata[24]),
    .A2(_02869_),
    .ZN(_02870_)
  );
  INV_X1 _07825_ (
    .A(_02870_),
    .ZN(_02871_)
  );
  AND2_X1 _07826_ (
    .A1(_02803_),
    .A2(_02871_),
    .ZN(_02872_)
  );
  INV_X1 _07827_ (
    .A(_02872_),
    .ZN(_02873_)
  );
  MUX2_X1 _07828_ (
    .A(reg_pmp_5_addr[24]),
    .B(_02873_),
    .S(_01525_),
    .Z(_00051_)
  );
  AND2_X1 _07829_ (
    .A1(io_rw_wdata[25]),
    .A2(_00903_),
    .ZN(_02874_)
  );
  INV_X1 _07830_ (
    .A(_02874_),
    .ZN(_02875_)
  );
  AND2_X1 _07831_ (
    .A1(reg_pmp_7_cfg_w),
    .A2(_00894_),
    .ZN(_02876_)
  );
  INV_X1 _07832_ (
    .A(_02876_),
    .ZN(_02877_)
  );
  AND2_X1 _07833_ (
    .A1(reg_pmp_4_addr[25]),
    .A2(_00968_),
    .ZN(_02878_)
  );
  INV_X1 _07834_ (
    .A(_02878_),
    .ZN(_02879_)
  );
  AND2_X1 _07835_ (
    .A1(_02877_),
    .A2(_02879_),
    .ZN(_02880_)
  );
  AND2_X1 _07836_ (
    .A1(reg_mtvec[25]),
    .A2(_00940_),
    .ZN(_02881_)
  );
  INV_X1 _07837_ (
    .A(_02881_),
    .ZN(_02882_)
  );
  AND2_X1 _07838_ (
    .A1(reg_pmp_5_addr[25]),
    .A2(_00948_),
    .ZN(_02883_)
  );
  INV_X1 _07839_ (
    .A(_02883_),
    .ZN(_02884_)
  );
  AND2_X1 _07840_ (
    .A1(_02882_),
    .A2(_02884_),
    .ZN(_02885_)
  );
  AND2_X1 _07841_ (
    .A1(_02880_),
    .A2(_02885_),
    .ZN(_02886_)
  );
  AND2_X1 _07842_ (
    .A1(reg_mepc[25]),
    .A2(_00943_),
    .ZN(_02887_)
  );
  INV_X1 _07843_ (
    .A(_02887_),
    .ZN(_02888_)
  );
  AND2_X1 _07844_ (
    .A1(reg_pmp_3_addr[25]),
    .A2(_01011_),
    .ZN(_02889_)
  );
  INV_X1 _07845_ (
    .A(_02889_),
    .ZN(_02890_)
  );
  AND2_X1 _07846_ (
    .A1(_02888_),
    .A2(_02890_),
    .ZN(_02891_)
  );
  AND2_X1 _07847_ (
    .A1(reg_mtval[25]),
    .A2(_00926_),
    .ZN(_02892_)
  );
  INV_X1 _07848_ (
    .A(_02892_),
    .ZN(_02893_)
  );
  AND2_X1 _07849_ (
    .A1(reg_pmp_0_addr[25]),
    .A2(_01004_),
    .ZN(_02894_)
  );
  INV_X1 _07850_ (
    .A(_02894_),
    .ZN(_02895_)
  );
  AND2_X1 _07851_ (
    .A1(_02893_),
    .A2(_02895_),
    .ZN(_02896_)
  );
  AND2_X1 _07852_ (
    .A1(_02891_),
    .A2(_02896_),
    .ZN(_02897_)
  );
  AND2_X1 _07853_ (
    .A1(reg_dscratch0[25]),
    .A2(_00958_),
    .ZN(_02898_)
  );
  INV_X1 _07854_ (
    .A(_02898_),
    .ZN(_02899_)
  );
  AND2_X1 _07855_ (
    .A1(reg_pmp_1_addr[25]),
    .A2(_01008_),
    .ZN(_02900_)
  );
  INV_X1 _07856_ (
    .A(_02900_),
    .ZN(_02901_)
  );
  AND2_X1 _07857_ (
    .A1(_02899_),
    .A2(_02901_),
    .ZN(_02902_)
  );
  AND2_X1 _07858_ (
    .A1(reg_mcause[25]),
    .A2(_01001_),
    .ZN(_02903_)
  );
  INV_X1 _07859_ (
    .A(_02903_),
    .ZN(_02904_)
  );
  AND2_X1 _07860_ (
    .A1(reg_bp_0_address[25]),
    .A2(_00962_),
    .ZN(_02905_)
  );
  INV_X1 _07861_ (
    .A(_02905_),
    .ZN(_02906_)
  );
  AND2_X1 _07862_ (
    .A1(_02904_),
    .A2(_02906_),
    .ZN(_02907_)
  );
  AND2_X1 _07863_ (
    .A1(_02902_),
    .A2(_02907_),
    .ZN(_02908_)
  );
  AND2_X1 _07864_ (
    .A1(_02897_),
    .A2(_02908_),
    .ZN(_02909_)
  );
  AND2_X1 _07865_ (
    .A1(_02886_),
    .A2(_02909_),
    .ZN(_02910_)
  );
  AND2_X1 _07866_ (
    .A1(reg_pmp_6_addr[25]),
    .A2(_00978_),
    .ZN(_02911_)
  );
  INV_X1 _07867_ (
    .A(_02911_),
    .ZN(_02912_)
  );
  AND2_X1 _07868_ (
    .A1(large_[19]),
    .A2(_00985_),
    .ZN(_02913_)
  );
  INV_X1 _07869_ (
    .A(_02913_),
    .ZN(_02914_)
  );
  AND2_X1 _07870_ (
    .A1(_02912_),
    .A2(_02914_),
    .ZN(_02915_)
  );
  AND2_X1 _07871_ (
    .A1(reg_pmp_7_addr[25]),
    .A2(_01016_),
    .ZN(_02916_)
  );
  INV_X1 _07872_ (
    .A(_02916_),
    .ZN(_02917_)
  );
  AND2_X1 _07873_ (
    .A1(large_1[51]),
    .A2(_01019_),
    .ZN(_02918_)
  );
  INV_X1 _07874_ (
    .A(_02918_),
    .ZN(_02919_)
  );
  AND2_X1 _07875_ (
    .A1(_02917_),
    .A2(_02919_),
    .ZN(_02920_)
  );
  AND2_X1 _07876_ (
    .A1(_02915_),
    .A2(_02920_),
    .ZN(_02921_)
  );
  AND2_X1 _07877_ (
    .A1(reg_mscratch[25]),
    .A2(_00929_),
    .ZN(_02922_)
  );
  INV_X1 _07878_ (
    .A(_02922_),
    .ZN(_02923_)
  );
  AND2_X1 _07879_ (
    .A1(reg_pmp_2_addr[25]),
    .A2(_00953_),
    .ZN(_02924_)
  );
  INV_X1 _07880_ (
    .A(_02924_),
    .ZN(_02925_)
  );
  AND2_X1 _07881_ (
    .A1(_02923_),
    .A2(_02925_),
    .ZN(_02926_)
  );
  AND2_X1 _07882_ (
    .A1(reg_dpc[25]),
    .A2(_00912_),
    .ZN(_02927_)
  );
  INV_X1 _07883_ (
    .A(_02927_),
    .ZN(_02928_)
  );
  AND2_X1 _07884_ (
    .A1(reg_pmp_3_cfg_w),
    .A2(_00916_),
    .ZN(_02929_)
  );
  INV_X1 _07885_ (
    .A(_02929_),
    .ZN(_02930_)
  );
  AND2_X1 _07886_ (
    .A1(_02928_),
    .A2(_02930_),
    .ZN(_02931_)
  );
  AND2_X1 _07887_ (
    .A1(_02926_),
    .A2(_02931_),
    .ZN(_02932_)
  );
  AND2_X1 _07888_ (
    .A1(large_[51]),
    .A2(_00991_),
    .ZN(_02933_)
  );
  INV_X1 _07889_ (
    .A(_02933_),
    .ZN(_02934_)
  );
  AND2_X1 _07890_ (
    .A1(large_1[19]),
    .A2(_00995_),
    .ZN(_02935_)
  );
  INV_X1 _07891_ (
    .A(_02935_),
    .ZN(_02936_)
  );
  AND2_X1 _07892_ (
    .A1(_02934_),
    .A2(_02936_),
    .ZN(_02937_)
  );
  AND2_X1 _07893_ (
    .A1(_02932_),
    .A2(_02937_),
    .ZN(_02938_)
  );
  AND2_X1 _07894_ (
    .A1(_02921_),
    .A2(_02938_),
    .ZN(_02939_)
  );
  AND2_X1 _07895_ (
    .A1(_02910_),
    .A2(_02939_),
    .ZN(_02940_)
  );
  INV_X1 _07896_ (
    .A(_02940_),
    .ZN(io_rw_rdata[25])
  );
  AND2_X1 _07897_ (
    .A1(io_rw_cmd[1]),
    .A2(_00860_),
    .ZN(_02941_)
  );
  AND2_X1 _07898_ (
    .A1(io_rw_rdata[25]),
    .A2(_02941_),
    .ZN(_02942_)
  );
  INV_X1 _07899_ (
    .A(_02942_),
    .ZN(_02943_)
  );
  AND2_X1 _07900_ (
    .A1(_02875_),
    .A2(_02943_),
    .ZN(_02944_)
  );
  INV_X1 _07901_ (
    .A(_02944_),
    .ZN(_02945_)
  );
  MUX2_X1 _07902_ (
    .A(reg_pmp_5_addr[25]),
    .B(_02945_),
    .S(_01525_),
    .Z(_00052_)
  );
  AND2_X1 _07903_ (
    .A1(io_rw_wdata[26]),
    .A2(_00903_),
    .ZN(_02946_)
  );
  INV_X1 _07904_ (
    .A(_02946_),
    .ZN(_02947_)
  );
  AND2_X1 _07905_ (
    .A1(reg_pmp_3_addr[26]),
    .A2(_01011_),
    .ZN(_02948_)
  );
  INV_X1 _07906_ (
    .A(_02948_),
    .ZN(_02949_)
  );
  AND2_X1 _07907_ (
    .A1(reg_mtval[26]),
    .A2(_00926_),
    .ZN(_02950_)
  );
  INV_X1 _07908_ (
    .A(_02950_),
    .ZN(_02951_)
  );
  AND2_X1 _07909_ (
    .A1(_02949_),
    .A2(_02951_),
    .ZN(_02952_)
  );
  AND2_X1 _07910_ (
    .A1(reg_pmp_1_addr[26]),
    .A2(_01008_),
    .ZN(_02953_)
  );
  INV_X1 _07911_ (
    .A(_02953_),
    .ZN(_02954_)
  );
  AND2_X1 _07912_ (
    .A1(reg_pmp_7_cfg_x),
    .A2(_00894_),
    .ZN(_02955_)
  );
  INV_X1 _07913_ (
    .A(_02955_),
    .ZN(_02956_)
  );
  AND2_X1 _07914_ (
    .A1(_02954_),
    .A2(_02956_),
    .ZN(_02957_)
  );
  AND2_X1 _07915_ (
    .A1(_02952_),
    .A2(_02957_),
    .ZN(_02958_)
  );
  AND2_X1 _07916_ (
    .A1(reg_mscratch[26]),
    .A2(_00929_),
    .ZN(_02959_)
  );
  INV_X1 _07917_ (
    .A(_02959_),
    .ZN(_02960_)
  );
  AND2_X1 _07918_ (
    .A1(reg_pmp_2_addr[26]),
    .A2(_00953_),
    .ZN(_02961_)
  );
  INV_X1 _07919_ (
    .A(_02961_),
    .ZN(_02962_)
  );
  AND2_X1 _07920_ (
    .A1(_02960_),
    .A2(_02962_),
    .ZN(_02963_)
  );
  AND2_X1 _07921_ (
    .A1(reg_pmp_3_cfg_x),
    .A2(_00916_),
    .ZN(_02964_)
  );
  INV_X1 _07922_ (
    .A(_02964_),
    .ZN(_02965_)
  );
  AND2_X1 _07923_ (
    .A1(reg_mtvec[26]),
    .A2(_00940_),
    .ZN(_02966_)
  );
  INV_X1 _07924_ (
    .A(_02966_),
    .ZN(_02967_)
  );
  AND2_X1 _07925_ (
    .A1(_02965_),
    .A2(_02967_),
    .ZN(_02968_)
  );
  AND2_X1 _07926_ (
    .A1(_02963_),
    .A2(_02968_),
    .ZN(_02969_)
  );
  AND2_X1 _07927_ (
    .A1(reg_pmp_4_addr[26]),
    .A2(_00968_),
    .ZN(_02970_)
  );
  INV_X1 _07928_ (
    .A(_02970_),
    .ZN(_02971_)
  );
  AND2_X1 _07929_ (
    .A1(reg_pmp_0_addr[26]),
    .A2(_01004_),
    .ZN(_02972_)
  );
  INV_X1 _07930_ (
    .A(_02972_),
    .ZN(_02973_)
  );
  AND2_X1 _07931_ (
    .A1(_02971_),
    .A2(_02973_),
    .ZN(_02974_)
  );
  AND2_X1 _07932_ (
    .A1(reg_bp_0_address[26]),
    .A2(_00962_),
    .ZN(_02975_)
  );
  INV_X1 _07933_ (
    .A(_02975_),
    .ZN(_02976_)
  );
  AND2_X1 _07934_ (
    .A1(reg_mepc[26]),
    .A2(_00943_),
    .ZN(_02977_)
  );
  INV_X1 _07935_ (
    .A(_02977_),
    .ZN(_02978_)
  );
  AND2_X1 _07936_ (
    .A1(_02976_),
    .A2(_02978_),
    .ZN(_02979_)
  );
  AND2_X1 _07937_ (
    .A1(_02974_),
    .A2(_02979_),
    .ZN(_02980_)
  );
  AND2_X1 _07938_ (
    .A1(_02969_),
    .A2(_02980_),
    .ZN(_02981_)
  );
  AND2_X1 _07939_ (
    .A1(_02958_),
    .A2(_02981_),
    .ZN(_02982_)
  );
  AND2_X1 _07940_ (
    .A1(large_1[52]),
    .A2(_01019_),
    .ZN(_02983_)
  );
  INV_X1 _07941_ (
    .A(_02983_),
    .ZN(_02984_)
  );
  AND2_X1 _07942_ (
    .A1(large_1[20]),
    .A2(_00995_),
    .ZN(_02985_)
  );
  INV_X1 _07943_ (
    .A(_02985_),
    .ZN(_02986_)
  );
  AND2_X1 _07944_ (
    .A1(_02984_),
    .A2(_02986_),
    .ZN(_02987_)
  );
  AND2_X1 _07945_ (
    .A1(large_[52]),
    .A2(_00991_),
    .ZN(_02988_)
  );
  INV_X1 _07946_ (
    .A(_02988_),
    .ZN(_02989_)
  );
  AND2_X1 _07947_ (
    .A1(large_[20]),
    .A2(_00985_),
    .ZN(_02990_)
  );
  INV_X1 _07948_ (
    .A(_02990_),
    .ZN(_02991_)
  );
  AND2_X1 _07949_ (
    .A1(_02989_),
    .A2(_02991_),
    .ZN(_02992_)
  );
  AND2_X1 _07950_ (
    .A1(_02987_),
    .A2(_02992_),
    .ZN(_02993_)
  );
  AND2_X1 _07951_ (
    .A1(reg_mcause[26]),
    .A2(_01001_),
    .ZN(_02994_)
  );
  INV_X1 _07952_ (
    .A(_02994_),
    .ZN(_02995_)
  );
  AND2_X1 _07953_ (
    .A1(reg_dscratch0[26]),
    .A2(_00958_),
    .ZN(_02996_)
  );
  INV_X1 _07954_ (
    .A(_02996_),
    .ZN(_02997_)
  );
  AND2_X1 _07955_ (
    .A1(_02995_),
    .A2(_02997_),
    .ZN(_02998_)
  );
  AND2_X1 _07956_ (
    .A1(reg_pmp_5_addr[26]),
    .A2(_00948_),
    .ZN(_02999_)
  );
  INV_X1 _07957_ (
    .A(_02999_),
    .ZN(_03000_)
  );
  AND2_X1 _07958_ (
    .A1(reg_dpc[26]),
    .A2(_00912_),
    .ZN(_03001_)
  );
  INV_X1 _07959_ (
    .A(_03001_),
    .ZN(_03002_)
  );
  AND2_X1 _07960_ (
    .A1(_03000_),
    .A2(_03002_),
    .ZN(_03003_)
  );
  AND2_X1 _07961_ (
    .A1(_02998_),
    .A2(_03003_),
    .ZN(_03004_)
  );
  AND2_X1 _07962_ (
    .A1(reg_pmp_6_addr[26]),
    .A2(_00978_),
    .ZN(_03005_)
  );
  INV_X1 _07963_ (
    .A(_03005_),
    .ZN(_03006_)
  );
  AND2_X1 _07964_ (
    .A1(reg_pmp_7_addr[26]),
    .A2(_01016_),
    .ZN(_03007_)
  );
  INV_X1 _07965_ (
    .A(_03007_),
    .ZN(_03008_)
  );
  AND2_X1 _07966_ (
    .A1(_03006_),
    .A2(_03008_),
    .ZN(_03009_)
  );
  AND2_X1 _07967_ (
    .A1(_03004_),
    .A2(_03009_),
    .ZN(_03010_)
  );
  AND2_X1 _07968_ (
    .A1(_02993_),
    .A2(_03010_),
    .ZN(_03011_)
  );
  AND2_X1 _07969_ (
    .A1(_02982_),
    .A2(_03011_),
    .ZN(_03012_)
  );
  INV_X1 _07970_ (
    .A(_03012_),
    .ZN(io_rw_rdata[26])
  );
  AND2_X1 _07971_ (
    .A1(io_rw_cmd[1]),
    .A2(_00861_),
    .ZN(_03013_)
  );
  AND2_X1 _07972_ (
    .A1(io_rw_rdata[26]),
    .A2(_03013_),
    .ZN(_03014_)
  );
  INV_X1 _07973_ (
    .A(_03014_),
    .ZN(_03015_)
  );
  AND2_X1 _07974_ (
    .A1(_02947_),
    .A2(_03015_),
    .ZN(_03016_)
  );
  INV_X1 _07975_ (
    .A(_03016_),
    .ZN(_03017_)
  );
  MUX2_X1 _07976_ (
    .A(reg_pmp_5_addr[26]),
    .B(_03017_),
    .S(_01525_),
    .Z(_00053_)
  );
  AND2_X1 _07977_ (
    .A1(reg_bp_0_control_dmode),
    .A2(_01341_),
    .ZN(_03018_)
  );
  INV_X1 _07978_ (
    .A(_03018_),
    .ZN(_03019_)
  );
  AND2_X1 _07979_ (
    .A1(reg_bp_0_address[27]),
    .A2(_00962_),
    .ZN(_03020_)
  );
  INV_X1 _07980_ (
    .A(_03020_),
    .ZN(_03021_)
  );
  AND2_X1 _07981_ (
    .A1(_03019_),
    .A2(_03021_),
    .ZN(_03022_)
  );
  AND2_X1 _07982_ (
    .A1(reg_pmp_3_cfg_a[0]),
    .A2(_00916_),
    .ZN(_03023_)
  );
  INV_X1 _07983_ (
    .A(_03023_),
    .ZN(_03024_)
  );
  AND2_X1 _07984_ (
    .A1(reg_mtval[27]),
    .A2(_00926_),
    .ZN(_03025_)
  );
  INV_X1 _07985_ (
    .A(_03025_),
    .ZN(_03026_)
  );
  AND2_X1 _07986_ (
    .A1(_03024_),
    .A2(_03026_),
    .ZN(_03027_)
  );
  AND2_X1 _07987_ (
    .A1(_03022_),
    .A2(_03027_),
    .ZN(_03028_)
  );
  AND2_X1 _07988_ (
    .A1(reg_dpc[27]),
    .A2(_00912_),
    .ZN(_03029_)
  );
  INV_X1 _07989_ (
    .A(_03029_),
    .ZN(_03030_)
  );
  AND2_X1 _07990_ (
    .A1(reg_pmp_4_addr[27]),
    .A2(_00968_),
    .ZN(_03031_)
  );
  INV_X1 _07991_ (
    .A(_03031_),
    .ZN(_03032_)
  );
  AND2_X1 _07992_ (
    .A1(_03030_),
    .A2(_03032_),
    .ZN(_03033_)
  );
  AND2_X1 _07993_ (
    .A1(reg_pmp_5_addr[27]),
    .A2(_00948_),
    .ZN(_03034_)
  );
  INV_X1 _07994_ (
    .A(_03034_),
    .ZN(_03035_)
  );
  AND2_X1 _07995_ (
    .A1(reg_pmp_0_addr[27]),
    .A2(_01004_),
    .ZN(_03036_)
  );
  INV_X1 _07996_ (
    .A(_03036_),
    .ZN(_03037_)
  );
  AND2_X1 _07997_ (
    .A1(_03035_),
    .A2(_03037_),
    .ZN(_03038_)
  );
  AND2_X1 _07998_ (
    .A1(_03033_),
    .A2(_03038_),
    .ZN(_03039_)
  );
  AND2_X1 _07999_ (
    .A1(_03028_),
    .A2(_03039_),
    .ZN(_03040_)
  );
  AND2_X1 _08000_ (
    .A1(reg_pmp_3_addr[27]),
    .A2(_01011_),
    .ZN(_03041_)
  );
  INV_X1 _08001_ (
    .A(_03041_),
    .ZN(_03042_)
  );
  AND2_X1 _08002_ (
    .A1(reg_pmp_1_addr[27]),
    .A2(_01008_),
    .ZN(_03043_)
  );
  INV_X1 _08003_ (
    .A(_03043_),
    .ZN(_03044_)
  );
  AND2_X1 _08004_ (
    .A1(reg_mepc[27]),
    .A2(_00943_),
    .ZN(_03045_)
  );
  INV_X1 _08005_ (
    .A(_03045_),
    .ZN(_03046_)
  );
  AND2_X1 _08006_ (
    .A1(_03044_),
    .A2(_03046_),
    .ZN(_03047_)
  );
  AND2_X1 _08007_ (
    .A1(_03042_),
    .A2(_03047_),
    .ZN(_03048_)
  );
  AND2_X1 _08008_ (
    .A1(reg_mtvec[27]),
    .A2(_00940_),
    .ZN(_03049_)
  );
  INV_X1 _08009_ (
    .A(_03049_),
    .ZN(_03050_)
  );
  AND2_X1 _08010_ (
    .A1(reg_mscratch[27]),
    .A2(_00929_),
    .ZN(_03051_)
  );
  INV_X1 _08011_ (
    .A(_03051_),
    .ZN(_03052_)
  );
  AND2_X1 _08012_ (
    .A1(_03050_),
    .A2(_03052_),
    .ZN(_03053_)
  );
  AND2_X1 _08013_ (
    .A1(reg_pmp_2_addr[27]),
    .A2(_00953_),
    .ZN(_03054_)
  );
  INV_X1 _08014_ (
    .A(_03054_),
    .ZN(_03055_)
  );
  AND2_X1 _08015_ (
    .A1(reg_mcause[27]),
    .A2(_01001_),
    .ZN(_03056_)
  );
  INV_X1 _08016_ (
    .A(_03056_),
    .ZN(_03057_)
  );
  AND2_X1 _08017_ (
    .A1(_03055_),
    .A2(_03057_),
    .ZN(_03058_)
  );
  AND2_X1 _08018_ (
    .A1(_03053_),
    .A2(_03058_),
    .ZN(_03059_)
  );
  AND2_X1 _08019_ (
    .A1(_03048_),
    .A2(_03059_),
    .ZN(_03060_)
  );
  AND2_X1 _08020_ (
    .A1(_03040_),
    .A2(_03060_),
    .ZN(_03061_)
  );
  AND2_X1 _08021_ (
    .A1(large_1[21]),
    .A2(_00995_),
    .ZN(_03062_)
  );
  INV_X1 _08022_ (
    .A(_03062_),
    .ZN(_03063_)
  );
  AND2_X1 _08023_ (
    .A1(large_[53]),
    .A2(_00991_),
    .ZN(_03064_)
  );
  INV_X1 _08024_ (
    .A(_03064_),
    .ZN(_03065_)
  );
  AND2_X1 _08025_ (
    .A1(large_1[53]),
    .A2(_01019_),
    .ZN(_03066_)
  );
  INV_X1 _08026_ (
    .A(_03066_),
    .ZN(_03067_)
  );
  AND2_X1 _08027_ (
    .A1(_03065_),
    .A2(_03067_),
    .ZN(_03068_)
  );
  AND2_X1 _08028_ (
    .A1(_03063_),
    .A2(_03068_),
    .ZN(_03069_)
  );
  AND2_X1 _08029_ (
    .A1(large_[21]),
    .A2(_00985_),
    .ZN(_03070_)
  );
  INV_X1 _08030_ (
    .A(_03070_),
    .ZN(_03071_)
  );
  AND2_X1 _08031_ (
    .A1(reg_dscratch0[27]),
    .A2(_00958_),
    .ZN(_03072_)
  );
  INV_X1 _08032_ (
    .A(_03072_),
    .ZN(_03073_)
  );
  AND2_X1 _08033_ (
    .A1(reg_pmp_7_cfg_a[0]),
    .A2(_00894_),
    .ZN(_03074_)
  );
  INV_X1 _08034_ (
    .A(_03074_),
    .ZN(_03075_)
  );
  AND2_X1 _08035_ (
    .A1(_03073_),
    .A2(_03075_),
    .ZN(_03076_)
  );
  AND2_X1 _08036_ (
    .A1(_03071_),
    .A2(_03076_),
    .ZN(_03077_)
  );
  AND2_X1 _08037_ (
    .A1(reg_pmp_7_addr[27]),
    .A2(_01016_),
    .ZN(_03078_)
  );
  INV_X1 _08038_ (
    .A(_03078_),
    .ZN(_03079_)
  );
  AND2_X1 _08039_ (
    .A1(reg_pmp_6_addr[27]),
    .A2(_00978_),
    .ZN(_03080_)
  );
  INV_X1 _08040_ (
    .A(_03080_),
    .ZN(_03081_)
  );
  AND2_X1 _08041_ (
    .A1(_03079_),
    .A2(_03081_),
    .ZN(_03082_)
  );
  AND2_X1 _08042_ (
    .A1(_03077_),
    .A2(_03082_),
    .ZN(_03083_)
  );
  AND2_X1 _08043_ (
    .A1(_03069_),
    .A2(_03083_),
    .ZN(_03084_)
  );
  AND2_X1 _08044_ (
    .A1(_03061_),
    .A2(_03084_),
    .ZN(_03085_)
  );
  INV_X1 _08045_ (
    .A(_03085_),
    .ZN(io_rw_rdata[27])
  );
  AND2_X1 _08046_ (
    .A1(io_rw_cmd[1]),
    .A2(io_rw_rdata[27]),
    .ZN(_03086_)
  );
  AND2_X1 _08047_ (
    .A1(io_rw_wdata[27]),
    .A2(_00902_),
    .ZN(_03087_)
  );
  INV_X1 _08048_ (
    .A(_03087_),
    .ZN(_03088_)
  );
  MUX2_X1 _08049_ (
    .A(_00903_),
    .B(_03086_),
    .S(_00862_),
    .Z(_03089_)
  );
  INV_X1 _08050_ (
    .A(_03089_),
    .ZN(_03090_)
  );
  MUX2_X1 _08051_ (
    .A(reg_pmp_5_addr[27]),
    .B(_03089_),
    .S(_01525_),
    .Z(_00054_)
  );
  AND2_X1 _08052_ (
    .A1(io_rw_wdata[28]),
    .A2(_00903_),
    .ZN(_03091_)
  );
  INV_X1 _08053_ (
    .A(_03091_),
    .ZN(_03092_)
  );
  AND2_X1 _08054_ (
    .A1(reg_dscratch0[28]),
    .A2(_00958_),
    .ZN(_03093_)
  );
  INV_X1 _08055_ (
    .A(_03093_),
    .ZN(_03094_)
  );
  AND2_X1 _08056_ (
    .A1(reg_mtval[28]),
    .A2(_00926_),
    .ZN(_03095_)
  );
  INV_X1 _08057_ (
    .A(_03095_),
    .ZN(_03096_)
  );
  AND2_X1 _08058_ (
    .A1(reg_mtvec[28]),
    .A2(_00940_),
    .ZN(_03097_)
  );
  INV_X1 _08059_ (
    .A(_03097_),
    .ZN(_03098_)
  );
  AND2_X1 _08060_ (
    .A1(reg_pmp_2_addr[28]),
    .A2(_00953_),
    .ZN(_03099_)
  );
  INV_X1 _08061_ (
    .A(_03099_),
    .ZN(_03100_)
  );
  AND2_X1 _08062_ (
    .A1(reg_pmp_7_cfg_a[1]),
    .A2(_00894_),
    .ZN(_03101_)
  );
  INV_X1 _08063_ (
    .A(_03101_),
    .ZN(_03102_)
  );
  AND2_X1 _08064_ (
    .A1(reg_pmp_3_addr[28]),
    .A2(_01011_),
    .ZN(_03103_)
  );
  INV_X1 _08065_ (
    .A(_03103_),
    .ZN(_03104_)
  );
  AND2_X1 _08066_ (
    .A1(reg_dpc[28]),
    .A2(_00912_),
    .ZN(_03105_)
  );
  INV_X1 _08067_ (
    .A(_03105_),
    .ZN(_03106_)
  );
  AND2_X1 _08068_ (
    .A1(reg_pmp_3_cfg_a[1]),
    .A2(_00916_),
    .ZN(_03107_)
  );
  INV_X1 _08069_ (
    .A(_03107_),
    .ZN(_03108_)
  );
  AND2_X1 _08070_ (
    .A1(reg_mepc[28]),
    .A2(_00943_),
    .ZN(_03109_)
  );
  INV_X1 _08071_ (
    .A(_03109_),
    .ZN(_03110_)
  );
  AND2_X1 _08072_ (
    .A1(reg_mscratch[28]),
    .A2(_00929_),
    .ZN(_03111_)
  );
  INV_X1 _08073_ (
    .A(_03111_),
    .ZN(_03112_)
  );
  AND2_X1 _08074_ (
    .A1(_03110_),
    .A2(_03112_),
    .ZN(_03113_)
  );
  AND2_X1 _08075_ (
    .A1(reg_pmp_4_addr[28]),
    .A2(_00968_),
    .ZN(_03114_)
  );
  INV_X1 _08076_ (
    .A(_03114_),
    .ZN(_03115_)
  );
  AND2_X1 _08077_ (
    .A1(reg_bp_0_address[28]),
    .A2(_00962_),
    .ZN(_03116_)
  );
  INV_X1 _08078_ (
    .A(_03116_),
    .ZN(_03117_)
  );
  AND2_X1 _08079_ (
    .A1(large_1[54]),
    .A2(_01019_),
    .ZN(_03118_)
  );
  INV_X1 _08080_ (
    .A(_03118_),
    .ZN(_03119_)
  );
  AND2_X1 _08081_ (
    .A1(large_[54]),
    .A2(_00991_),
    .ZN(_03120_)
  );
  INV_X1 _08082_ (
    .A(_03120_),
    .ZN(_03121_)
  );
  AND2_X1 _08083_ (
    .A1(reg_pmp_5_addr[28]),
    .A2(_00948_),
    .ZN(_03122_)
  );
  INV_X1 _08084_ (
    .A(_03122_),
    .ZN(_03123_)
  );
  AND2_X1 _08085_ (
    .A1(reg_mcause[28]),
    .A2(_01001_),
    .ZN(_03124_)
  );
  INV_X1 _08086_ (
    .A(_03124_),
    .ZN(_03125_)
  );
  AND2_X1 _08087_ (
    .A1(reg_pmp_1_addr[28]),
    .A2(_01008_),
    .ZN(_03126_)
  );
  INV_X1 _08088_ (
    .A(_03126_),
    .ZN(_03127_)
  );
  AND2_X1 _08089_ (
    .A1(reg_pmp_0_addr[28]),
    .A2(_01004_),
    .ZN(_03128_)
  );
  INV_X1 _08090_ (
    .A(_03128_),
    .ZN(_03129_)
  );
  AND2_X1 _08091_ (
    .A1(reg_pmp_7_addr[28]),
    .A2(_01016_),
    .ZN(_03130_)
  );
  INV_X1 _08092_ (
    .A(_03130_),
    .ZN(_03131_)
  );
  AND2_X1 _08093_ (
    .A1(reg_pmp_6_addr[28]),
    .A2(_00978_),
    .ZN(_03132_)
  );
  INV_X1 _08094_ (
    .A(_03132_),
    .ZN(_03133_)
  );
  AND2_X1 _08095_ (
    .A1(_03100_),
    .A2(_03104_),
    .ZN(_03134_)
  );
  AND2_X1 _08096_ (
    .A1(_03121_),
    .A2(_03134_),
    .ZN(_03135_)
  );
  AND2_X1 _08097_ (
    .A1(_03096_),
    .A2(_03098_),
    .ZN(_03136_)
  );
  AND2_X1 _08098_ (
    .A1(_03125_),
    .A2(_03129_),
    .ZN(_03137_)
  );
  AND2_X1 _08099_ (
    .A1(_03136_),
    .A2(_03137_),
    .ZN(_03138_)
  );
  AND2_X1 _08100_ (
    .A1(_03135_),
    .A2(_03138_),
    .ZN(_03139_)
  );
  AND2_X1 _08101_ (
    .A1(_03102_),
    .A2(_03108_),
    .ZN(_03140_)
  );
  AND2_X1 _08102_ (
    .A1(_03133_),
    .A2(_03140_),
    .ZN(_03141_)
  );
  AND2_X1 _08103_ (
    .A1(large_1[22]),
    .A2(_01029_),
    .ZN(_03142_)
  );
  INV_X1 _08104_ (
    .A(_03142_),
    .ZN(_03143_)
  );
  AND2_X1 _08105_ (
    .A1(_03115_),
    .A2(_03143_),
    .ZN(_03144_)
  );
  AND2_X1 _08106_ (
    .A1(large_[22]),
    .A2(_01027_),
    .ZN(_03145_)
  );
  INV_X1 _08107_ (
    .A(_03145_),
    .ZN(_03146_)
  );
  AND2_X1 _08108_ (
    .A1(_03123_),
    .A2(_03146_),
    .ZN(_03147_)
  );
  AND2_X1 _08109_ (
    .A1(_03144_),
    .A2(_03147_),
    .ZN(_03148_)
  );
  AND2_X1 _08110_ (
    .A1(_03141_),
    .A2(_03148_),
    .ZN(_03149_)
  );
  AND2_X1 _08111_ (
    .A1(_03139_),
    .A2(_03149_),
    .ZN(_03150_)
  );
  AND2_X1 _08112_ (
    .A1(_03113_),
    .A2(_03127_),
    .ZN(_03151_)
  );
  AND2_X1 _08113_ (
    .A1(_03119_),
    .A2(_03151_),
    .ZN(_03152_)
  );
  AND2_X1 _08114_ (
    .A1(_03106_),
    .A2(_03117_),
    .ZN(_03153_)
  );
  AND2_X1 _08115_ (
    .A1(_03131_),
    .A2(_03153_),
    .ZN(_03154_)
  );
  AND2_X1 _08116_ (
    .A1(_03094_),
    .A2(_03154_),
    .ZN(_03155_)
  );
  AND2_X1 _08117_ (
    .A1(_03152_),
    .A2(_03155_),
    .ZN(_03156_)
  );
  AND2_X1 _08118_ (
    .A1(_03150_),
    .A2(_03156_),
    .ZN(_03157_)
  );
  INV_X1 _08119_ (
    .A(_03157_),
    .ZN(io_rw_rdata[28])
  );
  AND2_X1 _08120_ (
    .A1(io_rw_cmd[1]),
    .A2(_00863_),
    .ZN(_03158_)
  );
  AND2_X1 _08121_ (
    .A1(io_rw_rdata[28]),
    .A2(_03158_),
    .ZN(_03159_)
  );
  INV_X1 _08122_ (
    .A(_03159_),
    .ZN(_03160_)
  );
  AND2_X1 _08123_ (
    .A1(_03092_),
    .A2(_03160_),
    .ZN(_03161_)
  );
  INV_X1 _08124_ (
    .A(_03161_),
    .ZN(_03162_)
  );
  MUX2_X1 _08125_ (
    .A(reg_pmp_5_addr[28]),
    .B(_03162_),
    .S(_01525_),
    .Z(_00055_)
  );
  AND2_X1 _08126_ (
    .A1(io_rw_wdata[29]),
    .A2(_00903_),
    .ZN(_03163_)
  );
  INV_X1 _08127_ (
    .A(_03163_),
    .ZN(_03164_)
  );
  AND2_X1 _08128_ (
    .A1(reg_pmp_1_addr[29]),
    .A2(_01008_),
    .ZN(_03165_)
  );
  INV_X1 _08129_ (
    .A(_03165_),
    .ZN(_03166_)
  );
  AND2_X1 _08130_ (
    .A1(reg_pmp_3_addr[29]),
    .A2(_01011_),
    .ZN(_03167_)
  );
  INV_X1 _08131_ (
    .A(_03167_),
    .ZN(_03168_)
  );
  AND2_X1 _08132_ (
    .A1(_03166_),
    .A2(_03168_),
    .ZN(_03169_)
  );
  AND2_X1 _08133_ (
    .A1(reg_mtvec[29]),
    .A2(_00940_),
    .ZN(_03170_)
  );
  INV_X1 _08134_ (
    .A(_03170_),
    .ZN(_03171_)
  );
  AND2_X1 _08135_ (
    .A1(reg_pmp_2_addr[29]),
    .A2(_00953_),
    .ZN(_03172_)
  );
  INV_X1 _08136_ (
    .A(_03172_),
    .ZN(_03173_)
  );
  AND2_X1 _08137_ (
    .A1(_03171_),
    .A2(_03173_),
    .ZN(_03174_)
  );
  AND2_X1 _08138_ (
    .A1(_03169_),
    .A2(_03174_),
    .ZN(_03175_)
  );
  AND2_X1 _08139_ (
    .A1(reg_mscratch[29]),
    .A2(_00929_),
    .ZN(_03176_)
  );
  INV_X1 _08140_ (
    .A(_03176_),
    .ZN(_03177_)
  );
  AND2_X1 _08141_ (
    .A1(reg_mepc[29]),
    .A2(_00943_),
    .ZN(_03178_)
  );
  INV_X1 _08142_ (
    .A(_03178_),
    .ZN(_03179_)
  );
  AND2_X1 _08143_ (
    .A1(_03177_),
    .A2(_03179_),
    .ZN(_03180_)
  );
  AND2_X1 _08144_ (
    .A1(reg_pmp_0_addr[29]),
    .A2(_01004_),
    .ZN(_03181_)
  );
  INV_X1 _08145_ (
    .A(_03181_),
    .ZN(_03182_)
  );
  AND2_X1 _08146_ (
    .A1(reg_pmp_4_addr[29]),
    .A2(_00968_),
    .ZN(_03183_)
  );
  INV_X1 _08147_ (
    .A(_03183_),
    .ZN(_03184_)
  );
  AND2_X1 _08148_ (
    .A1(_03182_),
    .A2(_03184_),
    .ZN(_03185_)
  );
  AND2_X1 _08149_ (
    .A1(_03180_),
    .A2(_03185_),
    .ZN(_03186_)
  );
  AND2_X1 _08150_ (
    .A1(reg_dscratch0[29]),
    .A2(_00958_),
    .ZN(_03187_)
  );
  INV_X1 _08151_ (
    .A(_03187_),
    .ZN(_03188_)
  );
  AND2_X1 _08152_ (
    .A1(reg_mtval[29]),
    .A2(_00926_),
    .ZN(_03189_)
  );
  INV_X1 _08153_ (
    .A(_03189_),
    .ZN(_03190_)
  );
  AND2_X1 _08154_ (
    .A1(_03188_),
    .A2(_03190_),
    .ZN(_03191_)
  );
  AND2_X1 _08155_ (
    .A1(reg_mcause[29]),
    .A2(_01001_),
    .ZN(_03192_)
  );
  INV_X1 _08156_ (
    .A(_03192_),
    .ZN(_03193_)
  );
  AND2_X1 _08157_ (
    .A1(reg_pmp_5_addr[29]),
    .A2(_00948_),
    .ZN(_03194_)
  );
  INV_X1 _08158_ (
    .A(_03194_),
    .ZN(_03195_)
  );
  AND2_X1 _08159_ (
    .A1(_03193_),
    .A2(_03195_),
    .ZN(_03196_)
  );
  AND2_X1 _08160_ (
    .A1(_03191_),
    .A2(_03196_),
    .ZN(_03197_)
  );
  AND2_X1 _08161_ (
    .A1(_03186_),
    .A2(_03197_),
    .ZN(_03198_)
  );
  AND2_X1 _08162_ (
    .A1(_03175_),
    .A2(_03198_),
    .ZN(_03199_)
  );
  AND2_X1 _08163_ (
    .A1(large_[55]),
    .A2(_00991_),
    .ZN(_03200_)
  );
  INV_X1 _08164_ (
    .A(_03200_),
    .ZN(_03201_)
  );
  AND2_X1 _08165_ (
    .A1(large_[23]),
    .A2(_00985_),
    .ZN(_03202_)
  );
  INV_X1 _08166_ (
    .A(_03202_),
    .ZN(_03203_)
  );
  AND2_X1 _08167_ (
    .A1(_03201_),
    .A2(_03203_),
    .ZN(_03204_)
  );
  AND2_X1 _08168_ (
    .A1(large_1[55]),
    .A2(_01019_),
    .ZN(_03205_)
  );
  INV_X1 _08169_ (
    .A(_03205_),
    .ZN(_03206_)
  );
  AND2_X1 _08170_ (
    .A1(large_1[23]),
    .A2(_00995_),
    .ZN(_03207_)
  );
  INV_X1 _08171_ (
    .A(_03207_),
    .ZN(_03208_)
  );
  AND2_X1 _08172_ (
    .A1(_03206_),
    .A2(_03208_),
    .ZN(_03209_)
  );
  AND2_X1 _08173_ (
    .A1(_03204_),
    .A2(_03209_),
    .ZN(_03210_)
  );
  AND2_X1 _08174_ (
    .A1(_01132_),
    .A2(_01342_),
    .ZN(_03211_)
  );
  AND2_X1 _08175_ (
    .A1(reg_dpc[29]),
    .A2(_00912_),
    .ZN(_03212_)
  );
  INV_X1 _08176_ (
    .A(_03212_),
    .ZN(_03213_)
  );
  AND2_X1 _08177_ (
    .A1(reg_bp_0_address[29]),
    .A2(_00962_),
    .ZN(_03214_)
  );
  INV_X1 _08178_ (
    .A(_03214_),
    .ZN(_03215_)
  );
  AND2_X1 _08179_ (
    .A1(_03213_),
    .A2(_03215_),
    .ZN(_03216_)
  );
  AND2_X1 _08180_ (
    .A1(_03211_),
    .A2(_03216_),
    .ZN(_03217_)
  );
  AND2_X1 _08181_ (
    .A1(reg_pmp_6_addr[29]),
    .A2(_00978_),
    .ZN(_03218_)
  );
  INV_X1 _08182_ (
    .A(_03218_),
    .ZN(_03219_)
  );
  AND2_X1 _08183_ (
    .A1(reg_pmp_7_addr[29]),
    .A2(_01016_),
    .ZN(_03220_)
  );
  INV_X1 _08184_ (
    .A(_03220_),
    .ZN(_03221_)
  );
  AND2_X1 _08185_ (
    .A1(_03219_),
    .A2(_03221_),
    .ZN(_03222_)
  );
  AND2_X1 _08186_ (
    .A1(_03217_),
    .A2(_03222_),
    .ZN(_03223_)
  );
  AND2_X1 _08187_ (
    .A1(_03210_),
    .A2(_03223_),
    .ZN(_03224_)
  );
  AND2_X1 _08188_ (
    .A1(_03199_),
    .A2(_03224_),
    .ZN(_03225_)
  );
  INV_X1 _08189_ (
    .A(_03225_),
    .ZN(io_rw_rdata[29])
  );
  AND2_X1 _08190_ (
    .A1(io_rw_cmd[1]),
    .A2(_00864_),
    .ZN(_03226_)
  );
  AND2_X1 _08191_ (
    .A1(io_rw_rdata[29]),
    .A2(_03226_),
    .ZN(_03227_)
  );
  INV_X1 _08192_ (
    .A(_03227_),
    .ZN(_03228_)
  );
  AND2_X1 _08193_ (
    .A1(_03164_),
    .A2(_03228_),
    .ZN(_03229_)
  );
  INV_X1 _08194_ (
    .A(_03229_),
    .ZN(_03230_)
  );
  MUX2_X1 _08195_ (
    .A(reg_pmp_5_addr[29]),
    .B(_03230_),
    .S(_01525_),
    .Z(_00056_)
  );
  AND2_X1 _08196_ (
    .A1(_00006_),
    .A2(_00916_),
    .ZN(_03231_)
  );
  AND2_X1 _08197_ (
    .A1(_00897_),
    .A2(_03231_),
    .ZN(_03232_)
  );
  INV_X1 _08198_ (
    .A(_03232_),
    .ZN(_03233_)
  );
  AND2_X1 _08199_ (
    .A1(_01613_),
    .A2(_01688_),
    .ZN(_03234_)
  );
  MUX2_X1 _08200_ (
    .A(reg_pmp_0_cfg_w),
    .B(_03234_),
    .S(_03232_),
    .Z(_00057_)
  );
  AND2_X1 _08201_ (
    .A1(_00807_),
    .A2(_01365_),
    .ZN(_03235_)
  );
  INV_X1 _08202_ (
    .A(_03235_),
    .ZN(_03236_)
  );
  AND2_X1 _08203_ (
    .A1(_00811_),
    .A2(_03236_),
    .ZN(_03237_)
  );
  AND2_X1 _08204_ (
    .A1(_01364_),
    .A2(_02313_),
    .ZN(_03238_)
  );
  INV_X1 _08205_ (
    .A(_03238_),
    .ZN(_03239_)
  );
  AND2_X1 _08206_ (
    .A1(_03237_),
    .A2(_03239_),
    .ZN(_00058_)
  );
  AND2_X1 _08207_ (
    .A1(_00806_),
    .A2(_01365_),
    .ZN(_03240_)
  );
  INV_X1 _08208_ (
    .A(_03240_),
    .ZN(_03241_)
  );
  AND2_X1 _08209_ (
    .A1(_00811_),
    .A2(_03241_),
    .ZN(_03242_)
  );
  AND2_X1 _08210_ (
    .A1(_01364_),
    .A2(_02390_),
    .ZN(_03243_)
  );
  INV_X1 _08211_ (
    .A(_03243_),
    .ZN(_03244_)
  );
  AND2_X1 _08212_ (
    .A1(_03242_),
    .A2(_03244_),
    .ZN(_00059_)
  );
  AND2_X1 _08213_ (
    .A1(_00805_),
    .A2(_01365_),
    .ZN(_03245_)
  );
  INV_X1 _08214_ (
    .A(_03245_),
    .ZN(_03246_)
  );
  AND2_X1 _08215_ (
    .A1(_00811_),
    .A2(_03246_),
    .ZN(_03247_)
  );
  AND2_X1 _08216_ (
    .A1(_01364_),
    .A2(_02596_),
    .ZN(_03248_)
  );
  INV_X1 _08217_ (
    .A(_03248_),
    .ZN(_03249_)
  );
  AND2_X1 _08218_ (
    .A1(_03247_),
    .A2(_03249_),
    .ZN(_00060_)
  );
  AND2_X1 _08219_ (
    .A1(reg_pmp_5_cfg_l),
    .A2(reg_pmp_5_cfg_a[0]),
    .ZN(_03250_)
  );
  AND2_X1 _08220_ (
    .A1(_00016_),
    .A2(_03250_),
    .ZN(_03251_)
  );
  INV_X1 _08221_ (
    .A(_03251_),
    .ZN(_03252_)
  );
  AND2_X1 _08222_ (
    .A1(_00802_),
    .A2(_03252_),
    .ZN(_03253_)
  );
  AND2_X1 _08223_ (
    .A1(_00897_),
    .A2(_03253_),
    .ZN(_03254_)
  );
  AND2_X1 _08224_ (
    .A1(_00968_),
    .A2(_03254_),
    .ZN(_03255_)
  );
  MUX2_X1 _08225_ (
    .A(reg_pmp_4_addr[0]),
    .B(_01613_),
    .S(_03255_),
    .Z(_00061_)
  );
  MUX2_X1 _08226_ (
    .A(reg_pmp_4_addr[1]),
    .B(_01688_),
    .S(_03255_),
    .Z(_00062_)
  );
  MUX2_X1 _08227_ (
    .A(reg_pmp_4_addr[2]),
    .B(_01774_),
    .S(_03255_),
    .Z(_00063_)
  );
  MUX2_X1 _08228_ (
    .A(reg_pmp_4_addr[3]),
    .B(_01865_),
    .S(_03255_),
    .Z(_00064_)
  );
  MUX2_X1 _08229_ (
    .A(reg_pmp_4_addr[4]),
    .B(_01938_),
    .S(_03255_),
    .Z(_00065_)
  );
  MUX2_X1 _08230_ (
    .A(reg_pmp_4_addr[5]),
    .B(_02005_),
    .S(_03255_),
    .Z(_00066_)
  );
  MUX2_X1 _08231_ (
    .A(reg_pmp_4_addr[6]),
    .B(_02076_),
    .S(_03255_),
    .Z(_00067_)
  );
  MUX2_X1 _08232_ (
    .A(reg_pmp_4_addr[7]),
    .B(_02163_),
    .S(_03255_),
    .Z(_00068_)
  );
  MUX2_X1 _08233_ (
    .A(reg_pmp_4_addr[8]),
    .B(_01446_),
    .S(_03255_),
    .Z(_00069_)
  );
  MUX2_X1 _08234_ (
    .A(reg_pmp_4_addr[9]),
    .B(_01518_),
    .S(_03255_),
    .Z(_00070_)
  );
  MUX2_X1 _08235_ (
    .A(reg_pmp_4_addr[10]),
    .B(_02235_),
    .S(_03255_),
    .Z(_00071_)
  );
  MUX2_X1 _08236_ (
    .A(reg_pmp_4_addr[11]),
    .B(_02314_),
    .S(_03255_),
    .Z(_00072_)
  );
  MUX2_X1 _08237_ (
    .A(reg_pmp_4_addr[12]),
    .B(_02389_),
    .S(_03255_),
    .Z(_00073_)
  );
  MUX2_X1 _08238_ (
    .A(reg_pmp_4_addr[13]),
    .B(_02456_),
    .S(_03255_),
    .Z(_00074_)
  );
  MUX2_X1 _08239_ (
    .A(reg_pmp_4_addr[14]),
    .B(_02522_),
    .S(_03255_),
    .Z(_00075_)
  );
  MUX2_X1 _08240_ (
    .A(reg_pmp_4_addr[15]),
    .B(_02597_),
    .S(_03255_),
    .Z(_00076_)
  );
  MUX2_X1 _08241_ (
    .A(reg_pmp_4_addr[16]),
    .B(_01035_),
    .S(_03255_),
    .Z(_00077_)
  );
  MUX2_X1 _08242_ (
    .A(reg_pmp_4_addr[17]),
    .B(_02669_),
    .S(_03255_),
    .Z(_00078_)
  );
  MUX2_X1 _08243_ (
    .A(reg_pmp_4_addr[18]),
    .B(_01107_),
    .S(_03255_),
    .Z(_00079_)
  );
  MUX2_X1 _08244_ (
    .A(reg_pmp_4_addr[19]),
    .B(_01199_),
    .S(_03255_),
    .Z(_00080_)
  );
  MUX2_X1 _08245_ (
    .A(reg_pmp_4_addr[20]),
    .B(_01277_),
    .S(_03255_),
    .Z(_00081_)
  );
  MUX2_X1 _08246_ (
    .A(reg_pmp_4_addr[21]),
    .B(_02735_),
    .S(_03255_),
    .Z(_00082_)
  );
  MUX2_X1 _08247_ (
    .A(reg_pmp_4_addr[22]),
    .B(_02801_),
    .S(_03255_),
    .Z(_00083_)
  );
  MUX2_X1 _08248_ (
    .A(reg_pmp_4_addr[23]),
    .B(_01360_),
    .S(_03255_),
    .Z(_00084_)
  );
  MUX2_X1 _08249_ (
    .A(reg_pmp_4_addr[24]),
    .B(_02873_),
    .S(_03255_),
    .Z(_00085_)
  );
  MUX2_X1 _08250_ (
    .A(reg_pmp_4_addr[25]),
    .B(_02945_),
    .S(_03255_),
    .Z(_00086_)
  );
  MUX2_X1 _08251_ (
    .A(reg_pmp_4_addr[26]),
    .B(_03017_),
    .S(_03255_),
    .Z(_00087_)
  );
  MUX2_X1 _08252_ (
    .A(reg_pmp_4_addr[27]),
    .B(_03089_),
    .S(_03255_),
    .Z(_00088_)
  );
  MUX2_X1 _08253_ (
    .A(reg_pmp_4_addr[28]),
    .B(_03162_),
    .S(_03255_),
    .Z(_00089_)
  );
  MUX2_X1 _08254_ (
    .A(reg_pmp_4_addr[29]),
    .B(_03230_),
    .S(_03255_),
    .Z(_00090_)
  );
  AND2_X1 _08255_ (
    .A1(_00013_),
    .A2(_00894_),
    .ZN(_03256_)
  );
  AND2_X1 _08256_ (
    .A1(_00897_),
    .A2(_03256_),
    .ZN(_03257_)
  );
  INV_X1 _08257_ (
    .A(_03257_),
    .ZN(_03258_)
  );
  MUX2_X1 _08258_ (
    .A(reg_pmp_4_cfg_w),
    .B(_03234_),
    .S(_03257_),
    .Z(_00091_)
  );
  MUX2_X1 _08259_ (
    .A(reg_pmp_4_cfg_x),
    .B(_01774_),
    .S(_03257_),
    .Z(_00092_)
  );
  AND2_X1 _08260_ (
    .A1(_00804_),
    .A2(_03258_),
    .ZN(_03259_)
  );
  INV_X1 _08261_ (
    .A(_03259_),
    .ZN(_03260_)
  );
  AND2_X1 _08262_ (
    .A1(_00811_),
    .A2(_03260_),
    .ZN(_03261_)
  );
  AND2_X1 _08263_ (
    .A1(_01864_),
    .A2(_03257_),
    .ZN(_03262_)
  );
  INV_X1 _08264_ (
    .A(_03262_),
    .ZN(_03263_)
  );
  AND2_X1 _08265_ (
    .A1(_03261_),
    .A2(_03263_),
    .ZN(_00093_)
  );
  AND2_X1 _08266_ (
    .A1(_00803_),
    .A2(_03258_),
    .ZN(_03264_)
  );
  INV_X1 _08267_ (
    .A(_03264_),
    .ZN(_03265_)
  );
  AND2_X1 _08268_ (
    .A1(_00811_),
    .A2(_03265_),
    .ZN(_03266_)
  );
  AND2_X1 _08269_ (
    .A1(_01937_),
    .A2(_03257_),
    .ZN(_03267_)
  );
  INV_X1 _08270_ (
    .A(_03267_),
    .ZN(_03268_)
  );
  AND2_X1 _08271_ (
    .A1(_03266_),
    .A2(_03268_),
    .ZN(_00094_)
  );
  AND2_X1 _08272_ (
    .A1(_00802_),
    .A2(_03258_),
    .ZN(_03269_)
  );
  INV_X1 _08273_ (
    .A(_03269_),
    .ZN(_03270_)
  );
  AND2_X1 _08274_ (
    .A1(_00811_),
    .A2(_03270_),
    .ZN(_03271_)
  );
  AND2_X1 _08275_ (
    .A1(_02162_),
    .A2(_03257_),
    .ZN(_03272_)
  );
  INV_X1 _08276_ (
    .A(_03272_),
    .ZN(_03273_)
  );
  AND2_X1 _08277_ (
    .A1(_03271_),
    .A2(_03273_),
    .ZN(_00095_)
  );
  AND2_X1 _08278_ (
    .A1(_00011_),
    .A2(_00916_),
    .ZN(_03274_)
  );
  AND2_X1 _08279_ (
    .A1(_00897_),
    .A2(_03274_),
    .ZN(_03275_)
  );
  INV_X1 _08280_ (
    .A(_03275_),
    .ZN(_03276_)
  );
  AND2_X1 _08281_ (
    .A1(_02873_),
    .A2(_02945_),
    .ZN(_03277_)
  );
  MUX2_X1 _08282_ (
    .A(reg_pmp_3_cfg_w),
    .B(_03277_),
    .S(_03275_),
    .Z(_00096_)
  );
  MUX2_X1 _08283_ (
    .A(reg_pmp_3_cfg_x),
    .B(_03017_),
    .S(_03275_),
    .Z(_00097_)
  );
  MUX2_X1 _08284_ (
    .A(reg_pmp_3_cfg_r),
    .B(_02873_),
    .S(_03275_),
    .Z(_00098_)
  );
  AND2_X1 _08285_ (
    .A1(_00009_),
    .A2(_00916_),
    .ZN(_03278_)
  );
  AND2_X1 _08286_ (
    .A1(_00897_),
    .A2(_03278_),
    .ZN(_03279_)
  );
  INV_X1 _08287_ (
    .A(_03279_),
    .ZN(_03280_)
  );
  AND2_X1 _08288_ (
    .A1(_01035_),
    .A2(_02669_),
    .ZN(_03281_)
  );
  MUX2_X1 _08289_ (
    .A(reg_pmp_2_cfg_w),
    .B(_03281_),
    .S(_03279_),
    .Z(_00099_)
  );
  AND2_X1 _08290_ (
    .A1(_00801_),
    .A2(_03276_),
    .ZN(_03282_)
  );
  INV_X1 _08291_ (
    .A(_03282_),
    .ZN(_03283_)
  );
  AND2_X1 _08292_ (
    .A1(_00811_),
    .A2(_03283_),
    .ZN(_03284_)
  );
  AND2_X1 _08293_ (
    .A1(_03090_),
    .A2(_03275_),
    .ZN(_03285_)
  );
  INV_X1 _08294_ (
    .A(_03285_),
    .ZN(_03286_)
  );
  AND2_X1 _08295_ (
    .A1(_03284_),
    .A2(_03286_),
    .ZN(_00100_)
  );
  AND2_X1 _08296_ (
    .A1(_00800_),
    .A2(_03276_),
    .ZN(_03287_)
  );
  INV_X1 _08297_ (
    .A(_03287_),
    .ZN(_03288_)
  );
  AND2_X1 _08298_ (
    .A1(_00811_),
    .A2(_03288_),
    .ZN(_03289_)
  );
  AND2_X1 _08299_ (
    .A1(_03161_),
    .A2(_03275_),
    .ZN(_03290_)
  );
  INV_X1 _08300_ (
    .A(_03290_),
    .ZN(_03291_)
  );
  AND2_X1 _08301_ (
    .A1(_03289_),
    .A2(_03291_),
    .ZN(_00101_)
  );
  AND2_X1 _08302_ (
    .A1(_00799_),
    .A2(_03276_),
    .ZN(_03292_)
  );
  INV_X1 _08303_ (
    .A(_03292_),
    .ZN(_03293_)
  );
  AND2_X1 _08304_ (
    .A1(_00811_),
    .A2(_03293_),
    .ZN(_03294_)
  );
  AND2_X1 _08305_ (
    .A1(io_rw_wdata[31]),
    .A2(_00903_),
    .ZN(_03295_)
  );
  INV_X1 _08306_ (
    .A(_03295_),
    .ZN(_03296_)
  );
  AND2_X1 _08307_ (
    .A1(large_1[57]),
    .A2(_01019_),
    .ZN(_03297_)
  );
  INV_X1 _08308_ (
    .A(_03297_),
    .ZN(_03298_)
  );
  AND2_X1 _08309_ (
    .A1(large_[57]),
    .A2(_00991_),
    .ZN(_03299_)
  );
  INV_X1 _08310_ (
    .A(_03299_),
    .ZN(_03300_)
  );
  AND2_X1 _08311_ (
    .A1(large_1[25]),
    .A2(_00995_),
    .ZN(_03301_)
  );
  INV_X1 _08312_ (
    .A(_03301_),
    .ZN(_03302_)
  );
  AND2_X1 _08313_ (
    .A1(_03300_),
    .A2(_03302_),
    .ZN(_03303_)
  );
  AND2_X1 _08314_ (
    .A1(_03298_),
    .A2(_03303_),
    .ZN(_03304_)
  );
  AND2_X1 _08315_ (
    .A1(reg_pmp_7_cfg_l),
    .A2(_00894_),
    .ZN(_03305_)
  );
  INV_X1 _08316_ (
    .A(_03305_),
    .ZN(_03306_)
  );
  AND2_X1 _08317_ (
    .A1(reg_pmp_3_cfg_l),
    .A2(_00916_),
    .ZN(_03307_)
  );
  INV_X1 _08318_ (
    .A(_03307_),
    .ZN(_03308_)
  );
  AND2_X1 _08319_ (
    .A1(_03306_),
    .A2(_03308_),
    .ZN(_03309_)
  );
  AND2_X1 _08320_ (
    .A1(reg_bp_0_address[31]),
    .A2(_00962_),
    .ZN(_03310_)
  );
  INV_X1 _08321_ (
    .A(_03310_),
    .ZN(_03311_)
  );
  AND2_X1 _08322_ (
    .A1(reg_mepc[31]),
    .A2(_00943_),
    .ZN(_03312_)
  );
  INV_X1 _08323_ (
    .A(_03312_),
    .ZN(_03313_)
  );
  AND2_X1 _08324_ (
    .A1(_03311_),
    .A2(_03313_),
    .ZN(_03314_)
  );
  AND2_X1 _08325_ (
    .A1(_03309_),
    .A2(_03314_),
    .ZN(_03315_)
  );
  AND2_X1 _08326_ (
    .A1(reg_mcause[31]),
    .A2(_01001_),
    .ZN(_03316_)
  );
  INV_X1 _08327_ (
    .A(_03316_),
    .ZN(_03317_)
  );
  AND2_X1 _08328_ (
    .A1(reg_dpc[31]),
    .A2(_00912_),
    .ZN(_03318_)
  );
  INV_X1 _08329_ (
    .A(_03318_),
    .ZN(_03319_)
  );
  AND2_X1 _08330_ (
    .A1(_03317_),
    .A2(_03319_),
    .ZN(_03320_)
  );
  AND2_X1 _08331_ (
    .A1(reg_dscratch0[31]),
    .A2(_00958_),
    .ZN(_03321_)
  );
  INV_X1 _08332_ (
    .A(_03321_),
    .ZN(_03322_)
  );
  AND2_X1 _08333_ (
    .A1(reg_mtvec[31]),
    .A2(_00940_),
    .ZN(_03323_)
  );
  INV_X1 _08334_ (
    .A(_03323_),
    .ZN(_03324_)
  );
  AND2_X1 _08335_ (
    .A1(_03322_),
    .A2(_03324_),
    .ZN(_03325_)
  );
  AND2_X1 _08336_ (
    .A1(_03320_),
    .A2(_03325_),
    .ZN(_03326_)
  );
  AND2_X1 _08337_ (
    .A1(large_[25]),
    .A2(_00985_),
    .ZN(_03327_)
  );
  INV_X1 _08338_ (
    .A(_03327_),
    .ZN(_03328_)
  );
  AND2_X1 _08339_ (
    .A1(reg_mtval[31]),
    .A2(_00926_),
    .ZN(_03329_)
  );
  INV_X1 _08340_ (
    .A(_03329_),
    .ZN(_03330_)
  );
  AND2_X1 _08341_ (
    .A1(reg_mscratch[31]),
    .A2(_00929_),
    .ZN(_03331_)
  );
  INV_X1 _08342_ (
    .A(_03331_),
    .ZN(_03332_)
  );
  AND2_X1 _08343_ (
    .A1(_03330_),
    .A2(_03332_),
    .ZN(_03333_)
  );
  AND2_X1 _08344_ (
    .A1(_03328_),
    .A2(_03333_),
    .ZN(_03334_)
  );
  AND2_X1 _08345_ (
    .A1(_03326_),
    .A2(_03334_),
    .ZN(_03335_)
  );
  AND2_X1 _08346_ (
    .A1(_03315_),
    .A2(_03335_),
    .ZN(_03336_)
  );
  AND2_X1 _08347_ (
    .A1(_03304_),
    .A2(_03336_),
    .ZN(_03337_)
  );
  INV_X1 _08348_ (
    .A(_03337_),
    .ZN(io_rw_rdata[31])
  );
  AND2_X1 _08349_ (
    .A1(io_rw_cmd[1]),
    .A2(_00866_),
    .ZN(_03338_)
  );
  AND2_X1 _08350_ (
    .A1(io_rw_rdata[31]),
    .A2(_03338_),
    .ZN(_03339_)
  );
  INV_X1 _08351_ (
    .A(_03339_),
    .ZN(_03340_)
  );
  AND2_X1 _08352_ (
    .A1(_03296_),
    .A2(_03340_),
    .ZN(_03341_)
  );
  INV_X1 _08353_ (
    .A(_03341_),
    .ZN(_03342_)
  );
  AND2_X1 _08354_ (
    .A1(_03275_),
    .A2(_03341_),
    .ZN(_03343_)
  );
  INV_X1 _08355_ (
    .A(_03343_),
    .ZN(_03344_)
  );
  AND2_X1 _08356_ (
    .A1(_03294_),
    .A2(_03344_),
    .ZN(_00102_)
  );
  AND2_X1 _08357_ (
    .A1(reg_pmp_3_cfg_l),
    .A2(reg_pmp_3_cfg_a[0]),
    .ZN(_03345_)
  );
  AND2_X1 _08358_ (
    .A1(_00012_),
    .A2(_03345_),
    .ZN(_03346_)
  );
  INV_X1 _08359_ (
    .A(_03346_),
    .ZN(_03347_)
  );
  AND2_X1 _08360_ (
    .A1(_00796_),
    .A2(_03347_),
    .ZN(_03348_)
  );
  AND2_X1 _08361_ (
    .A1(_00897_),
    .A2(_03348_),
    .ZN(_03349_)
  );
  AND2_X1 _08362_ (
    .A1(_00953_),
    .A2(_03349_),
    .ZN(_03350_)
  );
  MUX2_X1 _08363_ (
    .A(reg_pmp_2_addr[0]),
    .B(_01613_),
    .S(_03350_),
    .Z(_00103_)
  );
  MUX2_X1 _08364_ (
    .A(reg_pmp_2_addr[1]),
    .B(_01688_),
    .S(_03350_),
    .Z(_00104_)
  );
  MUX2_X1 _08365_ (
    .A(reg_pmp_2_addr[2]),
    .B(_01774_),
    .S(_03350_),
    .Z(_00105_)
  );
  MUX2_X1 _08366_ (
    .A(reg_pmp_2_addr[3]),
    .B(_01865_),
    .S(_03350_),
    .Z(_00106_)
  );
  MUX2_X1 _08367_ (
    .A(reg_pmp_2_addr[4]),
    .B(_01938_),
    .S(_03350_),
    .Z(_00107_)
  );
  MUX2_X1 _08368_ (
    .A(reg_pmp_2_addr[5]),
    .B(_02005_),
    .S(_03350_),
    .Z(_00108_)
  );
  MUX2_X1 _08369_ (
    .A(reg_pmp_2_addr[6]),
    .B(_02076_),
    .S(_03350_),
    .Z(_00109_)
  );
  MUX2_X1 _08370_ (
    .A(reg_pmp_2_addr[7]),
    .B(_02163_),
    .S(_03350_),
    .Z(_00110_)
  );
  MUX2_X1 _08371_ (
    .A(reg_pmp_2_addr[8]),
    .B(_01446_),
    .S(_03350_),
    .Z(_00111_)
  );
  MUX2_X1 _08372_ (
    .A(reg_pmp_2_addr[9]),
    .B(_01518_),
    .S(_03350_),
    .Z(_00112_)
  );
  MUX2_X1 _08373_ (
    .A(reg_pmp_2_addr[10]),
    .B(_02235_),
    .S(_03350_),
    .Z(_00113_)
  );
  MUX2_X1 _08374_ (
    .A(reg_pmp_2_addr[11]),
    .B(_02314_),
    .S(_03350_),
    .Z(_00114_)
  );
  MUX2_X1 _08375_ (
    .A(reg_pmp_2_addr[12]),
    .B(_02389_),
    .S(_03350_),
    .Z(_00115_)
  );
  MUX2_X1 _08376_ (
    .A(reg_pmp_2_addr[13]),
    .B(_02456_),
    .S(_03350_),
    .Z(_00116_)
  );
  MUX2_X1 _08377_ (
    .A(reg_pmp_2_addr[14]),
    .B(_02522_),
    .S(_03350_),
    .Z(_00117_)
  );
  MUX2_X1 _08378_ (
    .A(reg_pmp_2_addr[15]),
    .B(_02597_),
    .S(_03350_),
    .Z(_00118_)
  );
  MUX2_X1 _08379_ (
    .A(reg_pmp_2_addr[16]),
    .B(_01035_),
    .S(_03350_),
    .Z(_00119_)
  );
  MUX2_X1 _08380_ (
    .A(reg_pmp_2_addr[17]),
    .B(_02669_),
    .S(_03350_),
    .Z(_00120_)
  );
  MUX2_X1 _08381_ (
    .A(reg_pmp_2_addr[18]),
    .B(_01107_),
    .S(_03350_),
    .Z(_00121_)
  );
  MUX2_X1 _08382_ (
    .A(reg_pmp_2_addr[19]),
    .B(_01199_),
    .S(_03350_),
    .Z(_00122_)
  );
  MUX2_X1 _08383_ (
    .A(reg_pmp_2_addr[20]),
    .B(_01277_),
    .S(_03350_),
    .Z(_00123_)
  );
  MUX2_X1 _08384_ (
    .A(reg_pmp_2_addr[21]),
    .B(_02735_),
    .S(_03350_),
    .Z(_00124_)
  );
  MUX2_X1 _08385_ (
    .A(reg_pmp_2_addr[22]),
    .B(_02801_),
    .S(_03350_),
    .Z(_00125_)
  );
  MUX2_X1 _08386_ (
    .A(reg_pmp_2_addr[23]),
    .B(_01360_),
    .S(_03350_),
    .Z(_00126_)
  );
  MUX2_X1 _08387_ (
    .A(reg_pmp_2_addr[24]),
    .B(_02873_),
    .S(_03350_),
    .Z(_00127_)
  );
  MUX2_X1 _08388_ (
    .A(reg_pmp_2_addr[25]),
    .B(_02945_),
    .S(_03350_),
    .Z(_00128_)
  );
  MUX2_X1 _08389_ (
    .A(reg_pmp_2_addr[26]),
    .B(_03017_),
    .S(_03350_),
    .Z(_00129_)
  );
  MUX2_X1 _08390_ (
    .A(reg_pmp_2_addr[27]),
    .B(_03089_),
    .S(_03350_),
    .Z(_00130_)
  );
  MUX2_X1 _08391_ (
    .A(reg_pmp_2_addr[28]),
    .B(_03162_),
    .S(_03350_),
    .Z(_00131_)
  );
  MUX2_X1 _08392_ (
    .A(reg_pmp_2_addr[29]),
    .B(_03230_),
    .S(_03350_),
    .Z(_00132_)
  );
  AND2_X1 _08393_ (
    .A1(_00007_),
    .A2(_00916_),
    .ZN(_03351_)
  );
  AND2_X1 _08394_ (
    .A1(_00897_),
    .A2(_03351_),
    .ZN(_03352_)
  );
  INV_X1 _08395_ (
    .A(_03352_),
    .ZN(_03353_)
  );
  MUX2_X1 _08396_ (
    .A(reg_pmp_1_cfg_w),
    .B(_01519_),
    .S(_03352_),
    .Z(_00133_)
  );
  MUX2_X1 _08397_ (
    .A(reg_pmp_2_cfg_r),
    .B(_01035_),
    .S(_03279_),
    .Z(_00134_)
  );
  AND2_X1 _08398_ (
    .A1(reg_pmp_4_cfg_l),
    .A2(reg_pmp_4_cfg_a[0]),
    .ZN(_03354_)
  );
  AND2_X1 _08399_ (
    .A1(_00014_),
    .A2(_03354_),
    .ZN(_03355_)
  );
  INV_X1 _08400_ (
    .A(_03355_),
    .ZN(_03356_)
  );
  AND2_X1 _08401_ (
    .A1(_00799_),
    .A2(_03356_),
    .ZN(_03357_)
  );
  AND2_X1 _08402_ (
    .A1(_00897_),
    .A2(_03357_),
    .ZN(_03358_)
  );
  AND2_X1 _08403_ (
    .A1(_01011_),
    .A2(_03358_),
    .ZN(_03359_)
  );
  MUX2_X1 _08404_ (
    .A(reg_pmp_3_addr[0]),
    .B(_01613_),
    .S(_03359_),
    .Z(_00135_)
  );
  MUX2_X1 _08405_ (
    .A(reg_pmp_3_addr[1]),
    .B(_01688_),
    .S(_03359_),
    .Z(_00136_)
  );
  MUX2_X1 _08406_ (
    .A(reg_pmp_3_addr[2]),
    .B(_01774_),
    .S(_03359_),
    .Z(_00137_)
  );
  MUX2_X1 _08407_ (
    .A(reg_pmp_3_addr[3]),
    .B(_01865_),
    .S(_03359_),
    .Z(_00138_)
  );
  MUX2_X1 _08408_ (
    .A(reg_pmp_3_addr[4]),
    .B(_01938_),
    .S(_03359_),
    .Z(_00139_)
  );
  MUX2_X1 _08409_ (
    .A(reg_pmp_3_addr[5]),
    .B(_02005_),
    .S(_03359_),
    .Z(_00140_)
  );
  MUX2_X1 _08410_ (
    .A(reg_pmp_3_addr[6]),
    .B(_02076_),
    .S(_03359_),
    .Z(_00141_)
  );
  MUX2_X1 _08411_ (
    .A(reg_pmp_3_addr[7]),
    .B(_02163_),
    .S(_03359_),
    .Z(_00142_)
  );
  MUX2_X1 _08412_ (
    .A(reg_pmp_3_addr[8]),
    .B(_01446_),
    .S(_03359_),
    .Z(_00143_)
  );
  MUX2_X1 _08413_ (
    .A(reg_pmp_3_addr[9]),
    .B(_01518_),
    .S(_03359_),
    .Z(_00144_)
  );
  MUX2_X1 _08414_ (
    .A(reg_pmp_3_addr[10]),
    .B(_02235_),
    .S(_03359_),
    .Z(_00145_)
  );
  MUX2_X1 _08415_ (
    .A(reg_pmp_3_addr[11]),
    .B(_02314_),
    .S(_03359_),
    .Z(_00146_)
  );
  MUX2_X1 _08416_ (
    .A(reg_pmp_3_addr[12]),
    .B(_02389_),
    .S(_03359_),
    .Z(_00147_)
  );
  MUX2_X1 _08417_ (
    .A(reg_pmp_3_addr[13]),
    .B(_02456_),
    .S(_03359_),
    .Z(_00148_)
  );
  MUX2_X1 _08418_ (
    .A(reg_pmp_3_addr[14]),
    .B(_02522_),
    .S(_03359_),
    .Z(_00149_)
  );
  MUX2_X1 _08419_ (
    .A(reg_pmp_3_addr[15]),
    .B(_02597_),
    .S(_03359_),
    .Z(_00150_)
  );
  MUX2_X1 _08420_ (
    .A(reg_pmp_3_addr[16]),
    .B(_01035_),
    .S(_03359_),
    .Z(_00151_)
  );
  MUX2_X1 _08421_ (
    .A(reg_pmp_3_addr[17]),
    .B(_02669_),
    .S(_03359_),
    .Z(_00152_)
  );
  MUX2_X1 _08422_ (
    .A(reg_pmp_3_addr[18]),
    .B(_01107_),
    .S(_03359_),
    .Z(_00153_)
  );
  MUX2_X1 _08423_ (
    .A(reg_pmp_3_addr[19]),
    .B(_01199_),
    .S(_03359_),
    .Z(_00154_)
  );
  MUX2_X1 _08424_ (
    .A(reg_pmp_3_addr[20]),
    .B(_01277_),
    .S(_03359_),
    .Z(_00155_)
  );
  MUX2_X1 _08425_ (
    .A(reg_pmp_3_addr[21]),
    .B(_02735_),
    .S(_03359_),
    .Z(_00156_)
  );
  MUX2_X1 _08426_ (
    .A(reg_pmp_3_addr[22]),
    .B(_02801_),
    .S(_03359_),
    .Z(_00157_)
  );
  MUX2_X1 _08427_ (
    .A(reg_pmp_3_addr[23]),
    .B(_01360_),
    .S(_03359_),
    .Z(_00158_)
  );
  MUX2_X1 _08428_ (
    .A(reg_pmp_3_addr[24]),
    .B(_02873_),
    .S(_03359_),
    .Z(_00159_)
  );
  MUX2_X1 _08429_ (
    .A(reg_pmp_3_addr[25]),
    .B(_02945_),
    .S(_03359_),
    .Z(_00160_)
  );
  MUX2_X1 _08430_ (
    .A(reg_pmp_3_addr[26]),
    .B(_03017_),
    .S(_03359_),
    .Z(_00161_)
  );
  MUX2_X1 _08431_ (
    .A(reg_pmp_3_addr[27]),
    .B(_03089_),
    .S(_03359_),
    .Z(_00162_)
  );
  MUX2_X1 _08432_ (
    .A(reg_pmp_3_addr[28]),
    .B(_03162_),
    .S(_03359_),
    .Z(_00163_)
  );
  MUX2_X1 _08433_ (
    .A(reg_pmp_3_addr[29]),
    .B(_03230_),
    .S(_03359_),
    .Z(_00164_)
  );
  AND2_X1 _08434_ (
    .A1(_00798_),
    .A2(_03280_),
    .ZN(_03360_)
  );
  INV_X1 _08435_ (
    .A(_03360_),
    .ZN(_03361_)
  );
  AND2_X1 _08436_ (
    .A1(_00811_),
    .A2(_03361_),
    .ZN(_03362_)
  );
  AND2_X1 _08437_ (
    .A1(_01198_),
    .A2(_03279_),
    .ZN(_03363_)
  );
  INV_X1 _08438_ (
    .A(_03363_),
    .ZN(_03364_)
  );
  AND2_X1 _08439_ (
    .A1(_03362_),
    .A2(_03364_),
    .ZN(_00165_)
  );
  AND2_X1 _08440_ (
    .A1(_00797_),
    .A2(_03280_),
    .ZN(_03365_)
  );
  INV_X1 _08441_ (
    .A(_03365_),
    .ZN(_03366_)
  );
  AND2_X1 _08442_ (
    .A1(_00811_),
    .A2(_03366_),
    .ZN(_03367_)
  );
  AND2_X1 _08443_ (
    .A1(_01276_),
    .A2(_03279_),
    .ZN(_03368_)
  );
  INV_X1 _08444_ (
    .A(_03368_),
    .ZN(_03369_)
  );
  AND2_X1 _08445_ (
    .A1(_03367_),
    .A2(_03369_),
    .ZN(_00166_)
  );
  AND2_X1 _08446_ (
    .A1(_00796_),
    .A2(_03280_),
    .ZN(_03370_)
  );
  INV_X1 _08447_ (
    .A(_03370_),
    .ZN(_03371_)
  );
  AND2_X1 _08448_ (
    .A1(_00811_),
    .A2(_03371_),
    .ZN(_03372_)
  );
  AND2_X1 _08449_ (
    .A1(_01359_),
    .A2(_03279_),
    .ZN(_03373_)
  );
  INV_X1 _08450_ (
    .A(_03373_),
    .ZN(_03374_)
  );
  AND2_X1 _08451_ (
    .A1(_03372_),
    .A2(_03374_),
    .ZN(_00167_)
  );
  MUX2_X1 _08452_ (
    .A(reg_pmp_1_cfg_r),
    .B(_01446_),
    .S(_03352_),
    .Z(_00168_)
  );
  MUX2_X1 _08453_ (
    .A(reg_pmp_4_cfg_r),
    .B(_01613_),
    .S(_03257_),
    .Z(_00169_)
  );
  MUX2_X1 _08454_ (
    .A(reg_pmp_1_cfg_x),
    .B(_02235_),
    .S(_03352_),
    .Z(_00170_)
  );
  MUX2_X1 _08455_ (
    .A(reg_pmp_2_cfg_x),
    .B(_01107_),
    .S(_03279_),
    .Z(_00171_)
  );
  AND2_X1 _08456_ (
    .A1(_00795_),
    .A2(_03353_),
    .ZN(_03375_)
  );
  INV_X1 _08457_ (
    .A(_03375_),
    .ZN(_03376_)
  );
  AND2_X1 _08458_ (
    .A1(_00811_),
    .A2(_03376_),
    .ZN(_03377_)
  );
  AND2_X1 _08459_ (
    .A1(_02313_),
    .A2(_03352_),
    .ZN(_03378_)
  );
  INV_X1 _08460_ (
    .A(_03378_),
    .ZN(_03379_)
  );
  AND2_X1 _08461_ (
    .A1(_03377_),
    .A2(_03379_),
    .ZN(_00172_)
  );
  AND2_X1 _08462_ (
    .A1(_00794_),
    .A2(_03353_),
    .ZN(_03380_)
  );
  INV_X1 _08463_ (
    .A(_03380_),
    .ZN(_03381_)
  );
  AND2_X1 _08464_ (
    .A1(_00811_),
    .A2(_03381_),
    .ZN(_03382_)
  );
  AND2_X1 _08465_ (
    .A1(_02390_),
    .A2(_03352_),
    .ZN(_03383_)
  );
  INV_X1 _08466_ (
    .A(_03383_),
    .ZN(_03384_)
  );
  AND2_X1 _08467_ (
    .A1(_03382_),
    .A2(_03384_),
    .ZN(_00173_)
  );
  AND2_X1 _08468_ (
    .A1(_00793_),
    .A2(_03353_),
    .ZN(_03385_)
  );
  INV_X1 _08469_ (
    .A(_03385_),
    .ZN(_03386_)
  );
  AND2_X1 _08470_ (
    .A1(_00811_),
    .A2(_03386_),
    .ZN(_03387_)
  );
  AND2_X1 _08471_ (
    .A1(_02596_),
    .A2(_03352_),
    .ZN(_03388_)
  );
  INV_X1 _08472_ (
    .A(_03388_),
    .ZN(_03389_)
  );
  AND2_X1 _08473_ (
    .A1(_03387_),
    .A2(_03389_),
    .ZN(_00174_)
  );
  MUX2_X1 _08474_ (
    .A(reg_pmp_0_cfg_r),
    .B(_01613_),
    .S(_03232_),
    .Z(_00175_)
  );
  AND2_X1 _08475_ (
    .A1(reg_pmp_1_cfg_l),
    .A2(reg_pmp_1_cfg_a[0]),
    .ZN(_03390_)
  );
  AND2_X1 _08476_ (
    .A1(_00008_),
    .A2(_03390_),
    .ZN(_03391_)
  );
  INV_X1 _08477_ (
    .A(_03391_),
    .ZN(_03392_)
  );
  AND2_X1 _08478_ (
    .A1(_00790_),
    .A2(_03392_),
    .ZN(_03393_)
  );
  AND2_X1 _08479_ (
    .A1(_00897_),
    .A2(_03393_),
    .ZN(_03394_)
  );
  AND2_X1 _08480_ (
    .A1(_01004_),
    .A2(_03394_),
    .ZN(_03395_)
  );
  MUX2_X1 _08481_ (
    .A(reg_pmp_0_addr[0]),
    .B(_01613_),
    .S(_03395_),
    .Z(_00176_)
  );
  MUX2_X1 _08482_ (
    .A(reg_pmp_0_addr[1]),
    .B(_01688_),
    .S(_03395_),
    .Z(_00177_)
  );
  MUX2_X1 _08483_ (
    .A(reg_pmp_0_addr[2]),
    .B(_01774_),
    .S(_03395_),
    .Z(_00178_)
  );
  MUX2_X1 _08484_ (
    .A(reg_pmp_0_addr[3]),
    .B(_01865_),
    .S(_03395_),
    .Z(_00179_)
  );
  MUX2_X1 _08485_ (
    .A(reg_pmp_0_addr[4]),
    .B(_01938_),
    .S(_03395_),
    .Z(_00180_)
  );
  MUX2_X1 _08486_ (
    .A(reg_pmp_0_addr[5]),
    .B(_02005_),
    .S(_03395_),
    .Z(_00181_)
  );
  MUX2_X1 _08487_ (
    .A(reg_pmp_0_addr[6]),
    .B(_02076_),
    .S(_03395_),
    .Z(_00182_)
  );
  MUX2_X1 _08488_ (
    .A(reg_pmp_0_addr[7]),
    .B(_02163_),
    .S(_03395_),
    .Z(_00183_)
  );
  MUX2_X1 _08489_ (
    .A(reg_pmp_0_addr[8]),
    .B(_01446_),
    .S(_03395_),
    .Z(_00184_)
  );
  MUX2_X1 _08490_ (
    .A(reg_pmp_0_addr[9]),
    .B(_01518_),
    .S(_03395_),
    .Z(_00185_)
  );
  MUX2_X1 _08491_ (
    .A(reg_pmp_0_addr[10]),
    .B(_02235_),
    .S(_03395_),
    .Z(_00186_)
  );
  MUX2_X1 _08492_ (
    .A(reg_pmp_0_addr[11]),
    .B(_02314_),
    .S(_03395_),
    .Z(_00187_)
  );
  MUX2_X1 _08493_ (
    .A(reg_pmp_0_addr[12]),
    .B(_02389_),
    .S(_03395_),
    .Z(_00188_)
  );
  MUX2_X1 _08494_ (
    .A(reg_pmp_0_addr[13]),
    .B(_02456_),
    .S(_03395_),
    .Z(_00189_)
  );
  MUX2_X1 _08495_ (
    .A(reg_pmp_0_addr[14]),
    .B(_02522_),
    .S(_03395_),
    .Z(_00190_)
  );
  MUX2_X1 _08496_ (
    .A(reg_pmp_0_addr[15]),
    .B(_02597_),
    .S(_03395_),
    .Z(_00191_)
  );
  MUX2_X1 _08497_ (
    .A(reg_pmp_0_addr[16]),
    .B(_01035_),
    .S(_03395_),
    .Z(_00192_)
  );
  MUX2_X1 _08498_ (
    .A(reg_pmp_0_addr[17]),
    .B(_02669_),
    .S(_03395_),
    .Z(_00193_)
  );
  MUX2_X1 _08499_ (
    .A(reg_pmp_0_addr[18]),
    .B(_01107_),
    .S(_03395_),
    .Z(_00194_)
  );
  MUX2_X1 _08500_ (
    .A(reg_pmp_0_addr[19]),
    .B(_01199_),
    .S(_03395_),
    .Z(_00195_)
  );
  MUX2_X1 _08501_ (
    .A(reg_pmp_0_addr[20]),
    .B(_01277_),
    .S(_03395_),
    .Z(_00196_)
  );
  MUX2_X1 _08502_ (
    .A(reg_pmp_0_addr[21]),
    .B(_02735_),
    .S(_03395_),
    .Z(_00197_)
  );
  MUX2_X1 _08503_ (
    .A(reg_pmp_0_addr[22]),
    .B(_02801_),
    .S(_03395_),
    .Z(_00198_)
  );
  MUX2_X1 _08504_ (
    .A(reg_pmp_0_addr[23]),
    .B(_01360_),
    .S(_03395_),
    .Z(_00199_)
  );
  MUX2_X1 _08505_ (
    .A(reg_pmp_0_addr[24]),
    .B(_02873_),
    .S(_03395_),
    .Z(_00200_)
  );
  MUX2_X1 _08506_ (
    .A(reg_pmp_0_addr[25]),
    .B(_02945_),
    .S(_03395_),
    .Z(_00201_)
  );
  MUX2_X1 _08507_ (
    .A(reg_pmp_0_addr[26]),
    .B(_03017_),
    .S(_03395_),
    .Z(_00202_)
  );
  MUX2_X1 _08508_ (
    .A(reg_pmp_0_addr[27]),
    .B(_03089_),
    .S(_03395_),
    .Z(_00203_)
  );
  MUX2_X1 _08509_ (
    .A(reg_pmp_0_addr[28]),
    .B(_03162_),
    .S(_03395_),
    .Z(_00204_)
  );
  MUX2_X1 _08510_ (
    .A(reg_pmp_0_addr[29]),
    .B(_03230_),
    .S(_03395_),
    .Z(_00205_)
  );
  MUX2_X1 _08511_ (
    .A(reg_pmp_0_cfg_x),
    .B(_01774_),
    .S(_03232_),
    .Z(_00206_)
  );
  AND2_X1 _08512_ (
    .A1(_00870_),
    .A2(_00881_),
    .ZN(_03396_)
  );
  INV_X1 _08513_ (
    .A(_03396_),
    .ZN(_03397_)
  );
  AND2_X1 _08514_ (
    .A1(_00897_),
    .A2(_03397_),
    .ZN(_03398_)
  );
  AND2_X1 _08515_ (
    .A1(_00962_),
    .A2(_03398_),
    .ZN(_03399_)
  );
  MUX2_X1 _08516_ (
    .A(reg_bp_0_address[0]),
    .B(_01613_),
    .S(_03399_),
    .Z(_00207_)
  );
  MUX2_X1 _08517_ (
    .A(reg_bp_0_address[1]),
    .B(_01688_),
    .S(_03399_),
    .Z(_00208_)
  );
  MUX2_X1 _08518_ (
    .A(reg_bp_0_address[2]),
    .B(_01774_),
    .S(_03399_),
    .Z(_00209_)
  );
  MUX2_X1 _08519_ (
    .A(reg_bp_0_address[3]),
    .B(_01865_),
    .S(_03399_),
    .Z(_00210_)
  );
  MUX2_X1 _08520_ (
    .A(reg_bp_0_address[4]),
    .B(_01938_),
    .S(_03399_),
    .Z(_00211_)
  );
  MUX2_X1 _08521_ (
    .A(reg_bp_0_address[5]),
    .B(_02005_),
    .S(_03399_),
    .Z(_00212_)
  );
  MUX2_X1 _08522_ (
    .A(reg_bp_0_address[6]),
    .B(_02076_),
    .S(_03399_),
    .Z(_00213_)
  );
  MUX2_X1 _08523_ (
    .A(reg_bp_0_address[7]),
    .B(_02163_),
    .S(_03399_),
    .Z(_00214_)
  );
  MUX2_X1 _08524_ (
    .A(reg_bp_0_address[8]),
    .B(_01446_),
    .S(_03399_),
    .Z(_00215_)
  );
  MUX2_X1 _08525_ (
    .A(reg_bp_0_address[9]),
    .B(_01518_),
    .S(_03399_),
    .Z(_00216_)
  );
  MUX2_X1 _08526_ (
    .A(reg_bp_0_address[10]),
    .B(_02235_),
    .S(_03399_),
    .Z(_00217_)
  );
  MUX2_X1 _08527_ (
    .A(reg_bp_0_address[11]),
    .B(_02314_),
    .S(_03399_),
    .Z(_00218_)
  );
  MUX2_X1 _08528_ (
    .A(reg_bp_0_address[12]),
    .B(_02389_),
    .S(_03399_),
    .Z(_00219_)
  );
  MUX2_X1 _08529_ (
    .A(reg_bp_0_address[13]),
    .B(_02456_),
    .S(_03399_),
    .Z(_00220_)
  );
  MUX2_X1 _08530_ (
    .A(reg_bp_0_address[14]),
    .B(_02522_),
    .S(_03399_),
    .Z(_00221_)
  );
  MUX2_X1 _08531_ (
    .A(reg_bp_0_address[15]),
    .B(_02597_),
    .S(_03399_),
    .Z(_00222_)
  );
  MUX2_X1 _08532_ (
    .A(reg_bp_0_address[16]),
    .B(_01035_),
    .S(_03399_),
    .Z(_00223_)
  );
  MUX2_X1 _08533_ (
    .A(reg_bp_0_address[17]),
    .B(_02669_),
    .S(_03399_),
    .Z(_00224_)
  );
  MUX2_X1 _08534_ (
    .A(reg_bp_0_address[18]),
    .B(_01107_),
    .S(_03399_),
    .Z(_00225_)
  );
  MUX2_X1 _08535_ (
    .A(reg_bp_0_address[19]),
    .B(_01199_),
    .S(_03399_),
    .Z(_00226_)
  );
  MUX2_X1 _08536_ (
    .A(reg_bp_0_address[20]),
    .B(_01277_),
    .S(_03399_),
    .Z(_00227_)
  );
  MUX2_X1 _08537_ (
    .A(reg_bp_0_address[21]),
    .B(_02735_),
    .S(_03399_),
    .Z(_00228_)
  );
  MUX2_X1 _08538_ (
    .A(reg_bp_0_address[22]),
    .B(_02801_),
    .S(_03399_),
    .Z(_00229_)
  );
  MUX2_X1 _08539_ (
    .A(reg_bp_0_address[23]),
    .B(_01360_),
    .S(_03399_),
    .Z(_00230_)
  );
  MUX2_X1 _08540_ (
    .A(reg_bp_0_address[24]),
    .B(_02873_),
    .S(_03399_),
    .Z(_00231_)
  );
  MUX2_X1 _08541_ (
    .A(reg_bp_0_address[25]),
    .B(_02945_),
    .S(_03399_),
    .Z(_00232_)
  );
  MUX2_X1 _08542_ (
    .A(reg_bp_0_address[26]),
    .B(_03017_),
    .S(_03399_),
    .Z(_00233_)
  );
  MUX2_X1 _08543_ (
    .A(reg_bp_0_address[27]),
    .B(_03089_),
    .S(_03399_),
    .Z(_00234_)
  );
  MUX2_X1 _08544_ (
    .A(reg_bp_0_address[28]),
    .B(_03162_),
    .S(_03399_),
    .Z(_00235_)
  );
  MUX2_X1 _08545_ (
    .A(reg_bp_0_address[29]),
    .B(_03230_),
    .S(_03399_),
    .Z(_00236_)
  );
  AND2_X1 _08546_ (
    .A1(io_rw_wdata[30]),
    .A2(_00903_),
    .ZN(_03400_)
  );
  INV_X1 _08547_ (
    .A(_03400_),
    .ZN(_03401_)
  );
  AND2_X1 _08548_ (
    .A1(large_[56]),
    .A2(_00991_),
    .ZN(_03402_)
  );
  INV_X1 _08549_ (
    .A(_03402_),
    .ZN(_03403_)
  );
  AND2_X1 _08550_ (
    .A1(large_1[56]),
    .A2(_01019_),
    .ZN(_03404_)
  );
  INV_X1 _08551_ (
    .A(_03404_),
    .ZN(_03405_)
  );
  AND2_X1 _08552_ (
    .A1(reg_dscratch0[30]),
    .A2(_00958_),
    .ZN(_03406_)
  );
  INV_X1 _08553_ (
    .A(_03406_),
    .ZN(_03407_)
  );
  AND2_X1 _08554_ (
    .A1(reg_mtval[30]),
    .A2(_00926_),
    .ZN(_03408_)
  );
  INV_X1 _08555_ (
    .A(_03408_),
    .ZN(_03409_)
  );
  AND2_X1 _08556_ (
    .A1(reg_bp_0_address[30]),
    .A2(_00962_),
    .ZN(_03410_)
  );
  INV_X1 _08557_ (
    .A(_03410_),
    .ZN(_03411_)
  );
  AND2_X1 _08558_ (
    .A1(reg_mepc[30]),
    .A2(_00943_),
    .ZN(_03412_)
  );
  INV_X1 _08559_ (
    .A(_03412_),
    .ZN(_03413_)
  );
  AND2_X1 _08560_ (
    .A1(reg_dpc[30]),
    .A2(_00912_),
    .ZN(_03414_)
  );
  INV_X1 _08561_ (
    .A(_03414_),
    .ZN(_03415_)
  );
  AND2_X1 _08562_ (
    .A1(reg_mtvec[30]),
    .A2(_00940_),
    .ZN(_03416_)
  );
  INV_X1 _08563_ (
    .A(_03416_),
    .ZN(_03417_)
  );
  AND2_X1 _08564_ (
    .A1(reg_mcause[30]),
    .A2(_01001_),
    .ZN(_03418_)
  );
  INV_X1 _08565_ (
    .A(_03418_),
    .ZN(_03419_)
  );
  AND2_X1 _08566_ (
    .A1(reg_mscratch[30]),
    .A2(_00929_),
    .ZN(_03420_)
  );
  INV_X1 _08567_ (
    .A(_03420_),
    .ZN(_03421_)
  );
  AND2_X1 _08568_ (
    .A1(_01340_),
    .A2(_01382_),
    .ZN(_03422_)
  );
  AND2_X1 _08569_ (
    .A1(_03407_),
    .A2(_03415_),
    .ZN(_03423_)
  );
  AND2_X1 _08570_ (
    .A1(_03411_),
    .A2(_03423_),
    .ZN(_03424_)
  );
  AND2_X1 _08571_ (
    .A1(large_[24]),
    .A2(_01027_),
    .ZN(_03425_)
  );
  INV_X1 _08572_ (
    .A(_03425_),
    .ZN(_03426_)
  );
  AND2_X1 _08573_ (
    .A1(_03409_),
    .A2(_03413_),
    .ZN(_03427_)
  );
  AND2_X1 _08574_ (
    .A1(_03426_),
    .A2(_03427_),
    .ZN(_03428_)
  );
  AND2_X1 _08575_ (
    .A1(_03403_),
    .A2(_03428_),
    .ZN(_03429_)
  );
  AND2_X1 _08576_ (
    .A1(_03424_),
    .A2(_03429_),
    .ZN(_03430_)
  );
  AND2_X1 _08577_ (
    .A1(large_1[24]),
    .A2(_01029_),
    .ZN(_03431_)
  );
  INV_X1 _08578_ (
    .A(_03431_),
    .ZN(_03432_)
  );
  AND2_X1 _08579_ (
    .A1(_03419_),
    .A2(_03421_),
    .ZN(_03433_)
  );
  AND2_X1 _08580_ (
    .A1(_03432_),
    .A2(_03433_),
    .ZN(_03434_)
  );
  AND2_X1 _08581_ (
    .A1(_03417_),
    .A2(_03434_),
    .ZN(_03435_)
  );
  AND2_X1 _08582_ (
    .A1(_03405_),
    .A2(_03422_),
    .ZN(_03436_)
  );
  AND2_X1 _08583_ (
    .A1(_03435_),
    .A2(_03436_),
    .ZN(_03437_)
  );
  AND2_X1 _08584_ (
    .A1(_03430_),
    .A2(_03437_),
    .ZN(_03438_)
  );
  INV_X1 _08585_ (
    .A(_03438_),
    .ZN(io_rw_rdata[30])
  );
  AND2_X1 _08586_ (
    .A1(io_rw_cmd[1]),
    .A2(_00865_),
    .ZN(_03439_)
  );
  AND2_X1 _08587_ (
    .A1(io_rw_rdata[30]),
    .A2(_03439_),
    .ZN(_03440_)
  );
  INV_X1 _08588_ (
    .A(_03440_),
    .ZN(_03441_)
  );
  AND2_X1 _08589_ (
    .A1(_03401_),
    .A2(_03441_),
    .ZN(_03442_)
  );
  INV_X1 _08590_ (
    .A(_03442_),
    .ZN(_03443_)
  );
  MUX2_X1 _08591_ (
    .A(reg_bp_0_address[30]),
    .B(_03443_),
    .S(_03399_),
    .Z(_00237_)
  );
  MUX2_X1 _08592_ (
    .A(reg_bp_0_address[31]),
    .B(_03342_),
    .S(_03399_),
    .Z(_00238_)
  );
  AND2_X1 _08593_ (
    .A1(_00792_),
    .A2(_03233_),
    .ZN(_03444_)
  );
  INV_X1 _08594_ (
    .A(_03444_),
    .ZN(_03445_)
  );
  AND2_X1 _08595_ (
    .A1(_00811_),
    .A2(_03445_),
    .ZN(_03446_)
  );
  AND2_X1 _08596_ (
    .A1(_01864_),
    .A2(_03232_),
    .ZN(_03447_)
  );
  INV_X1 _08597_ (
    .A(_03447_),
    .ZN(_03448_)
  );
  AND2_X1 _08598_ (
    .A1(_03446_),
    .A2(_03448_),
    .ZN(_00239_)
  );
  AND2_X1 _08599_ (
    .A1(_00791_),
    .A2(_03233_),
    .ZN(_03449_)
  );
  INV_X1 _08600_ (
    .A(_03449_),
    .ZN(_03450_)
  );
  AND2_X1 _08601_ (
    .A1(_00811_),
    .A2(_03450_),
    .ZN(_03451_)
  );
  AND2_X1 _08602_ (
    .A1(_01937_),
    .A2(_03232_),
    .ZN(_03452_)
  );
  INV_X1 _08603_ (
    .A(_03452_),
    .ZN(_03453_)
  );
  AND2_X1 _08604_ (
    .A1(_03451_),
    .A2(_03453_),
    .ZN(_00240_)
  );
  AND2_X1 _08605_ (
    .A1(_00790_),
    .A2(_03233_),
    .ZN(_03454_)
  );
  INV_X1 _08606_ (
    .A(_03454_),
    .ZN(_03455_)
  );
  AND2_X1 _08607_ (
    .A1(_00811_),
    .A2(_03455_),
    .ZN(_03456_)
  );
  AND2_X1 _08608_ (
    .A1(_02162_),
    .A2(_03232_),
    .ZN(_03457_)
  );
  INV_X1 _08609_ (
    .A(_03457_),
    .ZN(_03458_)
  );
  AND2_X1 _08610_ (
    .A1(_03456_),
    .A2(_03458_),
    .ZN(_00241_)
  );
  AND2_X1 _08611_ (
    .A1(_01341_),
    .A2(_03398_),
    .ZN(_03459_)
  );
  INV_X1 _08612_ (
    .A(_03459_),
    .ZN(_03460_)
  );
  MUX2_X1 _08613_ (
    .A(reg_bp_0_control_tmatch[0]),
    .B(_02163_),
    .S(_03459_),
    .Z(_00242_)
  );
  MUX2_X1 _08614_ (
    .A(reg_bp_0_control_tmatch[1]),
    .B(_01446_),
    .S(_03459_),
    .Z(_00243_)
  );
  AND2_X1 _08615_ (
    .A1(_01612_),
    .A2(_03459_),
    .ZN(_03461_)
  );
  INV_X1 _08616_ (
    .A(_03461_),
    .ZN(_03462_)
  );
  AND2_X1 _08617_ (
    .A1(_00789_),
    .A2(_03460_),
    .ZN(_03463_)
  );
  INV_X1 _08618_ (
    .A(_03463_),
    .ZN(_03464_)
  );
  AND2_X1 _08619_ (
    .A1(_00811_),
    .A2(_03464_),
    .ZN(_03465_)
  );
  AND2_X1 _08620_ (
    .A1(_03462_),
    .A2(_03465_),
    .ZN(_00244_)
  );
  AND2_X1 _08621_ (
    .A1(_01687_),
    .A2(_03459_),
    .ZN(_03466_)
  );
  INV_X1 _08622_ (
    .A(_03466_),
    .ZN(_03467_)
  );
  AND2_X1 _08623_ (
    .A1(_00788_),
    .A2(_03460_),
    .ZN(_03468_)
  );
  INV_X1 _08624_ (
    .A(_03468_),
    .ZN(_03469_)
  );
  AND2_X1 _08625_ (
    .A1(_00811_),
    .A2(_03469_),
    .ZN(_03470_)
  );
  AND2_X1 _08626_ (
    .A1(_03467_),
    .A2(_03470_),
    .ZN(_00245_)
  );
  AND2_X1 _08627_ (
    .A1(_01773_),
    .A2(_03459_),
    .ZN(_03471_)
  );
  INV_X1 _08628_ (
    .A(_03471_),
    .ZN(_03472_)
  );
  AND2_X1 _08629_ (
    .A1(_00787_),
    .A2(_03460_),
    .ZN(_03473_)
  );
  INV_X1 _08630_ (
    .A(_03473_),
    .ZN(_03474_)
  );
  AND2_X1 _08631_ (
    .A1(_00811_),
    .A2(_03474_),
    .ZN(_03475_)
  );
  AND2_X1 _08632_ (
    .A1(_03472_),
    .A2(_03475_),
    .ZN(_00246_)
  );
  AND2_X1 _08633_ (
    .A1(reg_dcsr_step),
    .A2(_io_decode_0_read_illegal_T_15),
    .ZN(io_singleStep)
  );
  INV_X1 _08634_ (
    .A(io_singleStep),
    .ZN(_03476_)
  );
  AND2_X1 _08635_ (
    .A1(_00832_),
    .A2(_00833_),
    .ZN(_03477_)
  );
  AND2_X1 _08636_ (
    .A1(_00885_),
    .A2(_03477_),
    .ZN(_03478_)
  );
  AND2_X1 _08637_ (
    .A1(_00935_),
    .A2(_03478_),
    .ZN(_03479_)
  );
  AND2_X1 _08638_ (
    .A1(_00915_),
    .A2(_03479_),
    .ZN(_03480_)
  );
  AND2_X1 _08639_ (
    .A1(_01108_),
    .A2(_03480_),
    .ZN(_03481_)
  );
  INV_X1 _08640_ (
    .A(_03481_),
    .ZN(_03482_)
  );
  AND2_X1 _08641_ (
    .A1(_00884_),
    .A2(_03479_),
    .ZN(_03483_)
  );
  AND2_X1 _08642_ (
    .A1(_01108_),
    .A2(_03483_),
    .ZN(_03484_)
  );
  INV_X1 _08643_ (
    .A(_03484_),
    .ZN(_03485_)
  );
  AND2_X1 _08644_ (
    .A1(_03482_),
    .A2(_03485_),
    .ZN(_03486_)
  );
  AND2_X1 _08645_ (
    .A1(_00880_),
    .A2(_03486_),
    .ZN(_03487_)
  );
  INV_X1 _08646_ (
    .A(_03487_),
    .ZN(io_trace_0_exception)
  );
  AND2_X1 _08647_ (
    .A1(_00878_),
    .A2(_03487_),
    .ZN(_03488_)
  );
  INV_X1 _08648_ (
    .A(_03488_),
    .ZN(io_trace_0_valid)
  );
  AND2_X1 _08649_ (
    .A1(_00785_),
    .A2(_03488_),
    .ZN(_03489_)
  );
  INV_X1 _08650_ (
    .A(_03489_),
    .ZN(_03490_)
  );
  AND2_X1 _08651_ (
    .A1(io_singleStep),
    .A2(_03490_),
    .ZN(_00247_)
  );
  AND2_X1 _08652_ (
    .A1(reg_bp_0_control_action),
    .A2(_03460_),
    .ZN(_03491_)
  );
  INV_X1 _08653_ (
    .A(_03491_),
    .ZN(_03492_)
  );
  AND2_X1 _08654_ (
    .A1(reg_bp_0_control_dmode),
    .A2(io_rw_cmd[1]),
    .ZN(_03493_)
  );
  INV_X1 _08655_ (
    .A(_03493_),
    .ZN(_03494_)
  );
  AND2_X1 _08656_ (
    .A1(_00862_),
    .A2(_03494_),
    .ZN(_03495_)
  );
  INV_X1 _08657_ (
    .A(_03495_),
    .ZN(_03496_)
  );
  AND2_X1 _08658_ (
    .A1(reg_debug),
    .A2(_03088_),
    .ZN(_03497_)
  );
  AND2_X1 _08659_ (
    .A1(_03496_),
    .A2(_03497_),
    .ZN(_03498_)
  );
  AND2_X1 _08660_ (
    .A1(_03459_),
    .A2(_03498_),
    .ZN(_03499_)
  );
  AND2_X1 _08661_ (
    .A1(reg_bp_0_control_action),
    .A2(io_rw_cmd[1]),
    .ZN(_03500_)
  );
  MUX2_X1 _08662_ (
    .A(_03500_),
    .B(_00903_),
    .S(io_rw_wdata[12]),
    .Z(_03501_)
  );
  AND2_X1 _08663_ (
    .A1(_03499_),
    .A2(_03501_),
    .ZN(_03502_)
  );
  INV_X1 _08664_ (
    .A(_03502_),
    .ZN(_03503_)
  );
  AND2_X1 _08665_ (
    .A1(_03492_),
    .A2(_03503_),
    .ZN(_03504_)
  );
  INV_X1 _08666_ (
    .A(_03504_),
    .ZN(_03505_)
  );
  AND2_X1 _08667_ (
    .A1(_00811_),
    .A2(_03505_),
    .ZN(_00248_)
  );
  MUX2_X1 _08668_ (
    .A(reg_bp_0_control_dmode),
    .B(_03498_),
    .S(_03459_),
    .Z(_03506_)
  );
  AND2_X1 _08669_ (
    .A1(_00811_),
    .A2(_03506_),
    .ZN(_00249_)
  );
  AND2_X1 _08670_ (
    .A1(_00897_),
    .A2(_00958_),
    .ZN(_03507_)
  );
  MUX2_X1 _08671_ (
    .A(reg_dscratch0[0]),
    .B(_01613_),
    .S(_03507_),
    .Z(_00250_)
  );
  MUX2_X1 _08672_ (
    .A(reg_dscratch0[1]),
    .B(_01688_),
    .S(_03507_),
    .Z(_00251_)
  );
  MUX2_X1 _08673_ (
    .A(reg_dscratch0[2]),
    .B(_01774_),
    .S(_03507_),
    .Z(_00252_)
  );
  MUX2_X1 _08674_ (
    .A(reg_dscratch0[3]),
    .B(_01865_),
    .S(_03507_),
    .Z(_00253_)
  );
  MUX2_X1 _08675_ (
    .A(reg_dscratch0[4]),
    .B(_01938_),
    .S(_03507_),
    .Z(_00254_)
  );
  MUX2_X1 _08676_ (
    .A(reg_dscratch0[5]),
    .B(_02005_),
    .S(_03507_),
    .Z(_00255_)
  );
  MUX2_X1 _08677_ (
    .A(reg_dscratch0[6]),
    .B(_02076_),
    .S(_03507_),
    .Z(_00256_)
  );
  MUX2_X1 _08678_ (
    .A(reg_dscratch0[7]),
    .B(_02163_),
    .S(_03507_),
    .Z(_00257_)
  );
  MUX2_X1 _08679_ (
    .A(reg_dscratch0[8]),
    .B(_01446_),
    .S(_03507_),
    .Z(_00258_)
  );
  MUX2_X1 _08680_ (
    .A(reg_dscratch0[9]),
    .B(_01518_),
    .S(_03507_),
    .Z(_00259_)
  );
  MUX2_X1 _08681_ (
    .A(reg_dscratch0[10]),
    .B(_02235_),
    .S(_03507_),
    .Z(_00260_)
  );
  MUX2_X1 _08682_ (
    .A(reg_dscratch0[11]),
    .B(_02314_),
    .S(_03507_),
    .Z(_00261_)
  );
  MUX2_X1 _08683_ (
    .A(reg_dscratch0[12]),
    .B(_02389_),
    .S(_03507_),
    .Z(_00262_)
  );
  MUX2_X1 _08684_ (
    .A(reg_dscratch0[13]),
    .B(_02456_),
    .S(_03507_),
    .Z(_00263_)
  );
  MUX2_X1 _08685_ (
    .A(reg_dscratch0[14]),
    .B(_02522_),
    .S(_03507_),
    .Z(_00264_)
  );
  MUX2_X1 _08686_ (
    .A(reg_dscratch0[15]),
    .B(_02597_),
    .S(_03507_),
    .Z(_00265_)
  );
  MUX2_X1 _08687_ (
    .A(reg_dscratch0[16]),
    .B(_01035_),
    .S(_03507_),
    .Z(_00266_)
  );
  MUX2_X1 _08688_ (
    .A(reg_dscratch0[17]),
    .B(_02669_),
    .S(_03507_),
    .Z(_00267_)
  );
  MUX2_X1 _08689_ (
    .A(reg_dscratch0[18]),
    .B(_01107_),
    .S(_03507_),
    .Z(_00268_)
  );
  MUX2_X1 _08690_ (
    .A(reg_dscratch0[19]),
    .B(_01199_),
    .S(_03507_),
    .Z(_00269_)
  );
  MUX2_X1 _08691_ (
    .A(reg_dscratch0[20]),
    .B(_01277_),
    .S(_03507_),
    .Z(_00270_)
  );
  MUX2_X1 _08692_ (
    .A(reg_dscratch0[21]),
    .B(_02735_),
    .S(_03507_),
    .Z(_00271_)
  );
  MUX2_X1 _08693_ (
    .A(reg_dscratch0[22]),
    .B(_02801_),
    .S(_03507_),
    .Z(_00272_)
  );
  MUX2_X1 _08694_ (
    .A(reg_dscratch0[23]),
    .B(_01360_),
    .S(_03507_),
    .Z(_00273_)
  );
  MUX2_X1 _08695_ (
    .A(reg_dscratch0[24]),
    .B(_02873_),
    .S(_03507_),
    .Z(_00274_)
  );
  MUX2_X1 _08696_ (
    .A(reg_dscratch0[25]),
    .B(_02945_),
    .S(_03507_),
    .Z(_00275_)
  );
  MUX2_X1 _08697_ (
    .A(reg_dscratch0[26]),
    .B(_03017_),
    .S(_03507_),
    .Z(_00276_)
  );
  MUX2_X1 _08698_ (
    .A(reg_dscratch0[27]),
    .B(_03089_),
    .S(_03507_),
    .Z(_00277_)
  );
  MUX2_X1 _08699_ (
    .A(reg_dscratch0[28]),
    .B(_03162_),
    .S(_03507_),
    .Z(_00278_)
  );
  MUX2_X1 _08700_ (
    .A(reg_dscratch0[29]),
    .B(_03230_),
    .S(_03507_),
    .Z(_00279_)
  );
  MUX2_X1 _08701_ (
    .A(reg_dscratch0[30]),
    .B(_03443_),
    .S(_03507_),
    .Z(_00280_)
  );
  MUX2_X1 _08702_ (
    .A(reg_dscratch0[31]),
    .B(_03342_),
    .S(_03507_),
    .Z(_00281_)
  );
  AND2_X1 _08703_ (
    .A1(io_cause[5]),
    .A2(_03486_),
    .ZN(_03508_)
  );
  INV_X1 _08704_ (
    .A(_03508_),
    .ZN(_03509_)
  );
  AND2_X1 _08705_ (
    .A1(io_cause[7]),
    .A2(_03486_),
    .ZN(_03510_)
  );
  INV_X1 _08706_ (
    .A(_03510_),
    .ZN(_03511_)
  );
  AND2_X1 _08707_ (
    .A1(io_cause[6]),
    .A2(_03486_),
    .ZN(_03512_)
  );
  INV_X1 _08708_ (
    .A(_03512_),
    .ZN(_03513_)
  );
  AND2_X1 _08709_ (
    .A1(_03511_),
    .A2(_03513_),
    .ZN(_03514_)
  );
  AND2_X1 _08710_ (
    .A1(_03509_),
    .A2(_03514_),
    .ZN(_03515_)
  );
  AND2_X1 _08711_ (
    .A1(_00867_),
    .A2(_03486_),
    .ZN(_03516_)
  );
  INV_X1 _08712_ (
    .A(_03516_),
    .ZN(_03517_)
  );
  AND2_X1 _08713_ (
    .A1(io_cause[2]),
    .A2(_03486_),
    .ZN(_03518_)
  );
  AND2_X1 _08714_ (
    .A1(io_cause[3]),
    .A2(_03485_),
    .ZN(_03519_)
  );
  INV_X1 _08715_ (
    .A(_03519_),
    .ZN(_03520_)
  );
  AND2_X1 _08716_ (
    .A1(io_cause[1]),
    .A2(_00869_),
    .ZN(_03521_)
  );
  AND2_X1 _08717_ (
    .A1(_03519_),
    .A2(_03521_),
    .ZN(_03522_)
  );
  AND2_X1 _08718_ (
    .A1(_03518_),
    .A2(_03522_),
    .ZN(_03523_)
  );
  AND2_X1 _08719_ (
    .A1(_03482_),
    .A2(_03520_),
    .ZN(_03524_)
  );
  INV_X1 _08720_ (
    .A(_03524_),
    .ZN(_03525_)
  );
  AND2_X1 _08721_ (
    .A1(_03516_),
    .A2(_03523_),
    .ZN(_03526_)
  );
  AND2_X1 _08722_ (
    .A1(_03515_),
    .A2(_03526_),
    .ZN(_03527_)
  );
  INV_X1 _08723_ (
    .A(_03527_),
    .ZN(_03528_)
  );
  AND2_X1 _08724_ (
    .A1(_00785_),
    .A2(_00870_),
    .ZN(_03529_)
  );
  AND2_X1 _08725_ (
    .A1(reg_dcsr_ebreakm),
    .A2(_03484_),
    .ZN(_03530_)
  );
  INV_X1 _08726_ (
    .A(_03530_),
    .ZN(_03531_)
  );
  AND2_X1 _08727_ (
    .A1(_03529_),
    .A2(_03531_),
    .ZN(_03532_)
  );
  AND2_X1 _08728_ (
    .A1(_03528_),
    .A2(_03532_),
    .ZN(_03533_)
  );
  INV_X1 _08729_ (
    .A(_03533_),
    .ZN(_03534_)
  );
  AND2_X1 _08730_ (
    .A1(io_trace_0_exception),
    .A2(_03533_),
    .ZN(_03535_)
  );
  INV_X1 _08731_ (
    .A(_03535_),
    .ZN(_03536_)
  );
  AND2_X1 _08732_ (
    .A1(_00870_),
    .A2(_03487_),
    .ZN(_03537_)
  );
  INV_X1 _08733_ (
    .A(_03537_),
    .ZN(_03538_)
  );
  AND2_X1 _08734_ (
    .A1(_00882_),
    .A2(_00936_),
    .ZN(_03539_)
  );
  INV_X1 _08735_ (
    .A(_03539_),
    .ZN(_03540_)
  );
  AND2_X1 _08736_ (
    .A1(_00909_),
    .A2(_03540_),
    .ZN(_03541_)
  );
  INV_X1 _08737_ (
    .A(_03541_),
    .ZN(_03542_)
  );
  AND2_X1 _08738_ (
    .A1(_01108_),
    .A2(_03542_),
    .ZN(_03543_)
  );
  INV_X1 _08739_ (
    .A(_03543_),
    .ZN(_03544_)
  );
  AND2_X1 _08740_ (
    .A1(io_rw_addr[10]),
    .A2(io_rw_addr[7]),
    .ZN(_03545_)
  );
  INV_X1 _08741_ (
    .A(_03545_),
    .ZN(_03546_)
  );
  AND2_X1 _08742_ (
    .A1(_03543_),
    .A2(_03545_),
    .ZN(_03547_)
  );
  INV_X1 _08743_ (
    .A(_03547_),
    .ZN(_03548_)
  );
  AND2_X1 _08744_ (
    .A1(_03538_),
    .A2(_03548_),
    .ZN(_03549_)
  );
  AND2_X1 _08745_ (
    .A1(_00811_),
    .A2(_03549_),
    .ZN(_03550_)
  );
  AND2_X1 _08746_ (
    .A1(_03536_),
    .A2(_03550_),
    .ZN(_00282_)
  );
  AND2_X1 _08747_ (
    .A1(_03543_),
    .A2(_03546_),
    .ZN(_03551_)
  );
  INV_X1 _08748_ (
    .A(_03551_),
    .ZN(_03552_)
  );
  AND2_X1 _08749_ (
    .A1(reg_mstatus_mie),
    .A2(_03552_),
    .ZN(_03553_)
  );
  AND2_X1 _08750_ (
    .A1(_03536_),
    .A2(_03553_),
    .ZN(_03554_)
  );
  INV_X1 _08751_ (
    .A(_03554_),
    .ZN(_03555_)
  );
  AND2_X1 _08752_ (
    .A1(_00897_),
    .A2(_01813_),
    .ZN(_03556_)
  );
  INV_X1 _08753_ (
    .A(_03556_),
    .ZN(_03557_)
  );
  AND2_X1 _08754_ (
    .A1(reg_mstatus_mpie),
    .A2(_03551_),
    .ZN(_03558_)
  );
  INV_X1 _08755_ (
    .A(_03558_),
    .ZN(_03559_)
  );
  AND2_X1 _08756_ (
    .A1(_03552_),
    .A2(_03557_),
    .ZN(_03560_)
  );
  AND2_X1 _08757_ (
    .A1(_03557_),
    .A2(_03559_),
    .ZN(_03561_)
  );
  AND2_X1 _08758_ (
    .A1(_03555_),
    .A2(_03561_),
    .ZN(_03562_)
  );
  INV_X1 _08759_ (
    .A(_03562_),
    .ZN(_03563_)
  );
  AND2_X1 _08760_ (
    .A1(_01864_),
    .A2(_03556_),
    .ZN(_03564_)
  );
  INV_X1 _08761_ (
    .A(_03564_),
    .ZN(_03565_)
  );
  AND2_X1 _08762_ (
    .A1(_00811_),
    .A2(_03565_),
    .ZN(_03566_)
  );
  AND2_X1 _08763_ (
    .A1(_03563_),
    .A2(_03566_),
    .ZN(_00283_)
  );
  AND2_X1 _08764_ (
    .A1(_00897_),
    .A2(_01381_),
    .ZN(_03567_)
  );
  INV_X1 _08765_ (
    .A(_03567_),
    .ZN(_03568_)
  );
  AND2_X1 _08766_ (
    .A1(_01773_),
    .A2(_03567_),
    .ZN(_03569_)
  );
  INV_X1 _08767_ (
    .A(_03569_),
    .ZN(_03570_)
  );
  AND2_X1 _08768_ (
    .A1(_00786_),
    .A2(_03568_),
    .ZN(_03571_)
  );
  INV_X1 _08769_ (
    .A(_03571_),
    .ZN(_03572_)
  );
  AND2_X1 _08770_ (
    .A1(_00811_),
    .A2(_03572_),
    .ZN(_03573_)
  );
  AND2_X1 _08771_ (
    .A1(_03570_),
    .A2(_03573_),
    .ZN(_00284_)
  );
  AND2_X1 _08772_ (
    .A1(_io_decode_0_read_illegal_T_15),
    .A2(io_trace_0_exception),
    .ZN(_03574_)
  );
  AND2_X1 _08773_ (
    .A1(_03534_),
    .A2(_03574_),
    .ZN(_03575_)
  );
  INV_X1 _08774_ (
    .A(_03575_),
    .ZN(_03576_)
  );
  AND2_X1 _08775_ (
    .A1(io_cause[31]),
    .A2(_03486_),
    .ZN(_03577_)
  );
  INV_X1 _08776_ (
    .A(_03577_),
    .ZN(_03578_)
  );
  AND2_X1 _08777_ (
    .A1(_03527_),
    .A2(_03578_),
    .ZN(_03579_)
  );
  INV_X1 _08778_ (
    .A(_03579_),
    .ZN(_03580_)
  );
  AND2_X1 _08779_ (
    .A1(_00785_),
    .A2(_03580_),
    .ZN(_03581_)
  );
  MUX2_X1 _08780_ (
    .A(reg_dcsr_cause[0]),
    .B(_03581_),
    .S(_03575_),
    .Z(_03582_)
  );
  AND2_X1 _08781_ (
    .A1(_00811_),
    .A2(_03582_),
    .ZN(_00285_)
  );
  AND2_X1 _08782_ (
    .A1(reg_dcsr_cause[1]),
    .A2(_03576_),
    .ZN(_03583_)
  );
  INV_X1 _08783_ (
    .A(_03583_),
    .ZN(_03584_)
  );
  AND2_X1 _08784_ (
    .A1(_03527_),
    .A2(_03574_),
    .ZN(_03585_)
  );
  AND2_X1 _08785_ (
    .A1(_00785_),
    .A2(_03585_),
    .ZN(_03586_)
  );
  INV_X1 _08786_ (
    .A(_03586_),
    .ZN(_03587_)
  );
  AND2_X1 _08787_ (
    .A1(_03584_),
    .A2(_03587_),
    .ZN(_03588_)
  );
  INV_X1 _08788_ (
    .A(_03588_),
    .ZN(_03589_)
  );
  AND2_X1 _08789_ (
    .A1(_00811_),
    .A2(_03589_),
    .ZN(_00286_)
  );
  MUX2_X1 _08790_ (
    .A(reg_dcsr_cause[2]),
    .B(reg_singleStepped),
    .S(_03575_),
    .Z(_03590_)
  );
  AND2_X1 _08791_ (
    .A1(_00811_),
    .A2(_03590_),
    .ZN(_00287_)
  );
  AND2_X1 _08792_ (
    .A1(_02596_),
    .A2(_03567_),
    .ZN(_03591_)
  );
  INV_X1 _08793_ (
    .A(_03591_),
    .ZN(_03592_)
  );
  AND2_X1 _08794_ (
    .A1(_00784_),
    .A2(_03568_),
    .ZN(_03593_)
  );
  INV_X1 _08795_ (
    .A(_03593_),
    .ZN(_03594_)
  );
  AND2_X1 _08796_ (
    .A1(_00811_),
    .A2(_03594_),
    .ZN(_03595_)
  );
  AND2_X1 _08797_ (
    .A1(_03592_),
    .A2(_03595_),
    .ZN(_00288_)
  );
  MUX2_X1 _08798_ (
    .A(reg_mstatus_mpie),
    .B(reg_mstatus_mie),
    .S(_03535_),
    .Z(_03596_)
  );
  INV_X1 _08799_ (
    .A(_03596_),
    .ZN(_03597_)
  );
  AND2_X1 _08800_ (
    .A1(_03560_),
    .A2(_03597_),
    .ZN(_03598_)
  );
  INV_X1 _08801_ (
    .A(_03598_),
    .ZN(_03599_)
  );
  AND2_X1 _08802_ (
    .A1(_02162_),
    .A2(_03556_),
    .ZN(_03600_)
  );
  INV_X1 _08803_ (
    .A(_03600_),
    .ZN(_03601_)
  );
  AND2_X1 _08804_ (
    .A1(_00811_),
    .A2(_03601_),
    .ZN(_03602_)
  );
  AND2_X1 _08805_ (
    .A1(_03599_),
    .A2(_03602_),
    .ZN(_00289_)
  );
  AND2_X1 _08806_ (
    .A1(_00897_),
    .A2(_01607_),
    .ZN(_03603_)
  );
  INV_X1 _08807_ (
    .A(_03603_),
    .ZN(_03604_)
  );
  AND2_X1 _08808_ (
    .A1(_00783_),
    .A2(_03604_),
    .ZN(_03605_)
  );
  INV_X1 _08809_ (
    .A(_03605_),
    .ZN(_03606_)
  );
  AND2_X1 _08810_ (
    .A1(_00811_),
    .A2(_03606_),
    .ZN(_03607_)
  );
  AND2_X1 _08811_ (
    .A1(_01612_),
    .A2(_03603_),
    .ZN(_03608_)
  );
  INV_X1 _08812_ (
    .A(_03608_),
    .ZN(_03609_)
  );
  AND2_X1 _08813_ (
    .A1(_03607_),
    .A2(_03609_),
    .ZN(_00290_)
  );
  AND2_X1 _08814_ (
    .A1(_00782_),
    .A2(_03604_),
    .ZN(_03610_)
  );
  INV_X1 _08815_ (
    .A(_03610_),
    .ZN(_03611_)
  );
  AND2_X1 _08816_ (
    .A1(_00811_),
    .A2(_03611_),
    .ZN(_03612_)
  );
  AND2_X1 _08817_ (
    .A1(_01773_),
    .A2(_03603_),
    .ZN(_03613_)
  );
  INV_X1 _08818_ (
    .A(_03613_),
    .ZN(_03614_)
  );
  AND2_X1 _08819_ (
    .A1(_03612_),
    .A2(_03614_),
    .ZN(_00291_)
  );
  AND2_X1 _08820_ (
    .A1(_00786_),
    .A2(_00833_),
    .ZN(_03615_)
  );
  AND2_X1 _08821_ (
    .A1(_io_decode_0_read_illegal_T_15),
    .A2(_03615_),
    .ZN(_03616_)
  );
  AND2_X1 _08822_ (
    .A1(_01108_),
    .A2(_03616_),
    .ZN(_03617_)
  );
  AND2_X1 _08823_ (
    .A1(_00887_),
    .A2(_03617_),
    .ZN(_03618_)
  );
  INV_X1 _08824_ (
    .A(_03618_),
    .ZN(_03619_)
  );
  AND2_X1 _08825_ (
    .A1(_00877_),
    .A2(_03619_),
    .ZN(_03620_)
  );
  INV_X1 _08826_ (
    .A(_03620_),
    .ZN(_03621_)
  );
  AND2_X1 _08827_ (
    .A1(_00811_),
    .A2(_00835_),
    .ZN(_03622_)
  );
  AND2_X1 _08828_ (
    .A1(reg_mie[7]),
    .A2(io_interrupts_mtip),
    .ZN(_03623_)
  );
  INV_X1 _08829_ (
    .A(_03623_),
    .ZN(_03624_)
  );
  AND2_X1 _08830_ (
    .A1(reg_mie[3]),
    .A2(io_interrupts_msip),
    .ZN(_03625_)
  );
  INV_X1 _08831_ (
    .A(_03625_),
    .ZN(_03626_)
  );
  AND2_X1 _08832_ (
    .A1(reg_mie[11]),
    .A2(io_interrupts_meip),
    .ZN(_03627_)
  );
  INV_X1 _08833_ (
    .A(_03627_),
    .ZN(_03628_)
  );
  AND2_X1 _08834_ (
    .A1(_03626_),
    .A2(_03628_),
    .ZN(_03629_)
  );
  INV_X1 _08835_ (
    .A(_03629_),
    .ZN(_03630_)
  );
  AND2_X1 _08836_ (
    .A1(_03624_),
    .A2(_03629_),
    .ZN(_03631_)
  );
  INV_X1 _08837_ (
    .A(_03631_),
    .ZN(_03632_)
  );
  AND2_X1 _08838_ (
    .A1(_03622_),
    .A2(_03631_),
    .ZN(_03633_)
  );
  AND2_X1 _08839_ (
    .A1(_03621_),
    .A2(_03633_),
    .ZN(_03634_)
  );
  AND2_X1 _08840_ (
    .A1(_03487_),
    .A2(_03634_),
    .ZN(_00292_)
  );
  MUX2_X1 _08841_ (
    .A(reg_mstatus_gva),
    .B(io_gva),
    .S(_03535_),
    .Z(_03635_)
  );
  AND2_X1 _08842_ (
    .A1(_00811_),
    .A2(_03635_),
    .ZN(_00293_)
  );
  AND2_X1 _08843_ (
    .A1(large_1[17]),
    .A2(large_1[16]),
    .ZN(_03636_)
  );
  AND2_X1 _08844_ (
    .A1(large_1[15]),
    .A2(_03636_),
    .ZN(_03637_)
  );
  AND2_X1 _08845_ (
    .A1(large_1[20]),
    .A2(large_1[19]),
    .ZN(_03638_)
  );
  AND2_X1 _08846_ (
    .A1(large_1[23]),
    .A2(large_1[22]),
    .ZN(_03639_)
  );
  AND2_X1 _08847_ (
    .A1(large_1[21]),
    .A2(large_1[18]),
    .ZN(_03640_)
  );
  AND2_X1 _08848_ (
    .A1(_03639_),
    .A2(_03640_),
    .ZN(_03641_)
  );
  AND2_X1 _08849_ (
    .A1(_03638_),
    .A2(_03641_),
    .ZN(_03642_)
  );
  AND2_X1 _08850_ (
    .A1(_03637_),
    .A2(_03642_),
    .ZN(_03643_)
  );
  AND2_X1 _08851_ (
    .A1(large_1[13]),
    .A2(large_1[12]),
    .ZN(_03644_)
  );
  AND2_X1 _08852_ (
    .A1(large_1[14]),
    .A2(_03644_),
    .ZN(_03645_)
  );
  AND2_X1 _08853_ (
    .A1(large_1[8]),
    .A2(large_1[7]),
    .ZN(_03646_)
  );
  AND2_X1 _08854_ (
    .A1(large_1[9]),
    .A2(_03646_),
    .ZN(_03647_)
  );
  AND2_X1 _08855_ (
    .A1(large_1[4]),
    .A2(large_1[3]),
    .ZN(_03648_)
  );
  AND2_X1 _08856_ (
    .A1(large_1[3]),
    .A2(large_1[2]),
    .ZN(_03649_)
  );
  AND2_X1 _08857_ (
    .A1(large_1[5]),
    .A2(large_1[4]),
    .ZN(_03650_)
  );
  AND2_X1 _08858_ (
    .A1(_03649_),
    .A2(_03650_),
    .ZN(_03651_)
  );
  AND2_X1 _08859_ (
    .A1(large_1[6]),
    .A2(_03651_),
    .ZN(_03652_)
  );
  AND2_X1 _08860_ (
    .A1(_00877_),
    .A2(_00879_),
    .ZN(_03653_)
  );
  INV_X1 _08861_ (
    .A(_03653_),
    .ZN(io_csr_stall)
  );
  AND2_X1 _08862_ (
    .A1(small_1[0]),
    .A2(_03653_),
    .ZN(_03654_)
  );
  AND2_X1 _08863_ (
    .A1(small_1[1]),
    .A2(_03654_),
    .ZN(_03655_)
  );
  AND2_X1 _08864_ (
    .A1(small_1[2]),
    .A2(_03655_),
    .ZN(_03656_)
  );
  AND2_X1 _08865_ (
    .A1(small_1[3]),
    .A2(_03656_),
    .ZN(_03657_)
  );
  AND2_X1 _08866_ (
    .A1(small_1[4]),
    .A2(_03657_),
    .ZN(_03658_)
  );
  AND2_X1 _08867_ (
    .A1(small_1[5]),
    .A2(_T_15),
    .ZN(_03659_)
  );
  AND2_X1 _08868_ (
    .A1(_03658_),
    .A2(_03659_),
    .ZN(_03660_)
  );
  AND2_X1 _08869_ (
    .A1(large_1[0]),
    .A2(_03660_),
    .ZN(_03661_)
  );
  INV_X1 _08870_ (
    .A(_03661_),
    .ZN(_03662_)
  );
  AND2_X1 _08871_ (
    .A1(large_1[1]),
    .A2(_03661_),
    .ZN(_03663_)
  );
  AND2_X1 _08872_ (
    .A1(_03652_),
    .A2(_03663_),
    .ZN(_03664_)
  );
  AND2_X1 _08873_ (
    .A1(small_1[5]),
    .A2(_03658_),
    .ZN(_03665_)
  );
  AND2_X1 _08874_ (
    .A1(_T_15),
    .A2(_03665_),
    .ZN(_03666_)
  );
  AND2_X1 _08875_ (
    .A1(large_1[0]),
    .A2(_03666_),
    .ZN(_03667_)
  );
  AND2_X1 _08876_ (
    .A1(large_1[1]),
    .A2(_03667_),
    .ZN(_03668_)
  );
  INV_X1 _08877_ (
    .A(_03668_),
    .ZN(_03669_)
  );
  AND2_X1 _08878_ (
    .A1(_03652_),
    .A2(_03668_),
    .ZN(_03670_)
  );
  INV_X1 _08879_ (
    .A(_03670_),
    .ZN(_03671_)
  );
  AND2_X1 _08880_ (
    .A1(_03647_),
    .A2(_03670_),
    .ZN(_03672_)
  );
  INV_X1 _08881_ (
    .A(_03672_),
    .ZN(_03673_)
  );
  AND2_X1 _08882_ (
    .A1(large_1[10]),
    .A2(_03672_),
    .ZN(_03674_)
  );
  INV_X1 _08883_ (
    .A(_03674_),
    .ZN(_03675_)
  );
  AND2_X1 _08884_ (
    .A1(large_1[11]),
    .A2(_03674_),
    .ZN(_03676_)
  );
  INV_X1 _08885_ (
    .A(_03676_),
    .ZN(_03677_)
  );
  AND2_X1 _08886_ (
    .A1(_03645_),
    .A2(_03676_),
    .ZN(_03678_)
  );
  INV_X1 _08887_ (
    .A(_03678_),
    .ZN(_03679_)
  );
  AND2_X1 _08888_ (
    .A1(_03643_),
    .A2(_03678_),
    .ZN(_03680_)
  );
  AND2_X1 _08889_ (
    .A1(large_1[25]),
    .A2(large_1[24]),
    .ZN(_03681_)
  );
  AND2_X1 _08890_ (
    .A1(_03680_),
    .A2(_03681_),
    .ZN(_03682_)
  );
  AND2_X1 _08891_ (
    .A1(large_1[1]),
    .A2(large_1[0]),
    .ZN(_03683_)
  );
  AND2_X1 _08892_ (
    .A1(_03649_),
    .A2(_03683_),
    .ZN(_03684_)
  );
  AND2_X1 _08893_ (
    .A1(large_1[6]),
    .A2(_03650_),
    .ZN(_03685_)
  );
  AND2_X1 _08894_ (
    .A1(_03666_),
    .A2(_03685_),
    .ZN(_03686_)
  );
  AND2_X1 _08895_ (
    .A1(_03684_),
    .A2(_03686_),
    .ZN(_03687_)
  );
  AND2_X1 _08896_ (
    .A1(_03647_),
    .A2(_03687_),
    .ZN(_03688_)
  );
  AND2_X1 _08897_ (
    .A1(large_1[10]),
    .A2(_03688_),
    .ZN(_03689_)
  );
  AND2_X1 _08898_ (
    .A1(large_1[11]),
    .A2(_03689_),
    .ZN(_03690_)
  );
  AND2_X1 _08899_ (
    .A1(_03645_),
    .A2(_03690_),
    .ZN(_03691_)
  );
  AND2_X1 _08900_ (
    .A1(_03643_),
    .A2(_03691_),
    .ZN(_03692_)
  );
  INV_X1 _08901_ (
    .A(_03692_),
    .ZN(_03693_)
  );
  AND2_X1 _08902_ (
    .A1(large_1[24]),
    .A2(_03692_),
    .ZN(_03694_)
  );
  INV_X1 _08903_ (
    .A(_03694_),
    .ZN(_03695_)
  );
  AND2_X1 _08904_ (
    .A1(large_1[25]),
    .A2(_03694_),
    .ZN(_03696_)
  );
  INV_X1 _08905_ (
    .A(_03696_),
    .ZN(_03697_)
  );
  AND2_X1 _08906_ (
    .A1(_00781_),
    .A2(_03697_),
    .ZN(_03698_)
  );
  INV_X1 _08907_ (
    .A(_03698_),
    .ZN(_03699_)
  );
  AND2_X1 _08908_ (
    .A1(_00897_),
    .A2(_01019_),
    .ZN(_03700_)
  );
  INV_X1 _08909_ (
    .A(_03700_),
    .ZN(_03701_)
  );
  AND2_X1 _08910_ (
    .A1(_00897_),
    .A2(_00995_),
    .ZN(_03702_)
  );
  INV_X1 _08911_ (
    .A(_03702_),
    .ZN(_03703_)
  );
  AND2_X1 _08912_ (
    .A1(_00897_),
    .A2(_01020_),
    .ZN(_03704_)
  );
  AND2_X1 _08913_ (
    .A1(_00996_),
    .A2(_03704_),
    .ZN(_03705_)
  );
  AND2_X1 _08914_ (
    .A1(_03701_),
    .A2(_03703_),
    .ZN(_03706_)
  );
  AND2_X1 _08915_ (
    .A1(large_1[26]),
    .A2(_03682_),
    .ZN(_03707_)
  );
  AND2_X1 _08916_ (
    .A1(_00897_),
    .A2(_01029_),
    .ZN(_03708_)
  );
  INV_X1 _08917_ (
    .A(_03708_),
    .ZN(_03709_)
  );
  AND2_X1 _08918_ (
    .A1(_03701_),
    .A2(_03709_),
    .ZN(_03710_)
  );
  AND2_X1 _08919_ (
    .A1(large_1[26]),
    .A2(_03696_),
    .ZN(_03711_)
  );
  INV_X1 _08920_ (
    .A(_03711_),
    .ZN(_03712_)
  );
  AND2_X1 _08921_ (
    .A1(_03710_),
    .A2(_03712_),
    .ZN(_03713_)
  );
  AND2_X1 _08922_ (
    .A1(_03699_),
    .A2(_03713_),
    .ZN(_03714_)
  );
  INV_X1 _08923_ (
    .A(_03714_),
    .ZN(_03715_)
  );
  AND2_X1 _08924_ (
    .A1(_01613_),
    .A2(_03700_),
    .ZN(_03716_)
  );
  INV_X1 _08925_ (
    .A(_03716_),
    .ZN(_03717_)
  );
  AND2_X1 _08926_ (
    .A1(large_1[26]),
    .A2(_03702_),
    .ZN(_03718_)
  );
  INV_X1 _08927_ (
    .A(_03718_),
    .ZN(_03719_)
  );
  AND2_X1 _08928_ (
    .A1(_03717_),
    .A2(_03719_),
    .ZN(_03720_)
  );
  AND2_X1 _08929_ (
    .A1(_03715_),
    .A2(_03720_),
    .ZN(_03721_)
  );
  INV_X1 _08930_ (
    .A(_03721_),
    .ZN(_03722_)
  );
  AND2_X1 _08931_ (
    .A1(_00811_),
    .A2(_03722_),
    .ZN(_00294_)
  );
  AND2_X1 _08932_ (
    .A1(_00780_),
    .A2(_03712_),
    .ZN(_03723_)
  );
  INV_X1 _08933_ (
    .A(_03723_),
    .ZN(_03724_)
  );
  AND2_X1 _08934_ (
    .A1(large_1[27]),
    .A2(large_1[26]),
    .ZN(_03725_)
  );
  AND2_X1 _08935_ (
    .A1(large_1[27]),
    .A2(_03707_),
    .ZN(_03726_)
  );
  AND2_X1 _08936_ (
    .A1(_03681_),
    .A2(_03725_),
    .ZN(_03727_)
  );
  AND2_X1 _08937_ (
    .A1(_03692_),
    .A2(_03727_),
    .ZN(_03728_)
  );
  INV_X1 _08938_ (
    .A(_03728_),
    .ZN(_03729_)
  );
  AND2_X1 _08939_ (
    .A1(_03724_),
    .A2(_03729_),
    .ZN(_03730_)
  );
  AND2_X1 _08940_ (
    .A1(_03710_),
    .A2(_03730_),
    .ZN(_03731_)
  );
  INV_X1 _08941_ (
    .A(_03731_),
    .ZN(_03732_)
  );
  AND2_X1 _08942_ (
    .A1(_01688_),
    .A2(_03700_),
    .ZN(_03733_)
  );
  INV_X1 _08943_ (
    .A(_03733_),
    .ZN(_03734_)
  );
  AND2_X1 _08944_ (
    .A1(large_1[27]),
    .A2(_03702_),
    .ZN(_03735_)
  );
  INV_X1 _08945_ (
    .A(_03735_),
    .ZN(_03736_)
  );
  AND2_X1 _08946_ (
    .A1(_03734_),
    .A2(_03736_),
    .ZN(_03737_)
  );
  AND2_X1 _08947_ (
    .A1(_03732_),
    .A2(_03737_),
    .ZN(_03738_)
  );
  INV_X1 _08948_ (
    .A(_03738_),
    .ZN(_03739_)
  );
  AND2_X1 _08949_ (
    .A1(_00811_),
    .A2(_03739_),
    .ZN(_00295_)
  );
  AND2_X1 _08950_ (
    .A1(_00779_),
    .A2(_03729_),
    .ZN(_03740_)
  );
  INV_X1 _08951_ (
    .A(_03740_),
    .ZN(_03741_)
  );
  AND2_X1 _08952_ (
    .A1(_03710_),
    .A2(_03741_),
    .ZN(_03742_)
  );
  AND2_X1 _08953_ (
    .A1(large_1[28]),
    .A2(_03728_),
    .ZN(_03743_)
  );
  INV_X1 _08954_ (
    .A(_03743_),
    .ZN(_03744_)
  );
  AND2_X1 _08955_ (
    .A1(_03742_),
    .A2(_03744_),
    .ZN(_03745_)
  );
  INV_X1 _08956_ (
    .A(_03745_),
    .ZN(_03746_)
  );
  AND2_X1 _08957_ (
    .A1(_01774_),
    .A2(_03700_),
    .ZN(_03747_)
  );
  INV_X1 _08958_ (
    .A(_03747_),
    .ZN(_03748_)
  );
  AND2_X1 _08959_ (
    .A1(large_1[28]),
    .A2(_03702_),
    .ZN(_03749_)
  );
  INV_X1 _08960_ (
    .A(_03749_),
    .ZN(_03750_)
  );
  AND2_X1 _08961_ (
    .A1(_03748_),
    .A2(_03750_),
    .ZN(_03751_)
  );
  AND2_X1 _08962_ (
    .A1(_03746_),
    .A2(_03751_),
    .ZN(_03752_)
  );
  INV_X1 _08963_ (
    .A(_03752_),
    .ZN(_03753_)
  );
  AND2_X1 _08964_ (
    .A1(_00811_),
    .A2(_03753_),
    .ZN(_00296_)
  );
  AND2_X1 _08965_ (
    .A1(_00778_),
    .A2(_03744_),
    .ZN(_03754_)
  );
  INV_X1 _08966_ (
    .A(_03754_),
    .ZN(_03755_)
  );
  AND2_X1 _08967_ (
    .A1(large_1[29]),
    .A2(large_1[28]),
    .ZN(_03756_)
  );
  AND2_X1 _08968_ (
    .A1(_03726_),
    .A2(_03756_),
    .ZN(_03757_)
  );
  AND2_X1 _08969_ (
    .A1(large_1[29]),
    .A2(_03743_),
    .ZN(_03758_)
  );
  INV_X1 _08970_ (
    .A(_03758_),
    .ZN(_03759_)
  );
  AND2_X1 _08971_ (
    .A1(_03710_),
    .A2(_03759_),
    .ZN(_03760_)
  );
  AND2_X1 _08972_ (
    .A1(_03755_),
    .A2(_03760_),
    .ZN(_03761_)
  );
  INV_X1 _08973_ (
    .A(_03761_),
    .ZN(_03762_)
  );
  AND2_X1 _08974_ (
    .A1(_01865_),
    .A2(_03700_),
    .ZN(_03763_)
  );
  INV_X1 _08975_ (
    .A(_03763_),
    .ZN(_03764_)
  );
  AND2_X1 _08976_ (
    .A1(large_1[29]),
    .A2(_03708_),
    .ZN(_03765_)
  );
  INV_X1 _08977_ (
    .A(_03765_),
    .ZN(_03766_)
  );
  AND2_X1 _08978_ (
    .A1(_03764_),
    .A2(_03766_),
    .ZN(_03767_)
  );
  AND2_X1 _08979_ (
    .A1(_03762_),
    .A2(_03767_),
    .ZN(_03768_)
  );
  INV_X1 _08980_ (
    .A(_03768_),
    .ZN(_03769_)
  );
  AND2_X1 _08981_ (
    .A1(_00811_),
    .A2(_03769_),
    .ZN(_00297_)
  );
  AND2_X1 _08982_ (
    .A1(_00777_),
    .A2(_03759_),
    .ZN(_03770_)
  );
  INV_X1 _08983_ (
    .A(_03770_),
    .ZN(_03771_)
  );
  AND2_X1 _08984_ (
    .A1(large_1[30]),
    .A2(_03757_),
    .ZN(_03772_)
  );
  AND2_X1 _08985_ (
    .A1(large_1[30]),
    .A2(_03758_),
    .ZN(_03773_)
  );
  INV_X1 _08986_ (
    .A(_03773_),
    .ZN(_03774_)
  );
  AND2_X1 _08987_ (
    .A1(_03771_),
    .A2(_03774_),
    .ZN(_03775_)
  );
  AND2_X1 _08988_ (
    .A1(_03710_),
    .A2(_03775_),
    .ZN(_03776_)
  );
  INV_X1 _08989_ (
    .A(_03776_),
    .ZN(_03777_)
  );
  AND2_X1 _08990_ (
    .A1(_01938_),
    .A2(_03700_),
    .ZN(_03778_)
  );
  INV_X1 _08991_ (
    .A(_03778_),
    .ZN(_03779_)
  );
  AND2_X1 _08992_ (
    .A1(large_1[30]),
    .A2(_03702_),
    .ZN(_03780_)
  );
  INV_X1 _08993_ (
    .A(_03780_),
    .ZN(_03781_)
  );
  AND2_X1 _08994_ (
    .A1(_03779_),
    .A2(_03781_),
    .ZN(_03782_)
  );
  AND2_X1 _08995_ (
    .A1(_03777_),
    .A2(_03782_),
    .ZN(_03783_)
  );
  INV_X1 _08996_ (
    .A(_03783_),
    .ZN(_03784_)
  );
  AND2_X1 _08997_ (
    .A1(_00811_),
    .A2(_03784_),
    .ZN(_00298_)
  );
  AND2_X1 _08998_ (
    .A1(_00776_),
    .A2(_03774_),
    .ZN(_03785_)
  );
  INV_X1 _08999_ (
    .A(_03785_),
    .ZN(_03786_)
  );
  AND2_X1 _09000_ (
    .A1(large_1[31]),
    .A2(large_1[30]),
    .ZN(_03787_)
  );
  AND2_X1 _09001_ (
    .A1(large_1[31]),
    .A2(_03772_),
    .ZN(_03788_)
  );
  INV_X1 _09002_ (
    .A(_03788_),
    .ZN(_03789_)
  );
  AND2_X1 _09003_ (
    .A1(_03710_),
    .A2(_03789_),
    .ZN(_03790_)
  );
  AND2_X1 _09004_ (
    .A1(_03786_),
    .A2(_03790_),
    .ZN(_03791_)
  );
  INV_X1 _09005_ (
    .A(_03791_),
    .ZN(_03792_)
  );
  AND2_X1 _09006_ (
    .A1(_02005_),
    .A2(_03700_),
    .ZN(_03793_)
  );
  INV_X1 _09007_ (
    .A(_03793_),
    .ZN(_03794_)
  );
  AND2_X1 _09008_ (
    .A1(large_1[31]),
    .A2(_03702_),
    .ZN(_03795_)
  );
  INV_X1 _09009_ (
    .A(_03795_),
    .ZN(_03796_)
  );
  AND2_X1 _09010_ (
    .A1(_03794_),
    .A2(_03796_),
    .ZN(_03797_)
  );
  AND2_X1 _09011_ (
    .A1(_03792_),
    .A2(_03797_),
    .ZN(_03798_)
  );
  INV_X1 _09012_ (
    .A(_03798_),
    .ZN(_03799_)
  );
  AND2_X1 _09013_ (
    .A1(_00811_),
    .A2(_03799_),
    .ZN(_00299_)
  );
  AND2_X1 _09014_ (
    .A1(_03756_),
    .A2(_03787_),
    .ZN(_03800_)
  );
  AND2_X1 _09015_ (
    .A1(_00775_),
    .A2(_03789_),
    .ZN(_03801_)
  );
  INV_X1 _09016_ (
    .A(_03801_),
    .ZN(_03802_)
  );
  AND2_X1 _09017_ (
    .A1(large_1[32]),
    .A2(_03788_),
    .ZN(_03803_)
  );
  INV_X1 _09018_ (
    .A(_03803_),
    .ZN(_03804_)
  );
  AND2_X1 _09019_ (
    .A1(_03710_),
    .A2(_03804_),
    .ZN(_03805_)
  );
  AND2_X1 _09020_ (
    .A1(_03802_),
    .A2(_03805_),
    .ZN(_03806_)
  );
  INV_X1 _09021_ (
    .A(_03806_),
    .ZN(_03807_)
  );
  AND2_X1 _09022_ (
    .A1(_02076_),
    .A2(_03700_),
    .ZN(_03808_)
  );
  INV_X1 _09023_ (
    .A(_03808_),
    .ZN(_03809_)
  );
  AND2_X1 _09024_ (
    .A1(large_1[32]),
    .A2(_03702_),
    .ZN(_03810_)
  );
  INV_X1 _09025_ (
    .A(_03810_),
    .ZN(_03811_)
  );
  AND2_X1 _09026_ (
    .A1(_03809_),
    .A2(_03811_),
    .ZN(_03812_)
  );
  AND2_X1 _09027_ (
    .A1(_03807_),
    .A2(_03812_),
    .ZN(_03813_)
  );
  INV_X1 _09028_ (
    .A(_03813_),
    .ZN(_03814_)
  );
  AND2_X1 _09029_ (
    .A1(_00811_),
    .A2(_03814_),
    .ZN(_00300_)
  );
  AND2_X1 _09030_ (
    .A1(_00774_),
    .A2(_03804_),
    .ZN(_03815_)
  );
  INV_X1 _09031_ (
    .A(_03815_),
    .ZN(_03816_)
  );
  AND2_X1 _09032_ (
    .A1(_03710_),
    .A2(_03816_),
    .ZN(_03817_)
  );
  AND2_X1 _09033_ (
    .A1(large_1[33]),
    .A2(_03803_),
    .ZN(_03818_)
  );
  INV_X1 _09034_ (
    .A(_03818_),
    .ZN(_03819_)
  );
  AND2_X1 _09035_ (
    .A1(_03817_),
    .A2(_03819_),
    .ZN(_03820_)
  );
  INV_X1 _09036_ (
    .A(_03820_),
    .ZN(_03821_)
  );
  AND2_X1 _09037_ (
    .A1(_02163_),
    .A2(_03700_),
    .ZN(_03822_)
  );
  INV_X1 _09038_ (
    .A(_03822_),
    .ZN(_03823_)
  );
  AND2_X1 _09039_ (
    .A1(large_1[33]),
    .A2(_03708_),
    .ZN(_03824_)
  );
  INV_X1 _09040_ (
    .A(_03824_),
    .ZN(_03825_)
  );
  AND2_X1 _09041_ (
    .A1(_03823_),
    .A2(_03825_),
    .ZN(_03826_)
  );
  AND2_X1 _09042_ (
    .A1(_03821_),
    .A2(_03826_),
    .ZN(_03827_)
  );
  INV_X1 _09043_ (
    .A(_03827_),
    .ZN(_03828_)
  );
  AND2_X1 _09044_ (
    .A1(_00811_),
    .A2(_03828_),
    .ZN(_00301_)
  );
  AND2_X1 _09045_ (
    .A1(_00773_),
    .A2(_03819_),
    .ZN(_03829_)
  );
  INV_X1 _09046_ (
    .A(_03829_),
    .ZN(_03830_)
  );
  AND2_X1 _09047_ (
    .A1(large_1[34]),
    .A2(_03818_),
    .ZN(_03831_)
  );
  INV_X1 _09048_ (
    .A(_03831_),
    .ZN(_03832_)
  );
  AND2_X1 _09049_ (
    .A1(_03710_),
    .A2(_03832_),
    .ZN(_03833_)
  );
  AND2_X1 _09050_ (
    .A1(large_1[34]),
    .A2(large_1[33]),
    .ZN(_03834_)
  );
  AND2_X1 _09051_ (
    .A1(_03830_),
    .A2(_03833_),
    .ZN(_03835_)
  );
  INV_X1 _09052_ (
    .A(_03835_),
    .ZN(_03836_)
  );
  AND2_X1 _09053_ (
    .A1(_01446_),
    .A2(_03700_),
    .ZN(_03837_)
  );
  INV_X1 _09054_ (
    .A(_03837_),
    .ZN(_03838_)
  );
  AND2_X1 _09055_ (
    .A1(large_1[34]),
    .A2(_03702_),
    .ZN(_03839_)
  );
  INV_X1 _09056_ (
    .A(_03839_),
    .ZN(_03840_)
  );
  AND2_X1 _09057_ (
    .A1(_03838_),
    .A2(_03840_),
    .ZN(_03841_)
  );
  AND2_X1 _09058_ (
    .A1(_03836_),
    .A2(_03841_),
    .ZN(_03842_)
  );
  INV_X1 _09059_ (
    .A(_03842_),
    .ZN(_03843_)
  );
  AND2_X1 _09060_ (
    .A1(_00811_),
    .A2(_03843_),
    .ZN(_00302_)
  );
  AND2_X1 _09061_ (
    .A1(_00772_),
    .A2(_03832_),
    .ZN(_03844_)
  );
  INV_X1 _09062_ (
    .A(_03844_),
    .ZN(_03845_)
  );
  AND2_X1 _09063_ (
    .A1(large_1[35]),
    .A2(_03834_),
    .ZN(_03846_)
  );
  AND2_X1 _09064_ (
    .A1(_03803_),
    .A2(_03846_),
    .ZN(_03847_)
  );
  INV_X1 _09065_ (
    .A(_03847_),
    .ZN(_03848_)
  );
  AND2_X1 _09066_ (
    .A1(_03710_),
    .A2(_03848_),
    .ZN(_03849_)
  );
  AND2_X1 _09067_ (
    .A1(_03845_),
    .A2(_03849_),
    .ZN(_03850_)
  );
  INV_X1 _09068_ (
    .A(_03850_),
    .ZN(_03851_)
  );
  AND2_X1 _09069_ (
    .A1(_01518_),
    .A2(_03700_),
    .ZN(_03852_)
  );
  INV_X1 _09070_ (
    .A(_03852_),
    .ZN(_03853_)
  );
  AND2_X1 _09071_ (
    .A1(large_1[35]),
    .A2(_03702_),
    .ZN(_03854_)
  );
  INV_X1 _09072_ (
    .A(_03854_),
    .ZN(_03855_)
  );
  AND2_X1 _09073_ (
    .A1(_03853_),
    .A2(_03855_),
    .ZN(_03856_)
  );
  AND2_X1 _09074_ (
    .A1(_03851_),
    .A2(_03856_),
    .ZN(_03857_)
  );
  INV_X1 _09075_ (
    .A(_03857_),
    .ZN(_03858_)
  );
  AND2_X1 _09076_ (
    .A1(_00811_),
    .A2(_03858_),
    .ZN(_00303_)
  );
  AND2_X1 _09077_ (
    .A1(_00771_),
    .A2(_03848_),
    .ZN(_03859_)
  );
  INV_X1 _09078_ (
    .A(_03859_),
    .ZN(_03860_)
  );
  AND2_X1 _09079_ (
    .A1(large_1[36]),
    .A2(_03847_),
    .ZN(_03861_)
  );
  INV_X1 _09080_ (
    .A(_03861_),
    .ZN(_03862_)
  );
  AND2_X1 _09081_ (
    .A1(_03710_),
    .A2(_03862_),
    .ZN(_03863_)
  );
  AND2_X1 _09082_ (
    .A1(_03860_),
    .A2(_03863_),
    .ZN(_03864_)
  );
  INV_X1 _09083_ (
    .A(_03864_),
    .ZN(_03865_)
  );
  AND2_X1 _09084_ (
    .A1(_02235_),
    .A2(_03700_),
    .ZN(_03866_)
  );
  INV_X1 _09085_ (
    .A(_03866_),
    .ZN(_03867_)
  );
  AND2_X1 _09086_ (
    .A1(large_1[36]),
    .A2(_03702_),
    .ZN(_03868_)
  );
  INV_X1 _09087_ (
    .A(_03868_),
    .ZN(_03869_)
  );
  AND2_X1 _09088_ (
    .A1(_03867_),
    .A2(_03869_),
    .ZN(_03870_)
  );
  AND2_X1 _09089_ (
    .A1(_03865_),
    .A2(_03870_),
    .ZN(_03871_)
  );
  INV_X1 _09090_ (
    .A(_03871_),
    .ZN(_03872_)
  );
  AND2_X1 _09091_ (
    .A1(_00811_),
    .A2(_03872_),
    .ZN(_00304_)
  );
  AND2_X1 _09092_ (
    .A1(_00770_),
    .A2(_03862_),
    .ZN(_03873_)
  );
  INV_X1 _09093_ (
    .A(_03873_),
    .ZN(_03874_)
  );
  AND2_X1 _09094_ (
    .A1(_03710_),
    .A2(_03874_),
    .ZN(_03875_)
  );
  AND2_X1 _09095_ (
    .A1(large_1[37]),
    .A2(_03861_),
    .ZN(_03876_)
  );
  INV_X1 _09096_ (
    .A(_03876_),
    .ZN(_03877_)
  );
  AND2_X1 _09097_ (
    .A1(_03875_),
    .A2(_03877_),
    .ZN(_03878_)
  );
  INV_X1 _09098_ (
    .A(_03878_),
    .ZN(_03879_)
  );
  AND2_X1 _09099_ (
    .A1(_02314_),
    .A2(_03700_),
    .ZN(_03880_)
  );
  INV_X1 _09100_ (
    .A(_03880_),
    .ZN(_03881_)
  );
  AND2_X1 _09101_ (
    .A1(large_1[37]),
    .A2(_03702_),
    .ZN(_03882_)
  );
  INV_X1 _09102_ (
    .A(_03882_),
    .ZN(_03883_)
  );
  AND2_X1 _09103_ (
    .A1(_03881_),
    .A2(_03883_),
    .ZN(_03884_)
  );
  AND2_X1 _09104_ (
    .A1(_03879_),
    .A2(_03884_),
    .ZN(_03885_)
  );
  INV_X1 _09105_ (
    .A(_03885_),
    .ZN(_03886_)
  );
  AND2_X1 _09106_ (
    .A1(_00811_),
    .A2(_03886_),
    .ZN(_00305_)
  );
  AND2_X1 _09107_ (
    .A1(_00769_),
    .A2(_03877_),
    .ZN(_03887_)
  );
  INV_X1 _09108_ (
    .A(_03887_),
    .ZN(_03888_)
  );
  AND2_X1 _09109_ (
    .A1(large_1[38]),
    .A2(large_1[37]),
    .ZN(_03889_)
  );
  AND2_X1 _09110_ (
    .A1(large_1[36]),
    .A2(_03889_),
    .ZN(_03890_)
  );
  AND2_X1 _09111_ (
    .A1(_03847_),
    .A2(_03890_),
    .ZN(_03891_)
  );
  INV_X1 _09112_ (
    .A(_03891_),
    .ZN(_03892_)
  );
  AND2_X1 _09113_ (
    .A1(_03710_),
    .A2(_03892_),
    .ZN(_03893_)
  );
  AND2_X1 _09114_ (
    .A1(_03888_),
    .A2(_03893_),
    .ZN(_03894_)
  );
  INV_X1 _09115_ (
    .A(_03894_),
    .ZN(_03895_)
  );
  AND2_X1 _09116_ (
    .A1(_02389_),
    .A2(_03700_),
    .ZN(_03896_)
  );
  INV_X1 _09117_ (
    .A(_03896_),
    .ZN(_03897_)
  );
  AND2_X1 _09118_ (
    .A1(large_1[38]),
    .A2(_03702_),
    .ZN(_03898_)
  );
  INV_X1 _09119_ (
    .A(_03898_),
    .ZN(_03899_)
  );
  AND2_X1 _09120_ (
    .A1(_03897_),
    .A2(_03899_),
    .ZN(_03900_)
  );
  AND2_X1 _09121_ (
    .A1(_03895_),
    .A2(_03900_),
    .ZN(_03901_)
  );
  INV_X1 _09122_ (
    .A(_03901_),
    .ZN(_03902_)
  );
  AND2_X1 _09123_ (
    .A1(_00811_),
    .A2(_03902_),
    .ZN(_00306_)
  );
  AND2_X1 _09124_ (
    .A1(large_1[39]),
    .A2(_03891_),
    .ZN(_03903_)
  );
  INV_X1 _09125_ (
    .A(_03903_),
    .ZN(_03904_)
  );
  AND2_X1 _09126_ (
    .A1(_00768_),
    .A2(_03892_),
    .ZN(_03905_)
  );
  INV_X1 _09127_ (
    .A(_03905_),
    .ZN(_03906_)
  );
  AND2_X1 _09128_ (
    .A1(_03710_),
    .A2(_03906_),
    .ZN(_03907_)
  );
  AND2_X1 _09129_ (
    .A1(_03904_),
    .A2(_03907_),
    .ZN(_03908_)
  );
  INV_X1 _09130_ (
    .A(_03908_),
    .ZN(_03909_)
  );
  AND2_X1 _09131_ (
    .A1(_02456_),
    .A2(_03700_),
    .ZN(_03910_)
  );
  INV_X1 _09132_ (
    .A(_03910_),
    .ZN(_03911_)
  );
  AND2_X1 _09133_ (
    .A1(large_1[39]),
    .A2(_03702_),
    .ZN(_03912_)
  );
  INV_X1 _09134_ (
    .A(_03912_),
    .ZN(_03913_)
  );
  AND2_X1 _09135_ (
    .A1(_03911_),
    .A2(_03913_),
    .ZN(_03914_)
  );
  AND2_X1 _09136_ (
    .A1(_03909_),
    .A2(_03914_),
    .ZN(_03915_)
  );
  INV_X1 _09137_ (
    .A(_03915_),
    .ZN(_03916_)
  );
  AND2_X1 _09138_ (
    .A1(_00811_),
    .A2(_03916_),
    .ZN(_00307_)
  );
  AND2_X1 _09139_ (
    .A1(large_1[39]),
    .A2(large_1[32]),
    .ZN(_03917_)
  );
  AND2_X1 _09140_ (
    .A1(_03727_),
    .A2(_03917_),
    .ZN(_03918_)
  );
  AND2_X1 _09141_ (
    .A1(_03800_),
    .A2(_03846_),
    .ZN(_03919_)
  );
  AND2_X1 _09142_ (
    .A1(_03890_),
    .A2(_03918_),
    .ZN(_03920_)
  );
  AND2_X1 _09143_ (
    .A1(_03919_),
    .A2(_03920_),
    .ZN(_03921_)
  );
  AND2_X1 _09144_ (
    .A1(_03692_),
    .A2(_03921_),
    .ZN(_03922_)
  );
  INV_X1 _09145_ (
    .A(_03922_),
    .ZN(_03923_)
  );
  AND2_X1 _09146_ (
    .A1(_00767_),
    .A2(_03923_),
    .ZN(_03924_)
  );
  INV_X1 _09147_ (
    .A(_03924_),
    .ZN(_03925_)
  );
  AND2_X1 _09148_ (
    .A1(large_1[40]),
    .A2(_03922_),
    .ZN(_03926_)
  );
  INV_X1 _09149_ (
    .A(_03926_),
    .ZN(_03927_)
  );
  AND2_X1 _09150_ (
    .A1(_03925_),
    .A2(_03927_),
    .ZN(_03928_)
  );
  AND2_X1 _09151_ (
    .A1(_03710_),
    .A2(_03928_),
    .ZN(_03929_)
  );
  INV_X1 _09152_ (
    .A(_03929_),
    .ZN(_03930_)
  );
  AND2_X1 _09153_ (
    .A1(_02522_),
    .A2(_03700_),
    .ZN(_03931_)
  );
  INV_X1 _09154_ (
    .A(_03931_),
    .ZN(_03932_)
  );
  AND2_X1 _09155_ (
    .A1(large_1[40]),
    .A2(_03702_),
    .ZN(_03933_)
  );
  INV_X1 _09156_ (
    .A(_03933_),
    .ZN(_03934_)
  );
  AND2_X1 _09157_ (
    .A1(_03932_),
    .A2(_03934_),
    .ZN(_03935_)
  );
  AND2_X1 _09158_ (
    .A1(_03930_),
    .A2(_03935_),
    .ZN(_03936_)
  );
  INV_X1 _09159_ (
    .A(_03936_),
    .ZN(_03937_)
  );
  AND2_X1 _09160_ (
    .A1(_00811_),
    .A2(_03937_),
    .ZN(_00308_)
  );
  AND2_X1 _09161_ (
    .A1(_00766_),
    .A2(_03927_),
    .ZN(_03938_)
  );
  INV_X1 _09162_ (
    .A(_03938_),
    .ZN(_03939_)
  );
  AND2_X1 _09163_ (
    .A1(large_1[41]),
    .A2(large_1[40]),
    .ZN(_03940_)
  );
  AND2_X1 _09164_ (
    .A1(large_1[41]),
    .A2(_03926_),
    .ZN(_03941_)
  );
  INV_X1 _09165_ (
    .A(_03941_),
    .ZN(_03942_)
  );
  AND2_X1 _09166_ (
    .A1(_03710_),
    .A2(_03942_),
    .ZN(_03943_)
  );
  AND2_X1 _09167_ (
    .A1(_03939_),
    .A2(_03943_),
    .ZN(_03944_)
  );
  INV_X1 _09168_ (
    .A(_03944_),
    .ZN(_03945_)
  );
  AND2_X1 _09169_ (
    .A1(_02597_),
    .A2(_03700_),
    .ZN(_03946_)
  );
  INV_X1 _09170_ (
    .A(_03946_),
    .ZN(_03947_)
  );
  AND2_X1 _09171_ (
    .A1(large_1[41]),
    .A2(_03702_),
    .ZN(_03948_)
  );
  INV_X1 _09172_ (
    .A(_03948_),
    .ZN(_03949_)
  );
  AND2_X1 _09173_ (
    .A1(_03947_),
    .A2(_03949_),
    .ZN(_03950_)
  );
  AND2_X1 _09174_ (
    .A1(_03945_),
    .A2(_03950_),
    .ZN(_03951_)
  );
  INV_X1 _09175_ (
    .A(_03951_),
    .ZN(_03952_)
  );
  AND2_X1 _09176_ (
    .A1(_00811_),
    .A2(_03952_),
    .ZN(_00309_)
  );
  AND2_X1 _09177_ (
    .A1(_00765_),
    .A2(_03942_),
    .ZN(_03953_)
  );
  INV_X1 _09178_ (
    .A(_03953_),
    .ZN(_03954_)
  );
  AND2_X1 _09179_ (
    .A1(large_1[42]),
    .A2(_03941_),
    .ZN(_03955_)
  );
  INV_X1 _09180_ (
    .A(_03955_),
    .ZN(_03956_)
  );
  AND2_X1 _09181_ (
    .A1(_03954_),
    .A2(_03956_),
    .ZN(_03957_)
  );
  AND2_X1 _09182_ (
    .A1(_03710_),
    .A2(_03957_),
    .ZN(_03958_)
  );
  INV_X1 _09183_ (
    .A(_03958_),
    .ZN(_03959_)
  );
  AND2_X1 _09184_ (
    .A1(_01035_),
    .A2(_03700_),
    .ZN(_03960_)
  );
  INV_X1 _09185_ (
    .A(_03960_),
    .ZN(_03961_)
  );
  AND2_X1 _09186_ (
    .A1(large_1[42]),
    .A2(_03702_),
    .ZN(_03962_)
  );
  INV_X1 _09187_ (
    .A(_03962_),
    .ZN(_03963_)
  );
  AND2_X1 _09188_ (
    .A1(_03961_),
    .A2(_03963_),
    .ZN(_03964_)
  );
  AND2_X1 _09189_ (
    .A1(_03959_),
    .A2(_03964_),
    .ZN(_03965_)
  );
  INV_X1 _09190_ (
    .A(_03965_),
    .ZN(_03966_)
  );
  AND2_X1 _09191_ (
    .A1(_00811_),
    .A2(_03966_),
    .ZN(_00310_)
  );
  AND2_X1 _09192_ (
    .A1(_00764_),
    .A2(_03956_),
    .ZN(_03967_)
  );
  INV_X1 _09193_ (
    .A(_03967_),
    .ZN(_03968_)
  );
  AND2_X1 _09194_ (
    .A1(large_1[43]),
    .A2(large_1[42]),
    .ZN(_03969_)
  );
  AND2_X1 _09195_ (
    .A1(large_1[43]),
    .A2(_03955_),
    .ZN(_03970_)
  );
  INV_X1 _09196_ (
    .A(_03970_),
    .ZN(_03971_)
  );
  AND2_X1 _09197_ (
    .A1(_03710_),
    .A2(_03971_),
    .ZN(_03972_)
  );
  AND2_X1 _09198_ (
    .A1(_03968_),
    .A2(_03972_),
    .ZN(_03973_)
  );
  INV_X1 _09199_ (
    .A(_03973_),
    .ZN(_03974_)
  );
  AND2_X1 _09200_ (
    .A1(_02669_),
    .A2(_03700_),
    .ZN(_03975_)
  );
  INV_X1 _09201_ (
    .A(_03975_),
    .ZN(_03976_)
  );
  AND2_X1 _09202_ (
    .A1(large_1[43]),
    .A2(_03708_),
    .ZN(_03977_)
  );
  INV_X1 _09203_ (
    .A(_03977_),
    .ZN(_03978_)
  );
  AND2_X1 _09204_ (
    .A1(_03976_),
    .A2(_03978_),
    .ZN(_03979_)
  );
  AND2_X1 _09205_ (
    .A1(_03974_),
    .A2(_03979_),
    .ZN(_03980_)
  );
  INV_X1 _09206_ (
    .A(_03980_),
    .ZN(_03981_)
  );
  AND2_X1 _09207_ (
    .A1(_00811_),
    .A2(_03981_),
    .ZN(_00311_)
  );
  AND2_X1 _09208_ (
    .A1(_03940_),
    .A2(_03969_),
    .ZN(_03982_)
  );
  AND2_X1 _09209_ (
    .A1(_03922_),
    .A2(_03982_),
    .ZN(_03983_)
  );
  INV_X1 _09210_ (
    .A(_03983_),
    .ZN(_03984_)
  );
  AND2_X1 _09211_ (
    .A1(_00763_),
    .A2(_03984_),
    .ZN(_03985_)
  );
  INV_X1 _09212_ (
    .A(_03985_),
    .ZN(_03986_)
  );
  AND2_X1 _09213_ (
    .A1(large_1[44]),
    .A2(_03983_),
    .ZN(_03987_)
  );
  INV_X1 _09214_ (
    .A(_03987_),
    .ZN(_03988_)
  );
  AND2_X1 _09215_ (
    .A1(_03986_),
    .A2(_03988_),
    .ZN(_03989_)
  );
  AND2_X1 _09216_ (
    .A1(_03710_),
    .A2(_03989_),
    .ZN(_03990_)
  );
  INV_X1 _09217_ (
    .A(_03990_),
    .ZN(_03991_)
  );
  AND2_X1 _09218_ (
    .A1(_01107_),
    .A2(_03700_),
    .ZN(_03992_)
  );
  INV_X1 _09219_ (
    .A(_03992_),
    .ZN(_03993_)
  );
  AND2_X1 _09220_ (
    .A1(large_1[44]),
    .A2(_03702_),
    .ZN(_03994_)
  );
  INV_X1 _09221_ (
    .A(_03994_),
    .ZN(_03995_)
  );
  AND2_X1 _09222_ (
    .A1(_03993_),
    .A2(_03995_),
    .ZN(_03996_)
  );
  AND2_X1 _09223_ (
    .A1(_03991_),
    .A2(_03996_),
    .ZN(_03997_)
  );
  INV_X1 _09224_ (
    .A(_03997_),
    .ZN(_03998_)
  );
  AND2_X1 _09225_ (
    .A1(_00811_),
    .A2(_03998_),
    .ZN(_00312_)
  );
  AND2_X1 _09226_ (
    .A1(_00762_),
    .A2(_03988_),
    .ZN(_03999_)
  );
  INV_X1 _09227_ (
    .A(_03999_),
    .ZN(_04000_)
  );
  AND2_X1 _09228_ (
    .A1(large_1[45]),
    .A2(large_1[44]),
    .ZN(_04001_)
  );
  AND2_X1 _09229_ (
    .A1(large_1[45]),
    .A2(_03987_),
    .ZN(_04002_)
  );
  INV_X1 _09230_ (
    .A(_04002_),
    .ZN(_04003_)
  );
  AND2_X1 _09231_ (
    .A1(_03710_),
    .A2(_04003_),
    .ZN(_04004_)
  );
  AND2_X1 _09232_ (
    .A1(_04000_),
    .A2(_04004_),
    .ZN(_04005_)
  );
  INV_X1 _09233_ (
    .A(_04005_),
    .ZN(_04006_)
  );
  AND2_X1 _09234_ (
    .A1(_01199_),
    .A2(_03700_),
    .ZN(_04007_)
  );
  INV_X1 _09235_ (
    .A(_04007_),
    .ZN(_04008_)
  );
  AND2_X1 _09236_ (
    .A1(large_1[45]),
    .A2(_03702_),
    .ZN(_04009_)
  );
  INV_X1 _09237_ (
    .A(_04009_),
    .ZN(_04010_)
  );
  AND2_X1 _09238_ (
    .A1(_04008_),
    .A2(_04010_),
    .ZN(_04011_)
  );
  AND2_X1 _09239_ (
    .A1(_04006_),
    .A2(_04011_),
    .ZN(_04012_)
  );
  INV_X1 _09240_ (
    .A(_04012_),
    .ZN(_04013_)
  );
  AND2_X1 _09241_ (
    .A1(_00811_),
    .A2(_04013_),
    .ZN(_00313_)
  );
  AND2_X1 _09242_ (
    .A1(_00761_),
    .A2(_04003_),
    .ZN(_04014_)
  );
  INV_X1 _09243_ (
    .A(_04014_),
    .ZN(_04015_)
  );
  AND2_X1 _09244_ (
    .A1(large_1[46]),
    .A2(_04002_),
    .ZN(_04016_)
  );
  INV_X1 _09245_ (
    .A(_04016_),
    .ZN(_04017_)
  );
  AND2_X1 _09246_ (
    .A1(_04015_),
    .A2(_04017_),
    .ZN(_04018_)
  );
  AND2_X1 _09247_ (
    .A1(_03710_),
    .A2(_04018_),
    .ZN(_04019_)
  );
  INV_X1 _09248_ (
    .A(_04019_),
    .ZN(_04020_)
  );
  AND2_X1 _09249_ (
    .A1(_01277_),
    .A2(_03700_),
    .ZN(_04021_)
  );
  INV_X1 _09250_ (
    .A(_04021_),
    .ZN(_04022_)
  );
  AND2_X1 _09251_ (
    .A1(large_1[46]),
    .A2(_03702_),
    .ZN(_04023_)
  );
  INV_X1 _09252_ (
    .A(_04023_),
    .ZN(_04024_)
  );
  AND2_X1 _09253_ (
    .A1(_04022_),
    .A2(_04024_),
    .ZN(_04025_)
  );
  AND2_X1 _09254_ (
    .A1(_04020_),
    .A2(_04025_),
    .ZN(_04026_)
  );
  INV_X1 _09255_ (
    .A(_04026_),
    .ZN(_04027_)
  );
  AND2_X1 _09256_ (
    .A1(_00811_),
    .A2(_04027_),
    .ZN(_00314_)
  );
  AND2_X1 _09257_ (
    .A1(_00760_),
    .A2(_04017_),
    .ZN(_04028_)
  );
  INV_X1 _09258_ (
    .A(_04028_),
    .ZN(_04029_)
  );
  AND2_X1 _09259_ (
    .A1(large_1[47]),
    .A2(large_1[46]),
    .ZN(_04030_)
  );
  AND2_X1 _09260_ (
    .A1(_04001_),
    .A2(_04030_),
    .ZN(_04031_)
  );
  AND2_X1 _09261_ (
    .A1(large_1[47]),
    .A2(_04016_),
    .ZN(_04032_)
  );
  INV_X1 _09262_ (
    .A(_04032_),
    .ZN(_04033_)
  );
  AND2_X1 _09263_ (
    .A1(_03710_),
    .A2(_04033_),
    .ZN(_04034_)
  );
  AND2_X1 _09264_ (
    .A1(_04029_),
    .A2(_04034_),
    .ZN(_04035_)
  );
  INV_X1 _09265_ (
    .A(_04035_),
    .ZN(_04036_)
  );
  AND2_X1 _09266_ (
    .A1(_02735_),
    .A2(_03700_),
    .ZN(_04037_)
  );
  INV_X1 _09267_ (
    .A(_04037_),
    .ZN(_04038_)
  );
  AND2_X1 _09268_ (
    .A1(large_1[47]),
    .A2(_03702_),
    .ZN(_04039_)
  );
  INV_X1 _09269_ (
    .A(_04039_),
    .ZN(_04040_)
  );
  AND2_X1 _09270_ (
    .A1(_04038_),
    .A2(_04040_),
    .ZN(_04041_)
  );
  AND2_X1 _09271_ (
    .A1(_04036_),
    .A2(_04041_),
    .ZN(_04042_)
  );
  INV_X1 _09272_ (
    .A(_04042_),
    .ZN(_04043_)
  );
  AND2_X1 _09273_ (
    .A1(_00811_),
    .A2(_04043_),
    .ZN(_00315_)
  );
  AND2_X1 _09274_ (
    .A1(_03982_),
    .A2(_04031_),
    .ZN(_04044_)
  );
  AND2_X1 _09275_ (
    .A1(_03922_),
    .A2(_04044_),
    .ZN(_04045_)
  );
  INV_X1 _09276_ (
    .A(_04045_),
    .ZN(_04046_)
  );
  AND2_X1 _09277_ (
    .A1(_00759_),
    .A2(_04046_),
    .ZN(_04047_)
  );
  INV_X1 _09278_ (
    .A(_04047_),
    .ZN(_04048_)
  );
  AND2_X1 _09279_ (
    .A1(large_1[48]),
    .A2(_04045_),
    .ZN(_04049_)
  );
  INV_X1 _09280_ (
    .A(_04049_),
    .ZN(_04050_)
  );
  AND2_X1 _09281_ (
    .A1(_04048_),
    .A2(_04050_),
    .ZN(_04051_)
  );
  AND2_X1 _09282_ (
    .A1(_03710_),
    .A2(_04051_),
    .ZN(_04052_)
  );
  INV_X1 _09283_ (
    .A(_04052_),
    .ZN(_04053_)
  );
  AND2_X1 _09284_ (
    .A1(_02801_),
    .A2(_03700_),
    .ZN(_04054_)
  );
  INV_X1 _09285_ (
    .A(_04054_),
    .ZN(_04055_)
  );
  AND2_X1 _09286_ (
    .A1(large_1[48]),
    .A2(_03702_),
    .ZN(_04056_)
  );
  INV_X1 _09287_ (
    .A(_04056_),
    .ZN(_04057_)
  );
  AND2_X1 _09288_ (
    .A1(_04055_),
    .A2(_04057_),
    .ZN(_04058_)
  );
  AND2_X1 _09289_ (
    .A1(_04053_),
    .A2(_04058_),
    .ZN(_04059_)
  );
  INV_X1 _09290_ (
    .A(_04059_),
    .ZN(_04060_)
  );
  AND2_X1 _09291_ (
    .A1(_00811_),
    .A2(_04060_),
    .ZN(_00316_)
  );
  AND2_X1 _09292_ (
    .A1(_00758_),
    .A2(_04050_),
    .ZN(_04061_)
  );
  INV_X1 _09293_ (
    .A(_04061_),
    .ZN(_04062_)
  );
  AND2_X1 _09294_ (
    .A1(large_1[49]),
    .A2(_04049_),
    .ZN(_04063_)
  );
  INV_X1 _09295_ (
    .A(_04063_),
    .ZN(_04064_)
  );
  AND2_X1 _09296_ (
    .A1(_03710_),
    .A2(_04064_),
    .ZN(_04065_)
  );
  AND2_X1 _09297_ (
    .A1(_04062_),
    .A2(_04065_),
    .ZN(_04066_)
  );
  INV_X1 _09298_ (
    .A(_04066_),
    .ZN(_04067_)
  );
  AND2_X1 _09299_ (
    .A1(_01360_),
    .A2(_03700_),
    .ZN(_04068_)
  );
  INV_X1 _09300_ (
    .A(_04068_),
    .ZN(_04069_)
  );
  AND2_X1 _09301_ (
    .A1(large_1[49]),
    .A2(_03702_),
    .ZN(_04070_)
  );
  INV_X1 _09302_ (
    .A(_04070_),
    .ZN(_04071_)
  );
  AND2_X1 _09303_ (
    .A1(_04069_),
    .A2(_04071_),
    .ZN(_04072_)
  );
  AND2_X1 _09304_ (
    .A1(_04067_),
    .A2(_04072_),
    .ZN(_04073_)
  );
  INV_X1 _09305_ (
    .A(_04073_),
    .ZN(_04074_)
  );
  AND2_X1 _09306_ (
    .A1(_00811_),
    .A2(_04074_),
    .ZN(_00317_)
  );
  AND2_X1 _09307_ (
    .A1(_00757_),
    .A2(_04064_),
    .ZN(_04075_)
  );
  INV_X1 _09308_ (
    .A(_04075_),
    .ZN(_04076_)
  );
  AND2_X1 _09309_ (
    .A1(large_1[50]),
    .A2(large_1[49]),
    .ZN(_04077_)
  );
  AND2_X1 _09310_ (
    .A1(_04049_),
    .A2(_04077_),
    .ZN(_04078_)
  );
  INV_X1 _09311_ (
    .A(_04078_),
    .ZN(_04079_)
  );
  AND2_X1 _09312_ (
    .A1(_04076_),
    .A2(_04079_),
    .ZN(_04080_)
  );
  AND2_X1 _09313_ (
    .A1(_03710_),
    .A2(_04080_),
    .ZN(_04081_)
  );
  INV_X1 _09314_ (
    .A(_04081_),
    .ZN(_04082_)
  );
  AND2_X1 _09315_ (
    .A1(_02873_),
    .A2(_03700_),
    .ZN(_04083_)
  );
  INV_X1 _09316_ (
    .A(_04083_),
    .ZN(_04084_)
  );
  AND2_X1 _09317_ (
    .A1(large_1[50]),
    .A2(_03702_),
    .ZN(_04085_)
  );
  INV_X1 _09318_ (
    .A(_04085_),
    .ZN(_04086_)
  );
  AND2_X1 _09319_ (
    .A1(_04084_),
    .A2(_04086_),
    .ZN(_04087_)
  );
  AND2_X1 _09320_ (
    .A1(_04082_),
    .A2(_04087_),
    .ZN(_04088_)
  );
  INV_X1 _09321_ (
    .A(_04088_),
    .ZN(_04089_)
  );
  AND2_X1 _09322_ (
    .A1(_00811_),
    .A2(_04089_),
    .ZN(_00318_)
  );
  AND2_X1 _09323_ (
    .A1(_00756_),
    .A2(_04079_),
    .ZN(_04090_)
  );
  INV_X1 _09324_ (
    .A(_04090_),
    .ZN(_04091_)
  );
  AND2_X1 _09325_ (
    .A1(large_1[51]),
    .A2(_04078_),
    .ZN(_04092_)
  );
  INV_X1 _09326_ (
    .A(_04092_),
    .ZN(_04093_)
  );
  AND2_X1 _09327_ (
    .A1(_03710_),
    .A2(_04093_),
    .ZN(_04094_)
  );
  AND2_X1 _09328_ (
    .A1(_04091_),
    .A2(_04094_),
    .ZN(_04095_)
  );
  INV_X1 _09329_ (
    .A(_04095_),
    .ZN(_04096_)
  );
  AND2_X1 _09330_ (
    .A1(_02945_),
    .A2(_03700_),
    .ZN(_04097_)
  );
  INV_X1 _09331_ (
    .A(_04097_),
    .ZN(_04098_)
  );
  AND2_X1 _09332_ (
    .A1(large_1[51]),
    .A2(_03708_),
    .ZN(_04099_)
  );
  INV_X1 _09333_ (
    .A(_04099_),
    .ZN(_04100_)
  );
  AND2_X1 _09334_ (
    .A1(_04098_),
    .A2(_04100_),
    .ZN(_04101_)
  );
  AND2_X1 _09335_ (
    .A1(_04096_),
    .A2(_04101_),
    .ZN(_04102_)
  );
  INV_X1 _09336_ (
    .A(_04102_),
    .ZN(_04103_)
  );
  AND2_X1 _09337_ (
    .A1(_00811_),
    .A2(_04103_),
    .ZN(_00319_)
  );
  AND2_X1 _09338_ (
    .A1(_00755_),
    .A2(_04093_),
    .ZN(_04104_)
  );
  INV_X1 _09339_ (
    .A(_04104_),
    .ZN(_04105_)
  );
  AND2_X1 _09340_ (
    .A1(large_1[52]),
    .A2(_04092_),
    .ZN(_04106_)
  );
  INV_X1 _09341_ (
    .A(_04106_),
    .ZN(_04107_)
  );
  AND2_X1 _09342_ (
    .A1(_04105_),
    .A2(_04107_),
    .ZN(_04108_)
  );
  AND2_X1 _09343_ (
    .A1(_03710_),
    .A2(_04108_),
    .ZN(_04109_)
  );
  INV_X1 _09344_ (
    .A(_04109_),
    .ZN(_04110_)
  );
  AND2_X1 _09345_ (
    .A1(_03017_),
    .A2(_03700_),
    .ZN(_04111_)
  );
  INV_X1 _09346_ (
    .A(_04111_),
    .ZN(_04112_)
  );
  AND2_X1 _09347_ (
    .A1(large_1[52]),
    .A2(_03702_),
    .ZN(_04113_)
  );
  INV_X1 _09348_ (
    .A(_04113_),
    .ZN(_04114_)
  );
  AND2_X1 _09349_ (
    .A1(_04112_),
    .A2(_04114_),
    .ZN(_04115_)
  );
  AND2_X1 _09350_ (
    .A1(_04110_),
    .A2(_04115_),
    .ZN(_04116_)
  );
  INV_X1 _09351_ (
    .A(_04116_),
    .ZN(_04117_)
  );
  AND2_X1 _09352_ (
    .A1(_00811_),
    .A2(_04117_),
    .ZN(_00320_)
  );
  AND2_X1 _09353_ (
    .A1(_00754_),
    .A2(_04107_),
    .ZN(_04118_)
  );
  INV_X1 _09354_ (
    .A(_04118_),
    .ZN(_04119_)
  );
  AND2_X1 _09355_ (
    .A1(large_1[53]),
    .A2(_04106_),
    .ZN(_04120_)
  );
  INV_X1 _09356_ (
    .A(_04120_),
    .ZN(_04121_)
  );
  AND2_X1 _09357_ (
    .A1(_03710_),
    .A2(_04121_),
    .ZN(_04122_)
  );
  AND2_X1 _09358_ (
    .A1(_04119_),
    .A2(_04122_),
    .ZN(_04123_)
  );
  INV_X1 _09359_ (
    .A(_04123_),
    .ZN(_04124_)
  );
  AND2_X1 _09360_ (
    .A1(_03089_),
    .A2(_03700_),
    .ZN(_04125_)
  );
  INV_X1 _09361_ (
    .A(_04125_),
    .ZN(_04126_)
  );
  AND2_X1 _09362_ (
    .A1(large_1[53]),
    .A2(_03702_),
    .ZN(_04127_)
  );
  INV_X1 _09363_ (
    .A(_04127_),
    .ZN(_04128_)
  );
  AND2_X1 _09364_ (
    .A1(_04126_),
    .A2(_04128_),
    .ZN(_04129_)
  );
  AND2_X1 _09365_ (
    .A1(_04124_),
    .A2(_04129_),
    .ZN(_04130_)
  );
  INV_X1 _09366_ (
    .A(_04130_),
    .ZN(_04131_)
  );
  AND2_X1 _09367_ (
    .A1(_00811_),
    .A2(_04131_),
    .ZN(_00321_)
  );
  AND2_X1 _09368_ (
    .A1(_00753_),
    .A2(_04121_),
    .ZN(_04132_)
  );
  INV_X1 _09369_ (
    .A(_04132_),
    .ZN(_04133_)
  );
  AND2_X1 _09370_ (
    .A1(large_1[54]),
    .A2(_04120_),
    .ZN(_04134_)
  );
  INV_X1 _09371_ (
    .A(_04134_),
    .ZN(_04135_)
  );
  AND2_X1 _09372_ (
    .A1(_04133_),
    .A2(_04135_),
    .ZN(_04136_)
  );
  AND2_X1 _09373_ (
    .A1(_03710_),
    .A2(_04136_),
    .ZN(_04137_)
  );
  INV_X1 _09374_ (
    .A(_04137_),
    .ZN(_04138_)
  );
  AND2_X1 _09375_ (
    .A1(_03162_),
    .A2(_03700_),
    .ZN(_04139_)
  );
  INV_X1 _09376_ (
    .A(_04139_),
    .ZN(_04140_)
  );
  AND2_X1 _09377_ (
    .A1(large_1[54]),
    .A2(_03702_),
    .ZN(_04141_)
  );
  INV_X1 _09378_ (
    .A(_04141_),
    .ZN(_04142_)
  );
  AND2_X1 _09379_ (
    .A1(_04140_),
    .A2(_04142_),
    .ZN(_04143_)
  );
  AND2_X1 _09380_ (
    .A1(_04138_),
    .A2(_04143_),
    .ZN(_04144_)
  );
  INV_X1 _09381_ (
    .A(_04144_),
    .ZN(_04145_)
  );
  AND2_X1 _09382_ (
    .A1(_00811_),
    .A2(_04145_),
    .ZN(_00322_)
  );
  AND2_X1 _09383_ (
    .A1(_00752_),
    .A2(_04135_),
    .ZN(_04146_)
  );
  INV_X1 _09384_ (
    .A(_04146_),
    .ZN(_04147_)
  );
  AND2_X1 _09385_ (
    .A1(large_1[55]),
    .A2(_04134_),
    .ZN(_04148_)
  );
  INV_X1 _09386_ (
    .A(_04148_),
    .ZN(_04149_)
  );
  AND2_X1 _09387_ (
    .A1(_03710_),
    .A2(_04149_),
    .ZN(_04150_)
  );
  AND2_X1 _09388_ (
    .A1(_04147_),
    .A2(_04150_),
    .ZN(_04151_)
  );
  INV_X1 _09389_ (
    .A(_04151_),
    .ZN(_04152_)
  );
  AND2_X1 _09390_ (
    .A1(_03230_),
    .A2(_03700_),
    .ZN(_04153_)
  );
  INV_X1 _09391_ (
    .A(_04153_),
    .ZN(_04154_)
  );
  AND2_X1 _09392_ (
    .A1(large_1[55]),
    .A2(_03702_),
    .ZN(_04155_)
  );
  INV_X1 _09393_ (
    .A(_04155_),
    .ZN(_04156_)
  );
  AND2_X1 _09394_ (
    .A1(_04154_),
    .A2(_04156_),
    .ZN(_04157_)
  );
  AND2_X1 _09395_ (
    .A1(_04152_),
    .A2(_04157_),
    .ZN(_04158_)
  );
  INV_X1 _09396_ (
    .A(_04158_),
    .ZN(_04159_)
  );
  AND2_X1 _09397_ (
    .A1(_00811_),
    .A2(_04159_),
    .ZN(_00323_)
  );
  AND2_X1 _09398_ (
    .A1(_00751_),
    .A2(_04149_),
    .ZN(_04160_)
  );
  INV_X1 _09399_ (
    .A(_04160_),
    .ZN(_04161_)
  );
  AND2_X1 _09400_ (
    .A1(large_1[56]),
    .A2(_04148_),
    .ZN(_04162_)
  );
  INV_X1 _09401_ (
    .A(_04162_),
    .ZN(_04163_)
  );
  AND2_X1 _09402_ (
    .A1(_03710_),
    .A2(_04163_),
    .ZN(_04164_)
  );
  AND2_X1 _09403_ (
    .A1(_04161_),
    .A2(_04164_),
    .ZN(_04165_)
  );
  INV_X1 _09404_ (
    .A(_04165_),
    .ZN(_04166_)
  );
  AND2_X1 _09405_ (
    .A1(_03443_),
    .A2(_03700_),
    .ZN(_04167_)
  );
  INV_X1 _09406_ (
    .A(_04167_),
    .ZN(_04168_)
  );
  AND2_X1 _09407_ (
    .A1(large_1[56]),
    .A2(_03702_),
    .ZN(_04169_)
  );
  INV_X1 _09408_ (
    .A(_04169_),
    .ZN(_04170_)
  );
  AND2_X1 _09409_ (
    .A1(_04168_),
    .A2(_04170_),
    .ZN(_04171_)
  );
  AND2_X1 _09410_ (
    .A1(_04166_),
    .A2(_04171_),
    .ZN(_04172_)
  );
  INV_X1 _09411_ (
    .A(_04172_),
    .ZN(_04173_)
  );
  AND2_X1 _09412_ (
    .A1(_00811_),
    .A2(_04173_),
    .ZN(_00324_)
  );
  AND2_X1 _09413_ (
    .A1(large_1[57]),
    .A2(_04163_),
    .ZN(_04174_)
  );
  INV_X1 _09414_ (
    .A(_04174_),
    .ZN(_04175_)
  );
  AND2_X1 _09415_ (
    .A1(_00750_),
    .A2(_04162_),
    .ZN(_04176_)
  );
  INV_X1 _09416_ (
    .A(_04176_),
    .ZN(_04177_)
  );
  AND2_X1 _09417_ (
    .A1(_04175_),
    .A2(_04177_),
    .ZN(_04178_)
  );
  INV_X1 _09418_ (
    .A(_04178_),
    .ZN(_04179_)
  );
  AND2_X1 _09419_ (
    .A1(_03710_),
    .A2(_04179_),
    .ZN(_04180_)
  );
  INV_X1 _09420_ (
    .A(_04180_),
    .ZN(_04181_)
  );
  AND2_X1 _09421_ (
    .A1(_03342_),
    .A2(_03700_),
    .ZN(_04182_)
  );
  INV_X1 _09422_ (
    .A(_04182_),
    .ZN(_04183_)
  );
  AND2_X1 _09423_ (
    .A1(large_1[57]),
    .A2(_03708_),
    .ZN(_04184_)
  );
  INV_X1 _09424_ (
    .A(_04184_),
    .ZN(_04185_)
  );
  AND2_X1 _09425_ (
    .A1(_04183_),
    .A2(_04185_),
    .ZN(_04186_)
  );
  AND2_X1 _09426_ (
    .A1(_04181_),
    .A2(_04186_),
    .ZN(_04187_)
  );
  INV_X1 _09427_ (
    .A(_04187_),
    .ZN(_04188_)
  );
  AND2_X1 _09428_ (
    .A1(_00811_),
    .A2(_04188_),
    .ZN(_00325_)
  );
  AND2_X1 _09429_ (
    .A1(_00783_),
    .A2(_03653_),
    .ZN(_04189_)
  );
  INV_X1 _09430_ (
    .A(_04189_),
    .ZN(_04190_)
  );
  AND2_X1 _09431_ (
    .A1(small_1[0]),
    .A2(_04190_),
    .ZN(_04191_)
  );
  INV_X1 _09432_ (
    .A(_04191_),
    .ZN(_04192_)
  );
  AND2_X1 _09433_ (
    .A1(_00749_),
    .A2(_04189_),
    .ZN(_04193_)
  );
  INV_X1 _09434_ (
    .A(_04193_),
    .ZN(_04194_)
  );
  AND2_X1 _09435_ (
    .A1(_04192_),
    .A2(_04194_),
    .ZN(_04195_)
  );
  INV_X1 _09436_ (
    .A(_04195_),
    .ZN(_04196_)
  );
  AND2_X1 _09437_ (
    .A1(_03705_),
    .A2(_04196_),
    .ZN(_04197_)
  );
  INV_X1 _09438_ (
    .A(_04197_),
    .ZN(_04198_)
  );
  AND2_X1 _09439_ (
    .A1(small_1[0]),
    .A2(_03700_),
    .ZN(_04199_)
  );
  INV_X1 _09440_ (
    .A(_04199_),
    .ZN(_04200_)
  );
  AND2_X1 _09441_ (
    .A1(_00898_),
    .A2(_04196_),
    .ZN(_04201_)
  );
  INV_X1 _09442_ (
    .A(_04201_),
    .ZN(_04202_)
  );
  AND2_X1 _09443_ (
    .A1(_04200_),
    .A2(_04202_),
    .ZN(_04203_)
  );
  AND2_X1 _09444_ (
    .A1(_04198_),
    .A2(_04203_),
    .ZN(_04204_)
  );
  AND2_X1 _09445_ (
    .A1(_01613_),
    .A2(_03708_),
    .ZN(_04205_)
  );
  INV_X1 _09446_ (
    .A(_04205_),
    .ZN(_04206_)
  );
  AND2_X1 _09447_ (
    .A1(_04204_),
    .A2(_04206_),
    .ZN(_04207_)
  );
  INV_X1 _09448_ (
    .A(_04207_),
    .ZN(_04208_)
  );
  AND2_X1 _09449_ (
    .A1(_00811_),
    .A2(_04208_),
    .ZN(_00326_)
  );
  AND2_X1 _09450_ (
    .A1(small_1[1]),
    .A2(_03700_),
    .ZN(_04209_)
  );
  INV_X1 _09451_ (
    .A(_04209_),
    .ZN(_04210_)
  );
  AND2_X1 _09452_ (
    .A1(_00783_),
    .A2(_03654_),
    .ZN(_04211_)
  );
  INV_X1 _09453_ (
    .A(_04211_),
    .ZN(_04212_)
  );
  AND2_X1 _09454_ (
    .A1(small_1[1]),
    .A2(_04212_),
    .ZN(_04213_)
  );
  INV_X1 _09455_ (
    .A(_04213_),
    .ZN(_04214_)
  );
  AND2_X1 _09456_ (
    .A1(_00748_),
    .A2(_04211_),
    .ZN(_04215_)
  );
  INV_X1 _09457_ (
    .A(_04215_),
    .ZN(_04216_)
  );
  AND2_X1 _09458_ (
    .A1(_04214_),
    .A2(_04216_),
    .ZN(_04217_)
  );
  INV_X1 _09459_ (
    .A(_04217_),
    .ZN(_04218_)
  );
  AND2_X1 _09460_ (
    .A1(_03706_),
    .A2(_04218_),
    .ZN(_04219_)
  );
  INV_X1 _09461_ (
    .A(_04219_),
    .ZN(_04220_)
  );
  AND2_X1 _09462_ (
    .A1(_04210_),
    .A2(_04220_),
    .ZN(_04221_)
  );
  AND2_X1 _09463_ (
    .A1(_01688_),
    .A2(_03702_),
    .ZN(_04222_)
  );
  INV_X1 _09464_ (
    .A(_04222_),
    .ZN(_04223_)
  );
  AND2_X1 _09465_ (
    .A1(_04221_),
    .A2(_04223_),
    .ZN(_04224_)
  );
  INV_X1 _09466_ (
    .A(_04224_),
    .ZN(_04225_)
  );
  AND2_X1 _09467_ (
    .A1(_00811_),
    .A2(_04225_),
    .ZN(_00327_)
  );
  AND2_X1 _09468_ (
    .A1(small_1[2]),
    .A2(_03700_),
    .ZN(_04226_)
  );
  INV_X1 _09469_ (
    .A(_04226_),
    .ZN(_04227_)
  );
  AND2_X1 _09470_ (
    .A1(_00783_),
    .A2(_03655_),
    .ZN(_04228_)
  );
  INV_X1 _09471_ (
    .A(_04228_),
    .ZN(_04229_)
  );
  AND2_X1 _09472_ (
    .A1(small_1[2]),
    .A2(_04229_),
    .ZN(_04230_)
  );
  INV_X1 _09473_ (
    .A(_04230_),
    .ZN(_04231_)
  );
  AND2_X1 _09474_ (
    .A1(_00747_),
    .A2(_04228_),
    .ZN(_04232_)
  );
  INV_X1 _09475_ (
    .A(_04232_),
    .ZN(_04233_)
  );
  AND2_X1 _09476_ (
    .A1(_04231_),
    .A2(_04233_),
    .ZN(_04234_)
  );
  INV_X1 _09477_ (
    .A(_04234_),
    .ZN(_04235_)
  );
  AND2_X1 _09478_ (
    .A1(_03706_),
    .A2(_04235_),
    .ZN(_04236_)
  );
  INV_X1 _09479_ (
    .A(_04236_),
    .ZN(_04237_)
  );
  AND2_X1 _09480_ (
    .A1(_04227_),
    .A2(_04237_),
    .ZN(_04238_)
  );
  AND2_X1 _09481_ (
    .A1(_01774_),
    .A2(_03708_),
    .ZN(_04239_)
  );
  INV_X1 _09482_ (
    .A(_04239_),
    .ZN(_04240_)
  );
  AND2_X1 _09483_ (
    .A1(_04238_),
    .A2(_04240_),
    .ZN(_04241_)
  );
  INV_X1 _09484_ (
    .A(_04241_),
    .ZN(_04242_)
  );
  AND2_X1 _09485_ (
    .A1(_00811_),
    .A2(_04242_),
    .ZN(_00328_)
  );
  AND2_X1 _09486_ (
    .A1(small_1[3]),
    .A2(_03700_),
    .ZN(_04243_)
  );
  INV_X1 _09487_ (
    .A(_04243_),
    .ZN(_04244_)
  );
  AND2_X1 _09488_ (
    .A1(_00783_),
    .A2(_03656_),
    .ZN(_04245_)
  );
  INV_X1 _09489_ (
    .A(_04245_),
    .ZN(_04246_)
  );
  AND2_X1 _09490_ (
    .A1(_00746_),
    .A2(_04245_),
    .ZN(_04247_)
  );
  INV_X1 _09491_ (
    .A(_04247_),
    .ZN(_04248_)
  );
  AND2_X1 _09492_ (
    .A1(small_1[3]),
    .A2(_04246_),
    .ZN(_04249_)
  );
  INV_X1 _09493_ (
    .A(_04249_),
    .ZN(_04250_)
  );
  AND2_X1 _09494_ (
    .A1(_04248_),
    .A2(_04250_),
    .ZN(_04251_)
  );
  INV_X1 _09495_ (
    .A(_04251_),
    .ZN(_04252_)
  );
  AND2_X1 _09496_ (
    .A1(_03710_),
    .A2(_04252_),
    .ZN(_04253_)
  );
  INV_X1 _09497_ (
    .A(_04253_),
    .ZN(_04254_)
  );
  AND2_X1 _09498_ (
    .A1(_04244_),
    .A2(_04254_),
    .ZN(_04255_)
  );
  AND2_X1 _09499_ (
    .A1(_01865_),
    .A2(_03702_),
    .ZN(_04256_)
  );
  INV_X1 _09500_ (
    .A(_04256_),
    .ZN(_04257_)
  );
  AND2_X1 _09501_ (
    .A1(_04255_),
    .A2(_04257_),
    .ZN(_04258_)
  );
  INV_X1 _09502_ (
    .A(_04258_),
    .ZN(_04259_)
  );
  AND2_X1 _09503_ (
    .A1(_00811_),
    .A2(_04259_),
    .ZN(_00329_)
  );
  AND2_X1 _09504_ (
    .A1(_00783_),
    .A2(_03657_),
    .ZN(_04260_)
  );
  INV_X1 _09505_ (
    .A(_04260_),
    .ZN(_04261_)
  );
  AND2_X1 _09506_ (
    .A1(_00745_),
    .A2(_04261_),
    .ZN(_04262_)
  );
  INV_X1 _09507_ (
    .A(_04262_),
    .ZN(_04263_)
  );
  AND2_X1 _09508_ (
    .A1(small_1[4]),
    .A2(_04260_),
    .ZN(_04264_)
  );
  INV_X1 _09509_ (
    .A(_04264_),
    .ZN(_04265_)
  );
  AND2_X1 _09510_ (
    .A1(_03706_),
    .A2(_04265_),
    .ZN(_04266_)
  );
  AND2_X1 _09511_ (
    .A1(_04263_),
    .A2(_04266_),
    .ZN(_04267_)
  );
  INV_X1 _09512_ (
    .A(_04267_),
    .ZN(_04268_)
  );
  AND2_X1 _09513_ (
    .A1(small_1[4]),
    .A2(_03700_),
    .ZN(_04269_)
  );
  INV_X1 _09514_ (
    .A(_04269_),
    .ZN(_04270_)
  );
  AND2_X1 _09515_ (
    .A1(_04268_),
    .A2(_04270_),
    .ZN(_04271_)
  );
  AND2_X1 _09516_ (
    .A1(_01938_),
    .A2(_03702_),
    .ZN(_04272_)
  );
  INV_X1 _09517_ (
    .A(_04272_),
    .ZN(_04273_)
  );
  AND2_X1 _09518_ (
    .A1(_04271_),
    .A2(_04273_),
    .ZN(_04274_)
  );
  INV_X1 _09519_ (
    .A(_04274_),
    .ZN(_04275_)
  );
  AND2_X1 _09520_ (
    .A1(_00811_),
    .A2(_04275_),
    .ZN(_00330_)
  );
  AND2_X1 _09521_ (
    .A1(_02005_),
    .A2(_03702_),
    .ZN(_04276_)
  );
  INV_X1 _09522_ (
    .A(_04276_),
    .ZN(_04277_)
  );
  AND2_X1 _09523_ (
    .A1(small_1[5]),
    .A2(_03700_),
    .ZN(_04278_)
  );
  INV_X1 _09524_ (
    .A(_04278_),
    .ZN(_04279_)
  );
  AND2_X1 _09525_ (
    .A1(_00744_),
    .A2(_04265_),
    .ZN(_04280_)
  );
  INV_X1 _09526_ (
    .A(_04280_),
    .ZN(_04281_)
  );
  AND2_X1 _09527_ (
    .A1(small_1[5]),
    .A2(_04264_),
    .ZN(_04282_)
  );
  INV_X1 _09528_ (
    .A(_04282_),
    .ZN(_04283_)
  );
  AND2_X1 _09529_ (
    .A1(_03706_),
    .A2(_04283_),
    .ZN(_04284_)
  );
  AND2_X1 _09530_ (
    .A1(_04281_),
    .A2(_04284_),
    .ZN(_04285_)
  );
  INV_X1 _09531_ (
    .A(_04285_),
    .ZN(_04286_)
  );
  AND2_X1 _09532_ (
    .A1(_04279_),
    .A2(_04286_),
    .ZN(_04287_)
  );
  AND2_X1 _09533_ (
    .A1(_04277_),
    .A2(_04287_),
    .ZN(_04288_)
  );
  INV_X1 _09534_ (
    .A(_04288_),
    .ZN(_04289_)
  );
  AND2_X1 _09535_ (
    .A1(_00811_),
    .A2(_04289_),
    .ZN(_00331_)
  );
  AND2_X1 _09536_ (
    .A1(_00897_),
    .A2(_00929_),
    .ZN(_04290_)
  );
  MUX2_X1 _09537_ (
    .A(reg_mscratch[0]),
    .B(_01613_),
    .S(_04290_),
    .Z(_00332_)
  );
  MUX2_X1 _09538_ (
    .A(reg_mscratch[1]),
    .B(_01688_),
    .S(_04290_),
    .Z(_00333_)
  );
  MUX2_X1 _09539_ (
    .A(reg_mscratch[2]),
    .B(_01774_),
    .S(_04290_),
    .Z(_00334_)
  );
  MUX2_X1 _09540_ (
    .A(reg_mscratch[3]),
    .B(_01865_),
    .S(_04290_),
    .Z(_00335_)
  );
  MUX2_X1 _09541_ (
    .A(reg_mscratch[4]),
    .B(_01938_),
    .S(_04290_),
    .Z(_00336_)
  );
  MUX2_X1 _09542_ (
    .A(reg_mscratch[5]),
    .B(_02005_),
    .S(_04290_),
    .Z(_00337_)
  );
  MUX2_X1 _09543_ (
    .A(reg_mscratch[6]),
    .B(_02076_),
    .S(_04290_),
    .Z(_00338_)
  );
  MUX2_X1 _09544_ (
    .A(reg_mscratch[7]),
    .B(_02163_),
    .S(_04290_),
    .Z(_00339_)
  );
  MUX2_X1 _09545_ (
    .A(reg_mscratch[8]),
    .B(_01446_),
    .S(_04290_),
    .Z(_00340_)
  );
  MUX2_X1 _09546_ (
    .A(reg_mscratch[9]),
    .B(_01518_),
    .S(_04290_),
    .Z(_00341_)
  );
  MUX2_X1 _09547_ (
    .A(reg_mscratch[10]),
    .B(_02235_),
    .S(_04290_),
    .Z(_00342_)
  );
  MUX2_X1 _09548_ (
    .A(reg_mscratch[11]),
    .B(_02314_),
    .S(_04290_),
    .Z(_00343_)
  );
  MUX2_X1 _09549_ (
    .A(reg_mscratch[12]),
    .B(_02389_),
    .S(_04290_),
    .Z(_00344_)
  );
  MUX2_X1 _09550_ (
    .A(reg_mscratch[13]),
    .B(_02456_),
    .S(_04290_),
    .Z(_00345_)
  );
  MUX2_X1 _09551_ (
    .A(reg_mscratch[14]),
    .B(_02522_),
    .S(_04290_),
    .Z(_00346_)
  );
  MUX2_X1 _09552_ (
    .A(reg_mscratch[15]),
    .B(_02597_),
    .S(_04290_),
    .Z(_00347_)
  );
  MUX2_X1 _09553_ (
    .A(reg_mscratch[16]),
    .B(_01035_),
    .S(_04290_),
    .Z(_00348_)
  );
  MUX2_X1 _09554_ (
    .A(reg_mscratch[17]),
    .B(_02669_),
    .S(_04290_),
    .Z(_00349_)
  );
  MUX2_X1 _09555_ (
    .A(reg_mscratch[18]),
    .B(_01107_),
    .S(_04290_),
    .Z(_00350_)
  );
  MUX2_X1 _09556_ (
    .A(reg_mscratch[19]),
    .B(_01199_),
    .S(_04290_),
    .Z(_00351_)
  );
  MUX2_X1 _09557_ (
    .A(reg_mscratch[20]),
    .B(_01277_),
    .S(_04290_),
    .Z(_00352_)
  );
  MUX2_X1 _09558_ (
    .A(reg_mscratch[21]),
    .B(_02735_),
    .S(_04290_),
    .Z(_00353_)
  );
  MUX2_X1 _09559_ (
    .A(reg_mscratch[22]),
    .B(_02801_),
    .S(_04290_),
    .Z(_00354_)
  );
  MUX2_X1 _09560_ (
    .A(reg_mscratch[23]),
    .B(_01360_),
    .S(_04290_),
    .Z(_00355_)
  );
  MUX2_X1 _09561_ (
    .A(reg_mscratch[24]),
    .B(_02873_),
    .S(_04290_),
    .Z(_00356_)
  );
  MUX2_X1 _09562_ (
    .A(reg_mscratch[25]),
    .B(_02945_),
    .S(_04290_),
    .Z(_00357_)
  );
  MUX2_X1 _09563_ (
    .A(reg_mscratch[26]),
    .B(_03017_),
    .S(_04290_),
    .Z(_00358_)
  );
  MUX2_X1 _09564_ (
    .A(reg_mscratch[27]),
    .B(_03089_),
    .S(_04290_),
    .Z(_00359_)
  );
  MUX2_X1 _09565_ (
    .A(reg_mscratch[28]),
    .B(_03162_),
    .S(_04290_),
    .Z(_00360_)
  );
  MUX2_X1 _09566_ (
    .A(reg_mscratch[29]),
    .B(_03230_),
    .S(_04290_),
    .Z(_00361_)
  );
  MUX2_X1 _09567_ (
    .A(reg_mscratch[30]),
    .B(_03443_),
    .S(_04290_),
    .Z(_00362_)
  );
  MUX2_X1 _09568_ (
    .A(reg_mscratch[31]),
    .B(_03342_),
    .S(_04290_),
    .Z(_00363_)
  );
  MUX2_X1 _09569_ (
    .A(reg_pmp_5_cfg_x),
    .B(_02235_),
    .S(_01364_),
    .Z(_00364_)
  );
  AND2_X1 _09570_ (
    .A1(reg_pmp_2_cfg_l),
    .A2(reg_pmp_2_cfg_a[0]),
    .ZN(_04291_)
  );
  AND2_X1 _09571_ (
    .A1(_00010_),
    .A2(_04291_),
    .ZN(_04292_)
  );
  INV_X1 _09572_ (
    .A(_04292_),
    .ZN(_04293_)
  );
  AND2_X1 _09573_ (
    .A1(_00793_),
    .A2(_04293_),
    .ZN(_04294_)
  );
  AND2_X1 _09574_ (
    .A1(_00897_),
    .A2(_04294_),
    .ZN(_04295_)
  );
  AND2_X1 _09575_ (
    .A1(_01008_),
    .A2(_04295_),
    .ZN(_04296_)
  );
  MUX2_X1 _09576_ (
    .A(reg_pmp_1_addr[0]),
    .B(_01613_),
    .S(_04296_),
    .Z(_00365_)
  );
  MUX2_X1 _09577_ (
    .A(reg_pmp_1_addr[1]),
    .B(_01688_),
    .S(_04296_),
    .Z(_00366_)
  );
  MUX2_X1 _09578_ (
    .A(reg_pmp_1_addr[2]),
    .B(_01774_),
    .S(_04296_),
    .Z(_00367_)
  );
  MUX2_X1 _09579_ (
    .A(reg_pmp_1_addr[3]),
    .B(_01865_),
    .S(_04296_),
    .Z(_00368_)
  );
  MUX2_X1 _09580_ (
    .A(reg_pmp_1_addr[4]),
    .B(_01938_),
    .S(_04296_),
    .Z(_00369_)
  );
  MUX2_X1 _09581_ (
    .A(reg_pmp_1_addr[5]),
    .B(_02005_),
    .S(_04296_),
    .Z(_00370_)
  );
  MUX2_X1 _09582_ (
    .A(reg_pmp_1_addr[6]),
    .B(_02076_),
    .S(_04296_),
    .Z(_00371_)
  );
  MUX2_X1 _09583_ (
    .A(reg_pmp_1_addr[7]),
    .B(_02163_),
    .S(_04296_),
    .Z(_00372_)
  );
  MUX2_X1 _09584_ (
    .A(reg_pmp_1_addr[8]),
    .B(_01446_),
    .S(_04296_),
    .Z(_00373_)
  );
  MUX2_X1 _09585_ (
    .A(reg_pmp_1_addr[9]),
    .B(_01518_),
    .S(_04296_),
    .Z(_00374_)
  );
  MUX2_X1 _09586_ (
    .A(reg_pmp_1_addr[10]),
    .B(_02235_),
    .S(_04296_),
    .Z(_00375_)
  );
  MUX2_X1 _09587_ (
    .A(reg_pmp_1_addr[11]),
    .B(_02314_),
    .S(_04296_),
    .Z(_00376_)
  );
  MUX2_X1 _09588_ (
    .A(reg_pmp_1_addr[12]),
    .B(_02389_),
    .S(_04296_),
    .Z(_00377_)
  );
  MUX2_X1 _09589_ (
    .A(reg_pmp_1_addr[13]),
    .B(_02456_),
    .S(_04296_),
    .Z(_00378_)
  );
  MUX2_X1 _09590_ (
    .A(reg_pmp_1_addr[14]),
    .B(_02522_),
    .S(_04296_),
    .Z(_00379_)
  );
  MUX2_X1 _09591_ (
    .A(reg_pmp_1_addr[15]),
    .B(_02597_),
    .S(_04296_),
    .Z(_00380_)
  );
  MUX2_X1 _09592_ (
    .A(reg_pmp_1_addr[16]),
    .B(_01035_),
    .S(_04296_),
    .Z(_00381_)
  );
  MUX2_X1 _09593_ (
    .A(reg_pmp_1_addr[17]),
    .B(_02669_),
    .S(_04296_),
    .Z(_00382_)
  );
  MUX2_X1 _09594_ (
    .A(reg_pmp_1_addr[18]),
    .B(_01107_),
    .S(_04296_),
    .Z(_00383_)
  );
  MUX2_X1 _09595_ (
    .A(reg_pmp_1_addr[19]),
    .B(_01199_),
    .S(_04296_),
    .Z(_00384_)
  );
  MUX2_X1 _09596_ (
    .A(reg_pmp_1_addr[20]),
    .B(_01277_),
    .S(_04296_),
    .Z(_00385_)
  );
  MUX2_X1 _09597_ (
    .A(reg_pmp_1_addr[21]),
    .B(_02735_),
    .S(_04296_),
    .Z(_00386_)
  );
  MUX2_X1 _09598_ (
    .A(reg_pmp_1_addr[22]),
    .B(_02801_),
    .S(_04296_),
    .Z(_00387_)
  );
  MUX2_X1 _09599_ (
    .A(reg_pmp_1_addr[23]),
    .B(_01360_),
    .S(_04296_),
    .Z(_00388_)
  );
  MUX2_X1 _09600_ (
    .A(reg_pmp_1_addr[24]),
    .B(_02873_),
    .S(_04296_),
    .Z(_00389_)
  );
  MUX2_X1 _09601_ (
    .A(reg_pmp_1_addr[25]),
    .B(_02945_),
    .S(_04296_),
    .Z(_00390_)
  );
  MUX2_X1 _09602_ (
    .A(reg_pmp_1_addr[26]),
    .B(_03017_),
    .S(_04296_),
    .Z(_00391_)
  );
  MUX2_X1 _09603_ (
    .A(reg_pmp_1_addr[27]),
    .B(_03089_),
    .S(_04296_),
    .Z(_00392_)
  );
  MUX2_X1 _09604_ (
    .A(reg_pmp_1_addr[28]),
    .B(_03162_),
    .S(_04296_),
    .Z(_00393_)
  );
  MUX2_X1 _09605_ (
    .A(reg_pmp_1_addr[29]),
    .B(_03230_),
    .S(_04296_),
    .Z(_00394_)
  );
  AND2_X1 _09606_ (
    .A1(reg_pmp_7_cfg_l),
    .A2(reg_pmp_7_cfg_a[0]),
    .ZN(_04297_)
  );
  AND2_X1 _09607_ (
    .A1(_00004_),
    .A2(_04297_),
    .ZN(_04298_)
  );
  INV_X1 _09608_ (
    .A(_04298_),
    .ZN(_04299_)
  );
  AND2_X1 _09609_ (
    .A1(_00808_),
    .A2(_04299_),
    .ZN(_04300_)
  );
  AND2_X1 _09610_ (
    .A1(_00897_),
    .A2(_04300_),
    .ZN(_04301_)
  );
  AND2_X1 _09611_ (
    .A1(_00978_),
    .A2(_04301_),
    .ZN(_04302_)
  );
  MUX2_X1 _09612_ (
    .A(reg_pmp_6_addr[0]),
    .B(_01613_),
    .S(_04302_),
    .Z(_00395_)
  );
  MUX2_X1 _09613_ (
    .A(reg_pmp_6_addr[1]),
    .B(_01688_),
    .S(_04302_),
    .Z(_00396_)
  );
  MUX2_X1 _09614_ (
    .A(reg_pmp_6_addr[2]),
    .B(_01774_),
    .S(_04302_),
    .Z(_00397_)
  );
  MUX2_X1 _09615_ (
    .A(reg_pmp_6_addr[3]),
    .B(_01865_),
    .S(_04302_),
    .Z(_00398_)
  );
  MUX2_X1 _09616_ (
    .A(reg_pmp_6_addr[4]),
    .B(_01938_),
    .S(_04302_),
    .Z(_00399_)
  );
  MUX2_X1 _09617_ (
    .A(reg_pmp_6_addr[5]),
    .B(_02005_),
    .S(_04302_),
    .Z(_00400_)
  );
  MUX2_X1 _09618_ (
    .A(reg_pmp_6_addr[6]),
    .B(_02076_),
    .S(_04302_),
    .Z(_00401_)
  );
  MUX2_X1 _09619_ (
    .A(reg_pmp_6_addr[7]),
    .B(_02163_),
    .S(_04302_),
    .Z(_00402_)
  );
  MUX2_X1 _09620_ (
    .A(reg_pmp_6_addr[8]),
    .B(_01446_),
    .S(_04302_),
    .Z(_00403_)
  );
  MUX2_X1 _09621_ (
    .A(reg_pmp_6_addr[9]),
    .B(_01518_),
    .S(_04302_),
    .Z(_00404_)
  );
  MUX2_X1 _09622_ (
    .A(reg_pmp_6_addr[10]),
    .B(_02235_),
    .S(_04302_),
    .Z(_00405_)
  );
  MUX2_X1 _09623_ (
    .A(reg_pmp_6_addr[11]),
    .B(_02314_),
    .S(_04302_),
    .Z(_00406_)
  );
  MUX2_X1 _09624_ (
    .A(reg_pmp_6_addr[12]),
    .B(_02389_),
    .S(_04302_),
    .Z(_00407_)
  );
  MUX2_X1 _09625_ (
    .A(reg_pmp_6_addr[13]),
    .B(_02456_),
    .S(_04302_),
    .Z(_00408_)
  );
  MUX2_X1 _09626_ (
    .A(reg_pmp_6_addr[14]),
    .B(_02522_),
    .S(_04302_),
    .Z(_00409_)
  );
  MUX2_X1 _09627_ (
    .A(reg_pmp_6_addr[15]),
    .B(_02597_),
    .S(_04302_),
    .Z(_00410_)
  );
  MUX2_X1 _09628_ (
    .A(reg_pmp_6_addr[16]),
    .B(_01035_),
    .S(_04302_),
    .Z(_00411_)
  );
  MUX2_X1 _09629_ (
    .A(reg_pmp_6_addr[17]),
    .B(_02669_),
    .S(_04302_),
    .Z(_00412_)
  );
  MUX2_X1 _09630_ (
    .A(reg_pmp_6_addr[18]),
    .B(_01107_),
    .S(_04302_),
    .Z(_00413_)
  );
  MUX2_X1 _09631_ (
    .A(reg_pmp_6_addr[19]),
    .B(_01199_),
    .S(_04302_),
    .Z(_00414_)
  );
  MUX2_X1 _09632_ (
    .A(reg_pmp_6_addr[20]),
    .B(_01277_),
    .S(_04302_),
    .Z(_00415_)
  );
  MUX2_X1 _09633_ (
    .A(reg_pmp_6_addr[21]),
    .B(_02735_),
    .S(_04302_),
    .Z(_00416_)
  );
  MUX2_X1 _09634_ (
    .A(reg_pmp_6_addr[22]),
    .B(_02801_),
    .S(_04302_),
    .Z(_00417_)
  );
  MUX2_X1 _09635_ (
    .A(reg_pmp_6_addr[23]),
    .B(_01360_),
    .S(_04302_),
    .Z(_00418_)
  );
  MUX2_X1 _09636_ (
    .A(reg_pmp_6_addr[24]),
    .B(_02873_),
    .S(_04302_),
    .Z(_00419_)
  );
  MUX2_X1 _09637_ (
    .A(reg_pmp_6_addr[25]),
    .B(_02945_),
    .S(_04302_),
    .Z(_00420_)
  );
  MUX2_X1 _09638_ (
    .A(reg_pmp_6_addr[26]),
    .B(_03017_),
    .S(_04302_),
    .Z(_00421_)
  );
  MUX2_X1 _09639_ (
    .A(reg_pmp_6_addr[27]),
    .B(_03089_),
    .S(_04302_),
    .Z(_00422_)
  );
  MUX2_X1 _09640_ (
    .A(reg_pmp_6_addr[28]),
    .B(_03162_),
    .S(_04302_),
    .Z(_00423_)
  );
  MUX2_X1 _09641_ (
    .A(reg_pmp_6_addr[29]),
    .B(_03230_),
    .S(_04302_),
    .Z(_00424_)
  );
  AND2_X1 _09642_ (
    .A1(_00897_),
    .A2(_01842_),
    .ZN(_04303_)
  );
  INV_X1 _09643_ (
    .A(_04303_),
    .ZN(_04304_)
  );
  AND2_X1 _09644_ (
    .A1(_01865_),
    .A2(_04303_),
    .ZN(_04305_)
  );
  INV_X1 _09645_ (
    .A(_04305_),
    .ZN(_04306_)
  );
  AND2_X1 _09646_ (
    .A1(reg_custom_0[3]),
    .A2(_04304_),
    .ZN(_04307_)
  );
  INV_X1 _09647_ (
    .A(_04307_),
    .ZN(_04308_)
  );
  AND2_X1 _09648_ (
    .A1(_00811_),
    .A2(_04308_),
    .ZN(_04309_)
  );
  AND2_X1 _09649_ (
    .A1(_04306_),
    .A2(_04309_),
    .ZN(_04310_)
  );
  INV_X1 _09650_ (
    .A(_04310_),
    .ZN(_00425_)
  );
  AND2_X1 _09651_ (
    .A1(io_pc[1]),
    .A2(_01773_),
    .ZN(_04311_)
  );
  INV_X1 _09652_ (
    .A(_04311_),
    .ZN(_04312_)
  );
  AND2_X1 _09653_ (
    .A1(_00897_),
    .A2(_01339_),
    .ZN(_04313_)
  );
  AND2_X1 _09654_ (
    .A1(_04312_),
    .A2(_04313_),
    .ZN(_04314_)
  );
  MUX2_X1 _09655_ (
    .A(_00743_),
    .B(_01612_),
    .S(_04314_),
    .Z(_04315_)
  );
  AND2_X1 _09656_ (
    .A1(_00811_),
    .A2(_04315_),
    .ZN(_04316_)
  );
  INV_X1 _09657_ (
    .A(_04316_),
    .ZN(_00426_)
  );
  MUX2_X1 _09658_ (
    .A(_00742_),
    .B(_01773_),
    .S(_04314_),
    .Z(_04317_)
  );
  AND2_X1 _09659_ (
    .A1(_00811_),
    .A2(_04317_),
    .ZN(_04318_)
  );
  INV_X1 _09660_ (
    .A(_04318_),
    .ZN(_00427_)
  );
  MUX2_X1 _09661_ (
    .A(reg_misa[12]),
    .B(_02389_),
    .S(_04314_),
    .Z(_04319_)
  );
  INV_X1 _09662_ (
    .A(_04319_),
    .ZN(_04320_)
  );
  AND2_X1 _09663_ (
    .A1(_00811_),
    .A2(_04320_),
    .ZN(_04321_)
  );
  INV_X1 _09664_ (
    .A(_04321_),
    .ZN(_00428_)
  );
  AND2_X1 _09665_ (
    .A1(large_[16]),
    .A2(large_[15]),
    .ZN(_04322_)
  );
  AND2_X1 _09666_ (
    .A1(large_[17]),
    .A2(large_[14]),
    .ZN(_04323_)
  );
  AND2_X1 _09667_ (
    .A1(_04322_),
    .A2(_04323_),
    .ZN(_04324_)
  );
  AND2_X1 _09668_ (
    .A1(large_[19]),
    .A2(large_[18]),
    .ZN(_04325_)
  );
  AND2_X1 _09669_ (
    .A1(_04324_),
    .A2(_04325_),
    .ZN(_04326_)
  );
  AND2_X1 _09670_ (
    .A1(large_[11]),
    .A2(large_[10]),
    .ZN(_04327_)
  );
  AND2_X1 _09671_ (
    .A1(small_[4]),
    .A2(small_[3]),
    .ZN(_04328_)
  );
  AND2_X1 _09672_ (
    .A1(small_[5]),
    .A2(_T_14),
    .ZN(_04329_)
  );
  AND2_X1 _09673_ (
    .A1(_04328_),
    .A2(_04329_),
    .ZN(_04330_)
  );
  AND2_X1 _09674_ (
    .A1(small_[0]),
    .A2(io_retire),
    .ZN(_04331_)
  );
  AND2_X1 _09675_ (
    .A1(small_[2]),
    .A2(small_[1]),
    .ZN(_04332_)
  );
  AND2_X1 _09676_ (
    .A1(_04331_),
    .A2(_04332_),
    .ZN(_04333_)
  );
  AND2_X1 _09677_ (
    .A1(_04330_),
    .A2(_04333_),
    .ZN(_04334_)
  );
  AND2_X1 _09678_ (
    .A1(large_[1]),
    .A2(large_[0]),
    .ZN(_04335_)
  );
  AND2_X1 _09679_ (
    .A1(_04334_),
    .A2(_04335_),
    .ZN(_04336_)
  );
  INV_X1 _09680_ (
    .A(_04336_),
    .ZN(_04337_)
  );
  AND2_X1 _09681_ (
    .A1(large_[5]),
    .A2(large_[4]),
    .ZN(_04338_)
  );
  AND2_X1 _09682_ (
    .A1(large_[6]),
    .A2(large_[2]),
    .ZN(_04339_)
  );
  AND2_X1 _09683_ (
    .A1(_04338_),
    .A2(_04339_),
    .ZN(_04340_)
  );
  AND2_X1 _09684_ (
    .A1(large_[3]),
    .A2(_04340_),
    .ZN(_04341_)
  );
  AND2_X1 _09685_ (
    .A1(_04336_),
    .A2(_04341_),
    .ZN(_04342_)
  );
  AND2_X1 _09686_ (
    .A1(large_[7]),
    .A2(_04342_),
    .ZN(_04343_)
  );
  AND2_X1 _09687_ (
    .A1(large_[8]),
    .A2(_04343_),
    .ZN(_04344_)
  );
  AND2_X1 _09688_ (
    .A1(large_[9]),
    .A2(_04344_),
    .ZN(_04345_)
  );
  INV_X1 _09689_ (
    .A(_04345_),
    .ZN(_04346_)
  );
  AND2_X1 _09690_ (
    .A1(_04327_),
    .A2(_04345_),
    .ZN(_04347_)
  );
  INV_X1 _09691_ (
    .A(_04347_),
    .ZN(_04348_)
  );
  AND2_X1 _09692_ (
    .A1(large_[12]),
    .A2(_04347_),
    .ZN(_04349_)
  );
  AND2_X1 _09693_ (
    .A1(large_[13]),
    .A2(_04349_),
    .ZN(_04350_)
  );
  INV_X1 _09694_ (
    .A(_04350_),
    .ZN(_04351_)
  );
  AND2_X1 _09695_ (
    .A1(_04326_),
    .A2(_04350_),
    .ZN(_04352_)
  );
  INV_X1 _09696_ (
    .A(_04352_),
    .ZN(_04353_)
  );
  AND2_X1 _09697_ (
    .A1(large_[20]),
    .A2(_04352_),
    .ZN(_04354_)
  );
  INV_X1 _09698_ (
    .A(_04354_),
    .ZN(_04355_)
  );
  AND2_X1 _09699_ (
    .A1(large_[21]),
    .A2(_04354_),
    .ZN(_04356_)
  );
  INV_X1 _09700_ (
    .A(_04356_),
    .ZN(_04357_)
  );
  AND2_X1 _09701_ (
    .A1(large_[22]),
    .A2(_04356_),
    .ZN(_04358_)
  );
  INV_X1 _09702_ (
    .A(_04358_),
    .ZN(_04359_)
  );
  AND2_X1 _09703_ (
    .A1(large_[23]),
    .A2(_04358_),
    .ZN(_04360_)
  );
  INV_X1 _09704_ (
    .A(_04360_),
    .ZN(_04361_)
  );
  AND2_X1 _09705_ (
    .A1(large_[24]),
    .A2(_04360_),
    .ZN(_04362_)
  );
  INV_X1 _09706_ (
    .A(_04362_),
    .ZN(_04363_)
  );
  AND2_X1 _09707_ (
    .A1(large_[25]),
    .A2(_04362_),
    .ZN(_04364_)
  );
  INV_X1 _09708_ (
    .A(_04364_),
    .ZN(_04365_)
  );
  AND2_X1 _09709_ (
    .A1(large_[21]),
    .A2(large_[20]),
    .ZN(_04366_)
  );
  AND2_X1 _09710_ (
    .A1(large_[23]),
    .A2(large_[22]),
    .ZN(_04367_)
  );
  AND2_X1 _09711_ (
    .A1(large_[25]),
    .A2(large_[24]),
    .ZN(_04368_)
  );
  AND2_X1 _09712_ (
    .A1(_04367_),
    .A2(_04368_),
    .ZN(_04369_)
  );
  AND2_X1 _09713_ (
    .A1(large_[3]),
    .A2(large_[2]),
    .ZN(_04370_)
  );
  AND2_X1 _09714_ (
    .A1(_04335_),
    .A2(_04370_),
    .ZN(_04371_)
  );
  AND2_X1 _09715_ (
    .A1(large_[6]),
    .A2(_04338_),
    .ZN(_04372_)
  );
  AND2_X1 _09716_ (
    .A1(_04371_),
    .A2(_04372_),
    .ZN(_04373_)
  );
  AND2_X1 _09717_ (
    .A1(_04334_),
    .A2(_04373_),
    .ZN(_04374_)
  );
  INV_X1 _09718_ (
    .A(_04374_),
    .ZN(_04375_)
  );
  AND2_X1 _09719_ (
    .A1(large_[9]),
    .A2(large_[7]),
    .ZN(_04376_)
  );
  AND2_X1 _09720_ (
    .A1(large_[8]),
    .A2(_04376_),
    .ZN(_04377_)
  );
  AND2_X1 _09721_ (
    .A1(_04374_),
    .A2(_04377_),
    .ZN(_04378_)
  );
  AND2_X1 _09722_ (
    .A1(large_[12]),
    .A2(_04327_),
    .ZN(_04379_)
  );
  AND2_X1 _09723_ (
    .A1(_04378_),
    .A2(_04379_),
    .ZN(_04380_)
  );
  INV_X1 _09724_ (
    .A(_04380_),
    .ZN(_04381_)
  );
  AND2_X1 _09725_ (
    .A1(large_[13]),
    .A2(_04380_),
    .ZN(_04382_)
  );
  AND2_X1 _09726_ (
    .A1(_04326_),
    .A2(_04382_),
    .ZN(_04383_)
  );
  AND2_X1 _09727_ (
    .A1(_00741_),
    .A2(_04365_),
    .ZN(_04384_)
  );
  INV_X1 _09728_ (
    .A(_04384_),
    .ZN(_04385_)
  );
  AND2_X1 _09729_ (
    .A1(large_[26]),
    .A2(_04364_),
    .ZN(_04386_)
  );
  INV_X1 _09730_ (
    .A(_04386_),
    .ZN(_04387_)
  );
  AND2_X1 _09731_ (
    .A1(_00897_),
    .A2(_00991_),
    .ZN(_04388_)
  );
  INV_X1 _09732_ (
    .A(_04388_),
    .ZN(_04389_)
  );
  AND2_X1 _09733_ (
    .A1(_00897_),
    .A2(_00985_),
    .ZN(_04390_)
  );
  INV_X1 _09734_ (
    .A(_04390_),
    .ZN(_04391_)
  );
  AND2_X1 _09735_ (
    .A1(_00897_),
    .A2(_00992_),
    .ZN(_04392_)
  );
  AND2_X1 _09736_ (
    .A1(_01028_),
    .A2(_04392_),
    .ZN(_04393_)
  );
  AND2_X1 _09737_ (
    .A1(_04389_),
    .A2(_04391_),
    .ZN(_04394_)
  );
  AND2_X1 _09738_ (
    .A1(_04387_),
    .A2(_04394_),
    .ZN(_04395_)
  );
  AND2_X1 _09739_ (
    .A1(_00897_),
    .A2(_01027_),
    .ZN(_04396_)
  );
  INV_X1 _09740_ (
    .A(_04396_),
    .ZN(_04397_)
  );
  AND2_X1 _09741_ (
    .A1(_04389_),
    .A2(_04397_),
    .ZN(_04398_)
  );
  INV_X1 _09742_ (
    .A(_04398_),
    .ZN(_04399_)
  );
  AND2_X1 _09743_ (
    .A1(_04385_),
    .A2(_04395_),
    .ZN(_04400_)
  );
  INV_X1 _09744_ (
    .A(_04400_),
    .ZN(_04401_)
  );
  AND2_X1 _09745_ (
    .A1(_01613_),
    .A2(_04388_),
    .ZN(_04402_)
  );
  INV_X1 _09746_ (
    .A(_04402_),
    .ZN(_04403_)
  );
  AND2_X1 _09747_ (
    .A1(large_[26]),
    .A2(_04390_),
    .ZN(_04404_)
  );
  INV_X1 _09748_ (
    .A(_04404_),
    .ZN(_04405_)
  );
  AND2_X1 _09749_ (
    .A1(_04403_),
    .A2(_04405_),
    .ZN(_04406_)
  );
  AND2_X1 _09750_ (
    .A1(_04401_),
    .A2(_04406_),
    .ZN(_04407_)
  );
  INV_X1 _09751_ (
    .A(_04407_),
    .ZN(_04408_)
  );
  AND2_X1 _09752_ (
    .A1(_00811_),
    .A2(_04408_),
    .ZN(_00429_)
  );
  AND2_X1 _09753_ (
    .A1(large_[27]),
    .A2(_04386_),
    .ZN(_04409_)
  );
  INV_X1 _09754_ (
    .A(_04409_),
    .ZN(_04410_)
  );
  AND2_X1 _09755_ (
    .A1(_00740_),
    .A2(_04387_),
    .ZN(_04411_)
  );
  INV_X1 _09756_ (
    .A(_04411_),
    .ZN(_04412_)
  );
  AND2_X1 _09757_ (
    .A1(_04394_),
    .A2(_04412_),
    .ZN(_04413_)
  );
  AND2_X1 _09758_ (
    .A1(_04410_),
    .A2(_04413_),
    .ZN(_04414_)
  );
  INV_X1 _09759_ (
    .A(_04414_),
    .ZN(_04415_)
  );
  AND2_X1 _09760_ (
    .A1(_01688_),
    .A2(_04388_),
    .ZN(_04416_)
  );
  INV_X1 _09761_ (
    .A(_04416_),
    .ZN(_04417_)
  );
  AND2_X1 _09762_ (
    .A1(large_[27]),
    .A2(_04390_),
    .ZN(_04418_)
  );
  INV_X1 _09763_ (
    .A(_04418_),
    .ZN(_04419_)
  );
  AND2_X1 _09764_ (
    .A1(_04417_),
    .A2(_04419_),
    .ZN(_04420_)
  );
  AND2_X1 _09765_ (
    .A1(_04415_),
    .A2(_04420_),
    .ZN(_04421_)
  );
  INV_X1 _09766_ (
    .A(_04421_),
    .ZN(_04422_)
  );
  AND2_X1 _09767_ (
    .A1(_00811_),
    .A2(_04422_),
    .ZN(_00430_)
  );
  AND2_X1 _09768_ (
    .A1(large_[27]),
    .A2(large_[26]),
    .ZN(_04423_)
  );
  AND2_X1 _09769_ (
    .A1(_04366_),
    .A2(_04423_),
    .ZN(_04424_)
  );
  AND2_X1 _09770_ (
    .A1(_04369_),
    .A2(_04424_),
    .ZN(_04425_)
  );
  AND2_X1 _09771_ (
    .A1(_04383_),
    .A2(_04425_),
    .ZN(_04426_)
  );
  INV_X1 _09772_ (
    .A(_04426_),
    .ZN(_04427_)
  );
  AND2_X1 _09773_ (
    .A1(large_[28]),
    .A2(_04426_),
    .ZN(_04428_)
  );
  INV_X1 _09774_ (
    .A(_04428_),
    .ZN(_04429_)
  );
  AND2_X1 _09775_ (
    .A1(_00739_),
    .A2(_04427_),
    .ZN(_04430_)
  );
  INV_X1 _09776_ (
    .A(_04430_),
    .ZN(_04431_)
  );
  AND2_X1 _09777_ (
    .A1(_04398_),
    .A2(_04429_),
    .ZN(_04432_)
  );
  AND2_X1 _09778_ (
    .A1(_04431_),
    .A2(_04432_),
    .ZN(_04433_)
  );
  INV_X1 _09779_ (
    .A(_04433_),
    .ZN(_04434_)
  );
  AND2_X1 _09780_ (
    .A1(_01774_),
    .A2(_04388_),
    .ZN(_04435_)
  );
  INV_X1 _09781_ (
    .A(_04435_),
    .ZN(_04436_)
  );
  AND2_X1 _09782_ (
    .A1(large_[28]),
    .A2(_04396_),
    .ZN(_04437_)
  );
  INV_X1 _09783_ (
    .A(_04437_),
    .ZN(_04438_)
  );
  AND2_X1 _09784_ (
    .A1(_04434_),
    .A2(_04436_),
    .ZN(_04439_)
  );
  AND2_X1 _09785_ (
    .A1(_04438_),
    .A2(_04439_),
    .ZN(_04440_)
  );
  INV_X1 _09786_ (
    .A(_04440_),
    .ZN(_04441_)
  );
  AND2_X1 _09787_ (
    .A1(_00811_),
    .A2(_04441_),
    .ZN(_00431_)
  );
  AND2_X1 _09788_ (
    .A1(large_[29]),
    .A2(_04428_),
    .ZN(_04442_)
  );
  INV_X1 _09789_ (
    .A(_04442_),
    .ZN(_04443_)
  );
  AND2_X1 _09790_ (
    .A1(_00738_),
    .A2(_04429_),
    .ZN(_04444_)
  );
  INV_X1 _09791_ (
    .A(_04444_),
    .ZN(_04445_)
  );
  AND2_X1 _09792_ (
    .A1(large_[29]),
    .A2(large_[28]),
    .ZN(_04446_)
  );
  AND2_X1 _09793_ (
    .A1(_04426_),
    .A2(_04446_),
    .ZN(_04447_)
  );
  AND2_X1 _09794_ (
    .A1(_04398_),
    .A2(_04443_),
    .ZN(_04448_)
  );
  AND2_X1 _09795_ (
    .A1(_04445_),
    .A2(_04448_),
    .ZN(_04449_)
  );
  INV_X1 _09796_ (
    .A(_04449_),
    .ZN(_04450_)
  );
  AND2_X1 _09797_ (
    .A1(_01865_),
    .A2(_04388_),
    .ZN(_04451_)
  );
  INV_X1 _09798_ (
    .A(_04451_),
    .ZN(_04452_)
  );
  AND2_X1 _09799_ (
    .A1(large_[29]),
    .A2(_04396_),
    .ZN(_04453_)
  );
  INV_X1 _09800_ (
    .A(_04453_),
    .ZN(_04454_)
  );
  AND2_X1 _09801_ (
    .A1(_04450_),
    .A2(_04454_),
    .ZN(_04455_)
  );
  AND2_X1 _09802_ (
    .A1(_04452_),
    .A2(_04455_),
    .ZN(_04456_)
  );
  INV_X1 _09803_ (
    .A(_04456_),
    .ZN(_04457_)
  );
  AND2_X1 _09804_ (
    .A1(_00811_),
    .A2(_04457_),
    .ZN(_00432_)
  );
  AND2_X1 _09805_ (
    .A1(large_[30]),
    .A2(_04442_),
    .ZN(_04458_)
  );
  INV_X1 _09806_ (
    .A(_04458_),
    .ZN(_04459_)
  );
  AND2_X1 _09807_ (
    .A1(_00737_),
    .A2(_04443_),
    .ZN(_04460_)
  );
  INV_X1 _09808_ (
    .A(_04460_),
    .ZN(_04461_)
  );
  AND2_X1 _09809_ (
    .A1(large_[30]),
    .A2(_04447_),
    .ZN(_04462_)
  );
  AND2_X1 _09810_ (
    .A1(_04459_),
    .A2(_04461_),
    .ZN(_04463_)
  );
  AND2_X1 _09811_ (
    .A1(_04398_),
    .A2(_04463_),
    .ZN(_04464_)
  );
  INV_X1 _09812_ (
    .A(_04464_),
    .ZN(_04465_)
  );
  AND2_X1 _09813_ (
    .A1(_01938_),
    .A2(_04388_),
    .ZN(_04466_)
  );
  INV_X1 _09814_ (
    .A(_04466_),
    .ZN(_04467_)
  );
  AND2_X1 _09815_ (
    .A1(large_[30]),
    .A2(_04396_),
    .ZN(_04468_)
  );
  INV_X1 _09816_ (
    .A(_04468_),
    .ZN(_04469_)
  );
  AND2_X1 _09817_ (
    .A1(_04465_),
    .A2(_04467_),
    .ZN(_04470_)
  );
  AND2_X1 _09818_ (
    .A1(_04469_),
    .A2(_04470_),
    .ZN(_04471_)
  );
  INV_X1 _09819_ (
    .A(_04471_),
    .ZN(_04472_)
  );
  AND2_X1 _09820_ (
    .A1(_00811_),
    .A2(_04472_),
    .ZN(_00433_)
  );
  AND2_X1 _09821_ (
    .A1(_00736_),
    .A2(_04459_),
    .ZN(_04473_)
  );
  INV_X1 _09822_ (
    .A(_04473_),
    .ZN(_04474_)
  );
  AND2_X1 _09823_ (
    .A1(large_[31]),
    .A2(_04462_),
    .ZN(_04475_)
  );
  INV_X1 _09824_ (
    .A(_04475_),
    .ZN(_04476_)
  );
  AND2_X1 _09825_ (
    .A1(_04398_),
    .A2(_04476_),
    .ZN(_04477_)
  );
  AND2_X1 _09826_ (
    .A1(_04474_),
    .A2(_04477_),
    .ZN(_04478_)
  );
  INV_X1 _09827_ (
    .A(_04478_),
    .ZN(_04479_)
  );
  AND2_X1 _09828_ (
    .A1(_02005_),
    .A2(_04388_),
    .ZN(_04480_)
  );
  INV_X1 _09829_ (
    .A(_04480_),
    .ZN(_04481_)
  );
  AND2_X1 _09830_ (
    .A1(large_[31]),
    .A2(_04396_),
    .ZN(_04482_)
  );
  INV_X1 _09831_ (
    .A(_04482_),
    .ZN(_04483_)
  );
  AND2_X1 _09832_ (
    .A1(_04479_),
    .A2(_04483_),
    .ZN(_04484_)
  );
  AND2_X1 _09833_ (
    .A1(_04481_),
    .A2(_04484_),
    .ZN(_04485_)
  );
  INV_X1 _09834_ (
    .A(_04485_),
    .ZN(_04486_)
  );
  AND2_X1 _09835_ (
    .A1(_00811_),
    .A2(_04486_),
    .ZN(_00434_)
  );
  AND2_X1 _09836_ (
    .A1(large_[31]),
    .A2(_04446_),
    .ZN(_04487_)
  );
  AND2_X1 _09837_ (
    .A1(large_[30]),
    .A2(_04487_),
    .ZN(_04488_)
  );
  AND2_X1 _09838_ (
    .A1(_04426_),
    .A2(_04488_),
    .ZN(_04489_)
  );
  AND2_X1 _09839_ (
    .A1(_00735_),
    .A2(_04476_),
    .ZN(_04490_)
  );
  INV_X1 _09840_ (
    .A(_04490_),
    .ZN(_04491_)
  );
  AND2_X1 _09841_ (
    .A1(large_[32]),
    .A2(_04475_),
    .ZN(_04492_)
  );
  AND2_X1 _09842_ (
    .A1(large_[32]),
    .A2(_04489_),
    .ZN(_04493_)
  );
  INV_X1 _09843_ (
    .A(_04493_),
    .ZN(_04494_)
  );
  AND2_X1 _09844_ (
    .A1(_04491_),
    .A2(_04494_),
    .ZN(_04495_)
  );
  AND2_X1 _09845_ (
    .A1(_04398_),
    .A2(_04495_),
    .ZN(_04496_)
  );
  INV_X1 _09846_ (
    .A(_04496_),
    .ZN(_04497_)
  );
  AND2_X1 _09847_ (
    .A1(_02076_),
    .A2(_04388_),
    .ZN(_04498_)
  );
  INV_X1 _09848_ (
    .A(_04498_),
    .ZN(_04499_)
  );
  AND2_X1 _09849_ (
    .A1(large_[32]),
    .A2(_04396_),
    .ZN(_04500_)
  );
  INV_X1 _09850_ (
    .A(_04500_),
    .ZN(_04501_)
  );
  AND2_X1 _09851_ (
    .A1(_04497_),
    .A2(_04499_),
    .ZN(_04502_)
  );
  AND2_X1 _09852_ (
    .A1(_04501_),
    .A2(_04502_),
    .ZN(_04503_)
  );
  INV_X1 _09853_ (
    .A(_04503_),
    .ZN(_04504_)
  );
  AND2_X1 _09854_ (
    .A1(_00811_),
    .A2(_04504_),
    .ZN(_00435_)
  );
  AND2_X1 _09855_ (
    .A1(_00734_),
    .A2(_04494_),
    .ZN(_04505_)
  );
  INV_X1 _09856_ (
    .A(_04505_),
    .ZN(_04506_)
  );
  AND2_X1 _09857_ (
    .A1(large_[33]),
    .A2(_04492_),
    .ZN(_04507_)
  );
  INV_X1 _09858_ (
    .A(_04507_),
    .ZN(_04508_)
  );
  AND2_X1 _09859_ (
    .A1(_04398_),
    .A2(_04506_),
    .ZN(_04509_)
  );
  AND2_X1 _09860_ (
    .A1(_04508_),
    .A2(_04509_),
    .ZN(_04510_)
  );
  INV_X1 _09861_ (
    .A(_04510_),
    .ZN(_04511_)
  );
  AND2_X1 _09862_ (
    .A1(_02163_),
    .A2(_04388_),
    .ZN(_04512_)
  );
  INV_X1 _09863_ (
    .A(_04512_),
    .ZN(_04513_)
  );
  AND2_X1 _09864_ (
    .A1(large_[33]),
    .A2(_04396_),
    .ZN(_04514_)
  );
  INV_X1 _09865_ (
    .A(_04514_),
    .ZN(_04515_)
  );
  AND2_X1 _09866_ (
    .A1(_04511_),
    .A2(_04515_),
    .ZN(_04516_)
  );
  AND2_X1 _09867_ (
    .A1(_04513_),
    .A2(_04516_),
    .ZN(_04517_)
  );
  INV_X1 _09868_ (
    .A(_04517_),
    .ZN(_04518_)
  );
  AND2_X1 _09869_ (
    .A1(_00811_),
    .A2(_04518_),
    .ZN(_00436_)
  );
  AND2_X1 _09870_ (
    .A1(_00733_),
    .A2(_04508_),
    .ZN(_04519_)
  );
  INV_X1 _09871_ (
    .A(_04519_),
    .ZN(_04520_)
  );
  AND2_X1 _09872_ (
    .A1(large_[34]),
    .A2(_04507_),
    .ZN(_04521_)
  );
  INV_X1 _09873_ (
    .A(_04521_),
    .ZN(_04522_)
  );
  AND2_X1 _09874_ (
    .A1(_04398_),
    .A2(_04522_),
    .ZN(_04523_)
  );
  AND2_X1 _09875_ (
    .A1(large_[34]),
    .A2(large_[33]),
    .ZN(_04524_)
  );
  AND2_X1 _09876_ (
    .A1(_04520_),
    .A2(_04523_),
    .ZN(_04525_)
  );
  INV_X1 _09877_ (
    .A(_04525_),
    .ZN(_04526_)
  );
  AND2_X1 _09878_ (
    .A1(_01446_),
    .A2(_04388_),
    .ZN(_04527_)
  );
  INV_X1 _09879_ (
    .A(_04527_),
    .ZN(_04528_)
  );
  AND2_X1 _09880_ (
    .A1(large_[34]),
    .A2(_04396_),
    .ZN(_04529_)
  );
  INV_X1 _09881_ (
    .A(_04529_),
    .ZN(_04530_)
  );
  AND2_X1 _09882_ (
    .A1(_04526_),
    .A2(_04530_),
    .ZN(_04531_)
  );
  AND2_X1 _09883_ (
    .A1(_04528_),
    .A2(_04531_),
    .ZN(_04532_)
  );
  INV_X1 _09884_ (
    .A(_04532_),
    .ZN(_04533_)
  );
  AND2_X1 _09885_ (
    .A1(_00811_),
    .A2(_04533_),
    .ZN(_00437_)
  );
  AND2_X1 _09886_ (
    .A1(_00732_),
    .A2(_04522_),
    .ZN(_04534_)
  );
  INV_X1 _09887_ (
    .A(_04534_),
    .ZN(_04535_)
  );
  AND2_X1 _09888_ (
    .A1(large_[35]),
    .A2(_04521_),
    .ZN(_04536_)
  );
  AND2_X1 _09889_ (
    .A1(large_[35]),
    .A2(_04524_),
    .ZN(_04537_)
  );
  AND2_X1 _09890_ (
    .A1(_04493_),
    .A2(_04537_),
    .ZN(_04538_)
  );
  INV_X1 _09891_ (
    .A(_04538_),
    .ZN(_04539_)
  );
  AND2_X1 _09892_ (
    .A1(_04398_),
    .A2(_04539_),
    .ZN(_04540_)
  );
  AND2_X1 _09893_ (
    .A1(_04535_),
    .A2(_04540_),
    .ZN(_04541_)
  );
  INV_X1 _09894_ (
    .A(_04541_),
    .ZN(_04542_)
  );
  AND2_X1 _09895_ (
    .A1(_01518_),
    .A2(_04388_),
    .ZN(_04543_)
  );
  INV_X1 _09896_ (
    .A(_04543_),
    .ZN(_04544_)
  );
  AND2_X1 _09897_ (
    .A1(large_[35]),
    .A2(_04396_),
    .ZN(_04545_)
  );
  INV_X1 _09898_ (
    .A(_04545_),
    .ZN(_04546_)
  );
  AND2_X1 _09899_ (
    .A1(_04542_),
    .A2(_04544_),
    .ZN(_04547_)
  );
  AND2_X1 _09900_ (
    .A1(_04546_),
    .A2(_04547_),
    .ZN(_04548_)
  );
  INV_X1 _09901_ (
    .A(_04548_),
    .ZN(_04549_)
  );
  AND2_X1 _09902_ (
    .A1(_00811_),
    .A2(_04549_),
    .ZN(_00438_)
  );
  AND2_X1 _09903_ (
    .A1(_00731_),
    .A2(_04539_),
    .ZN(_04550_)
  );
  INV_X1 _09904_ (
    .A(_04550_),
    .ZN(_04551_)
  );
  AND2_X1 _09905_ (
    .A1(large_[36]),
    .A2(_04536_),
    .ZN(_04552_)
  );
  AND2_X1 _09906_ (
    .A1(large_[36]),
    .A2(_04538_),
    .ZN(_04553_)
  );
  INV_X1 _09907_ (
    .A(_04553_),
    .ZN(_04554_)
  );
  AND2_X1 _09908_ (
    .A1(_04551_),
    .A2(_04554_),
    .ZN(_04555_)
  );
  AND2_X1 _09909_ (
    .A1(_04398_),
    .A2(_04555_),
    .ZN(_04556_)
  );
  INV_X1 _09910_ (
    .A(_04556_),
    .ZN(_04557_)
  );
  AND2_X1 _09911_ (
    .A1(_02235_),
    .A2(_04388_),
    .ZN(_04558_)
  );
  INV_X1 _09912_ (
    .A(_04558_),
    .ZN(_04559_)
  );
  AND2_X1 _09913_ (
    .A1(large_[36]),
    .A2(_04396_),
    .ZN(_04560_)
  );
  INV_X1 _09914_ (
    .A(_04560_),
    .ZN(_04561_)
  );
  AND2_X1 _09915_ (
    .A1(_04557_),
    .A2(_04559_),
    .ZN(_04562_)
  );
  AND2_X1 _09916_ (
    .A1(_04561_),
    .A2(_04562_),
    .ZN(_04563_)
  );
  INV_X1 _09917_ (
    .A(_04563_),
    .ZN(_04564_)
  );
  AND2_X1 _09918_ (
    .A1(_00811_),
    .A2(_04564_),
    .ZN(_00439_)
  );
  AND2_X1 _09919_ (
    .A1(_00730_),
    .A2(_04554_),
    .ZN(_04565_)
  );
  INV_X1 _09920_ (
    .A(_04565_),
    .ZN(_04566_)
  );
  AND2_X1 _09921_ (
    .A1(large_[37]),
    .A2(large_[36]),
    .ZN(_04567_)
  );
  AND2_X1 _09922_ (
    .A1(large_[37]),
    .A2(_04552_),
    .ZN(_04568_)
  );
  INV_X1 _09923_ (
    .A(_04568_),
    .ZN(_04569_)
  );
  AND2_X1 _09924_ (
    .A1(_04398_),
    .A2(_04566_),
    .ZN(_04570_)
  );
  AND2_X1 _09925_ (
    .A1(_04569_),
    .A2(_04570_),
    .ZN(_04571_)
  );
  INV_X1 _09926_ (
    .A(_04571_),
    .ZN(_04572_)
  );
  AND2_X1 _09927_ (
    .A1(_02314_),
    .A2(_04388_),
    .ZN(_04573_)
  );
  INV_X1 _09928_ (
    .A(_04573_),
    .ZN(_04574_)
  );
  AND2_X1 _09929_ (
    .A1(large_[37]),
    .A2(_04390_),
    .ZN(_04575_)
  );
  INV_X1 _09930_ (
    .A(_04575_),
    .ZN(_04576_)
  );
  AND2_X1 _09931_ (
    .A1(_04574_),
    .A2(_04576_),
    .ZN(_04577_)
  );
  AND2_X1 _09932_ (
    .A1(_04572_),
    .A2(_04577_),
    .ZN(_04578_)
  );
  INV_X1 _09933_ (
    .A(_04578_),
    .ZN(_04579_)
  );
  AND2_X1 _09934_ (
    .A1(_00811_),
    .A2(_04579_),
    .ZN(_00440_)
  );
  AND2_X1 _09935_ (
    .A1(_00729_),
    .A2(_04569_),
    .ZN(_04580_)
  );
  INV_X1 _09936_ (
    .A(_04580_),
    .ZN(_04581_)
  );
  AND2_X1 _09937_ (
    .A1(large_[38]),
    .A2(_04568_),
    .ZN(_04582_)
  );
  INV_X1 _09938_ (
    .A(_04582_),
    .ZN(_04583_)
  );
  AND2_X1 _09939_ (
    .A1(_04398_),
    .A2(_04583_),
    .ZN(_04584_)
  );
  AND2_X1 _09940_ (
    .A1(large_[38]),
    .A2(_04567_),
    .ZN(_04585_)
  );
  AND2_X1 _09941_ (
    .A1(_04581_),
    .A2(_04584_),
    .ZN(_04586_)
  );
  INV_X1 _09942_ (
    .A(_04586_),
    .ZN(_04587_)
  );
  AND2_X1 _09943_ (
    .A1(_02389_),
    .A2(_04388_),
    .ZN(_04588_)
  );
  INV_X1 _09944_ (
    .A(_04588_),
    .ZN(_04589_)
  );
  AND2_X1 _09945_ (
    .A1(large_[38]),
    .A2(_04390_),
    .ZN(_04590_)
  );
  INV_X1 _09946_ (
    .A(_04590_),
    .ZN(_04591_)
  );
  AND2_X1 _09947_ (
    .A1(_04589_),
    .A2(_04591_),
    .ZN(_04592_)
  );
  AND2_X1 _09948_ (
    .A1(_04587_),
    .A2(_04592_),
    .ZN(_04593_)
  );
  INV_X1 _09949_ (
    .A(_04593_),
    .ZN(_04594_)
  );
  AND2_X1 _09950_ (
    .A1(_00811_),
    .A2(_04594_),
    .ZN(_00441_)
  );
  AND2_X1 _09951_ (
    .A1(_00728_),
    .A2(_04583_),
    .ZN(_04595_)
  );
  INV_X1 _09952_ (
    .A(_04595_),
    .ZN(_04596_)
  );
  AND2_X1 _09953_ (
    .A1(_04398_),
    .A2(_04596_),
    .ZN(_04597_)
  );
  AND2_X1 _09954_ (
    .A1(large_[39]),
    .A2(_04582_),
    .ZN(_04598_)
  );
  INV_X1 _09955_ (
    .A(_04598_),
    .ZN(_04599_)
  );
  AND2_X1 _09956_ (
    .A1(_04597_),
    .A2(_04599_),
    .ZN(_04600_)
  );
  INV_X1 _09957_ (
    .A(_04600_),
    .ZN(_04601_)
  );
  AND2_X1 _09958_ (
    .A1(_02456_),
    .A2(_04388_),
    .ZN(_04602_)
  );
  INV_X1 _09959_ (
    .A(_04602_),
    .ZN(_04603_)
  );
  AND2_X1 _09960_ (
    .A1(large_[39]),
    .A2(_04390_),
    .ZN(_04604_)
  );
  INV_X1 _09961_ (
    .A(_04604_),
    .ZN(_04605_)
  );
  AND2_X1 _09962_ (
    .A1(_04603_),
    .A2(_04605_),
    .ZN(_04606_)
  );
  AND2_X1 _09963_ (
    .A1(_04601_),
    .A2(_04606_),
    .ZN(_04607_)
  );
  INV_X1 _09964_ (
    .A(_04607_),
    .ZN(_04608_)
  );
  AND2_X1 _09965_ (
    .A1(_00811_),
    .A2(_04608_),
    .ZN(_00442_)
  );
  AND2_X1 _09966_ (
    .A1(large_[39]),
    .A2(large_[32]),
    .ZN(_04609_)
  );
  AND2_X1 _09967_ (
    .A1(large_[30]),
    .A2(_04609_),
    .ZN(_04610_)
  );
  AND2_X1 _09968_ (
    .A1(_04487_),
    .A2(_04610_),
    .ZN(_04611_)
  );
  AND2_X1 _09969_ (
    .A1(_04537_),
    .A2(_04585_),
    .ZN(_04612_)
  );
  AND2_X1 _09970_ (
    .A1(_04611_),
    .A2(_04612_),
    .ZN(_04613_)
  );
  AND2_X1 _09971_ (
    .A1(_04425_),
    .A2(_04613_),
    .ZN(_04614_)
  );
  AND2_X1 _09972_ (
    .A1(_04352_),
    .A2(_04614_),
    .ZN(_04615_)
  );
  AND2_X1 _09973_ (
    .A1(_04537_),
    .A2(_04609_),
    .ZN(_04616_)
  );
  AND2_X1 _09974_ (
    .A1(_04488_),
    .A2(_04616_),
    .ZN(_04617_)
  );
  AND2_X1 _09975_ (
    .A1(_04425_),
    .A2(_04585_),
    .ZN(_04618_)
  );
  AND2_X1 _09976_ (
    .A1(_04617_),
    .A2(_04618_),
    .ZN(_04619_)
  );
  AND2_X1 _09977_ (
    .A1(_04383_),
    .A2(_04619_),
    .ZN(_04620_)
  );
  INV_X1 _09978_ (
    .A(_04620_),
    .ZN(_04621_)
  );
  AND2_X1 _09979_ (
    .A1(_00727_),
    .A2(_04621_),
    .ZN(_04622_)
  );
  INV_X1 _09980_ (
    .A(_04622_),
    .ZN(_04623_)
  );
  AND2_X1 _09981_ (
    .A1(large_[40]),
    .A2(_04620_),
    .ZN(_04624_)
  );
  INV_X1 _09982_ (
    .A(_04624_),
    .ZN(_04625_)
  );
  AND2_X1 _09983_ (
    .A1(_04623_),
    .A2(_04625_),
    .ZN(_04626_)
  );
  AND2_X1 _09984_ (
    .A1(_04398_),
    .A2(_04626_),
    .ZN(_04627_)
  );
  INV_X1 _09985_ (
    .A(_04627_),
    .ZN(_04628_)
  );
  AND2_X1 _09986_ (
    .A1(_02522_),
    .A2(_04388_),
    .ZN(_04629_)
  );
  INV_X1 _09987_ (
    .A(_04629_),
    .ZN(_04630_)
  );
  AND2_X1 _09988_ (
    .A1(large_[40]),
    .A2(_04396_),
    .ZN(_04631_)
  );
  INV_X1 _09989_ (
    .A(_04631_),
    .ZN(_04632_)
  );
  AND2_X1 _09990_ (
    .A1(_04628_),
    .A2(_04630_),
    .ZN(_04633_)
  );
  AND2_X1 _09991_ (
    .A1(_04632_),
    .A2(_04633_),
    .ZN(_04634_)
  );
  INV_X1 _09992_ (
    .A(_04634_),
    .ZN(_04635_)
  );
  AND2_X1 _09993_ (
    .A1(_00811_),
    .A2(_04635_),
    .ZN(_00443_)
  );
  AND2_X1 _09994_ (
    .A1(_00726_),
    .A2(_04625_),
    .ZN(_04636_)
  );
  INV_X1 _09995_ (
    .A(_04636_),
    .ZN(_04637_)
  );
  AND2_X1 _09996_ (
    .A1(large_[41]),
    .A2(large_[40]),
    .ZN(_04638_)
  );
  AND2_X1 _09997_ (
    .A1(large_[41]),
    .A2(_04624_),
    .ZN(_04639_)
  );
  INV_X1 _09998_ (
    .A(_04639_),
    .ZN(_04640_)
  );
  AND2_X1 _09999_ (
    .A1(_04637_),
    .A2(_04640_),
    .ZN(_04641_)
  );
  AND2_X1 _10000_ (
    .A1(_04398_),
    .A2(_04641_),
    .ZN(_04642_)
  );
  INV_X1 _10001_ (
    .A(_04642_),
    .ZN(_04643_)
  );
  AND2_X1 _10002_ (
    .A1(_02597_),
    .A2(_04388_),
    .ZN(_04644_)
  );
  INV_X1 _10003_ (
    .A(_04644_),
    .ZN(_04645_)
  );
  AND2_X1 _10004_ (
    .A1(large_[41]),
    .A2(_04390_),
    .ZN(_04646_)
  );
  INV_X1 _10005_ (
    .A(_04646_),
    .ZN(_04647_)
  );
  AND2_X1 _10006_ (
    .A1(_04645_),
    .A2(_04647_),
    .ZN(_04648_)
  );
  AND2_X1 _10007_ (
    .A1(_04643_),
    .A2(_04648_),
    .ZN(_04649_)
  );
  INV_X1 _10008_ (
    .A(_04649_),
    .ZN(_04650_)
  );
  AND2_X1 _10009_ (
    .A1(_00811_),
    .A2(_04650_),
    .ZN(_00444_)
  );
  AND2_X1 _10010_ (
    .A1(_00725_),
    .A2(_04640_),
    .ZN(_04651_)
  );
  INV_X1 _10011_ (
    .A(_04651_),
    .ZN(_04652_)
  );
  AND2_X1 _10012_ (
    .A1(large_[42]),
    .A2(_04639_),
    .ZN(_04653_)
  );
  INV_X1 _10013_ (
    .A(_04653_),
    .ZN(_04654_)
  );
  AND2_X1 _10014_ (
    .A1(_04652_),
    .A2(_04654_),
    .ZN(_04655_)
  );
  AND2_X1 _10015_ (
    .A1(_04398_),
    .A2(_04655_),
    .ZN(_04656_)
  );
  INV_X1 _10016_ (
    .A(_04656_),
    .ZN(_04657_)
  );
  AND2_X1 _10017_ (
    .A1(_01035_),
    .A2(_04388_),
    .ZN(_04658_)
  );
  INV_X1 _10018_ (
    .A(_04658_),
    .ZN(_04659_)
  );
  AND2_X1 _10019_ (
    .A1(large_[42]),
    .A2(_04396_),
    .ZN(_04660_)
  );
  INV_X1 _10020_ (
    .A(_04660_),
    .ZN(_04661_)
  );
  AND2_X1 _10021_ (
    .A1(_04657_),
    .A2(_04659_),
    .ZN(_04662_)
  );
  AND2_X1 _10022_ (
    .A1(_04661_),
    .A2(_04662_),
    .ZN(_04663_)
  );
  INV_X1 _10023_ (
    .A(_04663_),
    .ZN(_04664_)
  );
  AND2_X1 _10024_ (
    .A1(_00811_),
    .A2(_04664_),
    .ZN(_00445_)
  );
  AND2_X1 _10025_ (
    .A1(_00724_),
    .A2(_04654_),
    .ZN(_04665_)
  );
  INV_X1 _10026_ (
    .A(_04665_),
    .ZN(_04666_)
  );
  AND2_X1 _10027_ (
    .A1(large_[43]),
    .A2(large_[42]),
    .ZN(_04667_)
  );
  AND2_X1 _10028_ (
    .A1(_04638_),
    .A2(_04667_),
    .ZN(_04668_)
  );
  AND2_X1 _10029_ (
    .A1(_04615_),
    .A2(_04668_),
    .ZN(_04669_)
  );
  INV_X1 _10030_ (
    .A(_04669_),
    .ZN(_04670_)
  );
  AND2_X1 _10031_ (
    .A1(_04398_),
    .A2(_04670_),
    .ZN(_04671_)
  );
  AND2_X1 _10032_ (
    .A1(_04666_),
    .A2(_04671_),
    .ZN(_04672_)
  );
  INV_X1 _10033_ (
    .A(_04672_),
    .ZN(_04673_)
  );
  AND2_X1 _10034_ (
    .A1(_02669_),
    .A2(_04388_),
    .ZN(_04674_)
  );
  INV_X1 _10035_ (
    .A(_04674_),
    .ZN(_04675_)
  );
  AND2_X1 _10036_ (
    .A1(large_[43]),
    .A2(_04390_),
    .ZN(_04676_)
  );
  INV_X1 _10037_ (
    .A(_04676_),
    .ZN(_04677_)
  );
  AND2_X1 _10038_ (
    .A1(_04675_),
    .A2(_04677_),
    .ZN(_04678_)
  );
  AND2_X1 _10039_ (
    .A1(_04673_),
    .A2(_04678_),
    .ZN(_04679_)
  );
  INV_X1 _10040_ (
    .A(_04679_),
    .ZN(_04680_)
  );
  AND2_X1 _10041_ (
    .A1(_00811_),
    .A2(_04680_),
    .ZN(_00446_)
  );
  AND2_X1 _10042_ (
    .A1(_04620_),
    .A2(_04668_),
    .ZN(_04681_)
  );
  AND2_X1 _10043_ (
    .A1(_00723_),
    .A2(_04670_),
    .ZN(_04682_)
  );
  INV_X1 _10044_ (
    .A(_04682_),
    .ZN(_04683_)
  );
  AND2_X1 _10045_ (
    .A1(large_[44]),
    .A2(_04669_),
    .ZN(_04684_)
  );
  INV_X1 _10046_ (
    .A(_04684_),
    .ZN(_04685_)
  );
  AND2_X1 _10047_ (
    .A1(_04398_),
    .A2(_04685_),
    .ZN(_04686_)
  );
  AND2_X1 _10048_ (
    .A1(large_[44]),
    .A2(_04681_),
    .ZN(_04687_)
  );
  AND2_X1 _10049_ (
    .A1(_04683_),
    .A2(_04686_),
    .ZN(_04688_)
  );
  INV_X1 _10050_ (
    .A(_04688_),
    .ZN(_04689_)
  );
  AND2_X1 _10051_ (
    .A1(_01107_),
    .A2(_04388_),
    .ZN(_04690_)
  );
  INV_X1 _10052_ (
    .A(_04690_),
    .ZN(_04691_)
  );
  AND2_X1 _10053_ (
    .A1(large_[44]),
    .A2(_04396_),
    .ZN(_04692_)
  );
  INV_X1 _10054_ (
    .A(_04692_),
    .ZN(_04693_)
  );
  AND2_X1 _10055_ (
    .A1(_04689_),
    .A2(_04691_),
    .ZN(_04694_)
  );
  AND2_X1 _10056_ (
    .A1(_04693_),
    .A2(_04694_),
    .ZN(_04695_)
  );
  INV_X1 _10057_ (
    .A(_04695_),
    .ZN(_04696_)
  );
  AND2_X1 _10058_ (
    .A1(_00811_),
    .A2(_04696_),
    .ZN(_00447_)
  );
  AND2_X1 _10059_ (
    .A1(_00722_),
    .A2(_04685_),
    .ZN(_04697_)
  );
  INV_X1 _10060_ (
    .A(_04697_),
    .ZN(_04698_)
  );
  AND2_X1 _10061_ (
    .A1(_04398_),
    .A2(_04698_),
    .ZN(_04699_)
  );
  AND2_X1 _10062_ (
    .A1(large_[45]),
    .A2(_04684_),
    .ZN(_04700_)
  );
  INV_X1 _10063_ (
    .A(_04700_),
    .ZN(_04701_)
  );
  AND2_X1 _10064_ (
    .A1(_04699_),
    .A2(_04701_),
    .ZN(_04702_)
  );
  INV_X1 _10065_ (
    .A(_04702_),
    .ZN(_04703_)
  );
  AND2_X1 _10066_ (
    .A1(_01199_),
    .A2(_04388_),
    .ZN(_04704_)
  );
  INV_X1 _10067_ (
    .A(_04704_),
    .ZN(_04705_)
  );
  AND2_X1 _10068_ (
    .A1(large_[45]),
    .A2(_04390_),
    .ZN(_04706_)
  );
  INV_X1 _10069_ (
    .A(_04706_),
    .ZN(_04707_)
  );
  AND2_X1 _10070_ (
    .A1(_04705_),
    .A2(_04707_),
    .ZN(_04708_)
  );
  AND2_X1 _10071_ (
    .A1(_04703_),
    .A2(_04708_),
    .ZN(_04709_)
  );
  INV_X1 _10072_ (
    .A(_04709_),
    .ZN(_04710_)
  );
  AND2_X1 _10073_ (
    .A1(_00811_),
    .A2(_04710_),
    .ZN(_00448_)
  );
  AND2_X1 _10074_ (
    .A1(_00721_),
    .A2(_04701_),
    .ZN(_04711_)
  );
  INV_X1 _10075_ (
    .A(_04711_),
    .ZN(_04712_)
  );
  AND2_X1 _10076_ (
    .A1(large_[46]),
    .A2(large_[45]),
    .ZN(_04713_)
  );
  AND2_X1 _10077_ (
    .A1(_04684_),
    .A2(_04713_),
    .ZN(_04714_)
  );
  INV_X1 _10078_ (
    .A(_04714_),
    .ZN(_04715_)
  );
  AND2_X1 _10079_ (
    .A1(_04398_),
    .A2(_04715_),
    .ZN(_04716_)
  );
  AND2_X1 _10080_ (
    .A1(_04687_),
    .A2(_04713_),
    .ZN(_04717_)
  );
  AND2_X1 _10081_ (
    .A1(_04712_),
    .A2(_04716_),
    .ZN(_04718_)
  );
  INV_X1 _10082_ (
    .A(_04718_),
    .ZN(_04719_)
  );
  AND2_X1 _10083_ (
    .A1(_01277_),
    .A2(_04388_),
    .ZN(_04720_)
  );
  INV_X1 _10084_ (
    .A(_04720_),
    .ZN(_04721_)
  );
  AND2_X1 _10085_ (
    .A1(large_[46]),
    .A2(_04390_),
    .ZN(_04722_)
  );
  INV_X1 _10086_ (
    .A(_04722_),
    .ZN(_04723_)
  );
  AND2_X1 _10087_ (
    .A1(_04721_),
    .A2(_04723_),
    .ZN(_04724_)
  );
  AND2_X1 _10088_ (
    .A1(_04719_),
    .A2(_04724_),
    .ZN(_04725_)
  );
  INV_X1 _10089_ (
    .A(_04725_),
    .ZN(_04726_)
  );
  AND2_X1 _10090_ (
    .A1(_00811_),
    .A2(_04726_),
    .ZN(_00449_)
  );
  AND2_X1 _10091_ (
    .A1(_00720_),
    .A2(_04715_),
    .ZN(_04727_)
  );
  INV_X1 _10092_ (
    .A(_04727_),
    .ZN(_04728_)
  );
  AND2_X1 _10093_ (
    .A1(_04398_),
    .A2(_04728_),
    .ZN(_04729_)
  );
  AND2_X1 _10094_ (
    .A1(large_[47]),
    .A2(_04714_),
    .ZN(_04730_)
  );
  INV_X1 _10095_ (
    .A(_04730_),
    .ZN(_04731_)
  );
  AND2_X1 _10096_ (
    .A1(large_[47]),
    .A2(_04717_),
    .ZN(_04732_)
  );
  AND2_X1 _10097_ (
    .A1(_04729_),
    .A2(_04731_),
    .ZN(_04733_)
  );
  INV_X1 _10098_ (
    .A(_04733_),
    .ZN(_04734_)
  );
  AND2_X1 _10099_ (
    .A1(_02735_),
    .A2(_04388_),
    .ZN(_04735_)
  );
  INV_X1 _10100_ (
    .A(_04735_),
    .ZN(_04736_)
  );
  AND2_X1 _10101_ (
    .A1(large_[47]),
    .A2(_04390_),
    .ZN(_04737_)
  );
  INV_X1 _10102_ (
    .A(_04737_),
    .ZN(_04738_)
  );
  AND2_X1 _10103_ (
    .A1(_04736_),
    .A2(_04738_),
    .ZN(_04739_)
  );
  AND2_X1 _10104_ (
    .A1(_04734_),
    .A2(_04739_),
    .ZN(_04740_)
  );
  INV_X1 _10105_ (
    .A(_04740_),
    .ZN(_04741_)
  );
  AND2_X1 _10106_ (
    .A1(_00811_),
    .A2(_04741_),
    .ZN(_00450_)
  );
  AND2_X1 _10107_ (
    .A1(_00719_),
    .A2(_04731_),
    .ZN(_04742_)
  );
  INV_X1 _10108_ (
    .A(_04742_),
    .ZN(_04743_)
  );
  AND2_X1 _10109_ (
    .A1(_04398_),
    .A2(_04743_),
    .ZN(_04744_)
  );
  AND2_X1 _10110_ (
    .A1(large_[48]),
    .A2(_04730_),
    .ZN(_04745_)
  );
  INV_X1 _10111_ (
    .A(_04745_),
    .ZN(_04746_)
  );
  AND2_X1 _10112_ (
    .A1(large_[48]),
    .A2(_04732_),
    .ZN(_04747_)
  );
  AND2_X1 _10113_ (
    .A1(_04744_),
    .A2(_04746_),
    .ZN(_04748_)
  );
  INV_X1 _10114_ (
    .A(_04748_),
    .ZN(_04749_)
  );
  AND2_X1 _10115_ (
    .A1(_02801_),
    .A2(_04388_),
    .ZN(_04750_)
  );
  INV_X1 _10116_ (
    .A(_04750_),
    .ZN(_04751_)
  );
  AND2_X1 _10117_ (
    .A1(large_[48]),
    .A2(_04396_),
    .ZN(_04752_)
  );
  INV_X1 _10118_ (
    .A(_04752_),
    .ZN(_04753_)
  );
  AND2_X1 _10119_ (
    .A1(_04751_),
    .A2(_04753_),
    .ZN(_04754_)
  );
  AND2_X1 _10120_ (
    .A1(_04749_),
    .A2(_04754_),
    .ZN(_04755_)
  );
  INV_X1 _10121_ (
    .A(_04755_),
    .ZN(_04756_)
  );
  AND2_X1 _10122_ (
    .A1(_00811_),
    .A2(_04756_),
    .ZN(_00451_)
  );
  AND2_X1 _10123_ (
    .A1(_00718_),
    .A2(_04746_),
    .ZN(_04757_)
  );
  INV_X1 _10124_ (
    .A(_04757_),
    .ZN(_04758_)
  );
  AND2_X1 _10125_ (
    .A1(_04398_),
    .A2(_04758_),
    .ZN(_04759_)
  );
  AND2_X1 _10126_ (
    .A1(large_[49]),
    .A2(_04745_),
    .ZN(_04760_)
  );
  INV_X1 _10127_ (
    .A(_04760_),
    .ZN(_04761_)
  );
  AND2_X1 _10128_ (
    .A1(large_[49]),
    .A2(_04747_),
    .ZN(_04762_)
  );
  AND2_X1 _10129_ (
    .A1(_04759_),
    .A2(_04761_),
    .ZN(_04763_)
  );
  INV_X1 _10130_ (
    .A(_04763_),
    .ZN(_04764_)
  );
  AND2_X1 _10131_ (
    .A1(_01360_),
    .A2(_04388_),
    .ZN(_04765_)
  );
  INV_X1 _10132_ (
    .A(_04765_),
    .ZN(_04766_)
  );
  AND2_X1 _10133_ (
    .A1(large_[49]),
    .A2(_04396_),
    .ZN(_04767_)
  );
  INV_X1 _10134_ (
    .A(_04767_),
    .ZN(_04768_)
  );
  AND2_X1 _10135_ (
    .A1(_04766_),
    .A2(_04768_),
    .ZN(_04769_)
  );
  AND2_X1 _10136_ (
    .A1(_04764_),
    .A2(_04769_),
    .ZN(_04770_)
  );
  INV_X1 _10137_ (
    .A(_04770_),
    .ZN(_04771_)
  );
  AND2_X1 _10138_ (
    .A1(_00811_),
    .A2(_04771_),
    .ZN(_00452_)
  );
  AND2_X1 _10139_ (
    .A1(_00717_),
    .A2(_04761_),
    .ZN(_04772_)
  );
  INV_X1 _10140_ (
    .A(_04772_),
    .ZN(_04773_)
  );
  AND2_X1 _10141_ (
    .A1(large_[50]),
    .A2(_04760_),
    .ZN(_04774_)
  );
  INV_X1 _10142_ (
    .A(_04774_),
    .ZN(_04775_)
  );
  AND2_X1 _10143_ (
    .A1(_04398_),
    .A2(_04775_),
    .ZN(_04776_)
  );
  AND2_X1 _10144_ (
    .A1(large_[50]),
    .A2(_04762_),
    .ZN(_04777_)
  );
  AND2_X1 _10145_ (
    .A1(_04773_),
    .A2(_04776_),
    .ZN(_04778_)
  );
  INV_X1 _10146_ (
    .A(_04778_),
    .ZN(_04779_)
  );
  AND2_X1 _10147_ (
    .A1(_02873_),
    .A2(_04388_),
    .ZN(_04780_)
  );
  INV_X1 _10148_ (
    .A(_04780_),
    .ZN(_04781_)
  );
  AND2_X1 _10149_ (
    .A1(large_[50]),
    .A2(_04390_),
    .ZN(_04782_)
  );
  INV_X1 _10150_ (
    .A(_04782_),
    .ZN(_04783_)
  );
  AND2_X1 _10151_ (
    .A1(_04781_),
    .A2(_04783_),
    .ZN(_04784_)
  );
  AND2_X1 _10152_ (
    .A1(_04779_),
    .A2(_04784_),
    .ZN(_04785_)
  );
  INV_X1 _10153_ (
    .A(_04785_),
    .ZN(_04786_)
  );
  AND2_X1 _10154_ (
    .A1(_00811_),
    .A2(_04786_),
    .ZN(_00453_)
  );
  AND2_X1 _10155_ (
    .A1(_00716_),
    .A2(_04775_),
    .ZN(_04787_)
  );
  INV_X1 _10156_ (
    .A(_04787_),
    .ZN(_04788_)
  );
  AND2_X1 _10157_ (
    .A1(_04398_),
    .A2(_04788_),
    .ZN(_04789_)
  );
  AND2_X1 _10158_ (
    .A1(large_[51]),
    .A2(_04774_),
    .ZN(_04790_)
  );
  INV_X1 _10159_ (
    .A(_04790_),
    .ZN(_04791_)
  );
  AND2_X1 _10160_ (
    .A1(large_[51]),
    .A2(_04777_),
    .ZN(_04792_)
  );
  AND2_X1 _10161_ (
    .A1(_04789_),
    .A2(_04791_),
    .ZN(_04793_)
  );
  INV_X1 _10162_ (
    .A(_04793_),
    .ZN(_04794_)
  );
  AND2_X1 _10163_ (
    .A1(_02945_),
    .A2(_04388_),
    .ZN(_04795_)
  );
  INV_X1 _10164_ (
    .A(_04795_),
    .ZN(_04796_)
  );
  AND2_X1 _10165_ (
    .A1(large_[51]),
    .A2(_04390_),
    .ZN(_04797_)
  );
  INV_X1 _10166_ (
    .A(_04797_),
    .ZN(_04798_)
  );
  AND2_X1 _10167_ (
    .A1(_04796_),
    .A2(_04798_),
    .ZN(_04799_)
  );
  AND2_X1 _10168_ (
    .A1(_04794_),
    .A2(_04799_),
    .ZN(_04800_)
  );
  INV_X1 _10169_ (
    .A(_04800_),
    .ZN(_04801_)
  );
  AND2_X1 _10170_ (
    .A1(_00811_),
    .A2(_04801_),
    .ZN(_00454_)
  );
  AND2_X1 _10171_ (
    .A1(_00715_),
    .A2(_04791_),
    .ZN(_04802_)
  );
  INV_X1 _10172_ (
    .A(_04802_),
    .ZN(_04803_)
  );
  AND2_X1 _10173_ (
    .A1(large_[52]),
    .A2(_04790_),
    .ZN(_04804_)
  );
  INV_X1 _10174_ (
    .A(_04804_),
    .ZN(_04805_)
  );
  AND2_X1 _10175_ (
    .A1(_04398_),
    .A2(_04805_),
    .ZN(_04806_)
  );
  AND2_X1 _10176_ (
    .A1(large_[52]),
    .A2(_04792_),
    .ZN(_04807_)
  );
  AND2_X1 _10177_ (
    .A1(_04803_),
    .A2(_04806_),
    .ZN(_04808_)
  );
  INV_X1 _10178_ (
    .A(_04808_),
    .ZN(_04809_)
  );
  AND2_X1 _10179_ (
    .A1(_03017_),
    .A2(_04388_),
    .ZN(_04810_)
  );
  INV_X1 _10180_ (
    .A(_04810_),
    .ZN(_04811_)
  );
  AND2_X1 _10181_ (
    .A1(large_[52]),
    .A2(_04390_),
    .ZN(_04812_)
  );
  INV_X1 _10182_ (
    .A(_04812_),
    .ZN(_04813_)
  );
  AND2_X1 _10183_ (
    .A1(_04811_),
    .A2(_04813_),
    .ZN(_04814_)
  );
  AND2_X1 _10184_ (
    .A1(_04809_),
    .A2(_04814_),
    .ZN(_04815_)
  );
  INV_X1 _10185_ (
    .A(_04815_),
    .ZN(_04816_)
  );
  AND2_X1 _10186_ (
    .A1(_00811_),
    .A2(_04816_),
    .ZN(_00455_)
  );
  AND2_X1 _10187_ (
    .A1(_00714_),
    .A2(_04805_),
    .ZN(_04817_)
  );
  INV_X1 _10188_ (
    .A(_04817_),
    .ZN(_04818_)
  );
  AND2_X1 _10189_ (
    .A1(_04398_),
    .A2(_04818_),
    .ZN(_04819_)
  );
  AND2_X1 _10190_ (
    .A1(large_[53]),
    .A2(_04804_),
    .ZN(_04820_)
  );
  INV_X1 _10191_ (
    .A(_04820_),
    .ZN(_04821_)
  );
  AND2_X1 _10192_ (
    .A1(large_[53]),
    .A2(_04807_),
    .ZN(_04822_)
  );
  AND2_X1 _10193_ (
    .A1(_04819_),
    .A2(_04821_),
    .ZN(_04823_)
  );
  INV_X1 _10194_ (
    .A(_04823_),
    .ZN(_04824_)
  );
  AND2_X1 _10195_ (
    .A1(_03089_),
    .A2(_04388_),
    .ZN(_04825_)
  );
  INV_X1 _10196_ (
    .A(_04825_),
    .ZN(_04826_)
  );
  AND2_X1 _10197_ (
    .A1(large_[53]),
    .A2(_04390_),
    .ZN(_04827_)
  );
  INV_X1 _10198_ (
    .A(_04827_),
    .ZN(_04828_)
  );
  AND2_X1 _10199_ (
    .A1(_04826_),
    .A2(_04828_),
    .ZN(_04829_)
  );
  AND2_X1 _10200_ (
    .A1(_04824_),
    .A2(_04829_),
    .ZN(_04830_)
  );
  INV_X1 _10201_ (
    .A(_04830_),
    .ZN(_04831_)
  );
  AND2_X1 _10202_ (
    .A1(_00811_),
    .A2(_04831_),
    .ZN(_00456_)
  );
  AND2_X1 _10203_ (
    .A1(_00713_),
    .A2(_04821_),
    .ZN(_04832_)
  );
  INV_X1 _10204_ (
    .A(_04832_),
    .ZN(_04833_)
  );
  AND2_X1 _10205_ (
    .A1(large_[54]),
    .A2(_04822_),
    .ZN(_04834_)
  );
  INV_X1 _10206_ (
    .A(_04834_),
    .ZN(_04835_)
  );
  AND2_X1 _10207_ (
    .A1(_04398_),
    .A2(_04835_),
    .ZN(_04836_)
  );
  AND2_X1 _10208_ (
    .A1(_04833_),
    .A2(_04836_),
    .ZN(_04837_)
  );
  INV_X1 _10209_ (
    .A(_04837_),
    .ZN(_04838_)
  );
  AND2_X1 _10210_ (
    .A1(_03162_),
    .A2(_04388_),
    .ZN(_04839_)
  );
  INV_X1 _10211_ (
    .A(_04839_),
    .ZN(_04840_)
  );
  AND2_X1 _10212_ (
    .A1(large_[54]),
    .A2(_04390_),
    .ZN(_04841_)
  );
  INV_X1 _10213_ (
    .A(_04841_),
    .ZN(_04842_)
  );
  AND2_X1 _10214_ (
    .A1(_04840_),
    .A2(_04842_),
    .ZN(_04843_)
  );
  AND2_X1 _10215_ (
    .A1(_04838_),
    .A2(_04843_),
    .ZN(_04844_)
  );
  INV_X1 _10216_ (
    .A(_04844_),
    .ZN(_04845_)
  );
  AND2_X1 _10217_ (
    .A1(_00811_),
    .A2(_04845_),
    .ZN(_00457_)
  );
  AND2_X1 _10218_ (
    .A1(_00712_),
    .A2(_04835_),
    .ZN(_04846_)
  );
  INV_X1 _10219_ (
    .A(_04846_),
    .ZN(_04847_)
  );
  AND2_X1 _10220_ (
    .A1(large_[55]),
    .A2(_04834_),
    .ZN(_04848_)
  );
  INV_X1 _10221_ (
    .A(_04848_),
    .ZN(_04849_)
  );
  AND2_X1 _10222_ (
    .A1(_04398_),
    .A2(_04849_),
    .ZN(_04850_)
  );
  AND2_X1 _10223_ (
    .A1(_04847_),
    .A2(_04850_),
    .ZN(_04851_)
  );
  INV_X1 _10224_ (
    .A(_04851_),
    .ZN(_04852_)
  );
  AND2_X1 _10225_ (
    .A1(_03230_),
    .A2(_04388_),
    .ZN(_04853_)
  );
  INV_X1 _10226_ (
    .A(_04853_),
    .ZN(_04854_)
  );
  AND2_X1 _10227_ (
    .A1(large_[55]),
    .A2(_04390_),
    .ZN(_04855_)
  );
  INV_X1 _10228_ (
    .A(_04855_),
    .ZN(_04856_)
  );
  AND2_X1 _10229_ (
    .A1(_04854_),
    .A2(_04856_),
    .ZN(_04857_)
  );
  AND2_X1 _10230_ (
    .A1(_04852_),
    .A2(_04857_),
    .ZN(_04858_)
  );
  INV_X1 _10231_ (
    .A(_04858_),
    .ZN(_04859_)
  );
  AND2_X1 _10232_ (
    .A1(_00811_),
    .A2(_04859_),
    .ZN(_00458_)
  );
  AND2_X1 _10233_ (
    .A1(_00711_),
    .A2(_04849_),
    .ZN(_04860_)
  );
  INV_X1 _10234_ (
    .A(_04860_),
    .ZN(_04861_)
  );
  AND2_X1 _10235_ (
    .A1(large_[56]),
    .A2(_04848_),
    .ZN(_04862_)
  );
  INV_X1 _10236_ (
    .A(_04862_),
    .ZN(_04863_)
  );
  AND2_X1 _10237_ (
    .A1(_04398_),
    .A2(_04863_),
    .ZN(_04864_)
  );
  AND2_X1 _10238_ (
    .A1(_04861_),
    .A2(_04864_),
    .ZN(_04865_)
  );
  INV_X1 _10239_ (
    .A(_04865_),
    .ZN(_04866_)
  );
  AND2_X1 _10240_ (
    .A1(_03443_),
    .A2(_04388_),
    .ZN(_04867_)
  );
  INV_X1 _10241_ (
    .A(_04867_),
    .ZN(_04868_)
  );
  AND2_X1 _10242_ (
    .A1(large_[56]),
    .A2(_04390_),
    .ZN(_04869_)
  );
  INV_X1 _10243_ (
    .A(_04869_),
    .ZN(_04870_)
  );
  AND2_X1 _10244_ (
    .A1(_04868_),
    .A2(_04870_),
    .ZN(_04871_)
  );
  AND2_X1 _10245_ (
    .A1(_04866_),
    .A2(_04871_),
    .ZN(_04872_)
  );
  INV_X1 _10246_ (
    .A(_04872_),
    .ZN(_04873_)
  );
  AND2_X1 _10247_ (
    .A1(_00811_),
    .A2(_04873_),
    .ZN(_00459_)
  );
  AND2_X1 _10248_ (
    .A1(large_[57]),
    .A2(_04863_),
    .ZN(_04874_)
  );
  INV_X1 _10249_ (
    .A(_04874_),
    .ZN(_04875_)
  );
  AND2_X1 _10250_ (
    .A1(_00710_),
    .A2(_04862_),
    .ZN(_04876_)
  );
  INV_X1 _10251_ (
    .A(_04876_),
    .ZN(_04877_)
  );
  AND2_X1 _10252_ (
    .A1(_04875_),
    .A2(_04877_),
    .ZN(_04878_)
  );
  INV_X1 _10253_ (
    .A(_04878_),
    .ZN(_04879_)
  );
  AND2_X1 _10254_ (
    .A1(_04398_),
    .A2(_04879_),
    .ZN(_04880_)
  );
  INV_X1 _10255_ (
    .A(_04880_),
    .ZN(_04881_)
  );
  AND2_X1 _10256_ (
    .A1(_03342_),
    .A2(_04388_),
    .ZN(_04882_)
  );
  INV_X1 _10257_ (
    .A(_04882_),
    .ZN(_04883_)
  );
  AND2_X1 _10258_ (
    .A1(large_[57]),
    .A2(_04390_),
    .ZN(_04884_)
  );
  INV_X1 _10259_ (
    .A(_04884_),
    .ZN(_04885_)
  );
  AND2_X1 _10260_ (
    .A1(_04883_),
    .A2(_04885_),
    .ZN(_04886_)
  );
  AND2_X1 _10261_ (
    .A1(_04881_),
    .A2(_04886_),
    .ZN(_04887_)
  );
  INV_X1 _10262_ (
    .A(_04887_),
    .ZN(_04888_)
  );
  AND2_X1 _10263_ (
    .A1(_00811_),
    .A2(_04888_),
    .ZN(_00460_)
  );
  AND2_X1 _10264_ (
    .A1(_00782_),
    .A2(io_retire),
    .ZN(_04889_)
  );
  INV_X1 _10265_ (
    .A(_04889_),
    .ZN(_04890_)
  );
  AND2_X1 _10266_ (
    .A1(_00782_),
    .A2(_04331_),
    .ZN(_04891_)
  );
  INV_X1 _10267_ (
    .A(_04891_),
    .ZN(_04892_)
  );
  AND2_X1 _10268_ (
    .A1(_00709_),
    .A2(_04890_),
    .ZN(_04893_)
  );
  INV_X1 _10269_ (
    .A(_04893_),
    .ZN(_04894_)
  );
  AND2_X1 _10270_ (
    .A1(_04892_),
    .A2(_04894_),
    .ZN(_04895_)
  );
  AND2_X1 _10271_ (
    .A1(_04393_),
    .A2(_04895_),
    .ZN(_04896_)
  );
  INV_X1 _10272_ (
    .A(_04896_),
    .ZN(_04897_)
  );
  AND2_X1 _10273_ (
    .A1(small_[0]),
    .A2(_04388_),
    .ZN(_04898_)
  );
  INV_X1 _10274_ (
    .A(_04898_),
    .ZN(_04899_)
  );
  AND2_X1 _10275_ (
    .A1(_00898_),
    .A2(_04895_),
    .ZN(_04900_)
  );
  INV_X1 _10276_ (
    .A(_04900_),
    .ZN(_04901_)
  );
  AND2_X1 _10277_ (
    .A1(_04899_),
    .A2(_04901_),
    .ZN(_04902_)
  );
  AND2_X1 _10278_ (
    .A1(_04897_),
    .A2(_04902_),
    .ZN(_04903_)
  );
  AND2_X1 _10279_ (
    .A1(_01613_),
    .A2(_04396_),
    .ZN(_04904_)
  );
  INV_X1 _10280_ (
    .A(_04904_),
    .ZN(_04905_)
  );
  AND2_X1 _10281_ (
    .A1(_04903_),
    .A2(_04905_),
    .ZN(_04906_)
  );
  INV_X1 _10282_ (
    .A(_04906_),
    .ZN(_04907_)
  );
  AND2_X1 _10283_ (
    .A1(_00811_),
    .A2(_04907_),
    .ZN(_00461_)
  );
  AND2_X1 _10284_ (
    .A1(_00708_),
    .A2(_04892_),
    .ZN(_04908_)
  );
  INV_X1 _10285_ (
    .A(_04908_),
    .ZN(_04909_)
  );
  AND2_X1 _10286_ (
    .A1(small_[1]),
    .A2(_04388_),
    .ZN(_04910_)
  );
  INV_X1 _10287_ (
    .A(_04910_),
    .ZN(_04911_)
  );
  AND2_X1 _10288_ (
    .A1(small_[1]),
    .A2(_04891_),
    .ZN(_04912_)
  );
  INV_X1 _10289_ (
    .A(_04912_),
    .ZN(_04913_)
  );
  AND2_X1 _10290_ (
    .A1(_04394_),
    .A2(_04913_),
    .ZN(_04914_)
  );
  INV_X1 _10291_ (
    .A(_04914_),
    .ZN(_04915_)
  );
  AND2_X1 _10292_ (
    .A1(_04911_),
    .A2(_04915_),
    .ZN(_04916_)
  );
  INV_X1 _10293_ (
    .A(_04916_),
    .ZN(_04917_)
  );
  AND2_X1 _10294_ (
    .A1(_04909_),
    .A2(_04917_),
    .ZN(_04918_)
  );
  INV_X1 _10295_ (
    .A(_04918_),
    .ZN(_04919_)
  );
  AND2_X1 _10296_ (
    .A1(_01688_),
    .A2(_04396_),
    .ZN(_04920_)
  );
  INV_X1 _10297_ (
    .A(_04920_),
    .ZN(_04921_)
  );
  AND2_X1 _10298_ (
    .A1(_04919_),
    .A2(_04921_),
    .ZN(_04922_)
  );
  INV_X1 _10299_ (
    .A(_04922_),
    .ZN(_04923_)
  );
  AND2_X1 _10300_ (
    .A1(_00811_),
    .A2(_04923_),
    .ZN(_00462_)
  );
  AND2_X1 _10301_ (
    .A1(small_[2]),
    .A2(_04388_),
    .ZN(_04924_)
  );
  INV_X1 _10302_ (
    .A(_04924_),
    .ZN(_04925_)
  );
  AND2_X1 _10303_ (
    .A1(_00782_),
    .A2(_04333_),
    .ZN(_04926_)
  );
  INV_X1 _10304_ (
    .A(_04926_),
    .ZN(_04927_)
  );
  AND2_X1 _10305_ (
    .A1(_00707_),
    .A2(_04913_),
    .ZN(_04928_)
  );
  INV_X1 _10306_ (
    .A(_04928_),
    .ZN(_04929_)
  );
  AND2_X1 _10307_ (
    .A1(_04927_),
    .A2(_04929_),
    .ZN(_04930_)
  );
  AND2_X1 _10308_ (
    .A1(_04394_),
    .A2(_04930_),
    .ZN(_04931_)
  );
  INV_X1 _10309_ (
    .A(_04931_),
    .ZN(_04932_)
  );
  AND2_X1 _10310_ (
    .A1(_04925_),
    .A2(_04932_),
    .ZN(_04933_)
  );
  AND2_X1 _10311_ (
    .A1(_01774_),
    .A2(_04390_),
    .ZN(_04934_)
  );
  INV_X1 _10312_ (
    .A(_04934_),
    .ZN(_04935_)
  );
  AND2_X1 _10313_ (
    .A1(_04933_),
    .A2(_04935_),
    .ZN(_04936_)
  );
  INV_X1 _10314_ (
    .A(_04936_),
    .ZN(_04937_)
  );
  AND2_X1 _10315_ (
    .A1(_00811_),
    .A2(_04937_),
    .ZN(_00463_)
  );
  AND2_X1 _10316_ (
    .A1(_00706_),
    .A2(_04927_),
    .ZN(_04938_)
  );
  INV_X1 _10317_ (
    .A(_04938_),
    .ZN(_04939_)
  );
  AND2_X1 _10318_ (
    .A1(small_[3]),
    .A2(_04388_),
    .ZN(_04940_)
  );
  INV_X1 _10319_ (
    .A(_04940_),
    .ZN(_04941_)
  );
  AND2_X1 _10320_ (
    .A1(small_[3]),
    .A2(_04926_),
    .ZN(_04942_)
  );
  INV_X1 _10321_ (
    .A(_04942_),
    .ZN(_04943_)
  );
  AND2_X1 _10322_ (
    .A1(_04398_),
    .A2(_04943_),
    .ZN(_04944_)
  );
  INV_X1 _10323_ (
    .A(_04944_),
    .ZN(_04945_)
  );
  AND2_X1 _10324_ (
    .A1(_04941_),
    .A2(_04945_),
    .ZN(_04946_)
  );
  INV_X1 _10325_ (
    .A(_04946_),
    .ZN(_04947_)
  );
  AND2_X1 _10326_ (
    .A1(_04939_),
    .A2(_04947_),
    .ZN(_04948_)
  );
  INV_X1 _10327_ (
    .A(_04948_),
    .ZN(_04949_)
  );
  AND2_X1 _10328_ (
    .A1(_01865_),
    .A2(_04390_),
    .ZN(_04950_)
  );
  INV_X1 _10329_ (
    .A(_04950_),
    .ZN(_04951_)
  );
  AND2_X1 _10330_ (
    .A1(_04949_),
    .A2(_04951_),
    .ZN(_04952_)
  );
  INV_X1 _10331_ (
    .A(_04952_),
    .ZN(_04953_)
  );
  AND2_X1 _10332_ (
    .A1(_00811_),
    .A2(_04953_),
    .ZN(_00464_)
  );
  AND2_X1 _10333_ (
    .A1(_00705_),
    .A2(_04943_),
    .ZN(_04954_)
  );
  INV_X1 _10334_ (
    .A(_04954_),
    .ZN(_04955_)
  );
  AND2_X1 _10335_ (
    .A1(small_[4]),
    .A2(_04388_),
    .ZN(_04956_)
  );
  INV_X1 _10336_ (
    .A(_04956_),
    .ZN(_04957_)
  );
  AND2_X1 _10337_ (
    .A1(_04328_),
    .A2(_04926_),
    .ZN(_04958_)
  );
  INV_X1 _10338_ (
    .A(_04958_),
    .ZN(_04959_)
  );
  AND2_X1 _10339_ (
    .A1(_04394_),
    .A2(_04959_),
    .ZN(_04960_)
  );
  INV_X1 _10340_ (
    .A(_04960_),
    .ZN(_04961_)
  );
  AND2_X1 _10341_ (
    .A1(_04957_),
    .A2(_04961_),
    .ZN(_04962_)
  );
  INV_X1 _10342_ (
    .A(_04962_),
    .ZN(_04963_)
  );
  AND2_X1 _10343_ (
    .A1(_04955_),
    .A2(_04963_),
    .ZN(_04964_)
  );
  INV_X1 _10344_ (
    .A(_04964_),
    .ZN(_04965_)
  );
  AND2_X1 _10345_ (
    .A1(_01938_),
    .A2(_04396_),
    .ZN(_04966_)
  );
  INV_X1 _10346_ (
    .A(_04966_),
    .ZN(_04967_)
  );
  AND2_X1 _10347_ (
    .A1(_04965_),
    .A2(_04967_),
    .ZN(_04968_)
  );
  INV_X1 _10348_ (
    .A(_04968_),
    .ZN(_04969_)
  );
  AND2_X1 _10349_ (
    .A1(_00811_),
    .A2(_04969_),
    .ZN(_00465_)
  );
  AND2_X1 _10350_ (
    .A1(small_[5]),
    .A2(_04958_),
    .ZN(_04970_)
  );
  INV_X1 _10351_ (
    .A(_04970_),
    .ZN(_04971_)
  );
  AND2_X1 _10352_ (
    .A1(small_[5]),
    .A2(_04388_),
    .ZN(_04972_)
  );
  INV_X1 _10353_ (
    .A(_04972_),
    .ZN(_04973_)
  );
  AND2_X1 _10354_ (
    .A1(_00704_),
    .A2(_04959_),
    .ZN(_04974_)
  );
  INV_X1 _10355_ (
    .A(_04974_),
    .ZN(_04975_)
  );
  AND2_X1 _10356_ (
    .A1(_04971_),
    .A2(_04975_),
    .ZN(_04976_)
  );
  AND2_X1 _10357_ (
    .A1(_04398_),
    .A2(_04976_),
    .ZN(_04977_)
  );
  INV_X1 _10358_ (
    .A(_04977_),
    .ZN(_04978_)
  );
  AND2_X1 _10359_ (
    .A1(_04973_),
    .A2(_04978_),
    .ZN(_04979_)
  );
  AND2_X1 _10360_ (
    .A1(_02005_),
    .A2(_04396_),
    .ZN(_04980_)
  );
  INV_X1 _10361_ (
    .A(_04980_),
    .ZN(_04981_)
  );
  AND2_X1 _10362_ (
    .A1(_04979_),
    .A2(_04981_),
    .ZN(_04982_)
  );
  INV_X1 _10363_ (
    .A(_04982_),
    .ZN(_04983_)
  );
  AND2_X1 _10364_ (
    .A1(_00811_),
    .A2(_04983_),
    .ZN(_00466_)
  );
  AND2_X1 _10365_ (
    .A1(_00897_),
    .A2(_00940_),
    .ZN(_04984_)
  );
  INV_X1 _10366_ (
    .A(_04984_),
    .ZN(_04985_)
  );
  AND2_X1 _10367_ (
    .A1(_01612_),
    .A2(_04984_),
    .ZN(_04986_)
  );
  INV_X1 _10368_ (
    .A(_04986_),
    .ZN(_04987_)
  );
  AND2_X1 _10369_ (
    .A1(_00703_),
    .A2(_04985_),
    .ZN(_04988_)
  );
  INV_X1 _10370_ (
    .A(_04988_),
    .ZN(_04989_)
  );
  AND2_X1 _10371_ (
    .A1(_00811_),
    .A2(_04989_),
    .ZN(_04990_)
  );
  AND2_X1 _10372_ (
    .A1(_04987_),
    .A2(_04990_),
    .ZN(_00467_)
  );
  AND2_X1 _10373_ (
    .A1(_01773_),
    .A2(_04984_),
    .ZN(_04991_)
  );
  INV_X1 _10374_ (
    .A(_04991_),
    .ZN(_04992_)
  );
  AND2_X1 _10375_ (
    .A1(_00702_),
    .A2(_04985_),
    .ZN(_04993_)
  );
  INV_X1 _10376_ (
    .A(_04993_),
    .ZN(_04994_)
  );
  AND2_X1 _10377_ (
    .A1(_00811_),
    .A2(_04994_),
    .ZN(_04995_)
  );
  AND2_X1 _10378_ (
    .A1(_04992_),
    .A2(_04995_),
    .ZN(_00468_)
  );
  AND2_X1 _10379_ (
    .A1(_01864_),
    .A2(_04984_),
    .ZN(_04996_)
  );
  INV_X1 _10380_ (
    .A(_04996_),
    .ZN(_04997_)
  );
  AND2_X1 _10381_ (
    .A1(_00701_),
    .A2(_04985_),
    .ZN(_04998_)
  );
  INV_X1 _10382_ (
    .A(_04998_),
    .ZN(_04999_)
  );
  AND2_X1 _10383_ (
    .A1(_00811_),
    .A2(_04999_),
    .ZN(_05000_)
  );
  AND2_X1 _10384_ (
    .A1(_04997_),
    .A2(_05000_),
    .ZN(_00469_)
  );
  AND2_X1 _10385_ (
    .A1(_01937_),
    .A2(_04984_),
    .ZN(_05001_)
  );
  INV_X1 _10386_ (
    .A(_05001_),
    .ZN(_05002_)
  );
  AND2_X1 _10387_ (
    .A1(_00700_),
    .A2(_04985_),
    .ZN(_05003_)
  );
  INV_X1 _10388_ (
    .A(_05003_),
    .ZN(_05004_)
  );
  AND2_X1 _10389_ (
    .A1(_00811_),
    .A2(_05004_),
    .ZN(_05005_)
  );
  AND2_X1 _10390_ (
    .A1(_05002_),
    .A2(_05005_),
    .ZN(_00470_)
  );
  AND2_X1 _10391_ (
    .A1(_02004_),
    .A2(_04984_),
    .ZN(_05006_)
  );
  INV_X1 _10392_ (
    .A(_05006_),
    .ZN(_05007_)
  );
  AND2_X1 _10393_ (
    .A1(_00699_),
    .A2(_04985_),
    .ZN(_05008_)
  );
  INV_X1 _10394_ (
    .A(_05008_),
    .ZN(_05009_)
  );
  AND2_X1 _10395_ (
    .A1(_00811_),
    .A2(_05009_),
    .ZN(_05010_)
  );
  AND2_X1 _10396_ (
    .A1(_05007_),
    .A2(_05010_),
    .ZN(_00471_)
  );
  AND2_X1 _10397_ (
    .A1(_02075_),
    .A2(_04984_),
    .ZN(_05011_)
  );
  INV_X1 _10398_ (
    .A(_05011_),
    .ZN(_05012_)
  );
  AND2_X1 _10399_ (
    .A1(_00698_),
    .A2(_04985_),
    .ZN(_05013_)
  );
  INV_X1 _10400_ (
    .A(_05013_),
    .ZN(_05014_)
  );
  AND2_X1 _10401_ (
    .A1(_00811_),
    .A2(_05014_),
    .ZN(_05015_)
  );
  AND2_X1 _10402_ (
    .A1(_05012_),
    .A2(_05015_),
    .ZN(_00472_)
  );
  AND2_X1 _10403_ (
    .A1(_02162_),
    .A2(_04984_),
    .ZN(_05016_)
  );
  INV_X1 _10404_ (
    .A(_05016_),
    .ZN(_05017_)
  );
  AND2_X1 _10405_ (
    .A1(_00697_),
    .A2(_04985_),
    .ZN(_05018_)
  );
  INV_X1 _10406_ (
    .A(_05018_),
    .ZN(_05019_)
  );
  AND2_X1 _10407_ (
    .A1(_00811_),
    .A2(_05019_),
    .ZN(_05020_)
  );
  AND2_X1 _10408_ (
    .A1(_05017_),
    .A2(_05020_),
    .ZN(_00473_)
  );
  AND2_X1 _10409_ (
    .A1(_01445_),
    .A2(_04984_),
    .ZN(_05021_)
  );
  INV_X1 _10410_ (
    .A(_05021_),
    .ZN(_05022_)
  );
  AND2_X1 _10411_ (
    .A1(_00696_),
    .A2(_04985_),
    .ZN(_05023_)
  );
  INV_X1 _10412_ (
    .A(_05023_),
    .ZN(_05024_)
  );
  AND2_X1 _10413_ (
    .A1(_00811_),
    .A2(_05024_),
    .ZN(_05025_)
  );
  AND2_X1 _10414_ (
    .A1(_05022_),
    .A2(_05025_),
    .ZN(_00474_)
  );
  AND2_X1 _10415_ (
    .A1(_01517_),
    .A2(_04984_),
    .ZN(_05026_)
  );
  INV_X1 _10416_ (
    .A(_05026_),
    .ZN(_05027_)
  );
  AND2_X1 _10417_ (
    .A1(_00695_),
    .A2(_04985_),
    .ZN(_05028_)
  );
  INV_X1 _10418_ (
    .A(_05028_),
    .ZN(_05029_)
  );
  AND2_X1 _10419_ (
    .A1(_00811_),
    .A2(_05029_),
    .ZN(_05030_)
  );
  AND2_X1 _10420_ (
    .A1(_05027_),
    .A2(_05030_),
    .ZN(_00475_)
  );
  AND2_X1 _10421_ (
    .A1(_02234_),
    .A2(_04984_),
    .ZN(_05031_)
  );
  INV_X1 _10422_ (
    .A(_05031_),
    .ZN(_05032_)
  );
  AND2_X1 _10423_ (
    .A1(_00694_),
    .A2(_04985_),
    .ZN(_05033_)
  );
  INV_X1 _10424_ (
    .A(_05033_),
    .ZN(_05034_)
  );
  AND2_X1 _10425_ (
    .A1(_00811_),
    .A2(_05034_),
    .ZN(_05035_)
  );
  AND2_X1 _10426_ (
    .A1(_05032_),
    .A2(_05035_),
    .ZN(_00476_)
  );
  AND2_X1 _10427_ (
    .A1(_02313_),
    .A2(_04984_),
    .ZN(_05036_)
  );
  INV_X1 _10428_ (
    .A(_05036_),
    .ZN(_05037_)
  );
  AND2_X1 _10429_ (
    .A1(_00693_),
    .A2(_04985_),
    .ZN(_05038_)
  );
  INV_X1 _10430_ (
    .A(_05038_),
    .ZN(_05039_)
  );
  AND2_X1 _10431_ (
    .A1(_00811_),
    .A2(_05039_),
    .ZN(_05040_)
  );
  AND2_X1 _10432_ (
    .A1(_05037_),
    .A2(_05040_),
    .ZN(_00477_)
  );
  AND2_X1 _10433_ (
    .A1(_02390_),
    .A2(_04984_),
    .ZN(_05041_)
  );
  INV_X1 _10434_ (
    .A(_05041_),
    .ZN(_05042_)
  );
  AND2_X1 _10435_ (
    .A1(_00692_),
    .A2(_04985_),
    .ZN(_05043_)
  );
  INV_X1 _10436_ (
    .A(_05043_),
    .ZN(_05044_)
  );
  AND2_X1 _10437_ (
    .A1(_00811_),
    .A2(_05044_),
    .ZN(_05045_)
  );
  AND2_X1 _10438_ (
    .A1(_05042_),
    .A2(_05045_),
    .ZN(_00478_)
  );
  AND2_X1 _10439_ (
    .A1(_02455_),
    .A2(_04984_),
    .ZN(_05046_)
  );
  INV_X1 _10440_ (
    .A(_05046_),
    .ZN(_05047_)
  );
  AND2_X1 _10441_ (
    .A1(_00691_),
    .A2(_04985_),
    .ZN(_05048_)
  );
  INV_X1 _10442_ (
    .A(_05048_),
    .ZN(_05049_)
  );
  AND2_X1 _10443_ (
    .A1(_00811_),
    .A2(_05049_),
    .ZN(_05050_)
  );
  AND2_X1 _10444_ (
    .A1(_05047_),
    .A2(_05050_),
    .ZN(_00479_)
  );
  AND2_X1 _10445_ (
    .A1(_02521_),
    .A2(_04984_),
    .ZN(_05051_)
  );
  INV_X1 _10446_ (
    .A(_05051_),
    .ZN(_05052_)
  );
  AND2_X1 _10447_ (
    .A1(_00690_),
    .A2(_04985_),
    .ZN(_05053_)
  );
  INV_X1 _10448_ (
    .A(_05053_),
    .ZN(_05054_)
  );
  AND2_X1 _10449_ (
    .A1(_00811_),
    .A2(_05054_),
    .ZN(_05055_)
  );
  AND2_X1 _10450_ (
    .A1(_05052_),
    .A2(_05055_),
    .ZN(_00480_)
  );
  AND2_X1 _10451_ (
    .A1(_02596_),
    .A2(_04984_),
    .ZN(_05056_)
  );
  INV_X1 _10452_ (
    .A(_05056_),
    .ZN(_05057_)
  );
  AND2_X1 _10453_ (
    .A1(_00689_),
    .A2(_04985_),
    .ZN(_05058_)
  );
  INV_X1 _10454_ (
    .A(_05058_),
    .ZN(_05059_)
  );
  AND2_X1 _10455_ (
    .A1(_00811_),
    .A2(_05059_),
    .ZN(_05060_)
  );
  AND2_X1 _10456_ (
    .A1(_05057_),
    .A2(_05060_),
    .ZN(_00481_)
  );
  AND2_X1 _10457_ (
    .A1(_01034_),
    .A2(_04984_),
    .ZN(_05061_)
  );
  INV_X1 _10458_ (
    .A(_05061_),
    .ZN(_05062_)
  );
  AND2_X1 _10459_ (
    .A1(_00688_),
    .A2(_04985_),
    .ZN(_05063_)
  );
  INV_X1 _10460_ (
    .A(_05063_),
    .ZN(_05064_)
  );
  AND2_X1 _10461_ (
    .A1(_00811_),
    .A2(_05064_),
    .ZN(_05065_)
  );
  AND2_X1 _10462_ (
    .A1(_05062_),
    .A2(_05065_),
    .ZN(_00482_)
  );
  AND2_X1 _10463_ (
    .A1(_02668_),
    .A2(_04984_),
    .ZN(_05066_)
  );
  INV_X1 _10464_ (
    .A(_05066_),
    .ZN(_05067_)
  );
  AND2_X1 _10465_ (
    .A1(_00687_),
    .A2(_04985_),
    .ZN(_05068_)
  );
  INV_X1 _10466_ (
    .A(_05068_),
    .ZN(_05069_)
  );
  AND2_X1 _10467_ (
    .A1(_00811_),
    .A2(_05069_),
    .ZN(_05070_)
  );
  AND2_X1 _10468_ (
    .A1(_05067_),
    .A2(_05070_),
    .ZN(_00483_)
  );
  AND2_X1 _10469_ (
    .A1(_01106_),
    .A2(_04984_),
    .ZN(_05071_)
  );
  INV_X1 _10470_ (
    .A(_05071_),
    .ZN(_05072_)
  );
  AND2_X1 _10471_ (
    .A1(_00686_),
    .A2(_04985_),
    .ZN(_05073_)
  );
  INV_X1 _10472_ (
    .A(_05073_),
    .ZN(_05074_)
  );
  AND2_X1 _10473_ (
    .A1(_00811_),
    .A2(_05074_),
    .ZN(_05075_)
  );
  AND2_X1 _10474_ (
    .A1(_05072_),
    .A2(_05075_),
    .ZN(_00484_)
  );
  AND2_X1 _10475_ (
    .A1(_01198_),
    .A2(_04984_),
    .ZN(_05076_)
  );
  INV_X1 _10476_ (
    .A(_05076_),
    .ZN(_05077_)
  );
  AND2_X1 _10477_ (
    .A1(_00685_),
    .A2(_04985_),
    .ZN(_05078_)
  );
  INV_X1 _10478_ (
    .A(_05078_),
    .ZN(_05079_)
  );
  AND2_X1 _10479_ (
    .A1(_00811_),
    .A2(_05079_),
    .ZN(_05080_)
  );
  AND2_X1 _10480_ (
    .A1(_05077_),
    .A2(_05080_),
    .ZN(_00485_)
  );
  AND2_X1 _10481_ (
    .A1(_01276_),
    .A2(_04984_),
    .ZN(_05081_)
  );
  INV_X1 _10482_ (
    .A(_05081_),
    .ZN(_05082_)
  );
  AND2_X1 _10483_ (
    .A1(_00684_),
    .A2(_04985_),
    .ZN(_05083_)
  );
  INV_X1 _10484_ (
    .A(_05083_),
    .ZN(_05084_)
  );
  AND2_X1 _10485_ (
    .A1(_00811_),
    .A2(_05084_),
    .ZN(_05085_)
  );
  AND2_X1 _10486_ (
    .A1(_05082_),
    .A2(_05085_),
    .ZN(_00486_)
  );
  AND2_X1 _10487_ (
    .A1(_02734_),
    .A2(_04984_),
    .ZN(_05086_)
  );
  INV_X1 _10488_ (
    .A(_05086_),
    .ZN(_05087_)
  );
  AND2_X1 _10489_ (
    .A1(_00683_),
    .A2(_04985_),
    .ZN(_05088_)
  );
  INV_X1 _10490_ (
    .A(_05088_),
    .ZN(_05089_)
  );
  AND2_X1 _10491_ (
    .A1(_00811_),
    .A2(_05089_),
    .ZN(_05090_)
  );
  AND2_X1 _10492_ (
    .A1(_05087_),
    .A2(_05090_),
    .ZN(_00487_)
  );
  AND2_X1 _10493_ (
    .A1(_02800_),
    .A2(_04984_),
    .ZN(_05091_)
  );
  INV_X1 _10494_ (
    .A(_05091_),
    .ZN(_05092_)
  );
  AND2_X1 _10495_ (
    .A1(_00682_),
    .A2(_04985_),
    .ZN(_05093_)
  );
  INV_X1 _10496_ (
    .A(_05093_),
    .ZN(_05094_)
  );
  AND2_X1 _10497_ (
    .A1(_00811_),
    .A2(_05094_),
    .ZN(_05095_)
  );
  AND2_X1 _10498_ (
    .A1(_05092_),
    .A2(_05095_),
    .ZN(_00488_)
  );
  AND2_X1 _10499_ (
    .A1(_01359_),
    .A2(_04984_),
    .ZN(_05096_)
  );
  INV_X1 _10500_ (
    .A(_05096_),
    .ZN(_05097_)
  );
  AND2_X1 _10501_ (
    .A1(_00681_),
    .A2(_04985_),
    .ZN(_05098_)
  );
  INV_X1 _10502_ (
    .A(_05098_),
    .ZN(_05099_)
  );
  AND2_X1 _10503_ (
    .A1(_00811_),
    .A2(_05099_),
    .ZN(_05100_)
  );
  AND2_X1 _10504_ (
    .A1(_05097_),
    .A2(_05100_),
    .ZN(_00489_)
  );
  AND2_X1 _10505_ (
    .A1(_02872_),
    .A2(_04984_),
    .ZN(_05101_)
  );
  INV_X1 _10506_ (
    .A(_05101_),
    .ZN(_05102_)
  );
  AND2_X1 _10507_ (
    .A1(_00680_),
    .A2(_04985_),
    .ZN(_05103_)
  );
  INV_X1 _10508_ (
    .A(_05103_),
    .ZN(_05104_)
  );
  AND2_X1 _10509_ (
    .A1(_00811_),
    .A2(_05104_),
    .ZN(_05105_)
  );
  AND2_X1 _10510_ (
    .A1(_05102_),
    .A2(_05105_),
    .ZN(_00490_)
  );
  AND2_X1 _10511_ (
    .A1(_02944_),
    .A2(_04984_),
    .ZN(_05106_)
  );
  INV_X1 _10512_ (
    .A(_05106_),
    .ZN(_05107_)
  );
  AND2_X1 _10513_ (
    .A1(_00679_),
    .A2(_04985_),
    .ZN(_05108_)
  );
  INV_X1 _10514_ (
    .A(_05108_),
    .ZN(_05109_)
  );
  AND2_X1 _10515_ (
    .A1(_00811_),
    .A2(_05109_),
    .ZN(_05110_)
  );
  AND2_X1 _10516_ (
    .A1(_05107_),
    .A2(_05110_),
    .ZN(_00491_)
  );
  AND2_X1 _10517_ (
    .A1(_03016_),
    .A2(_04984_),
    .ZN(_05111_)
  );
  INV_X1 _10518_ (
    .A(_05111_),
    .ZN(_05112_)
  );
  AND2_X1 _10519_ (
    .A1(_00678_),
    .A2(_04985_),
    .ZN(_05113_)
  );
  INV_X1 _10520_ (
    .A(_05113_),
    .ZN(_05114_)
  );
  AND2_X1 _10521_ (
    .A1(_00811_),
    .A2(_05114_),
    .ZN(_05115_)
  );
  AND2_X1 _10522_ (
    .A1(_05112_),
    .A2(_05115_),
    .ZN(_00492_)
  );
  AND2_X1 _10523_ (
    .A1(_03090_),
    .A2(_04984_),
    .ZN(_05116_)
  );
  INV_X1 _10524_ (
    .A(_05116_),
    .ZN(_05117_)
  );
  AND2_X1 _10525_ (
    .A1(_00677_),
    .A2(_04985_),
    .ZN(_05118_)
  );
  INV_X1 _10526_ (
    .A(_05118_),
    .ZN(_05119_)
  );
  AND2_X1 _10527_ (
    .A1(_00811_),
    .A2(_05119_),
    .ZN(_05120_)
  );
  AND2_X1 _10528_ (
    .A1(_05117_),
    .A2(_05120_),
    .ZN(_00493_)
  );
  AND2_X1 _10529_ (
    .A1(_03161_),
    .A2(_04984_),
    .ZN(_05121_)
  );
  INV_X1 _10530_ (
    .A(_05121_),
    .ZN(_05122_)
  );
  AND2_X1 _10531_ (
    .A1(_00676_),
    .A2(_04985_),
    .ZN(_05123_)
  );
  INV_X1 _10532_ (
    .A(_05123_),
    .ZN(_05124_)
  );
  AND2_X1 _10533_ (
    .A1(_00811_),
    .A2(_05124_),
    .ZN(_05125_)
  );
  AND2_X1 _10534_ (
    .A1(_05122_),
    .A2(_05125_),
    .ZN(_00494_)
  );
  AND2_X1 _10535_ (
    .A1(_03229_),
    .A2(_04984_),
    .ZN(_05126_)
  );
  INV_X1 _10536_ (
    .A(_05126_),
    .ZN(_05127_)
  );
  AND2_X1 _10537_ (
    .A1(_00675_),
    .A2(_04985_),
    .ZN(_05128_)
  );
  INV_X1 _10538_ (
    .A(_05128_),
    .ZN(_05129_)
  );
  AND2_X1 _10539_ (
    .A1(_00811_),
    .A2(_05129_),
    .ZN(_05130_)
  );
  AND2_X1 _10540_ (
    .A1(_05127_),
    .A2(_05130_),
    .ZN(_00495_)
  );
  AND2_X1 _10541_ (
    .A1(_03442_),
    .A2(_04984_),
    .ZN(_05131_)
  );
  INV_X1 _10542_ (
    .A(_05131_),
    .ZN(_05132_)
  );
  AND2_X1 _10543_ (
    .A1(_00674_),
    .A2(_04985_),
    .ZN(_05133_)
  );
  INV_X1 _10544_ (
    .A(_05133_),
    .ZN(_05134_)
  );
  AND2_X1 _10545_ (
    .A1(_00811_),
    .A2(_05134_),
    .ZN(_05135_)
  );
  AND2_X1 _10546_ (
    .A1(_05132_),
    .A2(_05135_),
    .ZN(_00496_)
  );
  AND2_X1 _10547_ (
    .A1(_03341_),
    .A2(_04984_),
    .ZN(_05136_)
  );
  INV_X1 _10548_ (
    .A(_05136_),
    .ZN(_05137_)
  );
  AND2_X1 _10549_ (
    .A1(_00673_),
    .A2(_04985_),
    .ZN(_05138_)
  );
  INV_X1 _10550_ (
    .A(_05138_),
    .ZN(_05139_)
  );
  AND2_X1 _10551_ (
    .A1(_00811_),
    .A2(_05139_),
    .ZN(_05140_)
  );
  AND2_X1 _10552_ (
    .A1(_05137_),
    .A2(_05140_),
    .ZN(_00497_)
  );
  AND2_X1 _10553_ (
    .A1(_00897_),
    .A2(_01001_),
    .ZN(_05141_)
  );
  INV_X1 _10554_ (
    .A(_05141_),
    .ZN(_05142_)
  );
  MUX2_X1 _10555_ (
    .A(reg_mcause[0]),
    .B(_03517_),
    .S(_03535_),
    .Z(_05143_)
  );
  MUX2_X1 _10556_ (
    .A(_01613_),
    .B(_05143_),
    .S(_05142_),
    .Z(_05144_)
  );
  AND2_X1 _10557_ (
    .A1(_00811_),
    .A2(_05144_),
    .ZN(_00498_)
  );
  AND2_X1 _10558_ (
    .A1(_00868_),
    .A2(_03486_),
    .ZN(_05145_)
  );
  MUX2_X1 _10559_ (
    .A(_00871_),
    .B(_05145_),
    .S(_03535_),
    .Z(_05146_)
  );
  AND2_X1 _10560_ (
    .A1(_05142_),
    .A2(_05146_),
    .ZN(_05147_)
  );
  INV_X1 _10561_ (
    .A(_05147_),
    .ZN(_05148_)
  );
  AND2_X1 _10562_ (
    .A1(_01687_),
    .A2(_05141_),
    .ZN(_05149_)
  );
  INV_X1 _10563_ (
    .A(_05149_),
    .ZN(_05150_)
  );
  AND2_X1 _10564_ (
    .A1(_00811_),
    .A2(_05150_),
    .ZN(_05151_)
  );
  AND2_X1 _10565_ (
    .A1(_05148_),
    .A2(_05151_),
    .ZN(_00499_)
  );
  MUX2_X1 _10566_ (
    .A(reg_mcause[2]),
    .B(_03518_),
    .S(_03535_),
    .Z(_05152_)
  );
  INV_X1 _10567_ (
    .A(_05152_),
    .ZN(_05153_)
  );
  AND2_X1 _10568_ (
    .A1(_05142_),
    .A2(_05153_),
    .ZN(_05154_)
  );
  INV_X1 _10569_ (
    .A(_05154_),
    .ZN(_05155_)
  );
  AND2_X1 _10570_ (
    .A1(_01773_),
    .A2(_05141_),
    .ZN(_05156_)
  );
  INV_X1 _10571_ (
    .A(_05156_),
    .ZN(_05157_)
  );
  AND2_X1 _10572_ (
    .A1(_00811_),
    .A2(_05157_),
    .ZN(_05158_)
  );
  AND2_X1 _10573_ (
    .A1(_05155_),
    .A2(_05158_),
    .ZN(_00500_)
  );
  MUX2_X1 _10574_ (
    .A(_00872_),
    .B(_03524_),
    .S(_03535_),
    .Z(_05159_)
  );
  AND2_X1 _10575_ (
    .A1(_05142_),
    .A2(_05159_),
    .ZN(_05160_)
  );
  INV_X1 _10576_ (
    .A(_05160_),
    .ZN(_05161_)
  );
  AND2_X1 _10577_ (
    .A1(_01864_),
    .A2(_05141_),
    .ZN(_05162_)
  );
  INV_X1 _10578_ (
    .A(_05162_),
    .ZN(_05163_)
  );
  AND2_X1 _10579_ (
    .A1(_00811_),
    .A2(_05163_),
    .ZN(_05164_)
  );
  AND2_X1 _10580_ (
    .A1(_05161_),
    .A2(_05164_),
    .ZN(_00501_)
  );
  AND2_X1 _10581_ (
    .A1(_00811_),
    .A2(_05142_),
    .ZN(_05165_)
  );
  AND2_X1 _10582_ (
    .A1(io_cause[4]),
    .A2(_03486_),
    .ZN(_05166_)
  );
  MUX2_X1 _10583_ (
    .A(reg_mcause[4]),
    .B(_05166_),
    .S(_03535_),
    .Z(_05167_)
  );
  AND2_X1 _10584_ (
    .A1(_05165_),
    .A2(_05167_),
    .ZN(_00502_)
  );
  MUX2_X1 _10585_ (
    .A(reg_mcause[5]),
    .B(_03508_),
    .S(_03535_),
    .Z(_05168_)
  );
  AND2_X1 _10586_ (
    .A1(_05165_),
    .A2(_05168_),
    .ZN(_00503_)
  );
  MUX2_X1 _10587_ (
    .A(reg_mcause[6]),
    .B(_03512_),
    .S(_03535_),
    .Z(_05169_)
  );
  AND2_X1 _10588_ (
    .A1(_05165_),
    .A2(_05169_),
    .ZN(_00504_)
  );
  MUX2_X1 _10589_ (
    .A(reg_mcause[7]),
    .B(_03510_),
    .S(_03535_),
    .Z(_05170_)
  );
  AND2_X1 _10590_ (
    .A1(_05165_),
    .A2(_05170_),
    .ZN(_00505_)
  );
  AND2_X1 _10591_ (
    .A1(io_cause[8]),
    .A2(_03486_),
    .ZN(_05171_)
  );
  MUX2_X1 _10592_ (
    .A(reg_mcause[8]),
    .B(_05171_),
    .S(_03535_),
    .Z(_05172_)
  );
  AND2_X1 _10593_ (
    .A1(_05165_),
    .A2(_05172_),
    .ZN(_00506_)
  );
  AND2_X1 _10594_ (
    .A1(io_cause[9]),
    .A2(_03486_),
    .ZN(_05173_)
  );
  MUX2_X1 _10595_ (
    .A(reg_mcause[9]),
    .B(_05173_),
    .S(_03535_),
    .Z(_05174_)
  );
  AND2_X1 _10596_ (
    .A1(_05165_),
    .A2(_05174_),
    .ZN(_00507_)
  );
  AND2_X1 _10597_ (
    .A1(io_cause[10]),
    .A2(_03486_),
    .ZN(_05175_)
  );
  MUX2_X1 _10598_ (
    .A(reg_mcause[10]),
    .B(_05175_),
    .S(_03535_),
    .Z(_05176_)
  );
  AND2_X1 _10599_ (
    .A1(_05165_),
    .A2(_05176_),
    .ZN(_00508_)
  );
  AND2_X1 _10600_ (
    .A1(io_cause[11]),
    .A2(_03486_),
    .ZN(_05177_)
  );
  MUX2_X1 _10601_ (
    .A(reg_mcause[11]),
    .B(_05177_),
    .S(_03535_),
    .Z(_05178_)
  );
  AND2_X1 _10602_ (
    .A1(_05165_),
    .A2(_05178_),
    .ZN(_00509_)
  );
  AND2_X1 _10603_ (
    .A1(io_cause[12]),
    .A2(_03486_),
    .ZN(_05179_)
  );
  MUX2_X1 _10604_ (
    .A(reg_mcause[12]),
    .B(_05179_),
    .S(_03535_),
    .Z(_05180_)
  );
  AND2_X1 _10605_ (
    .A1(_05165_),
    .A2(_05180_),
    .ZN(_00510_)
  );
  AND2_X1 _10606_ (
    .A1(io_cause[13]),
    .A2(_03486_),
    .ZN(_05181_)
  );
  MUX2_X1 _10607_ (
    .A(reg_mcause[13]),
    .B(_05181_),
    .S(_03535_),
    .Z(_05182_)
  );
  AND2_X1 _10608_ (
    .A1(_05165_),
    .A2(_05182_),
    .ZN(_00511_)
  );
  AND2_X1 _10609_ (
    .A1(io_cause[14]),
    .A2(_03486_),
    .ZN(_05183_)
  );
  MUX2_X1 _10610_ (
    .A(reg_mcause[14]),
    .B(_05183_),
    .S(_03535_),
    .Z(_05184_)
  );
  AND2_X1 _10611_ (
    .A1(_05165_),
    .A2(_05184_),
    .ZN(_00512_)
  );
  AND2_X1 _10612_ (
    .A1(io_cause[15]),
    .A2(_03486_),
    .ZN(_05185_)
  );
  MUX2_X1 _10613_ (
    .A(reg_mcause[15]),
    .B(_05185_),
    .S(_03535_),
    .Z(_05186_)
  );
  AND2_X1 _10614_ (
    .A1(_05165_),
    .A2(_05186_),
    .ZN(_00513_)
  );
  AND2_X1 _10615_ (
    .A1(io_cause[16]),
    .A2(_03486_),
    .ZN(_05187_)
  );
  MUX2_X1 _10616_ (
    .A(reg_mcause[16]),
    .B(_05187_),
    .S(_03535_),
    .Z(_05188_)
  );
  AND2_X1 _10617_ (
    .A1(_05165_),
    .A2(_05188_),
    .ZN(_00514_)
  );
  AND2_X1 _10618_ (
    .A1(io_cause[17]),
    .A2(_03486_),
    .ZN(_05189_)
  );
  MUX2_X1 _10619_ (
    .A(reg_mcause[17]),
    .B(_05189_),
    .S(_03535_),
    .Z(_05190_)
  );
  AND2_X1 _10620_ (
    .A1(_05165_),
    .A2(_05190_),
    .ZN(_00515_)
  );
  AND2_X1 _10621_ (
    .A1(io_cause[18]),
    .A2(_03486_),
    .ZN(_05191_)
  );
  MUX2_X1 _10622_ (
    .A(reg_mcause[18]),
    .B(_05191_),
    .S(_03535_),
    .Z(_05192_)
  );
  AND2_X1 _10623_ (
    .A1(_05165_),
    .A2(_05192_),
    .ZN(_00516_)
  );
  AND2_X1 _10624_ (
    .A1(io_cause[19]),
    .A2(_03486_),
    .ZN(_05193_)
  );
  MUX2_X1 _10625_ (
    .A(reg_mcause[19]),
    .B(_05193_),
    .S(_03535_),
    .Z(_05194_)
  );
  AND2_X1 _10626_ (
    .A1(_05165_),
    .A2(_05194_),
    .ZN(_00517_)
  );
  AND2_X1 _10627_ (
    .A1(io_cause[20]),
    .A2(_03486_),
    .ZN(_05195_)
  );
  MUX2_X1 _10628_ (
    .A(reg_mcause[20]),
    .B(_05195_),
    .S(_03535_),
    .Z(_05196_)
  );
  AND2_X1 _10629_ (
    .A1(_05165_),
    .A2(_05196_),
    .ZN(_00518_)
  );
  AND2_X1 _10630_ (
    .A1(io_cause[21]),
    .A2(_03486_),
    .ZN(_05197_)
  );
  MUX2_X1 _10631_ (
    .A(reg_mcause[21]),
    .B(_05197_),
    .S(_03535_),
    .Z(_05198_)
  );
  AND2_X1 _10632_ (
    .A1(_05165_),
    .A2(_05198_),
    .ZN(_00519_)
  );
  AND2_X1 _10633_ (
    .A1(io_cause[22]),
    .A2(_03486_),
    .ZN(_05199_)
  );
  MUX2_X1 _10634_ (
    .A(reg_mcause[22]),
    .B(_05199_),
    .S(_03535_),
    .Z(_05200_)
  );
  AND2_X1 _10635_ (
    .A1(_05165_),
    .A2(_05200_),
    .ZN(_00520_)
  );
  AND2_X1 _10636_ (
    .A1(io_cause[23]),
    .A2(_03486_),
    .ZN(_05201_)
  );
  MUX2_X1 _10637_ (
    .A(reg_mcause[23]),
    .B(_05201_),
    .S(_03535_),
    .Z(_05202_)
  );
  AND2_X1 _10638_ (
    .A1(_05165_),
    .A2(_05202_),
    .ZN(_00521_)
  );
  AND2_X1 _10639_ (
    .A1(io_cause[24]),
    .A2(_03486_),
    .ZN(_05203_)
  );
  MUX2_X1 _10640_ (
    .A(reg_mcause[24]),
    .B(_05203_),
    .S(_03535_),
    .Z(_05204_)
  );
  AND2_X1 _10641_ (
    .A1(_05165_),
    .A2(_05204_),
    .ZN(_00522_)
  );
  AND2_X1 _10642_ (
    .A1(io_cause[25]),
    .A2(_03486_),
    .ZN(_05205_)
  );
  MUX2_X1 _10643_ (
    .A(reg_mcause[25]),
    .B(_05205_),
    .S(_03535_),
    .Z(_05206_)
  );
  AND2_X1 _10644_ (
    .A1(_05165_),
    .A2(_05206_),
    .ZN(_00523_)
  );
  AND2_X1 _10645_ (
    .A1(io_cause[26]),
    .A2(_03486_),
    .ZN(_05207_)
  );
  MUX2_X1 _10646_ (
    .A(reg_mcause[26]),
    .B(_05207_),
    .S(_03535_),
    .Z(_05208_)
  );
  AND2_X1 _10647_ (
    .A1(_05165_),
    .A2(_05208_),
    .ZN(_00524_)
  );
  AND2_X1 _10648_ (
    .A1(io_cause[27]),
    .A2(_03486_),
    .ZN(_05209_)
  );
  MUX2_X1 _10649_ (
    .A(reg_mcause[27]),
    .B(_05209_),
    .S(_03535_),
    .Z(_05210_)
  );
  AND2_X1 _10650_ (
    .A1(_05165_),
    .A2(_05210_),
    .ZN(_00525_)
  );
  AND2_X1 _10651_ (
    .A1(io_cause[28]),
    .A2(_03486_),
    .ZN(_05211_)
  );
  MUX2_X1 _10652_ (
    .A(reg_mcause[28]),
    .B(_05211_),
    .S(_03535_),
    .Z(_05212_)
  );
  AND2_X1 _10653_ (
    .A1(_05165_),
    .A2(_05212_),
    .ZN(_00526_)
  );
  AND2_X1 _10654_ (
    .A1(io_cause[29]),
    .A2(_03486_),
    .ZN(_05213_)
  );
  MUX2_X1 _10655_ (
    .A(reg_mcause[29]),
    .B(_05213_),
    .S(_03535_),
    .Z(_05214_)
  );
  AND2_X1 _10656_ (
    .A1(_05165_),
    .A2(_05214_),
    .ZN(_00527_)
  );
  AND2_X1 _10657_ (
    .A1(io_cause[30]),
    .A2(_03486_),
    .ZN(_05215_)
  );
  MUX2_X1 _10658_ (
    .A(reg_mcause[30]),
    .B(_05215_),
    .S(_03535_),
    .Z(_05216_)
  );
  AND2_X1 _10659_ (
    .A1(_05165_),
    .A2(_05216_),
    .ZN(_00528_)
  );
  MUX2_X1 _10660_ (
    .A(reg_mcause[31]),
    .B(_03577_),
    .S(_03535_),
    .Z(_05217_)
  );
  INV_X1 _10661_ (
    .A(_05217_),
    .ZN(_05218_)
  );
  AND2_X1 _10662_ (
    .A1(_05142_),
    .A2(_05218_),
    .ZN(_05219_)
  );
  INV_X1 _10663_ (
    .A(_05219_),
    .ZN(_05220_)
  );
  AND2_X1 _10664_ (
    .A1(_03341_),
    .A2(_05141_),
    .ZN(_05221_)
  );
  INV_X1 _10665_ (
    .A(_05221_),
    .ZN(_05222_)
  );
  AND2_X1 _10666_ (
    .A1(_00811_),
    .A2(_05222_),
    .ZN(_05223_)
  );
  AND2_X1 _10667_ (
    .A1(_05220_),
    .A2(_05223_),
    .ZN(_00529_)
  );
  AND2_X1 _10668_ (
    .A1(_00897_),
    .A2(_01782_),
    .ZN(_05224_)
  );
  MUX2_X1 _10669_ (
    .A(reg_mie[3]),
    .B(_01865_),
    .S(_05224_),
    .Z(_00530_)
  );
  MUX2_X1 _10670_ (
    .A(reg_mie[7]),
    .B(_02163_),
    .S(_05224_),
    .Z(_00531_)
  );
  MUX2_X1 _10671_ (
    .A(reg_mie[11]),
    .B(_02314_),
    .S(_05224_),
    .Z(_00532_)
  );
  AND2_X1 _10672_ (
    .A1(_00003_),
    .A2(_00894_),
    .ZN(_05225_)
  );
  AND2_X1 _10673_ (
    .A1(_00897_),
    .A2(_05225_),
    .ZN(_05226_)
  );
  INV_X1 _10674_ (
    .A(_05226_),
    .ZN(_05227_)
  );
  MUX2_X1 _10675_ (
    .A(reg_pmp_7_cfg_r),
    .B(_02873_),
    .S(_05226_),
    .Z(_00533_)
  );
  MUX2_X1 _10676_ (
    .A(reg_pmp_7_cfg_w),
    .B(_03277_),
    .S(_05226_),
    .Z(_00534_)
  );
  MUX2_X1 _10677_ (
    .A(reg_pmp_7_cfg_x),
    .B(_03017_),
    .S(_05226_),
    .Z(_00535_)
  );
  AND2_X1 _10678_ (
    .A1(_00897_),
    .A2(_01016_),
    .ZN(_05228_)
  );
  AND2_X1 _10679_ (
    .A1(_00670_),
    .A2(_05228_),
    .ZN(_05229_)
  );
  MUX2_X1 _10680_ (
    .A(reg_pmp_7_addr[0]),
    .B(_01613_),
    .S(_05229_),
    .Z(_00536_)
  );
  MUX2_X1 _10681_ (
    .A(reg_pmp_7_addr[1]),
    .B(_01688_),
    .S(_05229_),
    .Z(_00537_)
  );
  MUX2_X1 _10682_ (
    .A(reg_pmp_7_addr[2]),
    .B(_01774_),
    .S(_05229_),
    .Z(_00538_)
  );
  MUX2_X1 _10683_ (
    .A(reg_pmp_7_addr[3]),
    .B(_01865_),
    .S(_05229_),
    .Z(_00539_)
  );
  MUX2_X1 _10684_ (
    .A(reg_pmp_7_addr[4]),
    .B(_01938_),
    .S(_05229_),
    .Z(_00540_)
  );
  MUX2_X1 _10685_ (
    .A(reg_pmp_7_addr[5]),
    .B(_02005_),
    .S(_05229_),
    .Z(_00541_)
  );
  MUX2_X1 _10686_ (
    .A(reg_pmp_7_addr[6]),
    .B(_02076_),
    .S(_05229_),
    .Z(_00542_)
  );
  MUX2_X1 _10687_ (
    .A(reg_pmp_7_addr[7]),
    .B(_02163_),
    .S(_05229_),
    .Z(_00543_)
  );
  MUX2_X1 _10688_ (
    .A(reg_pmp_7_addr[8]),
    .B(_01446_),
    .S(_05229_),
    .Z(_00544_)
  );
  MUX2_X1 _10689_ (
    .A(reg_pmp_7_addr[9]),
    .B(_01518_),
    .S(_05229_),
    .Z(_00545_)
  );
  MUX2_X1 _10690_ (
    .A(reg_pmp_7_addr[10]),
    .B(_02235_),
    .S(_05229_),
    .Z(_00546_)
  );
  MUX2_X1 _10691_ (
    .A(reg_pmp_7_addr[11]),
    .B(_02314_),
    .S(_05229_),
    .Z(_00547_)
  );
  MUX2_X1 _10692_ (
    .A(reg_pmp_7_addr[12]),
    .B(_02389_),
    .S(_05229_),
    .Z(_00548_)
  );
  MUX2_X1 _10693_ (
    .A(reg_pmp_7_addr[13]),
    .B(_02456_),
    .S(_05229_),
    .Z(_00549_)
  );
  MUX2_X1 _10694_ (
    .A(reg_pmp_7_addr[14]),
    .B(_02522_),
    .S(_05229_),
    .Z(_00550_)
  );
  MUX2_X1 _10695_ (
    .A(reg_pmp_7_addr[15]),
    .B(_02597_),
    .S(_05229_),
    .Z(_00551_)
  );
  MUX2_X1 _10696_ (
    .A(reg_pmp_7_addr[16]),
    .B(_01035_),
    .S(_05229_),
    .Z(_00552_)
  );
  MUX2_X1 _10697_ (
    .A(reg_pmp_7_addr[17]),
    .B(_02669_),
    .S(_05229_),
    .Z(_00553_)
  );
  MUX2_X1 _10698_ (
    .A(reg_pmp_7_addr[18]),
    .B(_01107_),
    .S(_05229_),
    .Z(_00554_)
  );
  MUX2_X1 _10699_ (
    .A(reg_pmp_7_addr[19]),
    .B(_01199_),
    .S(_05229_),
    .Z(_00555_)
  );
  MUX2_X1 _10700_ (
    .A(reg_pmp_7_addr[20]),
    .B(_01277_),
    .S(_05229_),
    .Z(_00556_)
  );
  MUX2_X1 _10701_ (
    .A(reg_pmp_7_addr[21]),
    .B(_02735_),
    .S(_05229_),
    .Z(_00557_)
  );
  MUX2_X1 _10702_ (
    .A(reg_pmp_7_addr[22]),
    .B(_02801_),
    .S(_05229_),
    .Z(_00558_)
  );
  MUX2_X1 _10703_ (
    .A(reg_pmp_7_addr[23]),
    .B(_01360_),
    .S(_05229_),
    .Z(_00559_)
  );
  MUX2_X1 _10704_ (
    .A(reg_pmp_7_addr[24]),
    .B(_02873_),
    .S(_05229_),
    .Z(_00560_)
  );
  MUX2_X1 _10705_ (
    .A(reg_pmp_7_addr[25]),
    .B(_02945_),
    .S(_05229_),
    .Z(_00561_)
  );
  MUX2_X1 _10706_ (
    .A(reg_pmp_7_addr[26]),
    .B(_03017_),
    .S(_05229_),
    .Z(_00562_)
  );
  MUX2_X1 _10707_ (
    .A(reg_pmp_7_addr[27]),
    .B(_03089_),
    .S(_05229_),
    .Z(_00563_)
  );
  MUX2_X1 _10708_ (
    .A(reg_pmp_7_addr[28]),
    .B(_03162_),
    .S(_05229_),
    .Z(_00564_)
  );
  MUX2_X1 _10709_ (
    .A(reg_pmp_7_addr[29]),
    .B(_03230_),
    .S(_05229_),
    .Z(_00565_)
  );
  AND2_X1 _10710_ (
    .A1(_00672_),
    .A2(_05227_),
    .ZN(_05230_)
  );
  INV_X1 _10711_ (
    .A(_05230_),
    .ZN(_05231_)
  );
  AND2_X1 _10712_ (
    .A1(_00811_),
    .A2(_05231_),
    .ZN(_05232_)
  );
  AND2_X1 _10713_ (
    .A1(_03090_),
    .A2(_05226_),
    .ZN(_05233_)
  );
  INV_X1 _10714_ (
    .A(_05233_),
    .ZN(_05234_)
  );
  AND2_X1 _10715_ (
    .A1(_05232_),
    .A2(_05234_),
    .ZN(_00566_)
  );
  AND2_X1 _10716_ (
    .A1(_00671_),
    .A2(_05227_),
    .ZN(_05235_)
  );
  INV_X1 _10717_ (
    .A(_05235_),
    .ZN(_05236_)
  );
  AND2_X1 _10718_ (
    .A1(_00811_),
    .A2(_05236_),
    .ZN(_05237_)
  );
  AND2_X1 _10719_ (
    .A1(_03161_),
    .A2(_05226_),
    .ZN(_05238_)
  );
  INV_X1 _10720_ (
    .A(_05238_),
    .ZN(_05239_)
  );
  AND2_X1 _10721_ (
    .A1(_05237_),
    .A2(_05239_),
    .ZN(_00567_)
  );
  AND2_X1 _10722_ (
    .A1(_00670_),
    .A2(_05227_),
    .ZN(_05240_)
  );
  INV_X1 _10723_ (
    .A(_05240_),
    .ZN(_05241_)
  );
  AND2_X1 _10724_ (
    .A1(_00811_),
    .A2(_05241_),
    .ZN(_05242_)
  );
  AND2_X1 _10725_ (
    .A1(_03341_),
    .A2(_05226_),
    .ZN(_05243_)
  );
  INV_X1 _10726_ (
    .A(_05243_),
    .ZN(_05244_)
  );
  AND2_X1 _10727_ (
    .A1(_05242_),
    .A2(_05244_),
    .ZN(_00568_)
  );
  AND2_X1 _10728_ (
    .A1(large_1[0]),
    .A2(_03700_),
    .ZN(_05245_)
  );
  INV_X1 _10729_ (
    .A(_05245_),
    .ZN(_05246_)
  );
  MUX2_X1 _10730_ (
    .A(large_1[0]),
    .B(_large_r_T_3[0]),
    .S(_03666_),
    .Z(_05247_)
  );
  AND2_X1 _10731_ (
    .A1(_03710_),
    .A2(_05247_),
    .ZN(_05248_)
  );
  INV_X1 _10732_ (
    .A(_05248_),
    .ZN(_05249_)
  );
  AND2_X1 _10733_ (
    .A1(_05246_),
    .A2(_05249_),
    .ZN(_05250_)
  );
  AND2_X1 _10734_ (
    .A1(_02076_),
    .A2(_03702_),
    .ZN(_05251_)
  );
  INV_X1 _10735_ (
    .A(_05251_),
    .ZN(_05252_)
  );
  AND2_X1 _10736_ (
    .A1(_05250_),
    .A2(_05252_),
    .ZN(_05253_)
  );
  INV_X1 _10737_ (
    .A(_05253_),
    .ZN(_05254_)
  );
  AND2_X1 _10738_ (
    .A1(_00811_),
    .A2(_05254_),
    .ZN(_00569_)
  );
  AND2_X1 _10739_ (
    .A1(_00669_),
    .A2(_03662_),
    .ZN(_05255_)
  );
  INV_X1 _10740_ (
    .A(_05255_),
    .ZN(_05256_)
  );
  AND2_X1 _10741_ (
    .A1(large_1[1]),
    .A2(_03700_),
    .ZN(_05257_)
  );
  INV_X1 _10742_ (
    .A(_05257_),
    .ZN(_05258_)
  );
  AND2_X1 _10743_ (
    .A1(_03710_),
    .A2(_05256_),
    .ZN(_05259_)
  );
  AND2_X1 _10744_ (
    .A1(_03666_),
    .A2(_03683_),
    .ZN(_05260_)
  );
  AND2_X1 _10745_ (
    .A1(_03669_),
    .A2(_05259_),
    .ZN(_05261_)
  );
  INV_X1 _10746_ (
    .A(_05261_),
    .ZN(_05262_)
  );
  AND2_X1 _10747_ (
    .A1(_05258_),
    .A2(_05262_),
    .ZN(_05263_)
  );
  AND2_X1 _10748_ (
    .A1(_02163_),
    .A2(_03702_),
    .ZN(_05264_)
  );
  INV_X1 _10749_ (
    .A(_05264_),
    .ZN(_05265_)
  );
  AND2_X1 _10750_ (
    .A1(_05263_),
    .A2(_05265_),
    .ZN(_05266_)
  );
  INV_X1 _10751_ (
    .A(_05266_),
    .ZN(_05267_)
  );
  AND2_X1 _10752_ (
    .A1(_00811_),
    .A2(_05267_),
    .ZN(_00570_)
  );
  AND2_X1 _10753_ (
    .A1(_00668_),
    .A2(_03669_),
    .ZN(_05268_)
  );
  INV_X1 _10754_ (
    .A(_05268_),
    .ZN(_05269_)
  );
  AND2_X1 _10755_ (
    .A1(large_1[2]),
    .A2(_03700_),
    .ZN(_05270_)
  );
  INV_X1 _10756_ (
    .A(_05270_),
    .ZN(_05271_)
  );
  AND2_X1 _10757_ (
    .A1(large_1[2]),
    .A2(_03663_),
    .ZN(_05272_)
  );
  AND2_X1 _10758_ (
    .A1(large_1[2]),
    .A2(_03668_),
    .ZN(_05273_)
  );
  INV_X1 _10759_ (
    .A(_05273_),
    .ZN(_05274_)
  );
  AND2_X1 _10760_ (
    .A1(_03710_),
    .A2(_05269_),
    .ZN(_05275_)
  );
  AND2_X1 _10761_ (
    .A1(_05274_),
    .A2(_05275_),
    .ZN(_05276_)
  );
  INV_X1 _10762_ (
    .A(_05276_),
    .ZN(_05277_)
  );
  AND2_X1 _10763_ (
    .A1(_01446_),
    .A2(_03708_),
    .ZN(_05278_)
  );
  INV_X1 _10764_ (
    .A(_05278_),
    .ZN(_05279_)
  );
  AND2_X1 _10765_ (
    .A1(_05277_),
    .A2(_05279_),
    .ZN(_05280_)
  );
  AND2_X1 _10766_ (
    .A1(_05271_),
    .A2(_05280_),
    .ZN(_05281_)
  );
  INV_X1 _10767_ (
    .A(_05281_),
    .ZN(_05282_)
  );
  AND2_X1 _10768_ (
    .A1(_00811_),
    .A2(_05282_),
    .ZN(_00571_)
  );
  AND2_X1 _10769_ (
    .A1(_00667_),
    .A2(_05274_),
    .ZN(_05283_)
  );
  INV_X1 _10770_ (
    .A(_05283_),
    .ZN(_05284_)
  );
  AND2_X1 _10771_ (
    .A1(large_1[3]),
    .A2(_03700_),
    .ZN(_05285_)
  );
  INV_X1 _10772_ (
    .A(_05285_),
    .ZN(_05286_)
  );
  AND2_X1 _10773_ (
    .A1(_03649_),
    .A2(_05260_),
    .ZN(_05287_)
  );
  INV_X1 _10774_ (
    .A(_05287_),
    .ZN(_05288_)
  );
  AND2_X1 _10775_ (
    .A1(_03710_),
    .A2(_05284_),
    .ZN(_05289_)
  );
  AND2_X1 _10776_ (
    .A1(_05288_),
    .A2(_05289_),
    .ZN(_05290_)
  );
  INV_X1 _10777_ (
    .A(_05290_),
    .ZN(_05291_)
  );
  AND2_X1 _10778_ (
    .A1(_01518_),
    .A2(_03708_),
    .ZN(_05292_)
  );
  INV_X1 _10779_ (
    .A(_05292_),
    .ZN(_05293_)
  );
  AND2_X1 _10780_ (
    .A1(_05286_),
    .A2(_05293_),
    .ZN(_05294_)
  );
  AND2_X1 _10781_ (
    .A1(_05291_),
    .A2(_05294_),
    .ZN(_05295_)
  );
  INV_X1 _10782_ (
    .A(_05295_),
    .ZN(_05296_)
  );
  AND2_X1 _10783_ (
    .A1(_00811_),
    .A2(_05296_),
    .ZN(_00572_)
  );
  AND2_X1 _10784_ (
    .A1(_00666_),
    .A2(_05288_),
    .ZN(_05297_)
  );
  INV_X1 _10785_ (
    .A(_05297_),
    .ZN(_05298_)
  );
  AND2_X1 _10786_ (
    .A1(_03648_),
    .A2(_05272_),
    .ZN(_05299_)
  );
  INV_X1 _10787_ (
    .A(_05299_),
    .ZN(_05300_)
  );
  AND2_X1 _10788_ (
    .A1(_03706_),
    .A2(_05300_),
    .ZN(_05301_)
  );
  AND2_X1 _10789_ (
    .A1(_05298_),
    .A2(_05301_),
    .ZN(_05302_)
  );
  INV_X1 _10790_ (
    .A(_05302_),
    .ZN(_05303_)
  );
  AND2_X1 _10791_ (
    .A1(large_1[4]),
    .A2(_03700_),
    .ZN(_05304_)
  );
  INV_X1 _10792_ (
    .A(_05304_),
    .ZN(_05305_)
  );
  AND2_X1 _10793_ (
    .A1(_05303_),
    .A2(_05305_),
    .ZN(_05306_)
  );
  AND2_X1 _10794_ (
    .A1(_02235_),
    .A2(_03702_),
    .ZN(_05307_)
  );
  INV_X1 _10795_ (
    .A(_05307_),
    .ZN(_05308_)
  );
  AND2_X1 _10796_ (
    .A1(_05306_),
    .A2(_05308_),
    .ZN(_05309_)
  );
  INV_X1 _10797_ (
    .A(_05309_),
    .ZN(_05310_)
  );
  AND2_X1 _10798_ (
    .A1(_00811_),
    .A2(_05310_),
    .ZN(_00573_)
  );
  AND2_X1 _10799_ (
    .A1(_00665_),
    .A2(_05300_),
    .ZN(_05311_)
  );
  INV_X1 _10800_ (
    .A(_05311_),
    .ZN(_05312_)
  );
  AND2_X1 _10801_ (
    .A1(large_1[5]),
    .A2(_03700_),
    .ZN(_05313_)
  );
  INV_X1 _10802_ (
    .A(_05313_),
    .ZN(_05314_)
  );
  AND2_X1 _10803_ (
    .A1(_03650_),
    .A2(_05287_),
    .ZN(_05315_)
  );
  INV_X1 _10804_ (
    .A(_05315_),
    .ZN(_05316_)
  );
  AND2_X1 _10805_ (
    .A1(_03710_),
    .A2(_05316_),
    .ZN(_05317_)
  );
  AND2_X1 _10806_ (
    .A1(_05312_),
    .A2(_05317_),
    .ZN(_05318_)
  );
  INV_X1 _10807_ (
    .A(_05318_),
    .ZN(_05319_)
  );
  AND2_X1 _10808_ (
    .A1(_02314_),
    .A2(_03708_),
    .ZN(_05320_)
  );
  INV_X1 _10809_ (
    .A(_05320_),
    .ZN(_05321_)
  );
  AND2_X1 _10810_ (
    .A1(_05314_),
    .A2(_05321_),
    .ZN(_05322_)
  );
  AND2_X1 _10811_ (
    .A1(_05319_),
    .A2(_05322_),
    .ZN(_05323_)
  );
  INV_X1 _10812_ (
    .A(_05323_),
    .ZN(_05324_)
  );
  AND2_X1 _10813_ (
    .A1(_00811_),
    .A2(_05324_),
    .ZN(_00574_)
  );
  AND2_X1 _10814_ (
    .A1(_00664_),
    .A2(_05316_),
    .ZN(_05325_)
  );
  INV_X1 _10815_ (
    .A(_05325_),
    .ZN(_05326_)
  );
  AND2_X1 _10816_ (
    .A1(large_1[6]),
    .A2(_03700_),
    .ZN(_05327_)
  );
  INV_X1 _10817_ (
    .A(_05327_),
    .ZN(_05328_)
  );
  AND2_X1 _10818_ (
    .A1(_03671_),
    .A2(_03710_),
    .ZN(_05329_)
  );
  AND2_X1 _10819_ (
    .A1(_05326_),
    .A2(_05329_),
    .ZN(_05330_)
  );
  INV_X1 _10820_ (
    .A(_05330_),
    .ZN(_05331_)
  );
  AND2_X1 _10821_ (
    .A1(_05328_),
    .A2(_05331_),
    .ZN(_05332_)
  );
  AND2_X1 _10822_ (
    .A1(_02389_),
    .A2(_03702_),
    .ZN(_05333_)
  );
  INV_X1 _10823_ (
    .A(_05333_),
    .ZN(_05334_)
  );
  AND2_X1 _10824_ (
    .A1(_05332_),
    .A2(_05334_),
    .ZN(_05335_)
  );
  INV_X1 _10825_ (
    .A(_05335_),
    .ZN(_05336_)
  );
  AND2_X1 _10826_ (
    .A1(_00811_),
    .A2(_05336_),
    .ZN(_00575_)
  );
  AND2_X1 _10827_ (
    .A1(_02456_),
    .A2(_03702_),
    .ZN(_05337_)
  );
  INV_X1 _10828_ (
    .A(_05337_),
    .ZN(_05338_)
  );
  AND2_X1 _10829_ (
    .A1(_00663_),
    .A2(_03671_),
    .ZN(_05339_)
  );
  INV_X1 _10830_ (
    .A(_05339_),
    .ZN(_05340_)
  );
  AND2_X1 _10831_ (
    .A1(_03710_),
    .A2(_05340_),
    .ZN(_05341_)
  );
  AND2_X1 _10832_ (
    .A1(large_1[7]),
    .A2(_03664_),
    .ZN(_05342_)
  );
  INV_X1 _10833_ (
    .A(_05342_),
    .ZN(_05343_)
  );
  AND2_X1 _10834_ (
    .A1(_05341_),
    .A2(_05343_),
    .ZN(_05344_)
  );
  INV_X1 _10835_ (
    .A(_05344_),
    .ZN(_05345_)
  );
  AND2_X1 _10836_ (
    .A1(large_1[7]),
    .A2(_03700_),
    .ZN(_05346_)
  );
  INV_X1 _10837_ (
    .A(_05346_),
    .ZN(_05347_)
  );
  AND2_X1 _10838_ (
    .A1(_05345_),
    .A2(_05347_),
    .ZN(_05348_)
  );
  AND2_X1 _10839_ (
    .A1(_05338_),
    .A2(_05348_),
    .ZN(_05349_)
  );
  INV_X1 _10840_ (
    .A(_05349_),
    .ZN(_05350_)
  );
  AND2_X1 _10841_ (
    .A1(_00811_),
    .A2(_05350_),
    .ZN(_00576_)
  );
  AND2_X1 _10842_ (
    .A1(_00662_),
    .A2(_05343_),
    .ZN(_05351_)
  );
  INV_X1 _10843_ (
    .A(_05351_),
    .ZN(_05352_)
  );
  AND2_X1 _10844_ (
    .A1(large_1[8]),
    .A2(_03700_),
    .ZN(_05353_)
  );
  INV_X1 _10845_ (
    .A(_05353_),
    .ZN(_05354_)
  );
  AND2_X1 _10846_ (
    .A1(_03646_),
    .A2(_03670_),
    .ZN(_05355_)
  );
  INV_X1 _10847_ (
    .A(_05355_),
    .ZN(_05356_)
  );
  AND2_X1 _10848_ (
    .A1(_03710_),
    .A2(_05356_),
    .ZN(_05357_)
  );
  AND2_X1 _10849_ (
    .A1(_05352_),
    .A2(_05357_),
    .ZN(_05358_)
  );
  INV_X1 _10850_ (
    .A(_05358_),
    .ZN(_05359_)
  );
  AND2_X1 _10851_ (
    .A1(_05354_),
    .A2(_05359_),
    .ZN(_05360_)
  );
  AND2_X1 _10852_ (
    .A1(_02522_),
    .A2(_03702_),
    .ZN(_05361_)
  );
  INV_X1 _10853_ (
    .A(_05361_),
    .ZN(_05362_)
  );
  AND2_X1 _10854_ (
    .A1(_05360_),
    .A2(_05362_),
    .ZN(_05363_)
  );
  INV_X1 _10855_ (
    .A(_05363_),
    .ZN(_05364_)
  );
  AND2_X1 _10856_ (
    .A1(_00811_),
    .A2(_05364_),
    .ZN(_00577_)
  );
  AND2_X1 _10857_ (
    .A1(_00661_),
    .A2(_05356_),
    .ZN(_05365_)
  );
  INV_X1 _10858_ (
    .A(_05365_),
    .ZN(_05366_)
  );
  AND2_X1 _10859_ (
    .A1(_03673_),
    .A2(_03710_),
    .ZN(_05367_)
  );
  AND2_X1 _10860_ (
    .A1(_05366_),
    .A2(_05367_),
    .ZN(_05368_)
  );
  INV_X1 _10861_ (
    .A(_05368_),
    .ZN(_05369_)
  );
  AND2_X1 _10862_ (
    .A1(large_1[9]),
    .A2(_03700_),
    .ZN(_05370_)
  );
  INV_X1 _10863_ (
    .A(_05370_),
    .ZN(_05371_)
  );
  AND2_X1 _10864_ (
    .A1(_02597_),
    .A2(_03708_),
    .ZN(_05372_)
  );
  INV_X1 _10865_ (
    .A(_05372_),
    .ZN(_05373_)
  );
  AND2_X1 _10866_ (
    .A1(_05369_),
    .A2(_05371_),
    .ZN(_05374_)
  );
  AND2_X1 _10867_ (
    .A1(_05373_),
    .A2(_05374_),
    .ZN(_05375_)
  );
  INV_X1 _10868_ (
    .A(_05375_),
    .ZN(_05376_)
  );
  AND2_X1 _10869_ (
    .A1(_00811_),
    .A2(_05376_),
    .ZN(_00578_)
  );
  AND2_X1 _10870_ (
    .A1(_00660_),
    .A2(_03673_),
    .ZN(_05377_)
  );
  INV_X1 _10871_ (
    .A(_05377_),
    .ZN(_05378_)
  );
  AND2_X1 _10872_ (
    .A1(large_1[10]),
    .A2(_03700_),
    .ZN(_05379_)
  );
  INV_X1 _10873_ (
    .A(_05379_),
    .ZN(_05380_)
  );
  AND2_X1 _10874_ (
    .A1(_03675_),
    .A2(_03710_),
    .ZN(_05381_)
  );
  AND2_X1 _10875_ (
    .A1(_05378_),
    .A2(_05381_),
    .ZN(_05382_)
  );
  INV_X1 _10876_ (
    .A(_05382_),
    .ZN(_05383_)
  );
  AND2_X1 _10877_ (
    .A1(_01035_),
    .A2(_03708_),
    .ZN(_05384_)
  );
  INV_X1 _10878_ (
    .A(_05384_),
    .ZN(_05385_)
  );
  AND2_X1 _10879_ (
    .A1(_05383_),
    .A2(_05385_),
    .ZN(_05386_)
  );
  AND2_X1 _10880_ (
    .A1(_05380_),
    .A2(_05386_),
    .ZN(_05387_)
  );
  INV_X1 _10881_ (
    .A(_05387_),
    .ZN(_05388_)
  );
  AND2_X1 _10882_ (
    .A1(_00811_),
    .A2(_05388_),
    .ZN(_00579_)
  );
  AND2_X1 _10883_ (
    .A1(_00659_),
    .A2(_03675_),
    .ZN(_05389_)
  );
  INV_X1 _10884_ (
    .A(_05389_),
    .ZN(_05390_)
  );
  AND2_X1 _10885_ (
    .A1(_03677_),
    .A2(_03710_),
    .ZN(_05391_)
  );
  AND2_X1 _10886_ (
    .A1(_05390_),
    .A2(_05391_),
    .ZN(_05392_)
  );
  INV_X1 _10887_ (
    .A(_05392_),
    .ZN(_05393_)
  );
  AND2_X1 _10888_ (
    .A1(large_1[11]),
    .A2(_03700_),
    .ZN(_05394_)
  );
  INV_X1 _10889_ (
    .A(_05394_),
    .ZN(_05395_)
  );
  AND2_X1 _10890_ (
    .A1(_02669_),
    .A2(_03708_),
    .ZN(_05396_)
  );
  INV_X1 _10891_ (
    .A(_05396_),
    .ZN(_05397_)
  );
  AND2_X1 _10892_ (
    .A1(_05393_),
    .A2(_05395_),
    .ZN(_05398_)
  );
  AND2_X1 _10893_ (
    .A1(_05397_),
    .A2(_05398_),
    .ZN(_05399_)
  );
  INV_X1 _10894_ (
    .A(_05399_),
    .ZN(_05400_)
  );
  AND2_X1 _10895_ (
    .A1(_00811_),
    .A2(_05400_),
    .ZN(_00580_)
  );
  AND2_X1 _10896_ (
    .A1(_00658_),
    .A2(_03677_),
    .ZN(_05401_)
  );
  INV_X1 _10897_ (
    .A(_05401_),
    .ZN(_05402_)
  );
  AND2_X1 _10898_ (
    .A1(_03710_),
    .A2(_05402_),
    .ZN(_05403_)
  );
  AND2_X1 _10899_ (
    .A1(large_1[12]),
    .A2(_03676_),
    .ZN(_05404_)
  );
  INV_X1 _10900_ (
    .A(_05404_),
    .ZN(_05405_)
  );
  AND2_X1 _10901_ (
    .A1(_05403_),
    .A2(_05405_),
    .ZN(_05406_)
  );
  INV_X1 _10902_ (
    .A(_05406_),
    .ZN(_05407_)
  );
  AND2_X1 _10903_ (
    .A1(large_1[12]),
    .A2(_03700_),
    .ZN(_05408_)
  );
  INV_X1 _10904_ (
    .A(_05408_),
    .ZN(_05409_)
  );
  AND2_X1 _10905_ (
    .A1(_01107_),
    .A2(_03708_),
    .ZN(_05410_)
  );
  INV_X1 _10906_ (
    .A(_05410_),
    .ZN(_05411_)
  );
  AND2_X1 _10907_ (
    .A1(_05409_),
    .A2(_05411_),
    .ZN(_05412_)
  );
  AND2_X1 _10908_ (
    .A1(_05407_),
    .A2(_05412_),
    .ZN(_05413_)
  );
  INV_X1 _10909_ (
    .A(_05413_),
    .ZN(_05414_)
  );
  AND2_X1 _10910_ (
    .A1(_00811_),
    .A2(_05414_),
    .ZN(_00581_)
  );
  AND2_X1 _10911_ (
    .A1(_00657_),
    .A2(_05405_),
    .ZN(_05415_)
  );
  INV_X1 _10912_ (
    .A(_05415_),
    .ZN(_05416_)
  );
  AND2_X1 _10913_ (
    .A1(large_1[13]),
    .A2(_05404_),
    .ZN(_05417_)
  );
  INV_X1 _10914_ (
    .A(_05417_),
    .ZN(_05418_)
  );
  AND2_X1 _10915_ (
    .A1(_03710_),
    .A2(_05418_),
    .ZN(_05419_)
  );
  AND2_X1 _10916_ (
    .A1(_05416_),
    .A2(_05419_),
    .ZN(_05420_)
  );
  INV_X1 _10917_ (
    .A(_05420_),
    .ZN(_05421_)
  );
  AND2_X1 _10918_ (
    .A1(large_1[13]),
    .A2(_03700_),
    .ZN(_05422_)
  );
  INV_X1 _10919_ (
    .A(_05422_),
    .ZN(_05423_)
  );
  AND2_X1 _10920_ (
    .A1(_01199_),
    .A2(_03708_),
    .ZN(_05424_)
  );
  INV_X1 _10921_ (
    .A(_05424_),
    .ZN(_05425_)
  );
  AND2_X1 _10922_ (
    .A1(_05423_),
    .A2(_05425_),
    .ZN(_05426_)
  );
  AND2_X1 _10923_ (
    .A1(_05421_),
    .A2(_05426_),
    .ZN(_05427_)
  );
  INV_X1 _10924_ (
    .A(_05427_),
    .ZN(_05428_)
  );
  AND2_X1 _10925_ (
    .A1(_00811_),
    .A2(_05428_),
    .ZN(_00582_)
  );
  AND2_X1 _10926_ (
    .A1(_00656_),
    .A2(_05418_),
    .ZN(_05429_)
  );
  INV_X1 _10927_ (
    .A(_05429_),
    .ZN(_05430_)
  );
  AND2_X1 _10928_ (
    .A1(_03679_),
    .A2(_03710_),
    .ZN(_05431_)
  );
  AND2_X1 _10929_ (
    .A1(_05430_),
    .A2(_05431_),
    .ZN(_05432_)
  );
  INV_X1 _10930_ (
    .A(_05432_),
    .ZN(_05433_)
  );
  AND2_X1 _10931_ (
    .A1(large_1[14]),
    .A2(_03700_),
    .ZN(_05434_)
  );
  INV_X1 _10932_ (
    .A(_05434_),
    .ZN(_05435_)
  );
  AND2_X1 _10933_ (
    .A1(_01277_),
    .A2(_03702_),
    .ZN(_05436_)
  );
  INV_X1 _10934_ (
    .A(_05436_),
    .ZN(_05437_)
  );
  AND2_X1 _10935_ (
    .A1(_05435_),
    .A2(_05437_),
    .ZN(_05438_)
  );
  AND2_X1 _10936_ (
    .A1(_05433_),
    .A2(_05438_),
    .ZN(_05439_)
  );
  INV_X1 _10937_ (
    .A(_05439_),
    .ZN(_05440_)
  );
  AND2_X1 _10938_ (
    .A1(_00811_),
    .A2(_05440_),
    .ZN(_00583_)
  );
  AND2_X1 _10939_ (
    .A1(_00655_),
    .A2(_03679_),
    .ZN(_05441_)
  );
  INV_X1 _10940_ (
    .A(_05441_),
    .ZN(_05442_)
  );
  AND2_X1 _10941_ (
    .A1(large_1[15]),
    .A2(_03678_),
    .ZN(_05443_)
  );
  INV_X1 _10942_ (
    .A(_05443_),
    .ZN(_05444_)
  );
  AND2_X1 _10943_ (
    .A1(_03710_),
    .A2(_05444_),
    .ZN(_05445_)
  );
  AND2_X1 _10944_ (
    .A1(large_1[15]),
    .A2(_03691_),
    .ZN(_05446_)
  );
  AND2_X1 _10945_ (
    .A1(_05442_),
    .A2(_05445_),
    .ZN(_05447_)
  );
  INV_X1 _10946_ (
    .A(_05447_),
    .ZN(_05448_)
  );
  AND2_X1 _10947_ (
    .A1(large_1[15]),
    .A2(_03700_),
    .ZN(_05449_)
  );
  INV_X1 _10948_ (
    .A(_05449_),
    .ZN(_05450_)
  );
  AND2_X1 _10949_ (
    .A1(_02735_),
    .A2(_03708_),
    .ZN(_05451_)
  );
  INV_X1 _10950_ (
    .A(_05451_),
    .ZN(_05452_)
  );
  AND2_X1 _10951_ (
    .A1(_05450_),
    .A2(_05452_),
    .ZN(_05453_)
  );
  AND2_X1 _10952_ (
    .A1(_05448_),
    .A2(_05453_),
    .ZN(_05454_)
  );
  INV_X1 _10953_ (
    .A(_05454_),
    .ZN(_05455_)
  );
  AND2_X1 _10954_ (
    .A1(_00811_),
    .A2(_05455_),
    .ZN(_00584_)
  );
  AND2_X1 _10955_ (
    .A1(_00654_),
    .A2(_05444_),
    .ZN(_05456_)
  );
  INV_X1 _10956_ (
    .A(_05456_),
    .ZN(_05457_)
  );
  AND2_X1 _10957_ (
    .A1(large_1[16]),
    .A2(_05443_),
    .ZN(_05458_)
  );
  INV_X1 _10958_ (
    .A(_05458_),
    .ZN(_05459_)
  );
  AND2_X1 _10959_ (
    .A1(_03710_),
    .A2(_05459_),
    .ZN(_05460_)
  );
  AND2_X1 _10960_ (
    .A1(_05457_),
    .A2(_05460_),
    .ZN(_05461_)
  );
  INV_X1 _10961_ (
    .A(_05461_),
    .ZN(_05462_)
  );
  AND2_X1 _10962_ (
    .A1(large_1[16]),
    .A2(_03700_),
    .ZN(_05463_)
  );
  INV_X1 _10963_ (
    .A(_05463_),
    .ZN(_05464_)
  );
  AND2_X1 _10964_ (
    .A1(_02801_),
    .A2(_03702_),
    .ZN(_05465_)
  );
  INV_X1 _10965_ (
    .A(_05465_),
    .ZN(_05466_)
  );
  AND2_X1 _10966_ (
    .A1(_05464_),
    .A2(_05466_),
    .ZN(_05467_)
  );
  AND2_X1 _10967_ (
    .A1(_05462_),
    .A2(_05467_),
    .ZN(_05468_)
  );
  INV_X1 _10968_ (
    .A(_05468_),
    .ZN(_05469_)
  );
  AND2_X1 _10969_ (
    .A1(_00811_),
    .A2(_05469_),
    .ZN(_00585_)
  );
  AND2_X1 _10970_ (
    .A1(_00653_),
    .A2(_05459_),
    .ZN(_05470_)
  );
  INV_X1 _10971_ (
    .A(_05470_),
    .ZN(_05471_)
  );
  AND2_X1 _10972_ (
    .A1(large_1[17]),
    .A2(_05458_),
    .ZN(_05472_)
  );
  AND2_X1 _10973_ (
    .A1(_03636_),
    .A2(_05446_),
    .ZN(_05473_)
  );
  INV_X1 _10974_ (
    .A(_05473_),
    .ZN(_05474_)
  );
  AND2_X1 _10975_ (
    .A1(_03710_),
    .A2(_05474_),
    .ZN(_05475_)
  );
  AND2_X1 _10976_ (
    .A1(_05471_),
    .A2(_05475_),
    .ZN(_05476_)
  );
  INV_X1 _10977_ (
    .A(_05476_),
    .ZN(_05477_)
  );
  AND2_X1 _10978_ (
    .A1(large_1[17]),
    .A2(_03700_),
    .ZN(_05478_)
  );
  INV_X1 _10979_ (
    .A(_05478_),
    .ZN(_05479_)
  );
  AND2_X1 _10980_ (
    .A1(_01360_),
    .A2(_03702_),
    .ZN(_05480_)
  );
  INV_X1 _10981_ (
    .A(_05480_),
    .ZN(_05481_)
  );
  AND2_X1 _10982_ (
    .A1(_05479_),
    .A2(_05481_),
    .ZN(_05482_)
  );
  AND2_X1 _10983_ (
    .A1(_05477_),
    .A2(_05482_),
    .ZN(_05483_)
  );
  INV_X1 _10984_ (
    .A(_05483_),
    .ZN(_05484_)
  );
  AND2_X1 _10985_ (
    .A1(_00811_),
    .A2(_05484_),
    .ZN(_00586_)
  );
  AND2_X1 _10986_ (
    .A1(_00652_),
    .A2(_05474_),
    .ZN(_05485_)
  );
  INV_X1 _10987_ (
    .A(_05485_),
    .ZN(_05486_)
  );
  AND2_X1 _10988_ (
    .A1(large_1[18]),
    .A2(_05472_),
    .ZN(_05487_)
  );
  AND2_X1 _10989_ (
    .A1(large_1[18]),
    .A2(_05473_),
    .ZN(_05488_)
  );
  INV_X1 _10990_ (
    .A(_05488_),
    .ZN(_05489_)
  );
  AND2_X1 _10991_ (
    .A1(_03710_),
    .A2(_05489_),
    .ZN(_05490_)
  );
  AND2_X1 _10992_ (
    .A1(_05486_),
    .A2(_05490_),
    .ZN(_05491_)
  );
  INV_X1 _10993_ (
    .A(_05491_),
    .ZN(_05492_)
  );
  AND2_X1 _10994_ (
    .A1(large_1[18]),
    .A2(_03700_),
    .ZN(_05493_)
  );
  INV_X1 _10995_ (
    .A(_05493_),
    .ZN(_05494_)
  );
  AND2_X1 _10996_ (
    .A1(_02873_),
    .A2(_03702_),
    .ZN(_05495_)
  );
  INV_X1 _10997_ (
    .A(_05495_),
    .ZN(_05496_)
  );
  AND2_X1 _10998_ (
    .A1(_05494_),
    .A2(_05496_),
    .ZN(_05497_)
  );
  AND2_X1 _10999_ (
    .A1(_05492_),
    .A2(_05497_),
    .ZN(_05498_)
  );
  INV_X1 _11000_ (
    .A(_05498_),
    .ZN(_05499_)
  );
  AND2_X1 _11001_ (
    .A1(_00811_),
    .A2(_05499_),
    .ZN(_00587_)
  );
  AND2_X1 _11002_ (
    .A1(_00651_),
    .A2(_05489_),
    .ZN(_05500_)
  );
  INV_X1 _11003_ (
    .A(_05500_),
    .ZN(_05501_)
  );
  AND2_X1 _11004_ (
    .A1(large_1[19]),
    .A2(_05487_),
    .ZN(_05502_)
  );
  INV_X1 _11005_ (
    .A(_05502_),
    .ZN(_05503_)
  );
  AND2_X1 _11006_ (
    .A1(_03710_),
    .A2(_05503_),
    .ZN(_05504_)
  );
  AND2_X1 _11007_ (
    .A1(_05501_),
    .A2(_05504_),
    .ZN(_05505_)
  );
  INV_X1 _11008_ (
    .A(_05505_),
    .ZN(_05506_)
  );
  AND2_X1 _11009_ (
    .A1(large_1[19]),
    .A2(_03700_),
    .ZN(_05507_)
  );
  INV_X1 _11010_ (
    .A(_05507_),
    .ZN(_05508_)
  );
  AND2_X1 _11011_ (
    .A1(_02945_),
    .A2(_03708_),
    .ZN(_05509_)
  );
  INV_X1 _11012_ (
    .A(_05509_),
    .ZN(_05510_)
  );
  AND2_X1 _11013_ (
    .A1(_05508_),
    .A2(_05510_),
    .ZN(_05511_)
  );
  AND2_X1 _11014_ (
    .A1(_05506_),
    .A2(_05511_),
    .ZN(_05512_)
  );
  INV_X1 _11015_ (
    .A(_05512_),
    .ZN(_05513_)
  );
  AND2_X1 _11016_ (
    .A1(_00811_),
    .A2(_05513_),
    .ZN(_00588_)
  );
  AND2_X1 _11017_ (
    .A1(_00650_),
    .A2(_05503_),
    .ZN(_05514_)
  );
  INV_X1 _11018_ (
    .A(_05514_),
    .ZN(_05515_)
  );
  AND2_X1 _11019_ (
    .A1(large_1[20]),
    .A2(_05502_),
    .ZN(_05516_)
  );
  INV_X1 _11020_ (
    .A(_05516_),
    .ZN(_05517_)
  );
  AND2_X1 _11021_ (
    .A1(_03710_),
    .A2(_05517_),
    .ZN(_05518_)
  );
  AND2_X1 _11022_ (
    .A1(_05515_),
    .A2(_05518_),
    .ZN(_05519_)
  );
  INV_X1 _11023_ (
    .A(_05519_),
    .ZN(_05520_)
  );
  AND2_X1 _11024_ (
    .A1(large_1[20]),
    .A2(_03700_),
    .ZN(_05521_)
  );
  INV_X1 _11025_ (
    .A(_05521_),
    .ZN(_05522_)
  );
  AND2_X1 _11026_ (
    .A1(_03017_),
    .A2(_03702_),
    .ZN(_05523_)
  );
  INV_X1 _11027_ (
    .A(_05523_),
    .ZN(_05524_)
  );
  AND2_X1 _11028_ (
    .A1(_05522_),
    .A2(_05524_),
    .ZN(_05525_)
  );
  AND2_X1 _11029_ (
    .A1(_05520_),
    .A2(_05525_),
    .ZN(_05526_)
  );
  INV_X1 _11030_ (
    .A(_05526_),
    .ZN(_05527_)
  );
  AND2_X1 _11031_ (
    .A1(_00811_),
    .A2(_05527_),
    .ZN(_00589_)
  );
  AND2_X1 _11032_ (
    .A1(_00649_),
    .A2(_05517_),
    .ZN(_05528_)
  );
  INV_X1 _11033_ (
    .A(_05528_),
    .ZN(_05529_)
  );
  AND2_X1 _11034_ (
    .A1(_03710_),
    .A2(_05529_),
    .ZN(_05530_)
  );
  AND2_X1 _11035_ (
    .A1(large_1[21]),
    .A2(_05516_),
    .ZN(_05531_)
  );
  INV_X1 _11036_ (
    .A(_05531_),
    .ZN(_05532_)
  );
  AND2_X1 _11037_ (
    .A1(_05530_),
    .A2(_05532_),
    .ZN(_05533_)
  );
  INV_X1 _11038_ (
    .A(_05533_),
    .ZN(_05534_)
  );
  AND2_X1 _11039_ (
    .A1(large_1[21]),
    .A2(_03700_),
    .ZN(_05535_)
  );
  INV_X1 _11040_ (
    .A(_05535_),
    .ZN(_05536_)
  );
  AND2_X1 _11041_ (
    .A1(_03089_),
    .A2(_03708_),
    .ZN(_05537_)
  );
  INV_X1 _11042_ (
    .A(_05537_),
    .ZN(_05538_)
  );
  AND2_X1 _11043_ (
    .A1(_05536_),
    .A2(_05538_),
    .ZN(_05539_)
  );
  AND2_X1 _11044_ (
    .A1(_05534_),
    .A2(_05539_),
    .ZN(_05540_)
  );
  INV_X1 _11045_ (
    .A(_05540_),
    .ZN(_05541_)
  );
  AND2_X1 _11046_ (
    .A1(_00811_),
    .A2(_05541_),
    .ZN(_00590_)
  );
  AND2_X1 _11047_ (
    .A1(_00648_),
    .A2(_05532_),
    .ZN(_05542_)
  );
  INV_X1 _11048_ (
    .A(_05542_),
    .ZN(_05543_)
  );
  AND2_X1 _11049_ (
    .A1(large_1[22]),
    .A2(_05531_),
    .ZN(_05544_)
  );
  INV_X1 _11050_ (
    .A(_05544_),
    .ZN(_05545_)
  );
  AND2_X1 _11051_ (
    .A1(_03710_),
    .A2(_05545_),
    .ZN(_05546_)
  );
  AND2_X1 _11052_ (
    .A1(_05543_),
    .A2(_05546_),
    .ZN(_05547_)
  );
  INV_X1 _11053_ (
    .A(_05547_),
    .ZN(_05548_)
  );
  AND2_X1 _11054_ (
    .A1(large_1[22]),
    .A2(_03700_),
    .ZN(_05549_)
  );
  INV_X1 _11055_ (
    .A(_05549_),
    .ZN(_05550_)
  );
  AND2_X1 _11056_ (
    .A1(_03162_),
    .A2(_03702_),
    .ZN(_05551_)
  );
  INV_X1 _11057_ (
    .A(_05551_),
    .ZN(_05552_)
  );
  AND2_X1 _11058_ (
    .A1(_05550_),
    .A2(_05552_),
    .ZN(_05553_)
  );
  AND2_X1 _11059_ (
    .A1(_05548_),
    .A2(_05553_),
    .ZN(_05554_)
  );
  INV_X1 _11060_ (
    .A(_05554_),
    .ZN(_05555_)
  );
  AND2_X1 _11061_ (
    .A1(_00811_),
    .A2(_05555_),
    .ZN(_00591_)
  );
  AND2_X1 _11062_ (
    .A1(_00647_),
    .A2(_05545_),
    .ZN(_05556_)
  );
  INV_X1 _11063_ (
    .A(_05556_),
    .ZN(_05557_)
  );
  AND2_X1 _11064_ (
    .A1(large_1[23]),
    .A2(_05544_),
    .ZN(_05558_)
  );
  INV_X1 _11065_ (
    .A(_05558_),
    .ZN(_05559_)
  );
  AND2_X1 _11066_ (
    .A1(_03710_),
    .A2(_05557_),
    .ZN(_05560_)
  );
  AND2_X1 _11067_ (
    .A1(_05559_),
    .A2(_05560_),
    .ZN(_05561_)
  );
  INV_X1 _11068_ (
    .A(_05561_),
    .ZN(_05562_)
  );
  AND2_X1 _11069_ (
    .A1(large_1[23]),
    .A2(_03700_),
    .ZN(_05563_)
  );
  INV_X1 _11070_ (
    .A(_05563_),
    .ZN(_05564_)
  );
  AND2_X1 _11071_ (
    .A1(_03230_),
    .A2(_03702_),
    .ZN(_05565_)
  );
  INV_X1 _11072_ (
    .A(_05565_),
    .ZN(_05566_)
  );
  AND2_X1 _11073_ (
    .A1(_05564_),
    .A2(_05566_),
    .ZN(_05567_)
  );
  AND2_X1 _11074_ (
    .A1(_05562_),
    .A2(_05567_),
    .ZN(_05568_)
  );
  INV_X1 _11075_ (
    .A(_05568_),
    .ZN(_05569_)
  );
  AND2_X1 _11076_ (
    .A1(_00811_),
    .A2(_05569_),
    .ZN(_00592_)
  );
  AND2_X1 _11077_ (
    .A1(_00646_),
    .A2(_03693_),
    .ZN(_05570_)
  );
  INV_X1 _11078_ (
    .A(_05570_),
    .ZN(_05571_)
  );
  AND2_X1 _11079_ (
    .A1(_03710_),
    .A2(_05571_),
    .ZN(_05572_)
  );
  AND2_X1 _11080_ (
    .A1(_03695_),
    .A2(_05572_),
    .ZN(_05573_)
  );
  INV_X1 _11081_ (
    .A(_05573_),
    .ZN(_05574_)
  );
  AND2_X1 _11082_ (
    .A1(large_1[24]),
    .A2(_03700_),
    .ZN(_05575_)
  );
  INV_X1 _11083_ (
    .A(_05575_),
    .ZN(_05576_)
  );
  AND2_X1 _11084_ (
    .A1(_03443_),
    .A2(_03702_),
    .ZN(_05577_)
  );
  INV_X1 _11085_ (
    .A(_05577_),
    .ZN(_05578_)
  );
  AND2_X1 _11086_ (
    .A1(_05576_),
    .A2(_05578_),
    .ZN(_05579_)
  );
  AND2_X1 _11087_ (
    .A1(_05574_),
    .A2(_05579_),
    .ZN(_05580_)
  );
  INV_X1 _11088_ (
    .A(_05580_),
    .ZN(_05581_)
  );
  AND2_X1 _11089_ (
    .A1(_00811_),
    .A2(_05581_),
    .ZN(_00593_)
  );
  AND2_X1 _11090_ (
    .A1(_00645_),
    .A2(_03695_),
    .ZN(_05582_)
  );
  INV_X1 _11091_ (
    .A(_05582_),
    .ZN(_05583_)
  );
  AND2_X1 _11092_ (
    .A1(_03710_),
    .A2(_05583_),
    .ZN(_05584_)
  );
  AND2_X1 _11093_ (
    .A1(_03697_),
    .A2(_05584_),
    .ZN(_05585_)
  );
  INV_X1 _11094_ (
    .A(_05585_),
    .ZN(_05586_)
  );
  AND2_X1 _11095_ (
    .A1(large_1[25]),
    .A2(_03700_),
    .ZN(_05587_)
  );
  INV_X1 _11096_ (
    .A(_05587_),
    .ZN(_05588_)
  );
  AND2_X1 _11097_ (
    .A1(_03342_),
    .A2(_03708_),
    .ZN(_05589_)
  );
  INV_X1 _11098_ (
    .A(_05589_),
    .ZN(_05590_)
  );
  AND2_X1 _11099_ (
    .A1(_05588_),
    .A2(_05590_),
    .ZN(_05591_)
  );
  AND2_X1 _11100_ (
    .A1(_05586_),
    .A2(_05591_),
    .ZN(_05592_)
  );
  INV_X1 _11101_ (
    .A(_05592_),
    .ZN(_05593_)
  );
  AND2_X1 _11102_ (
    .A1(_00811_),
    .A2(_05593_),
    .ZN(_00594_)
  );
  AND2_X1 _11103_ (
    .A1(large_[0]),
    .A2(_04388_),
    .ZN(_05594_)
  );
  INV_X1 _11104_ (
    .A(_05594_),
    .ZN(_05595_)
  );
  MUX2_X1 _11105_ (
    .A(large_[0]),
    .B(_large_r_T_1[0]),
    .S(_04334_),
    .Z(_05596_)
  );
  AND2_X1 _11106_ (
    .A1(_04398_),
    .A2(_05596_),
    .ZN(_05597_)
  );
  INV_X1 _11107_ (
    .A(_05597_),
    .ZN(_05598_)
  );
  AND2_X1 _11108_ (
    .A1(_05595_),
    .A2(_05598_),
    .ZN(_05599_)
  );
  AND2_X1 _11109_ (
    .A1(_02076_),
    .A2(_04396_),
    .ZN(_05600_)
  );
  INV_X1 _11110_ (
    .A(_05600_),
    .ZN(_05601_)
  );
  AND2_X1 _11111_ (
    .A1(_05599_),
    .A2(_05601_),
    .ZN(_05602_)
  );
  INV_X1 _11112_ (
    .A(_05602_),
    .ZN(_05603_)
  );
  AND2_X1 _11113_ (
    .A1(_00811_),
    .A2(_05603_),
    .ZN(_00595_)
  );
  AND2_X1 _11114_ (
    .A1(large_[0]),
    .A2(_04334_),
    .ZN(_05604_)
  );
  INV_X1 _11115_ (
    .A(_05604_),
    .ZN(_05605_)
  );
  AND2_X1 _11116_ (
    .A1(_00644_),
    .A2(_05605_),
    .ZN(_05606_)
  );
  INV_X1 _11117_ (
    .A(_05606_),
    .ZN(_05607_)
  );
  AND2_X1 _11118_ (
    .A1(large_[1]),
    .A2(_04388_),
    .ZN(_05608_)
  );
  INV_X1 _11119_ (
    .A(_05608_),
    .ZN(_05609_)
  );
  AND2_X1 _11120_ (
    .A1(_04337_),
    .A2(_04394_),
    .ZN(_05610_)
  );
  INV_X1 _11121_ (
    .A(_05610_),
    .ZN(_05611_)
  );
  AND2_X1 _11122_ (
    .A1(_05609_),
    .A2(_05611_),
    .ZN(_05612_)
  );
  INV_X1 _11123_ (
    .A(_05612_),
    .ZN(_05613_)
  );
  AND2_X1 _11124_ (
    .A1(_05607_),
    .A2(_05613_),
    .ZN(_05614_)
  );
  INV_X1 _11125_ (
    .A(_05614_),
    .ZN(_05615_)
  );
  AND2_X1 _11126_ (
    .A1(_02163_),
    .A2(_04396_),
    .ZN(_05616_)
  );
  INV_X1 _11127_ (
    .A(_05616_),
    .ZN(_05617_)
  );
  AND2_X1 _11128_ (
    .A1(_05615_),
    .A2(_05617_),
    .ZN(_05618_)
  );
  INV_X1 _11129_ (
    .A(_05618_),
    .ZN(_05619_)
  );
  AND2_X1 _11130_ (
    .A1(_00811_),
    .A2(_05619_),
    .ZN(_00596_)
  );
  AND2_X1 _11131_ (
    .A1(large_[2]),
    .A2(_04336_),
    .ZN(_05620_)
  );
  INV_X1 _11132_ (
    .A(_05620_),
    .ZN(_05621_)
  );
  AND2_X1 _11133_ (
    .A1(_00643_),
    .A2(_04337_),
    .ZN(_05622_)
  );
  INV_X1 _11134_ (
    .A(_05622_),
    .ZN(_05623_)
  );
  AND2_X1 _11135_ (
    .A1(_05621_),
    .A2(_05623_),
    .ZN(_05624_)
  );
  AND2_X1 _11136_ (
    .A1(_04393_),
    .A2(_05624_),
    .ZN(_05625_)
  );
  INV_X1 _11137_ (
    .A(_05625_),
    .ZN(_05626_)
  );
  AND2_X1 _11138_ (
    .A1(large_[2]),
    .A2(_04388_),
    .ZN(_05627_)
  );
  INV_X1 _11139_ (
    .A(_05627_),
    .ZN(_05628_)
  );
  AND2_X1 _11140_ (
    .A1(_00898_),
    .A2(_05624_),
    .ZN(_05629_)
  );
  INV_X1 _11141_ (
    .A(_05629_),
    .ZN(_05630_)
  );
  AND2_X1 _11142_ (
    .A1(_05628_),
    .A2(_05630_),
    .ZN(_05631_)
  );
  AND2_X1 _11143_ (
    .A1(_05626_),
    .A2(_05631_),
    .ZN(_05632_)
  );
  AND2_X1 _11144_ (
    .A1(_01446_),
    .A2(_04396_),
    .ZN(_05633_)
  );
  INV_X1 _11145_ (
    .A(_05633_),
    .ZN(_05634_)
  );
  AND2_X1 _11146_ (
    .A1(_05632_),
    .A2(_05634_),
    .ZN(_05635_)
  );
  INV_X1 _11147_ (
    .A(_05635_),
    .ZN(_05636_)
  );
  AND2_X1 _11148_ (
    .A1(_00811_),
    .A2(_05636_),
    .ZN(_00597_)
  );
  AND2_X1 _11149_ (
    .A1(_00642_),
    .A2(_05621_),
    .ZN(_05637_)
  );
  INV_X1 _11150_ (
    .A(_05637_),
    .ZN(_05638_)
  );
  AND2_X1 _11151_ (
    .A1(large_[3]),
    .A2(_04388_),
    .ZN(_05639_)
  );
  INV_X1 _11152_ (
    .A(_05639_),
    .ZN(_05640_)
  );
  AND2_X1 _11153_ (
    .A1(large_[3]),
    .A2(_05620_),
    .ZN(_05641_)
  );
  INV_X1 _11154_ (
    .A(_05641_),
    .ZN(_05642_)
  );
  AND2_X1 _11155_ (
    .A1(_01518_),
    .A2(_04396_),
    .ZN(_05643_)
  );
  INV_X1 _11156_ (
    .A(_05643_),
    .ZN(_05644_)
  );
  AND2_X1 _11157_ (
    .A1(_05638_),
    .A2(_05642_),
    .ZN(_05645_)
  );
  AND2_X1 _11158_ (
    .A1(_04398_),
    .A2(_05645_),
    .ZN(_05646_)
  );
  INV_X1 _11159_ (
    .A(_05646_),
    .ZN(_05647_)
  );
  AND2_X1 _11160_ (
    .A1(_05644_),
    .A2(_05647_),
    .ZN(_05648_)
  );
  AND2_X1 _11161_ (
    .A1(_05640_),
    .A2(_05648_),
    .ZN(_05649_)
  );
  INV_X1 _11162_ (
    .A(_05649_),
    .ZN(_05650_)
  );
  AND2_X1 _11163_ (
    .A1(_00811_),
    .A2(_05650_),
    .ZN(_00598_)
  );
  AND2_X1 _11164_ (
    .A1(_00641_),
    .A2(_05642_),
    .ZN(_05651_)
  );
  INV_X1 _11165_ (
    .A(_05651_),
    .ZN(_05652_)
  );
  AND2_X1 _11166_ (
    .A1(large_[4]),
    .A2(_04388_),
    .ZN(_05653_)
  );
  INV_X1 _11167_ (
    .A(_05653_),
    .ZN(_05654_)
  );
  AND2_X1 _11168_ (
    .A1(large_[4]),
    .A2(_05641_),
    .ZN(_05655_)
  );
  INV_X1 _11169_ (
    .A(_05655_),
    .ZN(_05656_)
  );
  AND2_X1 _11170_ (
    .A1(_05652_),
    .A2(_05656_),
    .ZN(_05657_)
  );
  AND2_X1 _11171_ (
    .A1(_04398_),
    .A2(_05657_),
    .ZN(_05658_)
  );
  INV_X1 _11172_ (
    .A(_05658_),
    .ZN(_05659_)
  );
  AND2_X1 _11173_ (
    .A1(_05654_),
    .A2(_05659_),
    .ZN(_05660_)
  );
  AND2_X1 _11174_ (
    .A1(_02235_),
    .A2(_04390_),
    .ZN(_05661_)
  );
  INV_X1 _11175_ (
    .A(_05661_),
    .ZN(_05662_)
  );
  AND2_X1 _11176_ (
    .A1(_05660_),
    .A2(_05662_),
    .ZN(_05663_)
  );
  INV_X1 _11177_ (
    .A(_05663_),
    .ZN(_05664_)
  );
  AND2_X1 _11178_ (
    .A1(_00811_),
    .A2(_05664_),
    .ZN(_00599_)
  );
  AND2_X1 _11179_ (
    .A1(large_[5]),
    .A2(_04388_),
    .ZN(_05665_)
  );
  INV_X1 _11180_ (
    .A(_05665_),
    .ZN(_05666_)
  );
  AND2_X1 _11181_ (
    .A1(_04338_),
    .A2(_05641_),
    .ZN(_05667_)
  );
  INV_X1 _11182_ (
    .A(_05667_),
    .ZN(_05668_)
  );
  AND2_X1 _11183_ (
    .A1(_00640_),
    .A2(_05656_),
    .ZN(_05669_)
  );
  INV_X1 _11184_ (
    .A(_05669_),
    .ZN(_05670_)
  );
  AND2_X1 _11185_ (
    .A1(_05668_),
    .A2(_05670_),
    .ZN(_05671_)
  );
  INV_X1 _11186_ (
    .A(_05671_),
    .ZN(_05672_)
  );
  AND2_X1 _11187_ (
    .A1(_02314_),
    .A2(_04390_),
    .ZN(_05673_)
  );
  INV_X1 _11188_ (
    .A(_05673_),
    .ZN(_05674_)
  );
  AND2_X1 _11189_ (
    .A1(_05672_),
    .A2(_05674_),
    .ZN(_05675_)
  );
  INV_X1 _11190_ (
    .A(_05675_),
    .ZN(_05676_)
  );
  AND2_X1 _11191_ (
    .A1(_02314_),
    .A2(_04389_),
    .ZN(_05677_)
  );
  INV_X1 _11192_ (
    .A(_05677_),
    .ZN(_05678_)
  );
  AND2_X1 _11193_ (
    .A1(_04399_),
    .A2(_05678_),
    .ZN(_05679_)
  );
  INV_X1 _11194_ (
    .A(_05679_),
    .ZN(_05680_)
  );
  AND2_X1 _11195_ (
    .A1(_05676_),
    .A2(_05680_),
    .ZN(_05681_)
  );
  INV_X1 _11196_ (
    .A(_05681_),
    .ZN(_05682_)
  );
  AND2_X1 _11197_ (
    .A1(_05666_),
    .A2(_05682_),
    .ZN(_05683_)
  );
  INV_X1 _11198_ (
    .A(_05683_),
    .ZN(_05684_)
  );
  AND2_X1 _11199_ (
    .A1(_00811_),
    .A2(_05684_),
    .ZN(_00600_)
  );
  AND2_X1 _11200_ (
    .A1(large_[6]),
    .A2(_04388_),
    .ZN(_05685_)
  );
  INV_X1 _11201_ (
    .A(_05685_),
    .ZN(_05686_)
  );
  AND2_X1 _11202_ (
    .A1(_00639_),
    .A2(_05668_),
    .ZN(_05687_)
  );
  INV_X1 _11203_ (
    .A(_05687_),
    .ZN(_05688_)
  );
  AND2_X1 _11204_ (
    .A1(large_[6]),
    .A2(_05667_),
    .ZN(_05689_)
  );
  INV_X1 _11205_ (
    .A(_05689_),
    .ZN(_05690_)
  );
  AND2_X1 _11206_ (
    .A1(_05688_),
    .A2(_05690_),
    .ZN(_05691_)
  );
  INV_X1 _11207_ (
    .A(_05691_),
    .ZN(_05692_)
  );
  AND2_X1 _11208_ (
    .A1(_02389_),
    .A2(_04390_),
    .ZN(_05693_)
  );
  INV_X1 _11209_ (
    .A(_05693_),
    .ZN(_05694_)
  );
  AND2_X1 _11210_ (
    .A1(_05692_),
    .A2(_05694_),
    .ZN(_05695_)
  );
  INV_X1 _11211_ (
    .A(_05695_),
    .ZN(_05696_)
  );
  AND2_X1 _11212_ (
    .A1(_02389_),
    .A2(_04389_),
    .ZN(_05697_)
  );
  INV_X1 _11213_ (
    .A(_05697_),
    .ZN(_05698_)
  );
  AND2_X1 _11214_ (
    .A1(_04399_),
    .A2(_05698_),
    .ZN(_05699_)
  );
  INV_X1 _11215_ (
    .A(_05699_),
    .ZN(_05700_)
  );
  AND2_X1 _11216_ (
    .A1(_05696_),
    .A2(_05700_),
    .ZN(_05701_)
  );
  INV_X1 _11217_ (
    .A(_05701_),
    .ZN(_05702_)
  );
  AND2_X1 _11218_ (
    .A1(_05686_),
    .A2(_05702_),
    .ZN(_05703_)
  );
  INV_X1 _11219_ (
    .A(_05703_),
    .ZN(_05704_)
  );
  AND2_X1 _11220_ (
    .A1(_00811_),
    .A2(_05704_),
    .ZN(_00601_)
  );
  AND2_X1 _11221_ (
    .A1(_00638_),
    .A2(_04375_),
    .ZN(_05705_)
  );
  INV_X1 _11222_ (
    .A(_05705_),
    .ZN(_05706_)
  );
  AND2_X1 _11223_ (
    .A1(large_[7]),
    .A2(_04374_),
    .ZN(_05707_)
  );
  INV_X1 _11224_ (
    .A(_05707_),
    .ZN(_05708_)
  );
  AND2_X1 _11225_ (
    .A1(_05706_),
    .A2(_05708_),
    .ZN(_05709_)
  );
  INV_X1 _11226_ (
    .A(_05709_),
    .ZN(_05710_)
  );
  AND2_X1 _11227_ (
    .A1(_01028_),
    .A2(_05710_),
    .ZN(_05711_)
  );
  INV_X1 _11228_ (
    .A(_05711_),
    .ZN(_05712_)
  );
  AND2_X1 _11229_ (
    .A1(_04392_),
    .A2(_05712_),
    .ZN(_05713_)
  );
  AND2_X1 _11230_ (
    .A1(_01027_),
    .A2(_02455_),
    .ZN(_05714_)
  );
  INV_X1 _11231_ (
    .A(_05714_),
    .ZN(_05715_)
  );
  AND2_X1 _11232_ (
    .A1(_05713_),
    .A2(_05715_),
    .ZN(_05716_)
  );
  INV_X1 _11233_ (
    .A(_05716_),
    .ZN(_05717_)
  );
  AND2_X1 _11234_ (
    .A1(_00898_),
    .A2(_05709_),
    .ZN(_05718_)
  );
  INV_X1 _11235_ (
    .A(_05718_),
    .ZN(_05719_)
  );
  AND2_X1 _11236_ (
    .A1(large_[7]),
    .A2(_04388_),
    .ZN(_05720_)
  );
  INV_X1 _11237_ (
    .A(_05720_),
    .ZN(_05721_)
  );
  AND2_X1 _11238_ (
    .A1(_05719_),
    .A2(_05721_),
    .ZN(_05722_)
  );
  AND2_X1 _11239_ (
    .A1(_05717_),
    .A2(_05722_),
    .ZN(_05723_)
  );
  INV_X1 _11240_ (
    .A(_05723_),
    .ZN(_05724_)
  );
  AND2_X1 _11241_ (
    .A1(_00811_),
    .A2(_05724_),
    .ZN(_00602_)
  );
  AND2_X1 _11242_ (
    .A1(large_[8]),
    .A2(_04388_),
    .ZN(_05725_)
  );
  INV_X1 _11243_ (
    .A(_05725_),
    .ZN(_05726_)
  );
  AND2_X1 _11244_ (
    .A1(_00637_),
    .A2(_05708_),
    .ZN(_05727_)
  );
  INV_X1 _11245_ (
    .A(_05727_),
    .ZN(_05728_)
  );
  AND2_X1 _11246_ (
    .A1(large_[8]),
    .A2(_05707_),
    .ZN(_05729_)
  );
  INV_X1 _11247_ (
    .A(_05729_),
    .ZN(_05730_)
  );
  AND2_X1 _11248_ (
    .A1(_05728_),
    .A2(_05730_),
    .ZN(_05731_)
  );
  INV_X1 _11249_ (
    .A(_05731_),
    .ZN(_05732_)
  );
  AND2_X1 _11250_ (
    .A1(_02522_),
    .A2(_04390_),
    .ZN(_05733_)
  );
  INV_X1 _11251_ (
    .A(_05733_),
    .ZN(_05734_)
  );
  AND2_X1 _11252_ (
    .A1(_05732_),
    .A2(_05734_),
    .ZN(_05735_)
  );
  INV_X1 _11253_ (
    .A(_05735_),
    .ZN(_05736_)
  );
  AND2_X1 _11254_ (
    .A1(_02522_),
    .A2(_04389_),
    .ZN(_05737_)
  );
  INV_X1 _11255_ (
    .A(_05737_),
    .ZN(_05738_)
  );
  AND2_X1 _11256_ (
    .A1(_04399_),
    .A2(_05738_),
    .ZN(_05739_)
  );
  INV_X1 _11257_ (
    .A(_05739_),
    .ZN(_05740_)
  );
  AND2_X1 _11258_ (
    .A1(_05736_),
    .A2(_05740_),
    .ZN(_05741_)
  );
  INV_X1 _11259_ (
    .A(_05741_),
    .ZN(_05742_)
  );
  AND2_X1 _11260_ (
    .A1(_05726_),
    .A2(_05742_),
    .ZN(_05743_)
  );
  INV_X1 _11261_ (
    .A(_05743_),
    .ZN(_05744_)
  );
  AND2_X1 _11262_ (
    .A1(_00811_),
    .A2(_05744_),
    .ZN(_00603_)
  );
  AND2_X1 _11263_ (
    .A1(_00636_),
    .A2(_05730_),
    .ZN(_05745_)
  );
  INV_X1 _11264_ (
    .A(_05745_),
    .ZN(_05746_)
  );
  AND2_X1 _11265_ (
    .A1(large_[9]),
    .A2(_04388_),
    .ZN(_05747_)
  );
  INV_X1 _11266_ (
    .A(_05747_),
    .ZN(_05748_)
  );
  AND2_X1 _11267_ (
    .A1(_04346_),
    .A2(_04398_),
    .ZN(_05749_)
  );
  AND2_X1 _11268_ (
    .A1(_05746_),
    .A2(_05749_),
    .ZN(_05750_)
  );
  INV_X1 _11269_ (
    .A(_05750_),
    .ZN(_05751_)
  );
  AND2_X1 _11270_ (
    .A1(_05748_),
    .A2(_05751_),
    .ZN(_05752_)
  );
  AND2_X1 _11271_ (
    .A1(_02597_),
    .A2(_04396_),
    .ZN(_05753_)
  );
  INV_X1 _11272_ (
    .A(_05753_),
    .ZN(_05754_)
  );
  AND2_X1 _11273_ (
    .A1(_05752_),
    .A2(_05754_),
    .ZN(_05755_)
  );
  INV_X1 _11274_ (
    .A(_05755_),
    .ZN(_05756_)
  );
  AND2_X1 _11275_ (
    .A1(_00811_),
    .A2(_05756_),
    .ZN(_00604_)
  );
  AND2_X1 _11276_ (
    .A1(_00635_),
    .A2(_04346_),
    .ZN(_05757_)
  );
  INV_X1 _11277_ (
    .A(_05757_),
    .ZN(_05758_)
  );
  AND2_X1 _11278_ (
    .A1(large_[10]),
    .A2(_04345_),
    .ZN(_05759_)
  );
  INV_X1 _11279_ (
    .A(_05759_),
    .ZN(_05760_)
  );
  AND2_X1 _11280_ (
    .A1(_04394_),
    .A2(_05760_),
    .ZN(_05761_)
  );
  AND2_X1 _11281_ (
    .A1(_05758_),
    .A2(_05761_),
    .ZN(_05762_)
  );
  INV_X1 _11282_ (
    .A(_05762_),
    .ZN(_05763_)
  );
  AND2_X1 _11283_ (
    .A1(large_[10]),
    .A2(_04388_),
    .ZN(_05764_)
  );
  INV_X1 _11284_ (
    .A(_05764_),
    .ZN(_05765_)
  );
  AND2_X1 _11285_ (
    .A1(_05763_),
    .A2(_05765_),
    .ZN(_05766_)
  );
  AND2_X1 _11286_ (
    .A1(_01035_),
    .A2(_04396_),
    .ZN(_05767_)
  );
  INV_X1 _11287_ (
    .A(_05767_),
    .ZN(_05768_)
  );
  AND2_X1 _11288_ (
    .A1(_05766_),
    .A2(_05768_),
    .ZN(_05769_)
  );
  INV_X1 _11289_ (
    .A(_05769_),
    .ZN(_05770_)
  );
  AND2_X1 _11290_ (
    .A1(_00811_),
    .A2(_05770_),
    .ZN(_00605_)
  );
  AND2_X1 _11291_ (
    .A1(_04348_),
    .A2(_04398_),
    .ZN(_05771_)
  );
  INV_X1 _11292_ (
    .A(_05771_),
    .ZN(_05772_)
  );
  AND2_X1 _11293_ (
    .A1(_05759_),
    .A2(_05771_),
    .ZN(_05773_)
  );
  INV_X1 _11294_ (
    .A(_05773_),
    .ZN(_05774_)
  );
  AND2_X1 _11295_ (
    .A1(_02669_),
    .A2(_04396_),
    .ZN(_05775_)
  );
  INV_X1 _11296_ (
    .A(_05775_),
    .ZN(_05776_)
  );
  AND2_X1 _11297_ (
    .A1(_04389_),
    .A2(_05772_),
    .ZN(_05777_)
  );
  INV_X1 _11298_ (
    .A(_05777_),
    .ZN(_05778_)
  );
  AND2_X1 _11299_ (
    .A1(large_[11]),
    .A2(_05778_),
    .ZN(_05779_)
  );
  INV_X1 _11300_ (
    .A(_05779_),
    .ZN(_05780_)
  );
  AND2_X1 _11301_ (
    .A1(_05776_),
    .A2(_05780_),
    .ZN(_05781_)
  );
  AND2_X1 _11302_ (
    .A1(_05774_),
    .A2(_05781_),
    .ZN(_05782_)
  );
  INV_X1 _11303_ (
    .A(_05782_),
    .ZN(_05783_)
  );
  AND2_X1 _11304_ (
    .A1(_00811_),
    .A2(_05783_),
    .ZN(_00606_)
  );
  AND2_X1 _11305_ (
    .A1(_04347_),
    .A2(_04398_),
    .ZN(_05784_)
  );
  INV_X1 _11306_ (
    .A(_05784_),
    .ZN(_05785_)
  );
  MUX2_X1 _11307_ (
    .A(_05785_),
    .B(_05777_),
    .S(large_[12]),
    .Z(_05786_)
  );
  AND2_X1 _11308_ (
    .A1(_01107_),
    .A2(_04390_),
    .ZN(_05787_)
  );
  INV_X1 _11309_ (
    .A(_05787_),
    .ZN(_05788_)
  );
  AND2_X1 _11310_ (
    .A1(_05786_),
    .A2(_05788_),
    .ZN(_05789_)
  );
  INV_X1 _11311_ (
    .A(_05789_),
    .ZN(_05790_)
  );
  AND2_X1 _11312_ (
    .A1(_00811_),
    .A2(_05790_),
    .ZN(_00607_)
  );
  AND2_X1 _11313_ (
    .A1(_00634_),
    .A2(_04381_),
    .ZN(_05791_)
  );
  INV_X1 _11314_ (
    .A(_05791_),
    .ZN(_05792_)
  );
  AND2_X1 _11315_ (
    .A1(large_[13]),
    .A2(_04388_),
    .ZN(_05793_)
  );
  INV_X1 _11316_ (
    .A(_05793_),
    .ZN(_05794_)
  );
  AND2_X1 _11317_ (
    .A1(_04351_),
    .A2(_04398_),
    .ZN(_05795_)
  );
  AND2_X1 _11318_ (
    .A1(_05792_),
    .A2(_05795_),
    .ZN(_05796_)
  );
  INV_X1 _11319_ (
    .A(_05796_),
    .ZN(_05797_)
  );
  AND2_X1 _11320_ (
    .A1(_05794_),
    .A2(_05797_),
    .ZN(_05798_)
  );
  AND2_X1 _11321_ (
    .A1(_01199_),
    .A2(_04396_),
    .ZN(_05799_)
  );
  INV_X1 _11322_ (
    .A(_05799_),
    .ZN(_05800_)
  );
  AND2_X1 _11323_ (
    .A1(_05798_),
    .A2(_05800_),
    .ZN(_05801_)
  );
  INV_X1 _11324_ (
    .A(_05801_),
    .ZN(_05802_)
  );
  AND2_X1 _11325_ (
    .A1(_00811_),
    .A2(_05802_),
    .ZN(_00608_)
  );
  AND2_X1 _11326_ (
    .A1(_00633_),
    .A2(_04351_),
    .ZN(_05803_)
  );
  INV_X1 _11327_ (
    .A(_05803_),
    .ZN(_05804_)
  );
  AND2_X1 _11328_ (
    .A1(large_[14]),
    .A2(_04388_),
    .ZN(_05805_)
  );
  INV_X1 _11329_ (
    .A(_05805_),
    .ZN(_05806_)
  );
  AND2_X1 _11330_ (
    .A1(large_[14]),
    .A2(_04350_),
    .ZN(_05807_)
  );
  INV_X1 _11331_ (
    .A(_05807_),
    .ZN(_05808_)
  );
  AND2_X1 _11332_ (
    .A1(_04398_),
    .A2(_05808_),
    .ZN(_05809_)
  );
  AND2_X1 _11333_ (
    .A1(_05804_),
    .A2(_05809_),
    .ZN(_05810_)
  );
  INV_X1 _11334_ (
    .A(_05810_),
    .ZN(_05811_)
  );
  AND2_X1 _11335_ (
    .A1(_05806_),
    .A2(_05811_),
    .ZN(_05812_)
  );
  AND2_X1 _11336_ (
    .A1(_01277_),
    .A2(_04390_),
    .ZN(_05813_)
  );
  INV_X1 _11337_ (
    .A(_05813_),
    .ZN(_05814_)
  );
  AND2_X1 _11338_ (
    .A1(_05812_),
    .A2(_05814_),
    .ZN(_05815_)
  );
  INV_X1 _11339_ (
    .A(_05815_),
    .ZN(_05816_)
  );
  AND2_X1 _11340_ (
    .A1(_00811_),
    .A2(_05816_),
    .ZN(_00609_)
  );
  AND2_X1 _11341_ (
    .A1(_00632_),
    .A2(_05808_),
    .ZN(_05817_)
  );
  INV_X1 _11342_ (
    .A(_05817_),
    .ZN(_05818_)
  );
  AND2_X1 _11343_ (
    .A1(large_[15]),
    .A2(_04388_),
    .ZN(_05819_)
  );
  INV_X1 _11344_ (
    .A(_05819_),
    .ZN(_05820_)
  );
  AND2_X1 _11345_ (
    .A1(large_[15]),
    .A2(_05807_),
    .ZN(_05821_)
  );
  INV_X1 _11346_ (
    .A(_05821_),
    .ZN(_05822_)
  );
  AND2_X1 _11347_ (
    .A1(_04398_),
    .A2(_05818_),
    .ZN(_05823_)
  );
  AND2_X1 _11348_ (
    .A1(_05822_),
    .A2(_05823_),
    .ZN(_05824_)
  );
  INV_X1 _11349_ (
    .A(_05824_),
    .ZN(_05825_)
  );
  AND2_X1 _11350_ (
    .A1(_05820_),
    .A2(_05825_),
    .ZN(_05826_)
  );
  AND2_X1 _11351_ (
    .A1(_02735_),
    .A2(_04390_),
    .ZN(_05827_)
  );
  INV_X1 _11352_ (
    .A(_05827_),
    .ZN(_05828_)
  );
  AND2_X1 _11353_ (
    .A1(_05826_),
    .A2(_05828_),
    .ZN(_05829_)
  );
  INV_X1 _11354_ (
    .A(_05829_),
    .ZN(_05830_)
  );
  AND2_X1 _11355_ (
    .A1(_00811_),
    .A2(_05830_),
    .ZN(_00610_)
  );
  AND2_X1 _11356_ (
    .A1(_00631_),
    .A2(_05822_),
    .ZN(_05831_)
  );
  INV_X1 _11357_ (
    .A(_05831_),
    .ZN(_05832_)
  );
  AND2_X1 _11358_ (
    .A1(large_[16]),
    .A2(_05821_),
    .ZN(_05833_)
  );
  INV_X1 _11359_ (
    .A(_05833_),
    .ZN(_05834_)
  );
  AND2_X1 _11360_ (
    .A1(_04398_),
    .A2(_05834_),
    .ZN(_05835_)
  );
  AND2_X1 _11361_ (
    .A1(_05832_),
    .A2(_05835_),
    .ZN(_05836_)
  );
  INV_X1 _11362_ (
    .A(_05836_),
    .ZN(_05837_)
  );
  AND2_X1 _11363_ (
    .A1(large_[16]),
    .A2(_04388_),
    .ZN(_05838_)
  );
  INV_X1 _11364_ (
    .A(_05838_),
    .ZN(_05839_)
  );
  AND2_X1 _11365_ (
    .A1(_02801_),
    .A2(_04396_),
    .ZN(_05840_)
  );
  INV_X1 _11366_ (
    .A(_05840_),
    .ZN(_05841_)
  );
  AND2_X1 _11367_ (
    .A1(_05837_),
    .A2(_05839_),
    .ZN(_05842_)
  );
  AND2_X1 _11368_ (
    .A1(_05841_),
    .A2(_05842_),
    .ZN(_05843_)
  );
  INV_X1 _11369_ (
    .A(_05843_),
    .ZN(_05844_)
  );
  AND2_X1 _11370_ (
    .A1(_00811_),
    .A2(_05844_),
    .ZN(_00611_)
  );
  AND2_X1 _11371_ (
    .A1(_00630_),
    .A2(_05834_),
    .ZN(_05845_)
  );
  INV_X1 _11372_ (
    .A(_05845_),
    .ZN(_05846_)
  );
  AND2_X1 _11373_ (
    .A1(large_[17]),
    .A2(_05833_),
    .ZN(_05847_)
  );
  INV_X1 _11374_ (
    .A(_05847_),
    .ZN(_05848_)
  );
  AND2_X1 _11375_ (
    .A1(_04398_),
    .A2(_05846_),
    .ZN(_05849_)
  );
  AND2_X1 _11376_ (
    .A1(_05848_),
    .A2(_05849_),
    .ZN(_05850_)
  );
  INV_X1 _11377_ (
    .A(_05850_),
    .ZN(_05851_)
  );
  AND2_X1 _11378_ (
    .A1(large_[17]),
    .A2(_04388_),
    .ZN(_05852_)
  );
  INV_X1 _11379_ (
    .A(_05852_),
    .ZN(_05853_)
  );
  AND2_X1 _11380_ (
    .A1(_01360_),
    .A2(_04396_),
    .ZN(_05854_)
  );
  INV_X1 _11381_ (
    .A(_05854_),
    .ZN(_05855_)
  );
  AND2_X1 _11382_ (
    .A1(_05851_),
    .A2(_05853_),
    .ZN(_05856_)
  );
  AND2_X1 _11383_ (
    .A1(_05855_),
    .A2(_05856_),
    .ZN(_05857_)
  );
  INV_X1 _11384_ (
    .A(_05857_),
    .ZN(_05858_)
  );
  AND2_X1 _11385_ (
    .A1(_00811_),
    .A2(_05858_),
    .ZN(_00612_)
  );
  AND2_X1 _11386_ (
    .A1(_00629_),
    .A2(_05848_),
    .ZN(_05859_)
  );
  INV_X1 _11387_ (
    .A(_05859_),
    .ZN(_05860_)
  );
  AND2_X1 _11388_ (
    .A1(large_[18]),
    .A2(_05847_),
    .ZN(_05861_)
  );
  INV_X1 _11389_ (
    .A(_05861_),
    .ZN(_05862_)
  );
  AND2_X1 _11390_ (
    .A1(_04398_),
    .A2(_05862_),
    .ZN(_05863_)
  );
  AND2_X1 _11391_ (
    .A1(_05860_),
    .A2(_05863_),
    .ZN(_05864_)
  );
  INV_X1 _11392_ (
    .A(_05864_),
    .ZN(_05865_)
  );
  AND2_X1 _11393_ (
    .A1(large_[18]),
    .A2(_04388_),
    .ZN(_05866_)
  );
  INV_X1 _11394_ (
    .A(_05866_),
    .ZN(_05867_)
  );
  AND2_X1 _11395_ (
    .A1(_02873_),
    .A2(_04390_),
    .ZN(_05868_)
  );
  INV_X1 _11396_ (
    .A(_05868_),
    .ZN(_05869_)
  );
  AND2_X1 _11397_ (
    .A1(_05867_),
    .A2(_05869_),
    .ZN(_05870_)
  );
  AND2_X1 _11398_ (
    .A1(_05865_),
    .A2(_05870_),
    .ZN(_05871_)
  );
  INV_X1 _11399_ (
    .A(_05871_),
    .ZN(_05872_)
  );
  AND2_X1 _11400_ (
    .A1(_00811_),
    .A2(_05872_),
    .ZN(_00613_)
  );
  AND2_X1 _11401_ (
    .A1(_00628_),
    .A2(_05862_),
    .ZN(_05873_)
  );
  INV_X1 _11402_ (
    .A(_05873_),
    .ZN(_05874_)
  );
  AND2_X1 _11403_ (
    .A1(_04353_),
    .A2(_04394_),
    .ZN(_05875_)
  );
  AND2_X1 _11404_ (
    .A1(_05874_),
    .A2(_05875_),
    .ZN(_05876_)
  );
  INV_X1 _11405_ (
    .A(_05876_),
    .ZN(_05877_)
  );
  AND2_X1 _11406_ (
    .A1(large_[19]),
    .A2(_04388_),
    .ZN(_05878_)
  );
  INV_X1 _11407_ (
    .A(_05878_),
    .ZN(_05879_)
  );
  AND2_X1 _11408_ (
    .A1(_02945_),
    .A2(_04396_),
    .ZN(_05880_)
  );
  INV_X1 _11409_ (
    .A(_05880_),
    .ZN(_05881_)
  );
  AND2_X1 _11410_ (
    .A1(_05879_),
    .A2(_05881_),
    .ZN(_05882_)
  );
  AND2_X1 _11411_ (
    .A1(_05877_),
    .A2(_05882_),
    .ZN(_05883_)
  );
  INV_X1 _11412_ (
    .A(_05883_),
    .ZN(_05884_)
  );
  AND2_X1 _11413_ (
    .A1(_00811_),
    .A2(_05884_),
    .ZN(_00614_)
  );
  AND2_X1 _11414_ (
    .A1(_00627_),
    .A2(_04353_),
    .ZN(_05885_)
  );
  INV_X1 _11415_ (
    .A(_05885_),
    .ZN(_05886_)
  );
  AND2_X1 _11416_ (
    .A1(_04355_),
    .A2(_04394_),
    .ZN(_05887_)
  );
  AND2_X1 _11417_ (
    .A1(_05886_),
    .A2(_05887_),
    .ZN(_05888_)
  );
  INV_X1 _11418_ (
    .A(_05888_),
    .ZN(_05889_)
  );
  AND2_X1 _11419_ (
    .A1(large_[20]),
    .A2(_04388_),
    .ZN(_05890_)
  );
  INV_X1 _11420_ (
    .A(_05890_),
    .ZN(_05891_)
  );
  AND2_X1 _11421_ (
    .A1(_03017_),
    .A2(_04396_),
    .ZN(_05892_)
  );
  INV_X1 _11422_ (
    .A(_05892_),
    .ZN(_05893_)
  );
  AND2_X1 _11423_ (
    .A1(_05889_),
    .A2(_05893_),
    .ZN(_05894_)
  );
  AND2_X1 _11424_ (
    .A1(_05891_),
    .A2(_05894_),
    .ZN(_05895_)
  );
  INV_X1 _11425_ (
    .A(_05895_),
    .ZN(_05896_)
  );
  AND2_X1 _11426_ (
    .A1(_00811_),
    .A2(_05896_),
    .ZN(_00615_)
  );
  AND2_X1 _11427_ (
    .A1(_00626_),
    .A2(_04355_),
    .ZN(_05897_)
  );
  INV_X1 _11428_ (
    .A(_05897_),
    .ZN(_05898_)
  );
  AND2_X1 _11429_ (
    .A1(_04357_),
    .A2(_04394_),
    .ZN(_05899_)
  );
  AND2_X1 _11430_ (
    .A1(_05898_),
    .A2(_05899_),
    .ZN(_05900_)
  );
  INV_X1 _11431_ (
    .A(_05900_),
    .ZN(_05901_)
  );
  AND2_X1 _11432_ (
    .A1(large_[21]),
    .A2(_04388_),
    .ZN(_05902_)
  );
  INV_X1 _11433_ (
    .A(_05902_),
    .ZN(_05903_)
  );
  AND2_X1 _11434_ (
    .A1(_03089_),
    .A2(_04396_),
    .ZN(_05904_)
  );
  INV_X1 _11435_ (
    .A(_05904_),
    .ZN(_05905_)
  );
  AND2_X1 _11436_ (
    .A1(_05901_),
    .A2(_05903_),
    .ZN(_05906_)
  );
  AND2_X1 _11437_ (
    .A1(_05905_),
    .A2(_05906_),
    .ZN(_05907_)
  );
  INV_X1 _11438_ (
    .A(_05907_),
    .ZN(_05908_)
  );
  AND2_X1 _11439_ (
    .A1(_00811_),
    .A2(_05908_),
    .ZN(_00616_)
  );
  AND2_X1 _11440_ (
    .A1(_00625_),
    .A2(_04357_),
    .ZN(_05909_)
  );
  INV_X1 _11441_ (
    .A(_05909_),
    .ZN(_05910_)
  );
  AND2_X1 _11442_ (
    .A1(_04359_),
    .A2(_04394_),
    .ZN(_05911_)
  );
  AND2_X1 _11443_ (
    .A1(_05910_),
    .A2(_05911_),
    .ZN(_05912_)
  );
  INV_X1 _11444_ (
    .A(_05912_),
    .ZN(_05913_)
  );
  AND2_X1 _11445_ (
    .A1(large_[22]),
    .A2(_04388_),
    .ZN(_05914_)
  );
  INV_X1 _11446_ (
    .A(_05914_),
    .ZN(_05915_)
  );
  AND2_X1 _11447_ (
    .A1(_03162_),
    .A2(_04396_),
    .ZN(_05916_)
  );
  INV_X1 _11448_ (
    .A(_05916_),
    .ZN(_05917_)
  );
  AND2_X1 _11449_ (
    .A1(_05913_),
    .A2(_05917_),
    .ZN(_05918_)
  );
  AND2_X1 _11450_ (
    .A1(_05915_),
    .A2(_05918_),
    .ZN(_05919_)
  );
  INV_X1 _11451_ (
    .A(_05919_),
    .ZN(_05920_)
  );
  AND2_X1 _11452_ (
    .A1(_00811_),
    .A2(_05920_),
    .ZN(_00617_)
  );
  AND2_X1 _11453_ (
    .A1(_00624_),
    .A2(_04359_),
    .ZN(_05921_)
  );
  INV_X1 _11454_ (
    .A(_05921_),
    .ZN(_05922_)
  );
  AND2_X1 _11455_ (
    .A1(_04361_),
    .A2(_04394_),
    .ZN(_05923_)
  );
  AND2_X1 _11456_ (
    .A1(_05922_),
    .A2(_05923_),
    .ZN(_05924_)
  );
  INV_X1 _11457_ (
    .A(_05924_),
    .ZN(_05925_)
  );
  AND2_X1 _11458_ (
    .A1(large_[23]),
    .A2(_04388_),
    .ZN(_05926_)
  );
  INV_X1 _11459_ (
    .A(_05926_),
    .ZN(_05927_)
  );
  AND2_X1 _11460_ (
    .A1(_03230_),
    .A2(_04396_),
    .ZN(_05928_)
  );
  INV_X1 _11461_ (
    .A(_05928_),
    .ZN(_05929_)
  );
  AND2_X1 _11462_ (
    .A1(_05927_),
    .A2(_05929_),
    .ZN(_05930_)
  );
  AND2_X1 _11463_ (
    .A1(_05925_),
    .A2(_05930_),
    .ZN(_05931_)
  );
  INV_X1 _11464_ (
    .A(_05931_),
    .ZN(_05932_)
  );
  AND2_X1 _11465_ (
    .A1(_00811_),
    .A2(_05932_),
    .ZN(_00618_)
  );
  AND2_X1 _11466_ (
    .A1(_00623_),
    .A2(_04361_),
    .ZN(_05933_)
  );
  INV_X1 _11467_ (
    .A(_05933_),
    .ZN(_05934_)
  );
  AND2_X1 _11468_ (
    .A1(_04363_),
    .A2(_04394_),
    .ZN(_05935_)
  );
  AND2_X1 _11469_ (
    .A1(_05934_),
    .A2(_05935_),
    .ZN(_05936_)
  );
  INV_X1 _11470_ (
    .A(_05936_),
    .ZN(_05937_)
  );
  AND2_X1 _11471_ (
    .A1(large_[24]),
    .A2(_04388_),
    .ZN(_05938_)
  );
  INV_X1 _11472_ (
    .A(_05938_),
    .ZN(_05939_)
  );
  AND2_X1 _11473_ (
    .A1(_03443_),
    .A2(_04390_),
    .ZN(_05940_)
  );
  INV_X1 _11474_ (
    .A(_05940_),
    .ZN(_05941_)
  );
  AND2_X1 _11475_ (
    .A1(_05939_),
    .A2(_05941_),
    .ZN(_05942_)
  );
  AND2_X1 _11476_ (
    .A1(_05937_),
    .A2(_05942_),
    .ZN(_05943_)
  );
  INV_X1 _11477_ (
    .A(_05943_),
    .ZN(_05944_)
  );
  AND2_X1 _11478_ (
    .A1(_00811_),
    .A2(_05944_),
    .ZN(_00619_)
  );
  AND2_X1 _11479_ (
    .A1(_00622_),
    .A2(_04363_),
    .ZN(_05945_)
  );
  INV_X1 _11480_ (
    .A(_05945_),
    .ZN(_05946_)
  );
  AND2_X1 _11481_ (
    .A1(_04365_),
    .A2(_04394_),
    .ZN(_05947_)
  );
  AND2_X1 _11482_ (
    .A1(_05946_),
    .A2(_05947_),
    .ZN(_05948_)
  );
  INV_X1 _11483_ (
    .A(_05948_),
    .ZN(_05949_)
  );
  AND2_X1 _11484_ (
    .A1(large_[25]),
    .A2(_04388_),
    .ZN(_05950_)
  );
  INV_X1 _11485_ (
    .A(_05950_),
    .ZN(_05951_)
  );
  AND2_X1 _11486_ (
    .A1(_03342_),
    .A2(_04390_),
    .ZN(_05952_)
  );
  INV_X1 _11487_ (
    .A(_05952_),
    .ZN(_05953_)
  );
  AND2_X1 _11488_ (
    .A1(_05951_),
    .A2(_05953_),
    .ZN(_05954_)
  );
  AND2_X1 _11489_ (
    .A1(_05949_),
    .A2(_05954_),
    .ZN(_05955_)
  );
  INV_X1 _11490_ (
    .A(_05955_),
    .ZN(_05956_)
  );
  AND2_X1 _11491_ (
    .A1(_00811_),
    .A2(_05956_),
    .ZN(_00620_)
  );
  MUX2_X1 _11492_ (
    .A(reg_pmp_6_cfg_w),
    .B(_03281_),
    .S(_00900_),
    .Z(_00621_)
  );
  AND2_X1 _11493_ (
    .A1(io_decode_0_inst[31]),
    .A2(io_decode_0_inst[30]),
    .ZN(io_decode_0_write_illegal)
  );
  AND2_X1 _11494_ (
    .A1(_00897_),
    .A2(_00912_),
    .ZN(_05957_)
  );
  AND2_X1 _11495_ (
    .A1(_00870_),
    .A2(io_trace_0_exception),
    .ZN(_05958_)
  );
  AND2_X1 _11496_ (
    .A1(_03534_),
    .A2(_05958_),
    .ZN(_05959_)
  );
  MUX2_X1 _11497_ (
    .A(reg_dpc[1]),
    .B(io_pc[1]),
    .S(_05959_),
    .Z(_05960_)
  );
  MUX2_X1 _11498_ (
    .A(_05960_),
    .B(_01688_),
    .S(_05957_),
    .Z(_00000_[1])
  );
  MUX2_X1 _11499_ (
    .A(reg_dpc[2]),
    .B(io_pc[2]),
    .S(_05959_),
    .Z(_05961_)
  );
  MUX2_X1 _11500_ (
    .A(_05961_),
    .B(_01774_),
    .S(_05957_),
    .Z(_00000_[2])
  );
  MUX2_X1 _11501_ (
    .A(reg_dpc[3]),
    .B(io_pc[3]),
    .S(_05959_),
    .Z(_05962_)
  );
  MUX2_X1 _11502_ (
    .A(_05962_),
    .B(_01865_),
    .S(_05957_),
    .Z(_00000_[3])
  );
  MUX2_X1 _11503_ (
    .A(reg_dpc[4]),
    .B(io_pc[4]),
    .S(_05959_),
    .Z(_05963_)
  );
  MUX2_X1 _11504_ (
    .A(_05963_),
    .B(_01938_),
    .S(_05957_),
    .Z(_00000_[4])
  );
  MUX2_X1 _11505_ (
    .A(reg_dpc[5]),
    .B(io_pc[5]),
    .S(_05959_),
    .Z(_05964_)
  );
  MUX2_X1 _11506_ (
    .A(_05964_),
    .B(_02005_),
    .S(_05957_),
    .Z(_00000_[5])
  );
  MUX2_X1 _11507_ (
    .A(reg_dpc[6]),
    .B(io_pc[6]),
    .S(_05959_),
    .Z(_05965_)
  );
  MUX2_X1 _11508_ (
    .A(_05965_),
    .B(_02076_),
    .S(_05957_),
    .Z(_00000_[6])
  );
  MUX2_X1 _11509_ (
    .A(reg_dpc[7]),
    .B(io_pc[7]),
    .S(_05959_),
    .Z(_05966_)
  );
  MUX2_X1 _11510_ (
    .A(_05966_),
    .B(_02163_),
    .S(_05957_),
    .Z(_00000_[7])
  );
  MUX2_X1 _11511_ (
    .A(reg_dpc[8]),
    .B(io_pc[8]),
    .S(_05959_),
    .Z(_05967_)
  );
  MUX2_X1 _11512_ (
    .A(_05967_),
    .B(_01446_),
    .S(_05957_),
    .Z(_00000_[8])
  );
  MUX2_X1 _11513_ (
    .A(reg_dpc[9]),
    .B(io_pc[9]),
    .S(_05959_),
    .Z(_05968_)
  );
  MUX2_X1 _11514_ (
    .A(_05968_),
    .B(_01518_),
    .S(_05957_),
    .Z(_00000_[9])
  );
  MUX2_X1 _11515_ (
    .A(reg_dpc[10]),
    .B(io_pc[10]),
    .S(_05959_),
    .Z(_05969_)
  );
  MUX2_X1 _11516_ (
    .A(_05969_),
    .B(_02235_),
    .S(_05957_),
    .Z(_00000_[10])
  );
  MUX2_X1 _11517_ (
    .A(reg_dpc[11]),
    .B(io_pc[11]),
    .S(_05959_),
    .Z(_05970_)
  );
  MUX2_X1 _11518_ (
    .A(_05970_),
    .B(_02314_),
    .S(_05957_),
    .Z(_00000_[11])
  );
  MUX2_X1 _11519_ (
    .A(reg_dpc[12]),
    .B(io_pc[12]),
    .S(_05959_),
    .Z(_05971_)
  );
  MUX2_X1 _11520_ (
    .A(_05971_),
    .B(_02389_),
    .S(_05957_),
    .Z(_00000_[12])
  );
  MUX2_X1 _11521_ (
    .A(reg_dpc[13]),
    .B(io_pc[13]),
    .S(_05959_),
    .Z(_05972_)
  );
  MUX2_X1 _11522_ (
    .A(_05972_),
    .B(_02456_),
    .S(_05957_),
    .Z(_00000_[13])
  );
  MUX2_X1 _11523_ (
    .A(reg_dpc[14]),
    .B(io_pc[14]),
    .S(_05959_),
    .Z(_05973_)
  );
  MUX2_X1 _11524_ (
    .A(_05973_),
    .B(_02522_),
    .S(_05957_),
    .Z(_00000_[14])
  );
  MUX2_X1 _11525_ (
    .A(reg_dpc[15]),
    .B(io_pc[15]),
    .S(_05959_),
    .Z(_05974_)
  );
  MUX2_X1 _11526_ (
    .A(_05974_),
    .B(_02597_),
    .S(_05957_),
    .Z(_00000_[15])
  );
  MUX2_X1 _11527_ (
    .A(reg_dpc[16]),
    .B(io_pc[16]),
    .S(_05959_),
    .Z(_05975_)
  );
  MUX2_X1 _11528_ (
    .A(_05975_),
    .B(_01035_),
    .S(_05957_),
    .Z(_00000_[16])
  );
  MUX2_X1 _11529_ (
    .A(reg_dpc[17]),
    .B(io_pc[17]),
    .S(_05959_),
    .Z(_05976_)
  );
  MUX2_X1 _11530_ (
    .A(_05976_),
    .B(_02669_),
    .S(_05957_),
    .Z(_00000_[17])
  );
  MUX2_X1 _11531_ (
    .A(reg_dpc[18]),
    .B(io_pc[18]),
    .S(_05959_),
    .Z(_05977_)
  );
  MUX2_X1 _11532_ (
    .A(_05977_),
    .B(_01107_),
    .S(_05957_),
    .Z(_00000_[18])
  );
  MUX2_X1 _11533_ (
    .A(reg_dpc[19]),
    .B(io_pc[19]),
    .S(_05959_),
    .Z(_05978_)
  );
  MUX2_X1 _11534_ (
    .A(_05978_),
    .B(_01199_),
    .S(_05957_),
    .Z(_00000_[19])
  );
  MUX2_X1 _11535_ (
    .A(reg_dpc[20]),
    .B(io_pc[20]),
    .S(_05959_),
    .Z(_05979_)
  );
  MUX2_X1 _11536_ (
    .A(_05979_),
    .B(_01277_),
    .S(_05957_),
    .Z(_00000_[20])
  );
  MUX2_X1 _11537_ (
    .A(reg_dpc[21]),
    .B(io_pc[21]),
    .S(_05959_),
    .Z(_05980_)
  );
  MUX2_X1 _11538_ (
    .A(_05980_),
    .B(_02735_),
    .S(_05957_),
    .Z(_00000_[21])
  );
  MUX2_X1 _11539_ (
    .A(reg_dpc[22]),
    .B(io_pc[22]),
    .S(_05959_),
    .Z(_05981_)
  );
  MUX2_X1 _11540_ (
    .A(_05981_),
    .B(_02801_),
    .S(_05957_),
    .Z(_00000_[22])
  );
  MUX2_X1 _11541_ (
    .A(reg_dpc[23]),
    .B(io_pc[23]),
    .S(_05959_),
    .Z(_05982_)
  );
  MUX2_X1 _11542_ (
    .A(_05982_),
    .B(_01360_),
    .S(_05957_),
    .Z(_00000_[23])
  );
  MUX2_X1 _11543_ (
    .A(reg_dpc[24]),
    .B(io_pc[24]),
    .S(_05959_),
    .Z(_05983_)
  );
  MUX2_X1 _11544_ (
    .A(_05983_),
    .B(_02873_),
    .S(_05957_),
    .Z(_00000_[24])
  );
  MUX2_X1 _11545_ (
    .A(reg_dpc[25]),
    .B(io_pc[25]),
    .S(_05959_),
    .Z(_05984_)
  );
  MUX2_X1 _11546_ (
    .A(_05984_),
    .B(_02945_),
    .S(_05957_),
    .Z(_00000_[25])
  );
  MUX2_X1 _11547_ (
    .A(reg_dpc[26]),
    .B(io_pc[26]),
    .S(_05959_),
    .Z(_05985_)
  );
  MUX2_X1 _11548_ (
    .A(_05985_),
    .B(_03017_),
    .S(_05957_),
    .Z(_00000_[26])
  );
  MUX2_X1 _11549_ (
    .A(reg_dpc[27]),
    .B(io_pc[27]),
    .S(_05959_),
    .Z(_05986_)
  );
  MUX2_X1 _11550_ (
    .A(_05986_),
    .B(_03089_),
    .S(_05957_),
    .Z(_00000_[27])
  );
  MUX2_X1 _11551_ (
    .A(reg_dpc[28]),
    .B(io_pc[28]),
    .S(_05959_),
    .Z(_05987_)
  );
  MUX2_X1 _11552_ (
    .A(_05987_),
    .B(_03162_),
    .S(_05957_),
    .Z(_00000_[28])
  );
  MUX2_X1 _11553_ (
    .A(reg_dpc[29]),
    .B(io_pc[29]),
    .S(_05959_),
    .Z(_05988_)
  );
  MUX2_X1 _11554_ (
    .A(_05988_),
    .B(_03230_),
    .S(_05957_),
    .Z(_00000_[29])
  );
  MUX2_X1 _11555_ (
    .A(reg_dpc[30]),
    .B(io_pc[30]),
    .S(_05959_),
    .Z(_05989_)
  );
  MUX2_X1 _11556_ (
    .A(_05989_),
    .B(_03443_),
    .S(_05957_),
    .Z(_00000_[30])
  );
  MUX2_X1 _11557_ (
    .A(reg_dpc[31]),
    .B(io_pc[31]),
    .S(_05959_),
    .Z(_05990_)
  );
  MUX2_X1 _11558_ (
    .A(_05990_),
    .B(_03342_),
    .S(_05957_),
    .Z(_00000_[31])
  );
  AND2_X1 _11559_ (
    .A1(_00897_),
    .A2(_00943_),
    .ZN(_05991_)
  );
  MUX2_X1 _11560_ (
    .A(reg_mepc[1]),
    .B(io_pc[1]),
    .S(_03535_),
    .Z(_05992_)
  );
  MUX2_X1 _11561_ (
    .A(_05992_),
    .B(_01688_),
    .S(_05991_),
    .Z(_00001_[1])
  );
  MUX2_X1 _11562_ (
    .A(reg_mepc[2]),
    .B(io_pc[2]),
    .S(_03535_),
    .Z(_05993_)
  );
  MUX2_X1 _11563_ (
    .A(_05993_),
    .B(_01774_),
    .S(_05991_),
    .Z(_00001_[2])
  );
  MUX2_X1 _11564_ (
    .A(reg_mepc[3]),
    .B(io_pc[3]),
    .S(_03535_),
    .Z(_05994_)
  );
  MUX2_X1 _11565_ (
    .A(_05994_),
    .B(_01865_),
    .S(_05991_),
    .Z(_00001_[3])
  );
  MUX2_X1 _11566_ (
    .A(reg_mepc[4]),
    .B(io_pc[4]),
    .S(_03535_),
    .Z(_05995_)
  );
  MUX2_X1 _11567_ (
    .A(_05995_),
    .B(_01938_),
    .S(_05991_),
    .Z(_00001_[4])
  );
  MUX2_X1 _11568_ (
    .A(reg_mepc[5]),
    .B(io_pc[5]),
    .S(_03535_),
    .Z(_05996_)
  );
  MUX2_X1 _11569_ (
    .A(_05996_),
    .B(_02005_),
    .S(_05991_),
    .Z(_00001_[5])
  );
  MUX2_X1 _11570_ (
    .A(reg_mepc[6]),
    .B(io_pc[6]),
    .S(_03535_),
    .Z(_05997_)
  );
  MUX2_X1 _11571_ (
    .A(_05997_),
    .B(_02076_),
    .S(_05991_),
    .Z(_00001_[6])
  );
  MUX2_X1 _11572_ (
    .A(reg_mepc[7]),
    .B(io_pc[7]),
    .S(_03535_),
    .Z(_05998_)
  );
  MUX2_X1 _11573_ (
    .A(_05998_),
    .B(_02163_),
    .S(_05991_),
    .Z(_00001_[7])
  );
  MUX2_X1 _11574_ (
    .A(reg_mepc[8]),
    .B(io_pc[8]),
    .S(_03535_),
    .Z(_05999_)
  );
  MUX2_X1 _11575_ (
    .A(_05999_),
    .B(_01446_),
    .S(_05991_),
    .Z(_00001_[8])
  );
  MUX2_X1 _11576_ (
    .A(reg_mepc[9]),
    .B(io_pc[9]),
    .S(_03535_),
    .Z(_06000_)
  );
  MUX2_X1 _11577_ (
    .A(_06000_),
    .B(_01518_),
    .S(_05991_),
    .Z(_00001_[9])
  );
  MUX2_X1 _11578_ (
    .A(reg_mepc[10]),
    .B(io_pc[10]),
    .S(_03535_),
    .Z(_06001_)
  );
  MUX2_X1 _11579_ (
    .A(_06001_),
    .B(_02235_),
    .S(_05991_),
    .Z(_00001_[10])
  );
  MUX2_X1 _11580_ (
    .A(reg_mepc[11]),
    .B(io_pc[11]),
    .S(_03535_),
    .Z(_06002_)
  );
  MUX2_X1 _11581_ (
    .A(_06002_),
    .B(_02314_),
    .S(_05991_),
    .Z(_00001_[11])
  );
  MUX2_X1 _11582_ (
    .A(reg_mepc[12]),
    .B(io_pc[12]),
    .S(_03535_),
    .Z(_06003_)
  );
  MUX2_X1 _11583_ (
    .A(_06003_),
    .B(_02389_),
    .S(_05991_),
    .Z(_00001_[12])
  );
  MUX2_X1 _11584_ (
    .A(reg_mepc[13]),
    .B(io_pc[13]),
    .S(_03535_),
    .Z(_06004_)
  );
  MUX2_X1 _11585_ (
    .A(_06004_),
    .B(_02456_),
    .S(_05991_),
    .Z(_00001_[13])
  );
  MUX2_X1 _11586_ (
    .A(reg_mepc[14]),
    .B(io_pc[14]),
    .S(_03535_),
    .Z(_06005_)
  );
  MUX2_X1 _11587_ (
    .A(_06005_),
    .B(_02522_),
    .S(_05991_),
    .Z(_00001_[14])
  );
  MUX2_X1 _11588_ (
    .A(reg_mepc[15]),
    .B(io_pc[15]),
    .S(_03535_),
    .Z(_06006_)
  );
  MUX2_X1 _11589_ (
    .A(_06006_),
    .B(_02597_),
    .S(_05991_),
    .Z(_00001_[15])
  );
  MUX2_X1 _11590_ (
    .A(reg_mepc[16]),
    .B(io_pc[16]),
    .S(_03535_),
    .Z(_06007_)
  );
  MUX2_X1 _11591_ (
    .A(_06007_),
    .B(_01035_),
    .S(_05991_),
    .Z(_00001_[16])
  );
  MUX2_X1 _11592_ (
    .A(reg_mepc[17]),
    .B(io_pc[17]),
    .S(_03535_),
    .Z(_06008_)
  );
  MUX2_X1 _11593_ (
    .A(_06008_),
    .B(_02669_),
    .S(_05991_),
    .Z(_00001_[17])
  );
  MUX2_X1 _11594_ (
    .A(reg_mepc[18]),
    .B(io_pc[18]),
    .S(_03535_),
    .Z(_06009_)
  );
  MUX2_X1 _11595_ (
    .A(_06009_),
    .B(_01107_),
    .S(_05991_),
    .Z(_00001_[18])
  );
  MUX2_X1 _11596_ (
    .A(reg_mepc[19]),
    .B(io_pc[19]),
    .S(_03535_),
    .Z(_06010_)
  );
  MUX2_X1 _11597_ (
    .A(_06010_),
    .B(_01199_),
    .S(_05991_),
    .Z(_00001_[19])
  );
  MUX2_X1 _11598_ (
    .A(reg_mepc[20]),
    .B(io_pc[20]),
    .S(_03535_),
    .Z(_06011_)
  );
  MUX2_X1 _11599_ (
    .A(_06011_),
    .B(_01277_),
    .S(_05991_),
    .Z(_00001_[20])
  );
  MUX2_X1 _11600_ (
    .A(reg_mepc[21]),
    .B(io_pc[21]),
    .S(_03535_),
    .Z(_06012_)
  );
  MUX2_X1 _11601_ (
    .A(_06012_),
    .B(_02735_),
    .S(_05991_),
    .Z(_00001_[21])
  );
  MUX2_X1 _11602_ (
    .A(reg_mepc[22]),
    .B(io_pc[22]),
    .S(_03535_),
    .Z(_06013_)
  );
  MUX2_X1 _11603_ (
    .A(_06013_),
    .B(_02801_),
    .S(_05991_),
    .Z(_00001_[22])
  );
  MUX2_X1 _11604_ (
    .A(reg_mepc[23]),
    .B(io_pc[23]),
    .S(_03535_),
    .Z(_06014_)
  );
  MUX2_X1 _11605_ (
    .A(_06014_),
    .B(_01360_),
    .S(_05991_),
    .Z(_00001_[23])
  );
  MUX2_X1 _11606_ (
    .A(reg_mepc[24]),
    .B(io_pc[24]),
    .S(_03535_),
    .Z(_06015_)
  );
  MUX2_X1 _11607_ (
    .A(_06015_),
    .B(_02873_),
    .S(_05991_),
    .Z(_00001_[24])
  );
  MUX2_X1 _11608_ (
    .A(reg_mepc[25]),
    .B(io_pc[25]),
    .S(_03535_),
    .Z(_06016_)
  );
  MUX2_X1 _11609_ (
    .A(_06016_),
    .B(_02945_),
    .S(_05991_),
    .Z(_00001_[25])
  );
  MUX2_X1 _11610_ (
    .A(reg_mepc[26]),
    .B(io_pc[26]),
    .S(_03535_),
    .Z(_06017_)
  );
  MUX2_X1 _11611_ (
    .A(_06017_),
    .B(_03017_),
    .S(_05991_),
    .Z(_00001_[26])
  );
  MUX2_X1 _11612_ (
    .A(reg_mepc[27]),
    .B(io_pc[27]),
    .S(_03535_),
    .Z(_06018_)
  );
  MUX2_X1 _11613_ (
    .A(_06018_),
    .B(_03089_),
    .S(_05991_),
    .Z(_00001_[27])
  );
  MUX2_X1 _11614_ (
    .A(reg_mepc[28]),
    .B(io_pc[28]),
    .S(_03535_),
    .Z(_06019_)
  );
  MUX2_X1 _11615_ (
    .A(_06019_),
    .B(_03162_),
    .S(_05991_),
    .Z(_00001_[28])
  );
  MUX2_X1 _11616_ (
    .A(reg_mepc[29]),
    .B(io_pc[29]),
    .S(_03535_),
    .Z(_06020_)
  );
  MUX2_X1 _11617_ (
    .A(_06020_),
    .B(_03230_),
    .S(_05991_),
    .Z(_00001_[29])
  );
  MUX2_X1 _11618_ (
    .A(reg_mepc[30]),
    .B(io_pc[30]),
    .S(_03535_),
    .Z(_06021_)
  );
  MUX2_X1 _11619_ (
    .A(_06021_),
    .B(_03443_),
    .S(_05991_),
    .Z(_00001_[30])
  );
  MUX2_X1 _11620_ (
    .A(reg_mepc[31]),
    .B(io_pc[31]),
    .S(_03535_),
    .Z(_06022_)
  );
  MUX2_X1 _11621_ (
    .A(_06022_),
    .B(_03342_),
    .S(_05991_),
    .Z(_00001_[31])
  );
  AND2_X1 _11622_ (
    .A1(_00897_),
    .A2(_00926_),
    .ZN(_06023_)
  );
  MUX2_X1 _11623_ (
    .A(reg_mtval[0]),
    .B(io_tval[0]),
    .S(_03535_),
    .Z(_06024_)
  );
  MUX2_X1 _11624_ (
    .A(_06024_),
    .B(_01613_),
    .S(_06023_),
    .Z(_00002_[0])
  );
  MUX2_X1 _11625_ (
    .A(reg_mtval[1]),
    .B(io_tval[1]),
    .S(_03535_),
    .Z(_06025_)
  );
  MUX2_X1 _11626_ (
    .A(_06025_),
    .B(_01688_),
    .S(_06023_),
    .Z(_00002_[1])
  );
  MUX2_X1 _11627_ (
    .A(reg_mtval[2]),
    .B(io_tval[2]),
    .S(_03535_),
    .Z(_06026_)
  );
  MUX2_X1 _11628_ (
    .A(_06026_),
    .B(_01774_),
    .S(_06023_),
    .Z(_00002_[2])
  );
  MUX2_X1 _11629_ (
    .A(reg_mtval[3]),
    .B(io_tval[3]),
    .S(_03535_),
    .Z(_06027_)
  );
  MUX2_X1 _11630_ (
    .A(_06027_),
    .B(_01865_),
    .S(_06023_),
    .Z(_00002_[3])
  );
  MUX2_X1 _11631_ (
    .A(reg_mtval[4]),
    .B(io_tval[4]),
    .S(_03535_),
    .Z(_06028_)
  );
  MUX2_X1 _11632_ (
    .A(_06028_),
    .B(_01938_),
    .S(_06023_),
    .Z(_00002_[4])
  );
  MUX2_X1 _11633_ (
    .A(reg_mtval[5]),
    .B(io_tval[5]),
    .S(_03535_),
    .Z(_06029_)
  );
  MUX2_X1 _11634_ (
    .A(_06029_),
    .B(_02005_),
    .S(_06023_),
    .Z(_00002_[5])
  );
  MUX2_X1 _11635_ (
    .A(reg_mtval[6]),
    .B(io_tval[6]),
    .S(_03535_),
    .Z(_06030_)
  );
  MUX2_X1 _11636_ (
    .A(_06030_),
    .B(_02076_),
    .S(_06023_),
    .Z(_00002_[6])
  );
  MUX2_X1 _11637_ (
    .A(reg_mtval[7]),
    .B(io_tval[7]),
    .S(_03535_),
    .Z(_06031_)
  );
  MUX2_X1 _11638_ (
    .A(_06031_),
    .B(_02163_),
    .S(_06023_),
    .Z(_00002_[7])
  );
  MUX2_X1 _11639_ (
    .A(reg_mtval[8]),
    .B(io_tval[8]),
    .S(_03535_),
    .Z(_06032_)
  );
  MUX2_X1 _11640_ (
    .A(_06032_),
    .B(_01446_),
    .S(_06023_),
    .Z(_00002_[8])
  );
  MUX2_X1 _11641_ (
    .A(reg_mtval[9]),
    .B(io_tval[9]),
    .S(_03535_),
    .Z(_06033_)
  );
  MUX2_X1 _11642_ (
    .A(_06033_),
    .B(_01518_),
    .S(_06023_),
    .Z(_00002_[9])
  );
  MUX2_X1 _11643_ (
    .A(reg_mtval[10]),
    .B(io_tval[10]),
    .S(_03535_),
    .Z(_06034_)
  );
  MUX2_X1 _11644_ (
    .A(_06034_),
    .B(_02235_),
    .S(_06023_),
    .Z(_00002_[10])
  );
  MUX2_X1 _11645_ (
    .A(reg_mtval[11]),
    .B(io_tval[11]),
    .S(_03535_),
    .Z(_06035_)
  );
  MUX2_X1 _11646_ (
    .A(_06035_),
    .B(_02314_),
    .S(_06023_),
    .Z(_00002_[11])
  );
  MUX2_X1 _11647_ (
    .A(reg_mtval[12]),
    .B(io_tval[12]),
    .S(_03535_),
    .Z(_06036_)
  );
  MUX2_X1 _11648_ (
    .A(_06036_),
    .B(_02389_),
    .S(_06023_),
    .Z(_00002_[12])
  );
  MUX2_X1 _11649_ (
    .A(reg_mtval[13]),
    .B(io_tval[13]),
    .S(_03535_),
    .Z(_06037_)
  );
  MUX2_X1 _11650_ (
    .A(_06037_),
    .B(_02456_),
    .S(_06023_),
    .Z(_00002_[13])
  );
  MUX2_X1 _11651_ (
    .A(reg_mtval[14]),
    .B(io_tval[14]),
    .S(_03535_),
    .Z(_06038_)
  );
  MUX2_X1 _11652_ (
    .A(_06038_),
    .B(_02522_),
    .S(_06023_),
    .Z(_00002_[14])
  );
  MUX2_X1 _11653_ (
    .A(reg_mtval[15]),
    .B(io_tval[15]),
    .S(_03535_),
    .Z(_06039_)
  );
  MUX2_X1 _11654_ (
    .A(_06039_),
    .B(_02597_),
    .S(_06023_),
    .Z(_00002_[15])
  );
  MUX2_X1 _11655_ (
    .A(reg_mtval[16]),
    .B(io_tval[16]),
    .S(_03535_),
    .Z(_06040_)
  );
  MUX2_X1 _11656_ (
    .A(_06040_),
    .B(_01035_),
    .S(_06023_),
    .Z(_00002_[16])
  );
  MUX2_X1 _11657_ (
    .A(reg_mtval[17]),
    .B(io_tval[17]),
    .S(_03535_),
    .Z(_06041_)
  );
  MUX2_X1 _11658_ (
    .A(_06041_),
    .B(_02669_),
    .S(_06023_),
    .Z(_00002_[17])
  );
  MUX2_X1 _11659_ (
    .A(reg_mtval[18]),
    .B(io_tval[18]),
    .S(_03535_),
    .Z(_06042_)
  );
  MUX2_X1 _11660_ (
    .A(_06042_),
    .B(_01107_),
    .S(_06023_),
    .Z(_00002_[18])
  );
  MUX2_X1 _11661_ (
    .A(reg_mtval[19]),
    .B(io_tval[19]),
    .S(_03535_),
    .Z(_06043_)
  );
  MUX2_X1 _11662_ (
    .A(_06043_),
    .B(_01199_),
    .S(_06023_),
    .Z(_00002_[19])
  );
  MUX2_X1 _11663_ (
    .A(reg_mtval[20]),
    .B(io_tval[20]),
    .S(_03535_),
    .Z(_06044_)
  );
  MUX2_X1 _11664_ (
    .A(_06044_),
    .B(_01277_),
    .S(_06023_),
    .Z(_00002_[20])
  );
  MUX2_X1 _11665_ (
    .A(reg_mtval[21]),
    .B(io_tval[21]),
    .S(_03535_),
    .Z(_06045_)
  );
  MUX2_X1 _11666_ (
    .A(_06045_),
    .B(_02735_),
    .S(_06023_),
    .Z(_00002_[21])
  );
  MUX2_X1 _11667_ (
    .A(reg_mtval[22]),
    .B(io_tval[22]),
    .S(_03535_),
    .Z(_06046_)
  );
  MUX2_X1 _11668_ (
    .A(_06046_),
    .B(_02801_),
    .S(_06023_),
    .Z(_00002_[22])
  );
  MUX2_X1 _11669_ (
    .A(reg_mtval[23]),
    .B(io_tval[23]),
    .S(_03535_),
    .Z(_06047_)
  );
  MUX2_X1 _11670_ (
    .A(_06047_),
    .B(_01360_),
    .S(_06023_),
    .Z(_00002_[23])
  );
  MUX2_X1 _11671_ (
    .A(reg_mtval[24]),
    .B(io_tval[24]),
    .S(_03535_),
    .Z(_06048_)
  );
  MUX2_X1 _11672_ (
    .A(_06048_),
    .B(_02873_),
    .S(_06023_),
    .Z(_00002_[24])
  );
  MUX2_X1 _11673_ (
    .A(reg_mtval[25]),
    .B(io_tval[25]),
    .S(_03535_),
    .Z(_06049_)
  );
  MUX2_X1 _11674_ (
    .A(_06049_),
    .B(_02945_),
    .S(_06023_),
    .Z(_00002_[25])
  );
  MUX2_X1 _11675_ (
    .A(reg_mtval[26]),
    .B(io_tval[26]),
    .S(_03535_),
    .Z(_06050_)
  );
  MUX2_X1 _11676_ (
    .A(_06050_),
    .B(_03017_),
    .S(_06023_),
    .Z(_00002_[26])
  );
  MUX2_X1 _11677_ (
    .A(reg_mtval[27]),
    .B(io_tval[27]),
    .S(_03535_),
    .Z(_06051_)
  );
  MUX2_X1 _11678_ (
    .A(_06051_),
    .B(_03089_),
    .S(_06023_),
    .Z(_00002_[27])
  );
  MUX2_X1 _11679_ (
    .A(reg_mtval[28]),
    .B(io_tval[28]),
    .S(_03535_),
    .Z(_06052_)
  );
  MUX2_X1 _11680_ (
    .A(_06052_),
    .B(_03162_),
    .S(_06023_),
    .Z(_00002_[28])
  );
  MUX2_X1 _11681_ (
    .A(reg_mtval[29]),
    .B(io_tval[29]),
    .S(_03535_),
    .Z(_06053_)
  );
  MUX2_X1 _11682_ (
    .A(_06053_),
    .B(_03230_),
    .S(_06023_),
    .Z(_00002_[29])
  );
  MUX2_X1 _11683_ (
    .A(reg_mtval[30]),
    .B(io_tval[30]),
    .S(_03535_),
    .Z(_06054_)
  );
  MUX2_X1 _11684_ (
    .A(_06054_),
    .B(_03443_),
    .S(_06023_),
    .Z(_00002_[30])
  );
  MUX2_X1 _11685_ (
    .A(reg_mtval[31]),
    .B(io_tval[31]),
    .S(_03535_),
    .Z(_06055_)
  );
  MUX2_X1 _11686_ (
    .A(_06055_),
    .B(_03342_),
    .S(_06023_),
    .Z(_00002_[31])
  );
  AND2_X1 _11687_ (
    .A1(reg_mstatus_mie),
    .A2(_00835_),
    .ZN(_06056_)
  );
  AND2_X1 _11688_ (
    .A1(_03632_),
    .A2(_06056_),
    .ZN(io_interrupt_cause[0])
  );
  INV_X1 _11689_ (
    .A(io_interrupt_cause[0]),
    .ZN(_06057_)
  );
  AND2_X1 _11690_ (
    .A1(_00835_),
    .A2(_06057_),
    .ZN(_06058_)
  );
  INV_X1 _11691_ (
    .A(_06058_),
    .ZN(io_interrupt_cause[1])
  );
  AND2_X1 _11692_ (
    .A1(_03630_),
    .A2(_06056_),
    .ZN(_06059_)
  );
  INV_X1 _11693_ (
    .A(_06059_),
    .ZN(io_interrupt_cause[2])
  );
  AND2_X1 _11694_ (
    .A1(reg_mstatus_mie),
    .A2(_03627_),
    .ZN(_06060_)
  );
  INV_X1 _11695_ (
    .A(_06060_),
    .ZN(_06061_)
  );
  AND2_X1 _11696_ (
    .A1(_00835_),
    .A2(_06061_),
    .ZN(_06062_)
  );
  INV_X1 _11697_ (
    .A(_06062_),
    .ZN(io_interrupt_cause[3])
  );
  AND2_X1 _11698_ (
    .A1(_01641_),
    .A2(_03551_),
    .ZN(_06063_)
  );
  INV_X1 _11699_ (
    .A(_06063_),
    .ZN(_06064_)
  );
  AND2_X1 _11700_ (
    .A1(_01630_),
    .A2(_03547_),
    .ZN(_06065_)
  );
  INV_X1 _11701_ (
    .A(_06065_),
    .ZN(_06066_)
  );
  AND2_X1 _11702_ (
    .A1(_06064_),
    .A2(_06066_),
    .ZN(_06067_)
  );
  INV_X1 _11703_ (
    .A(_06067_),
    .ZN(io_evec[1])
  );
  AND2_X1 _11704_ (
    .A1(_03533_),
    .A2(_03544_),
    .ZN(_06068_)
  );
  AND2_X1 _11705_ (
    .A1(reg_mtvec[0]),
    .A2(_03577_),
    .ZN(_06069_)
  );
  AND2_X1 _11706_ (
    .A1(_03515_),
    .A2(_06069_),
    .ZN(_06070_)
  );
  MUX2_X1 _11707_ (
    .A(_01717_),
    .B(io_cause[0]),
    .S(_06070_),
    .Z(_06071_)
  );
  AND2_X1 _11708_ (
    .A1(_06068_),
    .A2(_06071_),
    .ZN(_06072_)
  );
  INV_X1 _11709_ (
    .A(_06072_),
    .ZN(_06073_)
  );
  AND2_X1 _11710_ (
    .A1(reg_mepc[2]),
    .A2(_03551_),
    .ZN(_06074_)
  );
  INV_X1 _11711_ (
    .A(_06074_),
    .ZN(_06075_)
  );
  AND2_X1 _11712_ (
    .A1(reg_dpc[2]),
    .A2(_03547_),
    .ZN(_06076_)
  );
  INV_X1 _11713_ (
    .A(_06076_),
    .ZN(_06077_)
  );
  AND2_X1 _11714_ (
    .A1(_06075_),
    .A2(_06077_),
    .ZN(_06078_)
  );
  AND2_X1 _11715_ (
    .A1(_06073_),
    .A2(_06078_),
    .ZN(_06079_)
  );
  INV_X1 _11716_ (
    .A(_06079_),
    .ZN(io_evec[2])
  );
  AND2_X1 _11717_ (
    .A1(reg_debug),
    .A2(_03485_),
    .ZN(_06080_)
  );
  INV_X1 _11718_ (
    .A(_06080_),
    .ZN(_06081_)
  );
  MUX2_X1 _11719_ (
    .A(_01846_),
    .B(io_cause[1]),
    .S(_06070_),
    .Z(_06082_)
  );
  AND2_X1 _11720_ (
    .A1(_03533_),
    .A2(_06082_),
    .ZN(_06083_)
  );
  INV_X1 _11721_ (
    .A(_06083_),
    .ZN(_06084_)
  );
  AND2_X1 _11722_ (
    .A1(_06081_),
    .A2(_06084_),
    .ZN(_06085_)
  );
  INV_X1 _11723_ (
    .A(_06085_),
    .ZN(_06086_)
  );
  AND2_X1 _11724_ (
    .A1(_03544_),
    .A2(_06086_),
    .ZN(_06087_)
  );
  INV_X1 _11725_ (
    .A(_06087_),
    .ZN(_06088_)
  );
  AND2_X1 _11726_ (
    .A1(reg_dpc[3]),
    .A2(_03547_),
    .ZN(_06089_)
  );
  INV_X1 _11727_ (
    .A(_06089_),
    .ZN(_06090_)
  );
  AND2_X1 _11728_ (
    .A1(reg_mepc[3]),
    .A2(_03551_),
    .ZN(_06091_)
  );
  INV_X1 _11729_ (
    .A(_06091_),
    .ZN(_06092_)
  );
  AND2_X1 _11730_ (
    .A1(_06090_),
    .A2(_06092_),
    .ZN(_06093_)
  );
  AND2_X1 _11731_ (
    .A1(_06088_),
    .A2(_06093_),
    .ZN(_06094_)
  );
  INV_X1 _11732_ (
    .A(_06094_),
    .ZN(io_evec[3])
  );
  MUX2_X1 _11733_ (
    .A(_01879_),
    .B(io_cause[2]),
    .S(_06070_),
    .Z(_06095_)
  );
  AND2_X1 _11734_ (
    .A1(_06068_),
    .A2(_06095_),
    .ZN(_06096_)
  );
  INV_X1 _11735_ (
    .A(_06096_),
    .ZN(_06097_)
  );
  AND2_X1 _11736_ (
    .A1(reg_mepc[4]),
    .A2(_03551_),
    .ZN(_06098_)
  );
  INV_X1 _11737_ (
    .A(_06098_),
    .ZN(_06099_)
  );
  AND2_X1 _11738_ (
    .A1(reg_dpc[4]),
    .A2(_03547_),
    .ZN(_06100_)
  );
  INV_X1 _11739_ (
    .A(_06100_),
    .ZN(_06101_)
  );
  AND2_X1 _11740_ (
    .A1(_06099_),
    .A2(_06101_),
    .ZN(_06102_)
  );
  AND2_X1 _11741_ (
    .A1(_06097_),
    .A2(_06102_),
    .ZN(_06103_)
  );
  INV_X1 _11742_ (
    .A(_06103_),
    .ZN(io_evec[4])
  );
  MUX2_X1 _11743_ (
    .A(_01955_),
    .B(_03525_),
    .S(_06070_),
    .Z(_06104_)
  );
  AND2_X1 _11744_ (
    .A1(_06068_),
    .A2(_06104_),
    .ZN(_06105_)
  );
  INV_X1 _11745_ (
    .A(_06105_),
    .ZN(_06106_)
  );
  AND2_X1 _11746_ (
    .A1(reg_mepc[5]),
    .A2(_03551_),
    .ZN(_06107_)
  );
  INV_X1 _11747_ (
    .A(_06107_),
    .ZN(_06108_)
  );
  AND2_X1 _11748_ (
    .A1(reg_dpc[5]),
    .A2(_03547_),
    .ZN(_06109_)
  );
  INV_X1 _11749_ (
    .A(_06109_),
    .ZN(_06110_)
  );
  AND2_X1 _11750_ (
    .A1(_06108_),
    .A2(_06110_),
    .ZN(_06111_)
  );
  AND2_X1 _11751_ (
    .A1(_06106_),
    .A2(_06111_),
    .ZN(_06112_)
  );
  INV_X1 _11752_ (
    .A(_06112_),
    .ZN(io_evec[5])
  );
  MUX2_X1 _11753_ (
    .A(_02040_),
    .B(io_cause[4]),
    .S(_06070_),
    .Z(_06113_)
  );
  AND2_X1 _11754_ (
    .A1(_06068_),
    .A2(_06113_),
    .ZN(_06114_)
  );
  INV_X1 _11755_ (
    .A(_06114_),
    .ZN(_06115_)
  );
  AND2_X1 _11756_ (
    .A1(reg_mepc[6]),
    .A2(_03551_),
    .ZN(_06116_)
  );
  INV_X1 _11757_ (
    .A(_06116_),
    .ZN(_06117_)
  );
  AND2_X1 _11758_ (
    .A1(reg_dpc[6]),
    .A2(_03547_),
    .ZN(_06118_)
  );
  INV_X1 _11759_ (
    .A(_06118_),
    .ZN(_06119_)
  );
  AND2_X1 _11760_ (
    .A1(_06117_),
    .A2(_06119_),
    .ZN(_06120_)
  );
  AND2_X1 _11761_ (
    .A1(_06115_),
    .A2(_06120_),
    .ZN(_06121_)
  );
  INV_X1 _11762_ (
    .A(_06121_),
    .ZN(io_evec[6])
  );
  AND2_X1 _11763_ (
    .A1(reg_mtvec[7]),
    .A2(_06068_),
    .ZN(_06122_)
  );
  INV_X1 _11764_ (
    .A(_06122_),
    .ZN(_06123_)
  );
  AND2_X1 _11765_ (
    .A1(reg_mepc[7]),
    .A2(_03551_),
    .ZN(_06124_)
  );
  INV_X1 _11766_ (
    .A(_06124_),
    .ZN(_06125_)
  );
  AND2_X1 _11767_ (
    .A1(reg_dpc[7]),
    .A2(_03547_),
    .ZN(_06126_)
  );
  INV_X1 _11768_ (
    .A(_06126_),
    .ZN(_06127_)
  );
  AND2_X1 _11769_ (
    .A1(_06125_),
    .A2(_06127_),
    .ZN(_06128_)
  );
  AND2_X1 _11770_ (
    .A1(_06123_),
    .A2(_06128_),
    .ZN(_06129_)
  );
  INV_X1 _11771_ (
    .A(_06129_),
    .ZN(io_evec[7])
  );
  AND2_X1 _11772_ (
    .A1(reg_mtvec[8]),
    .A2(_06068_),
    .ZN(_06130_)
  );
  INV_X1 _11773_ (
    .A(_06130_),
    .ZN(_06131_)
  );
  AND2_X1 _11774_ (
    .A1(reg_mepc[8]),
    .A2(_03551_),
    .ZN(_06132_)
  );
  INV_X1 _11775_ (
    .A(_06132_),
    .ZN(_06133_)
  );
  AND2_X1 _11776_ (
    .A1(reg_dpc[8]),
    .A2(_03547_),
    .ZN(_06134_)
  );
  INV_X1 _11777_ (
    .A(_06134_),
    .ZN(_06135_)
  );
  AND2_X1 _11778_ (
    .A1(_06133_),
    .A2(_06135_),
    .ZN(_06136_)
  );
  AND2_X1 _11779_ (
    .A1(_06131_),
    .A2(_06136_),
    .ZN(_06137_)
  );
  INV_X1 _11780_ (
    .A(_06137_),
    .ZN(io_evec[8])
  );
  AND2_X1 _11781_ (
    .A1(reg_mtvec[9]),
    .A2(_06068_),
    .ZN(_06138_)
  );
  INV_X1 _11782_ (
    .A(_06138_),
    .ZN(_06139_)
  );
  AND2_X1 _11783_ (
    .A1(reg_dpc[9]),
    .A2(_03547_),
    .ZN(_06140_)
  );
  INV_X1 _11784_ (
    .A(_06140_),
    .ZN(_06141_)
  );
  AND2_X1 _11785_ (
    .A1(reg_mepc[9]),
    .A2(_03551_),
    .ZN(_06142_)
  );
  INV_X1 _11786_ (
    .A(_06142_),
    .ZN(_06143_)
  );
  AND2_X1 _11787_ (
    .A1(_06141_),
    .A2(_06143_),
    .ZN(_06144_)
  );
  AND2_X1 _11788_ (
    .A1(_06139_),
    .A2(_06144_),
    .ZN(_06145_)
  );
  INV_X1 _11789_ (
    .A(_06145_),
    .ZN(io_evec[9])
  );
  AND2_X1 _11790_ (
    .A1(reg_mtvec[10]),
    .A2(_06068_),
    .ZN(_06146_)
  );
  INV_X1 _11791_ (
    .A(_06146_),
    .ZN(_06147_)
  );
  AND2_X1 _11792_ (
    .A1(reg_mepc[10]),
    .A2(_03551_),
    .ZN(_06148_)
  );
  INV_X1 _11793_ (
    .A(_06148_),
    .ZN(_06149_)
  );
  AND2_X1 _11794_ (
    .A1(reg_dpc[10]),
    .A2(_03547_),
    .ZN(_06150_)
  );
  INV_X1 _11795_ (
    .A(_06150_),
    .ZN(_06151_)
  );
  AND2_X1 _11796_ (
    .A1(_06149_),
    .A2(_06151_),
    .ZN(_06152_)
  );
  AND2_X1 _11797_ (
    .A1(_06147_),
    .A2(_06152_),
    .ZN(_06153_)
  );
  INV_X1 _11798_ (
    .A(_06153_),
    .ZN(io_evec[10])
  );
  AND2_X1 _11799_ (
    .A1(_00693_),
    .A2(_03533_),
    .ZN(_06154_)
  );
  INV_X1 _11800_ (
    .A(_06154_),
    .ZN(_06155_)
  );
  AND2_X1 _11801_ (
    .A1(_03544_),
    .A2(_06155_),
    .ZN(_06156_)
  );
  INV_X1 _11802_ (
    .A(_06156_),
    .ZN(_06157_)
  );
  AND2_X1 _11803_ (
    .A1(reg_mepc[11]),
    .A2(_03551_),
    .ZN(_06158_)
  );
  INV_X1 _11804_ (
    .A(_06158_),
    .ZN(_06159_)
  );
  AND2_X1 _11805_ (
    .A1(reg_dpc[11]),
    .A2(_03547_),
    .ZN(_06160_)
  );
  INV_X1 _11806_ (
    .A(_06160_),
    .ZN(_06161_)
  );
  AND2_X1 _11807_ (
    .A1(_06159_),
    .A2(_06161_),
    .ZN(_06162_)
  );
  AND2_X1 _11808_ (
    .A1(_06157_),
    .A2(_06162_),
    .ZN(_06163_)
  );
  INV_X1 _11809_ (
    .A(_06163_),
    .ZN(io_evec[11])
  );
  AND2_X1 _11810_ (
    .A1(reg_mtvec[12]),
    .A2(_06068_),
    .ZN(_06164_)
  );
  INV_X1 _11811_ (
    .A(_06164_),
    .ZN(_06165_)
  );
  AND2_X1 _11812_ (
    .A1(reg_mepc[12]),
    .A2(_03551_),
    .ZN(_06166_)
  );
  INV_X1 _11813_ (
    .A(_06166_),
    .ZN(_06167_)
  );
  AND2_X1 _11814_ (
    .A1(reg_dpc[12]),
    .A2(_03547_),
    .ZN(_06168_)
  );
  INV_X1 _11815_ (
    .A(_06168_),
    .ZN(_06169_)
  );
  AND2_X1 _11816_ (
    .A1(_06167_),
    .A2(_06169_),
    .ZN(_06170_)
  );
  AND2_X1 _11817_ (
    .A1(_06165_),
    .A2(_06170_),
    .ZN(_06171_)
  );
  INV_X1 _11818_ (
    .A(_06171_),
    .ZN(io_evec[12])
  );
  AND2_X1 _11819_ (
    .A1(reg_mtvec[13]),
    .A2(_06068_),
    .ZN(_06172_)
  );
  INV_X1 _11820_ (
    .A(_06172_),
    .ZN(_06173_)
  );
  AND2_X1 _11821_ (
    .A1(reg_mepc[13]),
    .A2(_03551_),
    .ZN(_06174_)
  );
  INV_X1 _11822_ (
    .A(_06174_),
    .ZN(_06175_)
  );
  AND2_X1 _11823_ (
    .A1(reg_dpc[13]),
    .A2(_03547_),
    .ZN(_06176_)
  );
  INV_X1 _11824_ (
    .A(_06176_),
    .ZN(_06177_)
  );
  AND2_X1 _11825_ (
    .A1(_06175_),
    .A2(_06177_),
    .ZN(_06178_)
  );
  AND2_X1 _11826_ (
    .A1(_06173_),
    .A2(_06178_),
    .ZN(_06179_)
  );
  INV_X1 _11827_ (
    .A(_06179_),
    .ZN(io_evec[13])
  );
  AND2_X1 _11828_ (
    .A1(reg_mtvec[14]),
    .A2(_06068_),
    .ZN(_06180_)
  );
  INV_X1 _11829_ (
    .A(_06180_),
    .ZN(_06181_)
  );
  AND2_X1 _11830_ (
    .A1(reg_mepc[14]),
    .A2(_03551_),
    .ZN(_06182_)
  );
  INV_X1 _11831_ (
    .A(_06182_),
    .ZN(_06183_)
  );
  AND2_X1 _11832_ (
    .A1(reg_dpc[14]),
    .A2(_03547_),
    .ZN(_06184_)
  );
  INV_X1 _11833_ (
    .A(_06184_),
    .ZN(_06185_)
  );
  AND2_X1 _11834_ (
    .A1(_06183_),
    .A2(_06185_),
    .ZN(_06186_)
  );
  AND2_X1 _11835_ (
    .A1(_06181_),
    .A2(_06186_),
    .ZN(_06187_)
  );
  INV_X1 _11836_ (
    .A(_06187_),
    .ZN(io_evec[14])
  );
  AND2_X1 _11837_ (
    .A1(reg_mtvec[15]),
    .A2(_06068_),
    .ZN(_06188_)
  );
  INV_X1 _11838_ (
    .A(_06188_),
    .ZN(_06189_)
  );
  AND2_X1 _11839_ (
    .A1(reg_mepc[15]),
    .A2(_03551_),
    .ZN(_06190_)
  );
  INV_X1 _11840_ (
    .A(_06190_),
    .ZN(_06191_)
  );
  AND2_X1 _11841_ (
    .A1(reg_dpc[15]),
    .A2(_03547_),
    .ZN(_06192_)
  );
  INV_X1 _11842_ (
    .A(_06192_),
    .ZN(_06193_)
  );
  AND2_X1 _11843_ (
    .A1(_06191_),
    .A2(_06193_),
    .ZN(_06194_)
  );
  AND2_X1 _11844_ (
    .A1(_06189_),
    .A2(_06194_),
    .ZN(_06195_)
  );
  INV_X1 _11845_ (
    .A(_06195_),
    .ZN(io_evec[15])
  );
  AND2_X1 _11846_ (
    .A1(reg_mtvec[16]),
    .A2(_06068_),
    .ZN(_06196_)
  );
  INV_X1 _11847_ (
    .A(_06196_),
    .ZN(_06197_)
  );
  AND2_X1 _11848_ (
    .A1(reg_mepc[16]),
    .A2(_03551_),
    .ZN(_06198_)
  );
  INV_X1 _11849_ (
    .A(_06198_),
    .ZN(_06199_)
  );
  AND2_X1 _11850_ (
    .A1(reg_dpc[16]),
    .A2(_03547_),
    .ZN(_06200_)
  );
  INV_X1 _11851_ (
    .A(_06200_),
    .ZN(_06201_)
  );
  AND2_X1 _11852_ (
    .A1(_06199_),
    .A2(_06201_),
    .ZN(_06202_)
  );
  AND2_X1 _11853_ (
    .A1(_06197_),
    .A2(_06202_),
    .ZN(_06203_)
  );
  INV_X1 _11854_ (
    .A(_06203_),
    .ZN(io_evec[16])
  );
  AND2_X1 _11855_ (
    .A1(reg_mtvec[17]),
    .A2(_06068_),
    .ZN(_06204_)
  );
  INV_X1 _11856_ (
    .A(_06204_),
    .ZN(_06205_)
  );
  AND2_X1 _11857_ (
    .A1(reg_mepc[17]),
    .A2(_03551_),
    .ZN(_06206_)
  );
  INV_X1 _11858_ (
    .A(_06206_),
    .ZN(_06207_)
  );
  AND2_X1 _11859_ (
    .A1(reg_dpc[17]),
    .A2(_03547_),
    .ZN(_06208_)
  );
  INV_X1 _11860_ (
    .A(_06208_),
    .ZN(_06209_)
  );
  AND2_X1 _11861_ (
    .A1(_06207_),
    .A2(_06209_),
    .ZN(_06210_)
  );
  AND2_X1 _11862_ (
    .A1(_06205_),
    .A2(_06210_),
    .ZN(_06211_)
  );
  INV_X1 _11863_ (
    .A(_06211_),
    .ZN(io_evec[17])
  );
  AND2_X1 _11864_ (
    .A1(reg_mtvec[18]),
    .A2(_06068_),
    .ZN(_06212_)
  );
  INV_X1 _11865_ (
    .A(_06212_),
    .ZN(_06213_)
  );
  AND2_X1 _11866_ (
    .A1(reg_mepc[18]),
    .A2(_03551_),
    .ZN(_06214_)
  );
  INV_X1 _11867_ (
    .A(_06214_),
    .ZN(_06215_)
  );
  AND2_X1 _11868_ (
    .A1(reg_dpc[18]),
    .A2(_03547_),
    .ZN(_06216_)
  );
  INV_X1 _11869_ (
    .A(_06216_),
    .ZN(_06217_)
  );
  AND2_X1 _11870_ (
    .A1(_06215_),
    .A2(_06217_),
    .ZN(_06218_)
  );
  AND2_X1 _11871_ (
    .A1(_06213_),
    .A2(_06218_),
    .ZN(_06219_)
  );
  INV_X1 _11872_ (
    .A(_06219_),
    .ZN(io_evec[18])
  );
  AND2_X1 _11873_ (
    .A1(reg_mtvec[19]),
    .A2(_06068_),
    .ZN(_06220_)
  );
  INV_X1 _11874_ (
    .A(_06220_),
    .ZN(_06221_)
  );
  AND2_X1 _11875_ (
    .A1(reg_dpc[19]),
    .A2(_03547_),
    .ZN(_06222_)
  );
  INV_X1 _11876_ (
    .A(_06222_),
    .ZN(_06223_)
  );
  AND2_X1 _11877_ (
    .A1(reg_mepc[19]),
    .A2(_03551_),
    .ZN(_06224_)
  );
  INV_X1 _11878_ (
    .A(_06224_),
    .ZN(_06225_)
  );
  AND2_X1 _11879_ (
    .A1(_06223_),
    .A2(_06225_),
    .ZN(_06226_)
  );
  AND2_X1 _11880_ (
    .A1(_06221_),
    .A2(_06226_),
    .ZN(_06227_)
  );
  INV_X1 _11881_ (
    .A(_06227_),
    .ZN(io_evec[19])
  );
  AND2_X1 _11882_ (
    .A1(reg_mtvec[20]),
    .A2(_06068_),
    .ZN(_06228_)
  );
  INV_X1 _11883_ (
    .A(_06228_),
    .ZN(_06229_)
  );
  AND2_X1 _11884_ (
    .A1(reg_dpc[20]),
    .A2(_03547_),
    .ZN(_06230_)
  );
  INV_X1 _11885_ (
    .A(_06230_),
    .ZN(_06231_)
  );
  AND2_X1 _11886_ (
    .A1(reg_mepc[20]),
    .A2(_03551_),
    .ZN(_06232_)
  );
  INV_X1 _11887_ (
    .A(_06232_),
    .ZN(_06233_)
  );
  AND2_X1 _11888_ (
    .A1(_06231_),
    .A2(_06233_),
    .ZN(_06234_)
  );
  AND2_X1 _11889_ (
    .A1(_06229_),
    .A2(_06234_),
    .ZN(_06235_)
  );
  INV_X1 _11890_ (
    .A(_06235_),
    .ZN(io_evec[20])
  );
  AND2_X1 _11891_ (
    .A1(reg_mtvec[21]),
    .A2(_06068_),
    .ZN(_06236_)
  );
  INV_X1 _11892_ (
    .A(_06236_),
    .ZN(_06237_)
  );
  AND2_X1 _11893_ (
    .A1(reg_mepc[21]),
    .A2(_03551_),
    .ZN(_06238_)
  );
  INV_X1 _11894_ (
    .A(_06238_),
    .ZN(_06239_)
  );
  AND2_X1 _11895_ (
    .A1(reg_dpc[21]),
    .A2(_03547_),
    .ZN(_06240_)
  );
  INV_X1 _11896_ (
    .A(_06240_),
    .ZN(_06241_)
  );
  AND2_X1 _11897_ (
    .A1(_06239_),
    .A2(_06241_),
    .ZN(_06242_)
  );
  AND2_X1 _11898_ (
    .A1(_06237_),
    .A2(_06242_),
    .ZN(_06243_)
  );
  INV_X1 _11899_ (
    .A(_06243_),
    .ZN(io_evec[21])
  );
  AND2_X1 _11900_ (
    .A1(reg_mtvec[22]),
    .A2(_06068_),
    .ZN(_06244_)
  );
  INV_X1 _11901_ (
    .A(_06244_),
    .ZN(_06245_)
  );
  AND2_X1 _11902_ (
    .A1(reg_mepc[22]),
    .A2(_03551_),
    .ZN(_06246_)
  );
  INV_X1 _11903_ (
    .A(_06246_),
    .ZN(_06247_)
  );
  AND2_X1 _11904_ (
    .A1(reg_dpc[22]),
    .A2(_03547_),
    .ZN(_06248_)
  );
  INV_X1 _11905_ (
    .A(_06248_),
    .ZN(_06249_)
  );
  AND2_X1 _11906_ (
    .A1(_06247_),
    .A2(_06249_),
    .ZN(_06250_)
  );
  AND2_X1 _11907_ (
    .A1(_06245_),
    .A2(_06250_),
    .ZN(_06251_)
  );
  INV_X1 _11908_ (
    .A(_06251_),
    .ZN(io_evec[22])
  );
  AND2_X1 _11909_ (
    .A1(reg_mtvec[23]),
    .A2(_06068_),
    .ZN(_06252_)
  );
  INV_X1 _11910_ (
    .A(_06252_),
    .ZN(_06253_)
  );
  AND2_X1 _11911_ (
    .A1(reg_dpc[23]),
    .A2(_03547_),
    .ZN(_06254_)
  );
  INV_X1 _11912_ (
    .A(_06254_),
    .ZN(_06255_)
  );
  AND2_X1 _11913_ (
    .A1(reg_mepc[23]),
    .A2(_03551_),
    .ZN(_06256_)
  );
  INV_X1 _11914_ (
    .A(_06256_),
    .ZN(_06257_)
  );
  AND2_X1 _11915_ (
    .A1(_06255_),
    .A2(_06257_),
    .ZN(_06258_)
  );
  AND2_X1 _11916_ (
    .A1(_06253_),
    .A2(_06258_),
    .ZN(_06259_)
  );
  INV_X1 _11917_ (
    .A(_06259_),
    .ZN(io_evec[23])
  );
  AND2_X1 _11918_ (
    .A1(reg_mtvec[24]),
    .A2(_06068_),
    .ZN(_06260_)
  );
  INV_X1 _11919_ (
    .A(_06260_),
    .ZN(_06261_)
  );
  AND2_X1 _11920_ (
    .A1(reg_dpc[24]),
    .A2(_03547_),
    .ZN(_06262_)
  );
  INV_X1 _11921_ (
    .A(_06262_),
    .ZN(_06263_)
  );
  AND2_X1 _11922_ (
    .A1(reg_mepc[24]),
    .A2(_03551_),
    .ZN(_06264_)
  );
  INV_X1 _11923_ (
    .A(_06264_),
    .ZN(_06265_)
  );
  AND2_X1 _11924_ (
    .A1(_06263_),
    .A2(_06265_),
    .ZN(_06266_)
  );
  AND2_X1 _11925_ (
    .A1(_06261_),
    .A2(_06266_),
    .ZN(_06267_)
  );
  INV_X1 _11926_ (
    .A(_06267_),
    .ZN(io_evec[24])
  );
  AND2_X1 _11927_ (
    .A1(reg_mtvec[25]),
    .A2(_06068_),
    .ZN(_06268_)
  );
  INV_X1 _11928_ (
    .A(_06268_),
    .ZN(_06269_)
  );
  AND2_X1 _11929_ (
    .A1(reg_dpc[25]),
    .A2(_03547_),
    .ZN(_06270_)
  );
  INV_X1 _11930_ (
    .A(_06270_),
    .ZN(_06271_)
  );
  AND2_X1 _11931_ (
    .A1(reg_mepc[25]),
    .A2(_03551_),
    .ZN(_06272_)
  );
  INV_X1 _11932_ (
    .A(_06272_),
    .ZN(_06273_)
  );
  AND2_X1 _11933_ (
    .A1(_06271_),
    .A2(_06273_),
    .ZN(_06274_)
  );
  AND2_X1 _11934_ (
    .A1(_06269_),
    .A2(_06274_),
    .ZN(_06275_)
  );
  INV_X1 _11935_ (
    .A(_06275_),
    .ZN(io_evec[25])
  );
  AND2_X1 _11936_ (
    .A1(reg_mtvec[26]),
    .A2(_06068_),
    .ZN(_06276_)
  );
  INV_X1 _11937_ (
    .A(_06276_),
    .ZN(_06277_)
  );
  AND2_X1 _11938_ (
    .A1(reg_mepc[26]),
    .A2(_03551_),
    .ZN(_06278_)
  );
  INV_X1 _11939_ (
    .A(_06278_),
    .ZN(_06279_)
  );
  AND2_X1 _11940_ (
    .A1(reg_dpc[26]),
    .A2(_03547_),
    .ZN(_06280_)
  );
  INV_X1 _11941_ (
    .A(_06280_),
    .ZN(_06281_)
  );
  AND2_X1 _11942_ (
    .A1(_06279_),
    .A2(_06281_),
    .ZN(_06282_)
  );
  AND2_X1 _11943_ (
    .A1(_06277_),
    .A2(_06282_),
    .ZN(_06283_)
  );
  INV_X1 _11944_ (
    .A(_06283_),
    .ZN(io_evec[26])
  );
  AND2_X1 _11945_ (
    .A1(reg_mtvec[27]),
    .A2(_06068_),
    .ZN(_06284_)
  );
  INV_X1 _11946_ (
    .A(_06284_),
    .ZN(_06285_)
  );
  AND2_X1 _11947_ (
    .A1(reg_mepc[27]),
    .A2(_03551_),
    .ZN(_06286_)
  );
  INV_X1 _11948_ (
    .A(_06286_),
    .ZN(_06287_)
  );
  AND2_X1 _11949_ (
    .A1(reg_dpc[27]),
    .A2(_03547_),
    .ZN(_06288_)
  );
  INV_X1 _11950_ (
    .A(_06288_),
    .ZN(_06289_)
  );
  AND2_X1 _11951_ (
    .A1(_06287_),
    .A2(_06289_),
    .ZN(_06290_)
  );
  AND2_X1 _11952_ (
    .A1(_06285_),
    .A2(_06290_),
    .ZN(_06291_)
  );
  INV_X1 _11953_ (
    .A(_06291_),
    .ZN(io_evec[27])
  );
  AND2_X1 _11954_ (
    .A1(reg_mtvec[28]),
    .A2(_06068_),
    .ZN(_06292_)
  );
  INV_X1 _11955_ (
    .A(_06292_),
    .ZN(_06293_)
  );
  AND2_X1 _11956_ (
    .A1(reg_dpc[28]),
    .A2(_03547_),
    .ZN(_06294_)
  );
  INV_X1 _11957_ (
    .A(_06294_),
    .ZN(_06295_)
  );
  AND2_X1 _11958_ (
    .A1(reg_mepc[28]),
    .A2(_03551_),
    .ZN(_06296_)
  );
  INV_X1 _11959_ (
    .A(_06296_),
    .ZN(_06297_)
  );
  AND2_X1 _11960_ (
    .A1(_06295_),
    .A2(_06297_),
    .ZN(_06298_)
  );
  AND2_X1 _11961_ (
    .A1(_06293_),
    .A2(_06298_),
    .ZN(_06299_)
  );
  INV_X1 _11962_ (
    .A(_06299_),
    .ZN(io_evec[28])
  );
  AND2_X1 _11963_ (
    .A1(reg_mtvec[29]),
    .A2(_06068_),
    .ZN(_06300_)
  );
  INV_X1 _11964_ (
    .A(_06300_),
    .ZN(_06301_)
  );
  AND2_X1 _11965_ (
    .A1(reg_mepc[29]),
    .A2(_03551_),
    .ZN(_06302_)
  );
  INV_X1 _11966_ (
    .A(_06302_),
    .ZN(_06303_)
  );
  AND2_X1 _11967_ (
    .A1(reg_dpc[29]),
    .A2(_03547_),
    .ZN(_06304_)
  );
  INV_X1 _11968_ (
    .A(_06304_),
    .ZN(_06305_)
  );
  AND2_X1 _11969_ (
    .A1(_06303_),
    .A2(_06305_),
    .ZN(_06306_)
  );
  AND2_X1 _11970_ (
    .A1(_06301_),
    .A2(_06306_),
    .ZN(_06307_)
  );
  INV_X1 _11971_ (
    .A(_06307_),
    .ZN(io_evec[29])
  );
  AND2_X1 _11972_ (
    .A1(reg_mtvec[30]),
    .A2(_06068_),
    .ZN(_06308_)
  );
  INV_X1 _11973_ (
    .A(_06308_),
    .ZN(_06309_)
  );
  AND2_X1 _11974_ (
    .A1(reg_mepc[30]),
    .A2(_03551_),
    .ZN(_06310_)
  );
  INV_X1 _11975_ (
    .A(_06310_),
    .ZN(_06311_)
  );
  AND2_X1 _11976_ (
    .A1(reg_dpc[30]),
    .A2(_03547_),
    .ZN(_06312_)
  );
  INV_X1 _11977_ (
    .A(_06312_),
    .ZN(_06313_)
  );
  AND2_X1 _11978_ (
    .A1(_06311_),
    .A2(_06313_),
    .ZN(_06314_)
  );
  AND2_X1 _11979_ (
    .A1(_06309_),
    .A2(_06314_),
    .ZN(_06315_)
  );
  INV_X1 _11980_ (
    .A(_06315_),
    .ZN(io_evec[30])
  );
  AND2_X1 _11981_ (
    .A1(reg_mtvec[31]),
    .A2(_06068_),
    .ZN(_06316_)
  );
  INV_X1 _11982_ (
    .A(_06316_),
    .ZN(_06317_)
  );
  AND2_X1 _11983_ (
    .A1(reg_mepc[31]),
    .A2(_03551_),
    .ZN(_06318_)
  );
  INV_X1 _11984_ (
    .A(_06318_),
    .ZN(_06319_)
  );
  AND2_X1 _11985_ (
    .A1(reg_dpc[31]),
    .A2(_03547_),
    .ZN(_06320_)
  );
  INV_X1 _11986_ (
    .A(_06320_),
    .ZN(_06321_)
  );
  AND2_X1 _11987_ (
    .A1(_06319_),
    .A2(_06321_),
    .ZN(_06322_)
  );
  AND2_X1 _11988_ (
    .A1(_06317_),
    .A2(_06322_),
    .ZN(_06323_)
  );
  INV_X1 _11989_ (
    .A(_06323_),
    .ZN(io_evec[31])
  );
  AND2_X1 _11990_ (
    .A1(_00820_),
    .A2(_00821_),
    .ZN(_06324_)
  );
  AND2_X1 _11991_ (
    .A1(_00822_),
    .A2(_06324_),
    .ZN(_06325_)
  );
  AND2_X1 _11992_ (
    .A1(io_decode_0_inst[26]),
    .A2(_06325_),
    .ZN(_06326_)
  );
  AND2_X1 _11993_ (
    .A1(_00814_),
    .A2(_00819_),
    .ZN(_06327_)
  );
  INV_X1 _11994_ (
    .A(_06327_),
    .ZN(_06328_)
  );
  AND2_X1 _11995_ (
    .A1(_00816_),
    .A2(_00823_),
    .ZN(_06329_)
  );
  AND2_X1 _11996_ (
    .A1(_06327_),
    .A2(_06329_),
    .ZN(_06330_)
  );
  AND2_X1 _11997_ (
    .A1(io_decode_0_inst[21]),
    .A2(_06327_),
    .ZN(_06331_)
  );
  AND2_X1 _11998_ (
    .A1(_00815_),
    .A2(_00822_),
    .ZN(_06332_)
  );
  AND2_X1 _11999_ (
    .A1(_06326_),
    .A2(_06330_),
    .ZN(_06333_)
  );
  INV_X1 _12000_ (
    .A(_06333_),
    .ZN(io_decode_0_write_flush)
  );
  AND2_X1 _12001_ (
    .A1(reg_pmp_0_cfg_a[0]),
    .A2(reg_pmp_0_addr[0]),
    .ZN(io_pmp_0_mask[3])
  );
  AND2_X1 _12002_ (
    .A1(reg_pmp_0_addr[1]),
    .A2(io_pmp_0_mask[3]),
    .ZN(io_pmp_0_mask[4])
  );
  AND2_X1 _12003_ (
    .A1(reg_pmp_0_addr[2]),
    .A2(io_pmp_0_mask[4]),
    .ZN(io_pmp_0_mask[5])
  );
  AND2_X1 _12004_ (
    .A1(reg_pmp_0_addr[3]),
    .A2(io_pmp_0_mask[5]),
    .ZN(io_pmp_0_mask[6])
  );
  AND2_X1 _12005_ (
    .A1(reg_pmp_0_addr[4]),
    .A2(io_pmp_0_mask[6]),
    .ZN(io_pmp_0_mask[7])
  );
  AND2_X1 _12006_ (
    .A1(reg_pmp_0_addr[5]),
    .A2(io_pmp_0_mask[7]),
    .ZN(io_pmp_0_mask[8])
  );
  AND2_X1 _12007_ (
    .A1(reg_pmp_0_addr[6]),
    .A2(io_pmp_0_mask[8]),
    .ZN(io_pmp_0_mask[9])
  );
  AND2_X1 _12008_ (
    .A1(reg_pmp_0_addr[7]),
    .A2(io_pmp_0_mask[9]),
    .ZN(io_pmp_0_mask[10])
  );
  AND2_X1 _12009_ (
    .A1(reg_pmp_0_addr[8]),
    .A2(io_pmp_0_mask[10]),
    .ZN(io_pmp_0_mask[11])
  );
  AND2_X1 _12010_ (
    .A1(reg_pmp_0_addr[9]),
    .A2(io_pmp_0_mask[11]),
    .ZN(io_pmp_0_mask[12])
  );
  AND2_X1 _12011_ (
    .A1(reg_pmp_0_addr[10]),
    .A2(io_pmp_0_mask[12]),
    .ZN(io_pmp_0_mask[13])
  );
  AND2_X1 _12012_ (
    .A1(reg_pmp_0_addr[11]),
    .A2(io_pmp_0_mask[13]),
    .ZN(io_pmp_0_mask[14])
  );
  AND2_X1 _12013_ (
    .A1(reg_pmp_0_addr[12]),
    .A2(io_pmp_0_mask[14]),
    .ZN(io_pmp_0_mask[15])
  );
  AND2_X1 _12014_ (
    .A1(reg_pmp_0_addr[13]),
    .A2(io_pmp_0_mask[15]),
    .ZN(io_pmp_0_mask[16])
  );
  AND2_X1 _12015_ (
    .A1(reg_pmp_0_addr[14]),
    .A2(io_pmp_0_mask[16]),
    .ZN(io_pmp_0_mask[17])
  );
  AND2_X1 _12016_ (
    .A1(reg_pmp_0_addr[15]),
    .A2(io_pmp_0_mask[17]),
    .ZN(io_pmp_0_mask[18])
  );
  AND2_X1 _12017_ (
    .A1(reg_pmp_0_addr[16]),
    .A2(io_pmp_0_mask[18]),
    .ZN(io_pmp_0_mask[19])
  );
  AND2_X1 _12018_ (
    .A1(reg_pmp_0_addr[17]),
    .A2(io_pmp_0_mask[19]),
    .ZN(io_pmp_0_mask[20])
  );
  AND2_X1 _12019_ (
    .A1(reg_pmp_0_addr[18]),
    .A2(io_pmp_0_mask[20]),
    .ZN(io_pmp_0_mask[21])
  );
  AND2_X1 _12020_ (
    .A1(reg_pmp_0_addr[19]),
    .A2(io_pmp_0_mask[21]),
    .ZN(io_pmp_0_mask[22])
  );
  AND2_X1 _12021_ (
    .A1(reg_pmp_0_addr[20]),
    .A2(io_pmp_0_mask[22]),
    .ZN(io_pmp_0_mask[23])
  );
  AND2_X1 _12022_ (
    .A1(reg_pmp_0_addr[21]),
    .A2(io_pmp_0_mask[23]),
    .ZN(io_pmp_0_mask[24])
  );
  AND2_X1 _12023_ (
    .A1(reg_pmp_0_addr[22]),
    .A2(io_pmp_0_mask[24]),
    .ZN(io_pmp_0_mask[25])
  );
  AND2_X1 _12024_ (
    .A1(reg_pmp_0_addr[23]),
    .A2(io_pmp_0_mask[25]),
    .ZN(io_pmp_0_mask[26])
  );
  AND2_X1 _12025_ (
    .A1(reg_pmp_0_addr[24]),
    .A2(io_pmp_0_mask[26]),
    .ZN(io_pmp_0_mask[27])
  );
  AND2_X1 _12026_ (
    .A1(reg_pmp_0_addr[25]),
    .A2(io_pmp_0_mask[27]),
    .ZN(io_pmp_0_mask[28])
  );
  AND2_X1 _12027_ (
    .A1(reg_pmp_0_addr[26]),
    .A2(io_pmp_0_mask[28]),
    .ZN(io_pmp_0_mask[29])
  );
  AND2_X1 _12028_ (
    .A1(reg_pmp_0_addr[27]),
    .A2(io_pmp_0_mask[29]),
    .ZN(io_pmp_0_mask[30])
  );
  AND2_X1 _12029_ (
    .A1(reg_pmp_0_addr[28]),
    .A2(io_pmp_0_mask[30]),
    .ZN(io_pmp_0_mask[31])
  );
  AND2_X1 _12030_ (
    .A1(reg_pmp_1_cfg_a[0]),
    .A2(reg_pmp_1_addr[0]),
    .ZN(io_pmp_1_mask[3])
  );
  AND2_X1 _12031_ (
    .A1(reg_pmp_1_addr[1]),
    .A2(io_pmp_1_mask[3]),
    .ZN(io_pmp_1_mask[4])
  );
  AND2_X1 _12032_ (
    .A1(reg_pmp_1_addr[2]),
    .A2(io_pmp_1_mask[4]),
    .ZN(io_pmp_1_mask[5])
  );
  AND2_X1 _12033_ (
    .A1(reg_pmp_1_addr[3]),
    .A2(io_pmp_1_mask[5]),
    .ZN(io_pmp_1_mask[6])
  );
  AND2_X1 _12034_ (
    .A1(reg_pmp_1_addr[4]),
    .A2(io_pmp_1_mask[6]),
    .ZN(io_pmp_1_mask[7])
  );
  AND2_X1 _12035_ (
    .A1(reg_pmp_1_addr[5]),
    .A2(io_pmp_1_mask[7]),
    .ZN(io_pmp_1_mask[8])
  );
  AND2_X1 _12036_ (
    .A1(reg_pmp_1_addr[6]),
    .A2(io_pmp_1_mask[8]),
    .ZN(io_pmp_1_mask[9])
  );
  AND2_X1 _12037_ (
    .A1(reg_pmp_1_addr[7]),
    .A2(io_pmp_1_mask[9]),
    .ZN(io_pmp_1_mask[10])
  );
  AND2_X1 _12038_ (
    .A1(reg_pmp_1_addr[8]),
    .A2(io_pmp_1_mask[10]),
    .ZN(io_pmp_1_mask[11])
  );
  AND2_X1 _12039_ (
    .A1(reg_pmp_1_addr[9]),
    .A2(io_pmp_1_mask[11]),
    .ZN(io_pmp_1_mask[12])
  );
  AND2_X1 _12040_ (
    .A1(reg_pmp_1_addr[10]),
    .A2(io_pmp_1_mask[12]),
    .ZN(io_pmp_1_mask[13])
  );
  AND2_X1 _12041_ (
    .A1(reg_pmp_1_addr[11]),
    .A2(io_pmp_1_mask[13]),
    .ZN(io_pmp_1_mask[14])
  );
  AND2_X1 _12042_ (
    .A1(reg_pmp_1_addr[12]),
    .A2(io_pmp_1_mask[14]),
    .ZN(io_pmp_1_mask[15])
  );
  AND2_X1 _12043_ (
    .A1(reg_pmp_1_addr[13]),
    .A2(io_pmp_1_mask[15]),
    .ZN(io_pmp_1_mask[16])
  );
  AND2_X1 _12044_ (
    .A1(reg_pmp_1_addr[14]),
    .A2(io_pmp_1_mask[16]),
    .ZN(io_pmp_1_mask[17])
  );
  AND2_X1 _12045_ (
    .A1(reg_pmp_1_addr[15]),
    .A2(io_pmp_1_mask[17]),
    .ZN(io_pmp_1_mask[18])
  );
  AND2_X1 _12046_ (
    .A1(reg_pmp_1_addr[16]),
    .A2(io_pmp_1_mask[18]),
    .ZN(io_pmp_1_mask[19])
  );
  AND2_X1 _12047_ (
    .A1(reg_pmp_1_addr[17]),
    .A2(io_pmp_1_mask[19]),
    .ZN(io_pmp_1_mask[20])
  );
  AND2_X1 _12048_ (
    .A1(reg_pmp_1_addr[18]),
    .A2(io_pmp_1_mask[20]),
    .ZN(io_pmp_1_mask[21])
  );
  AND2_X1 _12049_ (
    .A1(reg_pmp_1_addr[19]),
    .A2(io_pmp_1_mask[21]),
    .ZN(io_pmp_1_mask[22])
  );
  AND2_X1 _12050_ (
    .A1(reg_pmp_1_addr[20]),
    .A2(io_pmp_1_mask[22]),
    .ZN(io_pmp_1_mask[23])
  );
  AND2_X1 _12051_ (
    .A1(reg_pmp_1_addr[21]),
    .A2(io_pmp_1_mask[23]),
    .ZN(io_pmp_1_mask[24])
  );
  AND2_X1 _12052_ (
    .A1(reg_pmp_1_addr[22]),
    .A2(io_pmp_1_mask[24]),
    .ZN(io_pmp_1_mask[25])
  );
  AND2_X1 _12053_ (
    .A1(reg_pmp_1_addr[23]),
    .A2(io_pmp_1_mask[25]),
    .ZN(io_pmp_1_mask[26])
  );
  AND2_X1 _12054_ (
    .A1(reg_pmp_1_addr[24]),
    .A2(io_pmp_1_mask[26]),
    .ZN(io_pmp_1_mask[27])
  );
  AND2_X1 _12055_ (
    .A1(reg_pmp_1_addr[25]),
    .A2(io_pmp_1_mask[27]),
    .ZN(io_pmp_1_mask[28])
  );
  AND2_X1 _12056_ (
    .A1(reg_pmp_1_addr[26]),
    .A2(io_pmp_1_mask[28]),
    .ZN(io_pmp_1_mask[29])
  );
  AND2_X1 _12057_ (
    .A1(reg_pmp_1_addr[27]),
    .A2(io_pmp_1_mask[29]),
    .ZN(io_pmp_1_mask[30])
  );
  AND2_X1 _12058_ (
    .A1(reg_pmp_1_addr[28]),
    .A2(io_pmp_1_mask[30]),
    .ZN(io_pmp_1_mask[31])
  );
  AND2_X1 _12059_ (
    .A1(reg_pmp_2_cfg_a[0]),
    .A2(reg_pmp_2_addr[0]),
    .ZN(io_pmp_2_mask[3])
  );
  AND2_X1 _12060_ (
    .A1(reg_pmp_2_addr[1]),
    .A2(io_pmp_2_mask[3]),
    .ZN(io_pmp_2_mask[4])
  );
  AND2_X1 _12061_ (
    .A1(reg_pmp_2_addr[2]),
    .A2(io_pmp_2_mask[4]),
    .ZN(io_pmp_2_mask[5])
  );
  AND2_X1 _12062_ (
    .A1(reg_pmp_2_addr[3]),
    .A2(io_pmp_2_mask[5]),
    .ZN(io_pmp_2_mask[6])
  );
  AND2_X1 _12063_ (
    .A1(reg_pmp_2_addr[4]),
    .A2(io_pmp_2_mask[6]),
    .ZN(io_pmp_2_mask[7])
  );
  AND2_X1 _12064_ (
    .A1(reg_pmp_2_addr[5]),
    .A2(io_pmp_2_mask[7]),
    .ZN(io_pmp_2_mask[8])
  );
  AND2_X1 _12065_ (
    .A1(reg_pmp_2_addr[6]),
    .A2(io_pmp_2_mask[8]),
    .ZN(io_pmp_2_mask[9])
  );
  AND2_X1 _12066_ (
    .A1(reg_pmp_2_addr[7]),
    .A2(io_pmp_2_mask[9]),
    .ZN(io_pmp_2_mask[10])
  );
  AND2_X1 _12067_ (
    .A1(reg_pmp_2_addr[8]),
    .A2(io_pmp_2_mask[10]),
    .ZN(io_pmp_2_mask[11])
  );
  AND2_X1 _12068_ (
    .A1(reg_pmp_2_addr[9]),
    .A2(io_pmp_2_mask[11]),
    .ZN(io_pmp_2_mask[12])
  );
  AND2_X1 _12069_ (
    .A1(reg_pmp_2_addr[10]),
    .A2(io_pmp_2_mask[12]),
    .ZN(io_pmp_2_mask[13])
  );
  AND2_X1 _12070_ (
    .A1(reg_pmp_2_addr[11]),
    .A2(io_pmp_2_mask[13]),
    .ZN(io_pmp_2_mask[14])
  );
  AND2_X1 _12071_ (
    .A1(reg_pmp_2_addr[12]),
    .A2(io_pmp_2_mask[14]),
    .ZN(io_pmp_2_mask[15])
  );
  AND2_X1 _12072_ (
    .A1(reg_pmp_2_addr[13]),
    .A2(io_pmp_2_mask[15]),
    .ZN(io_pmp_2_mask[16])
  );
  AND2_X1 _12073_ (
    .A1(reg_pmp_2_addr[14]),
    .A2(io_pmp_2_mask[16]),
    .ZN(io_pmp_2_mask[17])
  );
  AND2_X1 _12074_ (
    .A1(reg_pmp_2_addr[15]),
    .A2(io_pmp_2_mask[17]),
    .ZN(io_pmp_2_mask[18])
  );
  AND2_X1 _12075_ (
    .A1(reg_pmp_2_addr[16]),
    .A2(io_pmp_2_mask[18]),
    .ZN(io_pmp_2_mask[19])
  );
  AND2_X1 _12076_ (
    .A1(reg_pmp_2_addr[17]),
    .A2(io_pmp_2_mask[19]),
    .ZN(io_pmp_2_mask[20])
  );
  AND2_X1 _12077_ (
    .A1(reg_pmp_2_addr[18]),
    .A2(io_pmp_2_mask[20]),
    .ZN(io_pmp_2_mask[21])
  );
  AND2_X1 _12078_ (
    .A1(reg_pmp_2_addr[19]),
    .A2(io_pmp_2_mask[21]),
    .ZN(io_pmp_2_mask[22])
  );
  AND2_X1 _12079_ (
    .A1(reg_pmp_2_addr[20]),
    .A2(io_pmp_2_mask[22]),
    .ZN(io_pmp_2_mask[23])
  );
  AND2_X1 _12080_ (
    .A1(reg_pmp_2_addr[21]),
    .A2(io_pmp_2_mask[23]),
    .ZN(io_pmp_2_mask[24])
  );
  AND2_X1 _12081_ (
    .A1(reg_pmp_2_addr[22]),
    .A2(io_pmp_2_mask[24]),
    .ZN(io_pmp_2_mask[25])
  );
  AND2_X1 _12082_ (
    .A1(reg_pmp_2_addr[23]),
    .A2(io_pmp_2_mask[25]),
    .ZN(io_pmp_2_mask[26])
  );
  AND2_X1 _12083_ (
    .A1(reg_pmp_2_addr[24]),
    .A2(io_pmp_2_mask[26]),
    .ZN(io_pmp_2_mask[27])
  );
  AND2_X1 _12084_ (
    .A1(reg_pmp_2_addr[25]),
    .A2(io_pmp_2_mask[27]),
    .ZN(io_pmp_2_mask[28])
  );
  AND2_X1 _12085_ (
    .A1(reg_pmp_2_addr[26]),
    .A2(io_pmp_2_mask[28]),
    .ZN(io_pmp_2_mask[29])
  );
  AND2_X1 _12086_ (
    .A1(reg_pmp_2_addr[27]),
    .A2(io_pmp_2_mask[29]),
    .ZN(io_pmp_2_mask[30])
  );
  AND2_X1 _12087_ (
    .A1(reg_pmp_2_addr[28]),
    .A2(io_pmp_2_mask[30]),
    .ZN(io_pmp_2_mask[31])
  );
  AND2_X1 _12088_ (
    .A1(reg_pmp_3_cfg_a[0]),
    .A2(reg_pmp_3_addr[0]),
    .ZN(io_pmp_3_mask[3])
  );
  AND2_X1 _12089_ (
    .A1(reg_pmp_3_addr[1]),
    .A2(io_pmp_3_mask[3]),
    .ZN(io_pmp_3_mask[4])
  );
  AND2_X1 _12090_ (
    .A1(reg_pmp_3_addr[2]),
    .A2(io_pmp_3_mask[4]),
    .ZN(io_pmp_3_mask[5])
  );
  AND2_X1 _12091_ (
    .A1(reg_pmp_3_addr[3]),
    .A2(io_pmp_3_mask[5]),
    .ZN(io_pmp_3_mask[6])
  );
  AND2_X1 _12092_ (
    .A1(reg_pmp_3_addr[4]),
    .A2(io_pmp_3_mask[6]),
    .ZN(io_pmp_3_mask[7])
  );
  AND2_X1 _12093_ (
    .A1(reg_pmp_3_addr[5]),
    .A2(io_pmp_3_mask[7]),
    .ZN(io_pmp_3_mask[8])
  );
  AND2_X1 _12094_ (
    .A1(reg_pmp_3_addr[6]),
    .A2(io_pmp_3_mask[8]),
    .ZN(io_pmp_3_mask[9])
  );
  AND2_X1 _12095_ (
    .A1(reg_pmp_3_addr[7]),
    .A2(io_pmp_3_mask[9]),
    .ZN(io_pmp_3_mask[10])
  );
  AND2_X1 _12096_ (
    .A1(reg_pmp_3_addr[8]),
    .A2(io_pmp_3_mask[10]),
    .ZN(io_pmp_3_mask[11])
  );
  AND2_X1 _12097_ (
    .A1(reg_pmp_3_addr[9]),
    .A2(io_pmp_3_mask[11]),
    .ZN(io_pmp_3_mask[12])
  );
  AND2_X1 _12098_ (
    .A1(reg_pmp_3_addr[10]),
    .A2(io_pmp_3_mask[12]),
    .ZN(io_pmp_3_mask[13])
  );
  AND2_X1 _12099_ (
    .A1(reg_pmp_3_addr[11]),
    .A2(io_pmp_3_mask[13]),
    .ZN(io_pmp_3_mask[14])
  );
  AND2_X1 _12100_ (
    .A1(reg_pmp_3_addr[12]),
    .A2(io_pmp_3_mask[14]),
    .ZN(io_pmp_3_mask[15])
  );
  AND2_X1 _12101_ (
    .A1(reg_pmp_3_addr[13]),
    .A2(io_pmp_3_mask[15]),
    .ZN(io_pmp_3_mask[16])
  );
  AND2_X1 _12102_ (
    .A1(reg_pmp_3_addr[14]),
    .A2(io_pmp_3_mask[16]),
    .ZN(io_pmp_3_mask[17])
  );
  AND2_X1 _12103_ (
    .A1(reg_pmp_3_addr[15]),
    .A2(io_pmp_3_mask[17]),
    .ZN(io_pmp_3_mask[18])
  );
  AND2_X1 _12104_ (
    .A1(reg_pmp_3_addr[16]),
    .A2(io_pmp_3_mask[18]),
    .ZN(io_pmp_3_mask[19])
  );
  AND2_X1 _12105_ (
    .A1(reg_pmp_3_addr[17]),
    .A2(io_pmp_3_mask[19]),
    .ZN(io_pmp_3_mask[20])
  );
  AND2_X1 _12106_ (
    .A1(reg_pmp_3_addr[18]),
    .A2(io_pmp_3_mask[20]),
    .ZN(io_pmp_3_mask[21])
  );
  AND2_X1 _12107_ (
    .A1(reg_pmp_3_addr[19]),
    .A2(io_pmp_3_mask[21]),
    .ZN(io_pmp_3_mask[22])
  );
  AND2_X1 _12108_ (
    .A1(reg_pmp_3_addr[20]),
    .A2(io_pmp_3_mask[22]),
    .ZN(io_pmp_3_mask[23])
  );
  AND2_X1 _12109_ (
    .A1(reg_pmp_3_addr[21]),
    .A2(io_pmp_3_mask[23]),
    .ZN(io_pmp_3_mask[24])
  );
  AND2_X1 _12110_ (
    .A1(reg_pmp_3_addr[22]),
    .A2(io_pmp_3_mask[24]),
    .ZN(io_pmp_3_mask[25])
  );
  AND2_X1 _12111_ (
    .A1(reg_pmp_3_addr[23]),
    .A2(io_pmp_3_mask[25]),
    .ZN(io_pmp_3_mask[26])
  );
  AND2_X1 _12112_ (
    .A1(reg_pmp_3_addr[24]),
    .A2(io_pmp_3_mask[26]),
    .ZN(io_pmp_3_mask[27])
  );
  AND2_X1 _12113_ (
    .A1(reg_pmp_3_addr[25]),
    .A2(io_pmp_3_mask[27]),
    .ZN(io_pmp_3_mask[28])
  );
  AND2_X1 _12114_ (
    .A1(reg_pmp_3_addr[26]),
    .A2(io_pmp_3_mask[28]),
    .ZN(io_pmp_3_mask[29])
  );
  AND2_X1 _12115_ (
    .A1(reg_pmp_3_addr[27]),
    .A2(io_pmp_3_mask[29]),
    .ZN(io_pmp_3_mask[30])
  );
  AND2_X1 _12116_ (
    .A1(reg_pmp_3_addr[28]),
    .A2(io_pmp_3_mask[30]),
    .ZN(io_pmp_3_mask[31])
  );
  AND2_X1 _12117_ (
    .A1(reg_pmp_4_cfg_a[0]),
    .A2(reg_pmp_4_addr[0]),
    .ZN(io_pmp_4_mask[3])
  );
  AND2_X1 _12118_ (
    .A1(reg_pmp_4_addr[1]),
    .A2(io_pmp_4_mask[3]),
    .ZN(io_pmp_4_mask[4])
  );
  AND2_X1 _12119_ (
    .A1(reg_pmp_4_addr[2]),
    .A2(io_pmp_4_mask[4]),
    .ZN(io_pmp_4_mask[5])
  );
  AND2_X1 _12120_ (
    .A1(reg_pmp_4_addr[3]),
    .A2(io_pmp_4_mask[5]),
    .ZN(io_pmp_4_mask[6])
  );
  AND2_X1 _12121_ (
    .A1(reg_pmp_4_addr[4]),
    .A2(io_pmp_4_mask[6]),
    .ZN(io_pmp_4_mask[7])
  );
  AND2_X1 _12122_ (
    .A1(reg_pmp_4_addr[5]),
    .A2(io_pmp_4_mask[7]),
    .ZN(io_pmp_4_mask[8])
  );
  AND2_X1 _12123_ (
    .A1(reg_pmp_4_addr[6]),
    .A2(io_pmp_4_mask[8]),
    .ZN(io_pmp_4_mask[9])
  );
  AND2_X1 _12124_ (
    .A1(reg_pmp_4_addr[7]),
    .A2(io_pmp_4_mask[9]),
    .ZN(io_pmp_4_mask[10])
  );
  AND2_X1 _12125_ (
    .A1(reg_pmp_4_addr[8]),
    .A2(io_pmp_4_mask[10]),
    .ZN(io_pmp_4_mask[11])
  );
  AND2_X1 _12126_ (
    .A1(reg_pmp_4_addr[9]),
    .A2(io_pmp_4_mask[11]),
    .ZN(io_pmp_4_mask[12])
  );
  AND2_X1 _12127_ (
    .A1(reg_pmp_4_addr[10]),
    .A2(io_pmp_4_mask[12]),
    .ZN(io_pmp_4_mask[13])
  );
  AND2_X1 _12128_ (
    .A1(reg_pmp_4_addr[11]),
    .A2(io_pmp_4_mask[13]),
    .ZN(io_pmp_4_mask[14])
  );
  AND2_X1 _12129_ (
    .A1(reg_pmp_4_addr[12]),
    .A2(io_pmp_4_mask[14]),
    .ZN(io_pmp_4_mask[15])
  );
  AND2_X1 _12130_ (
    .A1(reg_pmp_4_addr[13]),
    .A2(io_pmp_4_mask[15]),
    .ZN(io_pmp_4_mask[16])
  );
  AND2_X1 _12131_ (
    .A1(reg_pmp_4_addr[14]),
    .A2(io_pmp_4_mask[16]),
    .ZN(io_pmp_4_mask[17])
  );
  AND2_X1 _12132_ (
    .A1(reg_pmp_4_addr[15]),
    .A2(io_pmp_4_mask[17]),
    .ZN(io_pmp_4_mask[18])
  );
  AND2_X1 _12133_ (
    .A1(reg_pmp_4_addr[16]),
    .A2(io_pmp_4_mask[18]),
    .ZN(io_pmp_4_mask[19])
  );
  AND2_X1 _12134_ (
    .A1(reg_pmp_4_addr[17]),
    .A2(io_pmp_4_mask[19]),
    .ZN(io_pmp_4_mask[20])
  );
  AND2_X1 _12135_ (
    .A1(reg_pmp_4_addr[18]),
    .A2(io_pmp_4_mask[20]),
    .ZN(io_pmp_4_mask[21])
  );
  AND2_X1 _12136_ (
    .A1(reg_pmp_4_addr[19]),
    .A2(io_pmp_4_mask[21]),
    .ZN(io_pmp_4_mask[22])
  );
  AND2_X1 _12137_ (
    .A1(reg_pmp_4_addr[20]),
    .A2(io_pmp_4_mask[22]),
    .ZN(io_pmp_4_mask[23])
  );
  AND2_X1 _12138_ (
    .A1(reg_pmp_4_addr[21]),
    .A2(io_pmp_4_mask[23]),
    .ZN(io_pmp_4_mask[24])
  );
  AND2_X1 _12139_ (
    .A1(reg_pmp_4_addr[22]),
    .A2(io_pmp_4_mask[24]),
    .ZN(io_pmp_4_mask[25])
  );
  AND2_X1 _12140_ (
    .A1(reg_pmp_4_addr[23]),
    .A2(io_pmp_4_mask[25]),
    .ZN(io_pmp_4_mask[26])
  );
  AND2_X1 _12141_ (
    .A1(reg_pmp_4_addr[24]),
    .A2(io_pmp_4_mask[26]),
    .ZN(io_pmp_4_mask[27])
  );
  AND2_X1 _12142_ (
    .A1(reg_pmp_4_addr[25]),
    .A2(io_pmp_4_mask[27]),
    .ZN(io_pmp_4_mask[28])
  );
  AND2_X1 _12143_ (
    .A1(reg_pmp_4_addr[26]),
    .A2(io_pmp_4_mask[28]),
    .ZN(io_pmp_4_mask[29])
  );
  AND2_X1 _12144_ (
    .A1(reg_pmp_4_addr[27]),
    .A2(io_pmp_4_mask[29]),
    .ZN(io_pmp_4_mask[30])
  );
  AND2_X1 _12145_ (
    .A1(reg_pmp_4_addr[28]),
    .A2(io_pmp_4_mask[30]),
    .ZN(io_pmp_4_mask[31])
  );
  AND2_X1 _12146_ (
    .A1(reg_pmp_5_cfg_a[0]),
    .A2(reg_pmp_5_addr[0]),
    .ZN(io_pmp_5_mask[3])
  );
  AND2_X1 _12147_ (
    .A1(reg_pmp_5_addr[1]),
    .A2(io_pmp_5_mask[3]),
    .ZN(io_pmp_5_mask[4])
  );
  AND2_X1 _12148_ (
    .A1(reg_pmp_5_addr[2]),
    .A2(io_pmp_5_mask[4]),
    .ZN(io_pmp_5_mask[5])
  );
  AND2_X1 _12149_ (
    .A1(reg_pmp_5_addr[3]),
    .A2(io_pmp_5_mask[5]),
    .ZN(io_pmp_5_mask[6])
  );
  AND2_X1 _12150_ (
    .A1(reg_pmp_5_addr[4]),
    .A2(io_pmp_5_mask[6]),
    .ZN(io_pmp_5_mask[7])
  );
  AND2_X1 _12151_ (
    .A1(reg_pmp_5_addr[5]),
    .A2(io_pmp_5_mask[7]),
    .ZN(io_pmp_5_mask[8])
  );
  AND2_X1 _12152_ (
    .A1(reg_pmp_5_addr[6]),
    .A2(io_pmp_5_mask[8]),
    .ZN(io_pmp_5_mask[9])
  );
  AND2_X1 _12153_ (
    .A1(reg_pmp_5_addr[7]),
    .A2(io_pmp_5_mask[9]),
    .ZN(io_pmp_5_mask[10])
  );
  AND2_X1 _12154_ (
    .A1(reg_pmp_5_addr[8]),
    .A2(io_pmp_5_mask[10]),
    .ZN(io_pmp_5_mask[11])
  );
  AND2_X1 _12155_ (
    .A1(reg_pmp_5_addr[9]),
    .A2(io_pmp_5_mask[11]),
    .ZN(io_pmp_5_mask[12])
  );
  AND2_X1 _12156_ (
    .A1(reg_pmp_5_addr[10]),
    .A2(io_pmp_5_mask[12]),
    .ZN(io_pmp_5_mask[13])
  );
  AND2_X1 _12157_ (
    .A1(reg_pmp_5_addr[11]),
    .A2(io_pmp_5_mask[13]),
    .ZN(io_pmp_5_mask[14])
  );
  AND2_X1 _12158_ (
    .A1(reg_pmp_5_addr[12]),
    .A2(io_pmp_5_mask[14]),
    .ZN(io_pmp_5_mask[15])
  );
  AND2_X1 _12159_ (
    .A1(reg_pmp_5_addr[13]),
    .A2(io_pmp_5_mask[15]),
    .ZN(io_pmp_5_mask[16])
  );
  AND2_X1 _12160_ (
    .A1(reg_pmp_5_addr[14]),
    .A2(io_pmp_5_mask[16]),
    .ZN(io_pmp_5_mask[17])
  );
  AND2_X1 _12161_ (
    .A1(reg_pmp_5_addr[15]),
    .A2(io_pmp_5_mask[17]),
    .ZN(io_pmp_5_mask[18])
  );
  AND2_X1 _12162_ (
    .A1(reg_pmp_5_addr[16]),
    .A2(io_pmp_5_mask[18]),
    .ZN(io_pmp_5_mask[19])
  );
  AND2_X1 _12163_ (
    .A1(reg_pmp_5_addr[17]),
    .A2(io_pmp_5_mask[19]),
    .ZN(io_pmp_5_mask[20])
  );
  AND2_X1 _12164_ (
    .A1(reg_pmp_5_addr[18]),
    .A2(io_pmp_5_mask[20]),
    .ZN(io_pmp_5_mask[21])
  );
  AND2_X1 _12165_ (
    .A1(reg_pmp_5_addr[19]),
    .A2(io_pmp_5_mask[21]),
    .ZN(io_pmp_5_mask[22])
  );
  AND2_X1 _12166_ (
    .A1(reg_pmp_5_addr[20]),
    .A2(io_pmp_5_mask[22]),
    .ZN(io_pmp_5_mask[23])
  );
  AND2_X1 _12167_ (
    .A1(reg_pmp_5_addr[21]),
    .A2(io_pmp_5_mask[23]),
    .ZN(io_pmp_5_mask[24])
  );
  AND2_X1 _12168_ (
    .A1(reg_pmp_5_addr[22]),
    .A2(io_pmp_5_mask[24]),
    .ZN(io_pmp_5_mask[25])
  );
  AND2_X1 _12169_ (
    .A1(reg_pmp_5_addr[23]),
    .A2(io_pmp_5_mask[25]),
    .ZN(io_pmp_5_mask[26])
  );
  AND2_X1 _12170_ (
    .A1(reg_pmp_5_addr[24]),
    .A2(io_pmp_5_mask[26]),
    .ZN(io_pmp_5_mask[27])
  );
  AND2_X1 _12171_ (
    .A1(reg_pmp_5_addr[25]),
    .A2(io_pmp_5_mask[27]),
    .ZN(io_pmp_5_mask[28])
  );
  AND2_X1 _12172_ (
    .A1(reg_pmp_5_addr[26]),
    .A2(io_pmp_5_mask[28]),
    .ZN(io_pmp_5_mask[29])
  );
  AND2_X1 _12173_ (
    .A1(reg_pmp_5_addr[27]),
    .A2(io_pmp_5_mask[29]),
    .ZN(io_pmp_5_mask[30])
  );
  AND2_X1 _12174_ (
    .A1(reg_pmp_5_addr[28]),
    .A2(io_pmp_5_mask[30]),
    .ZN(io_pmp_5_mask[31])
  );
  AND2_X1 _12175_ (
    .A1(reg_pmp_6_cfg_a[0]),
    .A2(reg_pmp_6_addr[0]),
    .ZN(io_pmp_6_mask[3])
  );
  AND2_X1 _12176_ (
    .A1(reg_pmp_6_addr[1]),
    .A2(io_pmp_6_mask[3]),
    .ZN(io_pmp_6_mask[4])
  );
  AND2_X1 _12177_ (
    .A1(reg_pmp_6_addr[2]),
    .A2(io_pmp_6_mask[4]),
    .ZN(io_pmp_6_mask[5])
  );
  AND2_X1 _12178_ (
    .A1(reg_pmp_6_addr[3]),
    .A2(io_pmp_6_mask[5]),
    .ZN(io_pmp_6_mask[6])
  );
  AND2_X1 _12179_ (
    .A1(reg_pmp_6_addr[4]),
    .A2(io_pmp_6_mask[6]),
    .ZN(io_pmp_6_mask[7])
  );
  AND2_X1 _12180_ (
    .A1(reg_pmp_6_addr[5]),
    .A2(io_pmp_6_mask[7]),
    .ZN(io_pmp_6_mask[8])
  );
  AND2_X1 _12181_ (
    .A1(reg_pmp_6_addr[6]),
    .A2(io_pmp_6_mask[8]),
    .ZN(io_pmp_6_mask[9])
  );
  AND2_X1 _12182_ (
    .A1(reg_pmp_6_addr[7]),
    .A2(io_pmp_6_mask[9]),
    .ZN(io_pmp_6_mask[10])
  );
  AND2_X1 _12183_ (
    .A1(reg_pmp_6_addr[8]),
    .A2(io_pmp_6_mask[10]),
    .ZN(io_pmp_6_mask[11])
  );
  AND2_X1 _12184_ (
    .A1(reg_pmp_6_addr[9]),
    .A2(io_pmp_6_mask[11]),
    .ZN(io_pmp_6_mask[12])
  );
  AND2_X1 _12185_ (
    .A1(reg_pmp_6_addr[10]),
    .A2(io_pmp_6_mask[12]),
    .ZN(io_pmp_6_mask[13])
  );
  AND2_X1 _12186_ (
    .A1(reg_pmp_6_addr[11]),
    .A2(io_pmp_6_mask[13]),
    .ZN(io_pmp_6_mask[14])
  );
  AND2_X1 _12187_ (
    .A1(reg_pmp_6_addr[12]),
    .A2(io_pmp_6_mask[14]),
    .ZN(io_pmp_6_mask[15])
  );
  AND2_X1 _12188_ (
    .A1(reg_pmp_6_addr[13]),
    .A2(io_pmp_6_mask[15]),
    .ZN(io_pmp_6_mask[16])
  );
  AND2_X1 _12189_ (
    .A1(reg_pmp_6_addr[14]),
    .A2(io_pmp_6_mask[16]),
    .ZN(io_pmp_6_mask[17])
  );
  AND2_X1 _12190_ (
    .A1(reg_pmp_6_addr[15]),
    .A2(io_pmp_6_mask[17]),
    .ZN(io_pmp_6_mask[18])
  );
  AND2_X1 _12191_ (
    .A1(reg_pmp_6_addr[16]),
    .A2(io_pmp_6_mask[18]),
    .ZN(io_pmp_6_mask[19])
  );
  AND2_X1 _12192_ (
    .A1(reg_pmp_6_addr[17]),
    .A2(io_pmp_6_mask[19]),
    .ZN(io_pmp_6_mask[20])
  );
  AND2_X1 _12193_ (
    .A1(reg_pmp_6_addr[18]),
    .A2(io_pmp_6_mask[20]),
    .ZN(io_pmp_6_mask[21])
  );
  AND2_X1 _12194_ (
    .A1(reg_pmp_6_addr[19]),
    .A2(io_pmp_6_mask[21]),
    .ZN(io_pmp_6_mask[22])
  );
  AND2_X1 _12195_ (
    .A1(reg_pmp_6_addr[20]),
    .A2(io_pmp_6_mask[22]),
    .ZN(io_pmp_6_mask[23])
  );
  AND2_X1 _12196_ (
    .A1(reg_pmp_6_addr[21]),
    .A2(io_pmp_6_mask[23]),
    .ZN(io_pmp_6_mask[24])
  );
  AND2_X1 _12197_ (
    .A1(reg_pmp_6_addr[22]),
    .A2(io_pmp_6_mask[24]),
    .ZN(io_pmp_6_mask[25])
  );
  AND2_X1 _12198_ (
    .A1(reg_pmp_6_addr[23]),
    .A2(io_pmp_6_mask[25]),
    .ZN(io_pmp_6_mask[26])
  );
  AND2_X1 _12199_ (
    .A1(reg_pmp_6_addr[24]),
    .A2(io_pmp_6_mask[26]),
    .ZN(io_pmp_6_mask[27])
  );
  AND2_X1 _12200_ (
    .A1(reg_pmp_6_addr[25]),
    .A2(io_pmp_6_mask[27]),
    .ZN(io_pmp_6_mask[28])
  );
  AND2_X1 _12201_ (
    .A1(reg_pmp_6_addr[26]),
    .A2(io_pmp_6_mask[28]),
    .ZN(io_pmp_6_mask[29])
  );
  AND2_X1 _12202_ (
    .A1(reg_pmp_6_addr[27]),
    .A2(io_pmp_6_mask[29]),
    .ZN(io_pmp_6_mask[30])
  );
  AND2_X1 _12203_ (
    .A1(reg_pmp_6_addr[28]),
    .A2(io_pmp_6_mask[30]),
    .ZN(io_pmp_6_mask[31])
  );
  AND2_X1 _12204_ (
    .A1(reg_pmp_7_cfg_a[0]),
    .A2(reg_pmp_7_addr[0]),
    .ZN(io_pmp_7_mask[3])
  );
  AND2_X1 _12205_ (
    .A1(reg_pmp_7_addr[1]),
    .A2(io_pmp_7_mask[3]),
    .ZN(io_pmp_7_mask[4])
  );
  AND2_X1 _12206_ (
    .A1(reg_pmp_7_addr[2]),
    .A2(io_pmp_7_mask[4]),
    .ZN(io_pmp_7_mask[5])
  );
  AND2_X1 _12207_ (
    .A1(reg_pmp_7_addr[3]),
    .A2(io_pmp_7_mask[5]),
    .ZN(io_pmp_7_mask[6])
  );
  AND2_X1 _12208_ (
    .A1(reg_pmp_7_addr[4]),
    .A2(io_pmp_7_mask[6]),
    .ZN(io_pmp_7_mask[7])
  );
  AND2_X1 _12209_ (
    .A1(reg_pmp_7_addr[5]),
    .A2(io_pmp_7_mask[7]),
    .ZN(io_pmp_7_mask[8])
  );
  AND2_X1 _12210_ (
    .A1(reg_pmp_7_addr[6]),
    .A2(io_pmp_7_mask[8]),
    .ZN(io_pmp_7_mask[9])
  );
  AND2_X1 _12211_ (
    .A1(reg_pmp_7_addr[7]),
    .A2(io_pmp_7_mask[9]),
    .ZN(io_pmp_7_mask[10])
  );
  AND2_X1 _12212_ (
    .A1(reg_pmp_7_addr[8]),
    .A2(io_pmp_7_mask[10]),
    .ZN(io_pmp_7_mask[11])
  );
  AND2_X1 _12213_ (
    .A1(reg_pmp_7_addr[9]),
    .A2(io_pmp_7_mask[11]),
    .ZN(io_pmp_7_mask[12])
  );
  AND2_X1 _12214_ (
    .A1(reg_pmp_7_addr[10]),
    .A2(io_pmp_7_mask[12]),
    .ZN(io_pmp_7_mask[13])
  );
  AND2_X1 _12215_ (
    .A1(reg_pmp_7_addr[11]),
    .A2(io_pmp_7_mask[13]),
    .ZN(io_pmp_7_mask[14])
  );
  AND2_X1 _12216_ (
    .A1(reg_pmp_7_addr[12]),
    .A2(io_pmp_7_mask[14]),
    .ZN(io_pmp_7_mask[15])
  );
  AND2_X1 _12217_ (
    .A1(reg_pmp_7_addr[13]),
    .A2(io_pmp_7_mask[15]),
    .ZN(io_pmp_7_mask[16])
  );
  AND2_X1 _12218_ (
    .A1(reg_pmp_7_addr[14]),
    .A2(io_pmp_7_mask[16]),
    .ZN(io_pmp_7_mask[17])
  );
  AND2_X1 _12219_ (
    .A1(reg_pmp_7_addr[15]),
    .A2(io_pmp_7_mask[17]),
    .ZN(io_pmp_7_mask[18])
  );
  AND2_X1 _12220_ (
    .A1(reg_pmp_7_addr[16]),
    .A2(io_pmp_7_mask[18]),
    .ZN(io_pmp_7_mask[19])
  );
  AND2_X1 _12221_ (
    .A1(reg_pmp_7_addr[17]),
    .A2(io_pmp_7_mask[19]),
    .ZN(io_pmp_7_mask[20])
  );
  AND2_X1 _12222_ (
    .A1(reg_pmp_7_addr[18]),
    .A2(io_pmp_7_mask[20]),
    .ZN(io_pmp_7_mask[21])
  );
  AND2_X1 _12223_ (
    .A1(reg_pmp_7_addr[19]),
    .A2(io_pmp_7_mask[21]),
    .ZN(io_pmp_7_mask[22])
  );
  AND2_X1 _12224_ (
    .A1(reg_pmp_7_addr[20]),
    .A2(io_pmp_7_mask[22]),
    .ZN(io_pmp_7_mask[23])
  );
  AND2_X1 _12225_ (
    .A1(reg_pmp_7_addr[21]),
    .A2(io_pmp_7_mask[23]),
    .ZN(io_pmp_7_mask[24])
  );
  AND2_X1 _12226_ (
    .A1(reg_pmp_7_addr[22]),
    .A2(io_pmp_7_mask[24]),
    .ZN(io_pmp_7_mask[25])
  );
  AND2_X1 _12227_ (
    .A1(reg_pmp_7_addr[23]),
    .A2(io_pmp_7_mask[25]),
    .ZN(io_pmp_7_mask[26])
  );
  AND2_X1 _12228_ (
    .A1(reg_pmp_7_addr[24]),
    .A2(io_pmp_7_mask[26]),
    .ZN(io_pmp_7_mask[27])
  );
  AND2_X1 _12229_ (
    .A1(reg_pmp_7_addr[25]),
    .A2(io_pmp_7_mask[27]),
    .ZN(io_pmp_7_mask[28])
  );
  AND2_X1 _12230_ (
    .A1(reg_pmp_7_addr[26]),
    .A2(io_pmp_7_mask[28]),
    .ZN(io_pmp_7_mask[29])
  );
  AND2_X1 _12231_ (
    .A1(reg_pmp_7_addr[27]),
    .A2(io_pmp_7_mask[29]),
    .ZN(io_pmp_7_mask[30])
  );
  AND2_X1 _12232_ (
    .A1(reg_pmp_7_addr[28]),
    .A2(io_pmp_7_mask[30]),
    .ZN(io_pmp_7_mask[31])
  );
  AND2_X1 _12233_ (
    .A1(_00815_),
    .A2(io_decode_0_inst[27]),
    .ZN(_06334_)
  );
  AND2_X1 _12234_ (
    .A1(io_decode_0_inst[25]),
    .A2(_06334_),
    .ZN(_06335_)
  );
  AND2_X1 _12235_ (
    .A1(_06327_),
    .A2(_06335_),
    .ZN(_06336_)
  );
  INV_X1 _12236_ (
    .A(_06336_),
    .ZN(_06337_)
  );
  AND2_X1 _12237_ (
    .A1(io_decode_0_inst[21]),
    .A2(io_decode_0_inst[20]),
    .ZN(_06338_)
  );
  INV_X1 _12238_ (
    .A(_06338_),
    .ZN(_06339_)
  );
  AND2_X1 _12239_ (
    .A1(io_decode_0_inst[24]),
    .A2(_06338_),
    .ZN(_06340_)
  );
  INV_X1 _12240_ (
    .A(_06340_),
    .ZN(_06341_)
  );
  AND2_X1 _12241_ (
    .A1(_06336_),
    .A2(_06341_),
    .ZN(_06342_)
  );
  INV_X1 _12242_ (
    .A(_06342_),
    .ZN(_06343_)
  );
  AND2_X1 _12243_ (
    .A1(_00817_),
    .A2(io_decode_0_inst[20]),
    .ZN(_06344_)
  );
  AND2_X1 _12244_ (
    .A1(_06327_),
    .A2(_06344_),
    .ZN(_06345_)
  );
  AND2_X1 _12245_ (
    .A1(io_decode_0_inst[26]),
    .A2(io_decode_0_inst[27]),
    .ZN(_06346_)
  );
  AND2_X1 _12246_ (
    .A1(_06324_),
    .A2(_06346_),
    .ZN(_06347_)
  );
  AND2_X1 _12247_ (
    .A1(_06345_),
    .A2(_06347_),
    .ZN(_06348_)
  );
  INV_X1 _12248_ (
    .A(_06348_),
    .ZN(_06349_)
  );
  AND2_X1 _12249_ (
    .A1(io_decode_0_inst[30]),
    .A2(_06349_),
    .ZN(_06350_)
  );
  AND2_X1 _12250_ (
    .A1(_06343_),
    .A2(_06350_),
    .ZN(_06351_)
  );
  INV_X1 _12251_ (
    .A(_06351_),
    .ZN(_06352_)
  );
  AND2_X1 _12252_ (
    .A1(io_decode_0_inst[22]),
    .A2(_00819_),
    .ZN(_06353_)
  );
  MUX2_X1 _12253_ (
    .A(_00821_),
    .B(_06353_),
    .S(_00818_),
    .Z(_06354_)
  );
  AND2_X1 _12254_ (
    .A1(io_decode_0_inst[21]),
    .A2(_06354_),
    .ZN(_06355_)
  );
  INV_X1 _12255_ (
    .A(_06355_),
    .ZN(_06356_)
  );
  AND2_X1 _12256_ (
    .A1(_00821_),
    .A2(_06328_),
    .ZN(_06357_)
  );
  INV_X1 _12257_ (
    .A(_06357_),
    .ZN(_06358_)
  );
  AND2_X1 _12258_ (
    .A1(io_decode_0_inst[22]),
    .A2(io_decode_0_inst[23]),
    .ZN(_06359_)
  );
  AND2_X1 _12259_ (
    .A1(_06344_),
    .A2(_06359_),
    .ZN(_06360_)
  );
  INV_X1 _12260_ (
    .A(_06360_),
    .ZN(_06361_)
  );
  AND2_X1 _12261_ (
    .A1(_06358_),
    .A2(_06361_),
    .ZN(_06362_)
  );
  AND2_X1 _12262_ (
    .A1(_06356_),
    .A2(_06362_),
    .ZN(_06363_)
  );
  INV_X1 _12263_ (
    .A(_06363_),
    .ZN(_06364_)
  );
  AND2_X1 _12264_ (
    .A1(io_decode_0_inst[25]),
    .A2(_06364_),
    .ZN(_06365_)
  );
  INV_X1 _12265_ (
    .A(_06365_),
    .ZN(_06366_)
  );
  AND2_X1 _12266_ (
    .A1(_00817_),
    .A2(_00818_),
    .ZN(_06367_)
  );
  INV_X1 _12267_ (
    .A(_06367_),
    .ZN(_06368_)
  );
  AND2_X1 _12268_ (
    .A1(_00819_),
    .A2(_00821_),
    .ZN(_06369_)
  );
  AND2_X1 _12269_ (
    .A1(_06367_),
    .A2(_06369_),
    .ZN(_06370_)
  );
  INV_X1 _12270_ (
    .A(_06370_),
    .ZN(_06371_)
  );
  AND2_X1 _12271_ (
    .A1(_06366_),
    .A2(_06371_),
    .ZN(_06372_)
  );
  INV_X1 _12272_ (
    .A(_06372_),
    .ZN(_06373_)
  );
  AND2_X1 _12273_ (
    .A1(_00815_),
    .A2(_06373_),
    .ZN(_06374_)
  );
  INV_X1 _12274_ (
    .A(_06374_),
    .ZN(_06375_)
  );
  AND2_X1 _12275_ (
    .A1(io_decode_0_inst[22]),
    .A2(io_decode_0_inst[20]),
    .ZN(_06376_)
  );
  INV_X1 _12276_ (
    .A(_06376_),
    .ZN(_06377_)
  );
  AND2_X1 _12277_ (
    .A1(_00817_),
    .A2(_00819_),
    .ZN(_06378_)
  );
  AND2_X1 _12278_ (
    .A1(_06324_),
    .A2(_06378_),
    .ZN(_06379_)
  );
  AND2_X1 _12279_ (
    .A1(_06377_),
    .A2(_06379_),
    .ZN(_06380_)
  );
  INV_X1 _12280_ (
    .A(_06380_),
    .ZN(_06381_)
  );
  AND2_X1 _12281_ (
    .A1(_06375_),
    .A2(_06381_),
    .ZN(_06382_)
  );
  INV_X1 _12282_ (
    .A(_06382_),
    .ZN(_06383_)
  );
  AND2_X1 _12283_ (
    .A1(_00822_),
    .A2(_06383_),
    .ZN(_06384_)
  );
  INV_X1 _12284_ (
    .A(_06384_),
    .ZN(_06385_)
  );
  AND2_X1 _12285_ (
    .A1(io_decode_0_inst[25]),
    .A2(io_decode_0_inst[24]),
    .ZN(_06386_)
  );
  AND2_X1 _12286_ (
    .A1(_06334_),
    .A2(_06386_),
    .ZN(_06387_)
  );
  INV_X1 _12287_ (
    .A(_06387_),
    .ZN(_06388_)
  );
  AND2_X1 _12288_ (
    .A1(_06344_),
    .A2(_06353_),
    .ZN(_06389_)
  );
  AND2_X1 _12289_ (
    .A1(_06324_),
    .A2(_06332_),
    .ZN(_06390_)
  );
  AND2_X1 _12290_ (
    .A1(_06389_),
    .A2(_06390_),
    .ZN(_06391_)
  );
  INV_X1 _12291_ (
    .A(_06391_),
    .ZN(_06392_)
  );
  AND2_X1 _12292_ (
    .A1(_06332_),
    .A2(_06386_),
    .ZN(_06393_)
  );
  AND2_X1 _12293_ (
    .A1(_00817_),
    .A2(_06353_),
    .ZN(_06394_)
  );
  AND2_X1 _12294_ (
    .A1(_06393_),
    .A2(_06394_),
    .ZN(_06395_)
  );
  INV_X1 _12295_ (
    .A(_06395_),
    .ZN(_06396_)
  );
  AND2_X1 _12296_ (
    .A1(_06392_),
    .A2(_06396_),
    .ZN(_06397_)
  );
  AND2_X1 _12297_ (
    .A1(_06388_),
    .A2(_06397_),
    .ZN(_06398_)
  );
  AND2_X1 _12298_ (
    .A1(_00818_),
    .A2(io_decode_0_inst[23]),
    .ZN(_06399_)
  );
  INV_X1 _12299_ (
    .A(_06399_),
    .ZN(_06400_)
  );
  AND2_X1 _12300_ (
    .A1(io_decode_0_inst[22]),
    .A2(_06339_),
    .ZN(_06401_)
  );
  AND2_X1 _12301_ (
    .A1(_06400_),
    .A2(_06401_),
    .ZN(_06402_)
  );
  INV_X1 _12302_ (
    .A(_06402_),
    .ZN(_06403_)
  );
  AND2_X1 _12303_ (
    .A1(_06393_),
    .A2(_06403_),
    .ZN(_06404_)
  );
  INV_X1 _12304_ (
    .A(_06404_),
    .ZN(_06405_)
  );
  AND2_X1 _12305_ (
    .A1(_06326_),
    .A2(_06331_),
    .ZN(_06406_)
  );
  INV_X1 _12306_ (
    .A(_06406_),
    .ZN(_06407_)
  );
  AND2_X1 _12307_ (
    .A1(_00823_),
    .A2(_06337_),
    .ZN(_06408_)
  );
  AND2_X1 _12308_ (
    .A1(_06407_),
    .A2(_06408_),
    .ZN(_06409_)
  );
  AND2_X1 _12309_ (
    .A1(_06405_),
    .A2(_06409_),
    .ZN(_06410_)
  );
  AND2_X1 _12310_ (
    .A1(_06398_),
    .A2(_06410_),
    .ZN(_06411_)
  );
  AND2_X1 _12311_ (
    .A1(_06385_),
    .A2(_06411_),
    .ZN(_06412_)
  );
  INV_X1 _12312_ (
    .A(_06412_),
    .ZN(_06413_)
  );
  AND2_X1 _12313_ (
    .A1(_06352_),
    .A2(_06413_),
    .ZN(_06414_)
  );
  INV_X1 _12314_ (
    .A(_06414_),
    .ZN(_06415_)
  );
  AND2_X1 _12315_ (
    .A1(_00816_),
    .A2(_06415_),
    .ZN(_06416_)
  );
  INV_X1 _12316_ (
    .A(_06416_),
    .ZN(_06417_)
  );
  AND2_X1 _12317_ (
    .A1(_06353_),
    .A2(_06367_),
    .ZN(_06418_)
  );
  AND2_X1 _12318_ (
    .A1(_00820_),
    .A2(io_decode_0_inst[24]),
    .ZN(_06419_)
  );
  AND2_X1 _12319_ (
    .A1(_00815_),
    .A2(_06419_),
    .ZN(_06420_)
  );
  AND2_X1 _12320_ (
    .A1(_06332_),
    .A2(_06419_),
    .ZN(_06421_)
  );
  AND2_X1 _12321_ (
    .A1(_06418_),
    .A2(_06421_),
    .ZN(_06422_)
  );
  INV_X1 _12322_ (
    .A(_06422_),
    .ZN(_06423_)
  );
  AND2_X1 _12323_ (
    .A1(io_decode_0_inst[30]),
    .A2(_06423_),
    .ZN(_06424_)
  );
  INV_X1 _12324_ (
    .A(_06424_),
    .ZN(_06425_)
  );
  AND2_X1 _12325_ (
    .A1(_06327_),
    .A2(_06368_),
    .ZN(_06426_)
  );
  MUX2_X1 _12326_ (
    .A(_06327_),
    .B(_06353_),
    .S(_06367_),
    .Z(_06427_)
  );
  AND2_X1 _12327_ (
    .A1(io_decode_0_inst[27]),
    .A2(_06427_),
    .ZN(_06428_)
  );
  INV_X1 _12328_ (
    .A(_06428_),
    .ZN(_06429_)
  );
  AND2_X1 _12329_ (
    .A1(_06327_),
    .A2(_06367_),
    .ZN(_06430_)
  );
  INV_X1 _12330_ (
    .A(_06430_),
    .ZN(_06431_)
  );
  AND2_X1 _12331_ (
    .A1(io_decode_0_inst[22]),
    .A2(_06338_),
    .ZN(_06432_)
  );
  INV_X1 _12332_ (
    .A(_06432_),
    .ZN(_06433_)
  );
  AND2_X1 _12333_ (
    .A1(io_decode_0_inst[23]),
    .A2(_06433_),
    .ZN(_06434_)
  );
  INV_X1 _12334_ (
    .A(_06434_),
    .ZN(_06435_)
  );
  AND2_X1 _12335_ (
    .A1(_06431_),
    .A2(_06435_),
    .ZN(_06436_)
  );
  AND2_X1 _12336_ (
    .A1(_06429_),
    .A2(_06436_),
    .ZN(_06437_)
  );
  INV_X1 _12337_ (
    .A(_06437_),
    .ZN(_06438_)
  );
  AND2_X1 _12338_ (
    .A1(_06419_),
    .A2(_06438_),
    .ZN(_06439_)
  );
  INV_X1 _12339_ (
    .A(_06439_),
    .ZN(_06440_)
  );
  AND2_X1 _12340_ (
    .A1(_06353_),
    .A2(_06368_),
    .ZN(_06441_)
  );
  INV_X1 _12341_ (
    .A(_06441_),
    .ZN(_06442_)
  );
  AND2_X1 _12342_ (
    .A1(_06327_),
    .A2(_06339_),
    .ZN(_06443_)
  );
  INV_X1 _12343_ (
    .A(_06443_),
    .ZN(_06444_)
  );
  AND2_X1 _12344_ (
    .A1(_06324_),
    .A2(_06444_),
    .ZN(_06445_)
  );
  AND2_X1 _12345_ (
    .A1(_06442_),
    .A2(_06445_),
    .ZN(_06446_)
  );
  INV_X1 _12346_ (
    .A(_06446_),
    .ZN(_06447_)
  );
  AND2_X1 _12347_ (
    .A1(_00820_),
    .A2(_06389_),
    .ZN(_06448_)
  );
  INV_X1 _12348_ (
    .A(_06448_),
    .ZN(_06449_)
  );
  AND2_X1 _12349_ (
    .A1(_00818_),
    .A2(_06324_),
    .ZN(_06450_)
  );
  AND2_X1 _12350_ (
    .A1(_06327_),
    .A2(_06450_),
    .ZN(_06451_)
  );
  INV_X1 _12351_ (
    .A(_06451_),
    .ZN(_06452_)
  );
  AND2_X1 _12352_ (
    .A1(_06449_),
    .A2(_06452_),
    .ZN(_06453_)
  );
  AND2_X1 _12353_ (
    .A1(_06447_),
    .A2(_06453_),
    .ZN(_06454_)
  );
  AND2_X1 _12354_ (
    .A1(_06440_),
    .A2(_06454_),
    .ZN(_06455_)
  );
  INV_X1 _12355_ (
    .A(_06455_),
    .ZN(_06456_)
  );
  AND2_X1 _12356_ (
    .A1(_00815_),
    .A2(_06456_),
    .ZN(_06457_)
  );
  INV_X1 _12357_ (
    .A(_06457_),
    .ZN(_06458_)
  );
  AND2_X1 _12358_ (
    .A1(_00815_),
    .A2(_00820_),
    .ZN(_06459_)
  );
  AND2_X1 _12359_ (
    .A1(_06353_),
    .A2(_06459_),
    .ZN(_06460_)
  );
  AND2_X1 _12360_ (
    .A1(io_decode_0_inst[21]),
    .A2(_06460_),
    .ZN(_06461_)
  );
  INV_X1 _12361_ (
    .A(_06461_),
    .ZN(_06462_)
  );
  AND2_X1 _12362_ (
    .A1(_06338_),
    .A2(_06359_),
    .ZN(_06463_)
  );
  AND2_X1 _12363_ (
    .A1(_06420_),
    .A2(_06463_),
    .ZN(_06464_)
  );
  INV_X1 _12364_ (
    .A(_06464_),
    .ZN(_06465_)
  );
  AND2_X1 _12365_ (
    .A1(_06423_),
    .A2(_06465_),
    .ZN(_06466_)
  );
  AND2_X1 _12366_ (
    .A1(_06462_),
    .A2(_06466_),
    .ZN(_06467_)
  );
  AND2_X1 _12367_ (
    .A1(_06458_),
    .A2(_06467_),
    .ZN(_06468_)
  );
  INV_X1 _12368_ (
    .A(_06468_),
    .ZN(_06469_)
  );
  AND2_X1 _12369_ (
    .A1(_06425_),
    .A2(_06469_),
    .ZN(_06470_)
  );
  INV_X1 _12370_ (
    .A(_06470_),
    .ZN(_06471_)
  );
  AND2_X1 _12371_ (
    .A1(_06421_),
    .A2(_06426_),
    .ZN(_06472_)
  );
  INV_X1 _12372_ (
    .A(_06472_),
    .ZN(_06473_)
  );
  AND2_X1 _12373_ (
    .A1(io_decode_0_inst[31]),
    .A2(_06473_),
    .ZN(_06474_)
  );
  AND2_X1 _12374_ (
    .A1(_06471_),
    .A2(_06474_),
    .ZN(_06475_)
  );
  INV_X1 _12375_ (
    .A(_06475_),
    .ZN(_06476_)
  );
  AND2_X1 _12376_ (
    .A1(io_decode_0_inst[29]),
    .A2(io_decode_0_inst[28]),
    .ZN(_06477_)
  );
  AND2_X1 _12377_ (
    .A1(_00816_),
    .A2(io_decode_0_inst[30]),
    .ZN(_06478_)
  );
  AND2_X1 _12378_ (
    .A1(_io_decode_0_read_illegal_T_15),
    .A2(_06477_),
    .ZN(_06479_)
  );
  AND2_X1 _12379_ (
    .A1(_06478_),
    .A2(_06479_),
    .ZN(_06480_)
  );
  AND2_X1 _12380_ (
    .A1(_06387_),
    .A2(_06480_),
    .ZN(_06481_)
  );
  INV_X1 _12381_ (
    .A(_06481_),
    .ZN(_06482_)
  );
  AND2_X1 _12382_ (
    .A1(_06477_),
    .A2(_06482_),
    .ZN(_06483_)
  );
  AND2_X1 _12383_ (
    .A1(_06476_),
    .A2(_06483_),
    .ZN(_06484_)
  );
  AND2_X1 _12384_ (
    .A1(_06417_),
    .A2(_06484_),
    .ZN(_06485_)
  );
  INV_X1 _12385_ (
    .A(_06485_),
    .ZN(io_decode_0_read_illegal)
  );
  AND2_X1 _12386_ (
    .A1(io_decode_0_inst[27]),
    .A2(_io_decode_0_read_illegal_T_15),
    .ZN(_06486_)
  );
  AND2_X1 _12387_ (
    .A1(_06478_),
    .A2(_06486_),
    .ZN(io_decode_0_system_illegal)
  );
  AND2_X1 _12388_ (
    .A1(_03486_),
    .A2(_03544_),
    .ZN(_06487_)
  );
  INV_X1 _12389_ (
    .A(_06487_),
    .ZN(io_eret)
  );
  AND2_X1 _12390_ (
    .A1(_03476_),
    .A2(io_interrupt_cause[1]),
    .ZN(_06488_)
  );
  INV_X1 _12391_ (
    .A(_06488_),
    .ZN(_06489_)
  );
  AND2_X1 _12392_ (
    .A1(_00785_),
    .A2(_06489_),
    .ZN(_06490_)
  );
  INV_X1 _12393_ (
    .A(_06490_),
    .ZN(_06491_)
  );
  AND2_X1 _12394_ (
    .A1(_00870_),
    .A2(_00879_),
    .ZN(_06492_)
  );
  AND2_X1 _12395_ (
    .A1(_06491_),
    .A2(_06492_),
    .ZN(io_interrupt)
  );
  INV_X1 _12396_ (
    .A(large_[25]),
    .ZN(_00622_)
  );
  INV_X1 _12397_ (
    .A(large_[24]),
    .ZN(_00623_)
  );
  INV_X1 _12398_ (
    .A(large_[23]),
    .ZN(_00624_)
  );
  INV_X1 _12399_ (
    .A(large_[22]),
    .ZN(_00625_)
  );
  INV_X1 _12400_ (
    .A(large_[21]),
    .ZN(_00626_)
  );
  INV_X1 _12401_ (
    .A(large_[20]),
    .ZN(_00627_)
  );
  INV_X1 _12402_ (
    .A(large_[19]),
    .ZN(_00628_)
  );
  INV_X1 _12403_ (
    .A(large_[18]),
    .ZN(_00629_)
  );
  INV_X1 _12404_ (
    .A(large_[17]),
    .ZN(_00630_)
  );
  INV_X1 _12405_ (
    .A(large_[16]),
    .ZN(_00631_)
  );
  INV_X1 _12406_ (
    .A(large_[15]),
    .ZN(_00632_)
  );
  INV_X1 _12407_ (
    .A(large_[14]),
    .ZN(_00633_)
  );
  INV_X1 _12408_ (
    .A(large_[13]),
    .ZN(_00634_)
  );
  INV_X1 _12409_ (
    .A(large_[10]),
    .ZN(_00635_)
  );
  INV_X1 _12410_ (
    .A(large_[9]),
    .ZN(_00636_)
  );
  INV_X1 _12411_ (
    .A(large_[8]),
    .ZN(_00637_)
  );
  INV_X1 _12412_ (
    .A(large_[7]),
    .ZN(_00638_)
  );
  INV_X1 _12413_ (
    .A(large_[6]),
    .ZN(_00639_)
  );
  INV_X1 _12414_ (
    .A(large_[5]),
    .ZN(_00640_)
  );
  INV_X1 _12415_ (
    .A(large_[4]),
    .ZN(_00641_)
  );
  INV_X1 _12416_ (
    .A(large_[3]),
    .ZN(_00642_)
  );
  INV_X1 _12417_ (
    .A(large_[2]),
    .ZN(_00643_)
  );
  INV_X1 _12418_ (
    .A(large_[1]),
    .ZN(_00644_)
  );
  INV_X1 _12419_ (
    .A(large_1[25]),
    .ZN(_00645_)
  );
  INV_X1 _12420_ (
    .A(large_1[24]),
    .ZN(_00646_)
  );
  INV_X1 _12421_ (
    .A(large_1[23]),
    .ZN(_00647_)
  );
  INV_X1 _12422_ (
    .A(large_1[22]),
    .ZN(_00648_)
  );
  INV_X1 _12423_ (
    .A(large_1[21]),
    .ZN(_00649_)
  );
  INV_X1 _12424_ (
    .A(large_1[20]),
    .ZN(_00650_)
  );
  INV_X1 _12425_ (
    .A(large_1[19]),
    .ZN(_00651_)
  );
  INV_X1 _12426_ (
    .A(large_1[18]),
    .ZN(_00652_)
  );
  INV_X1 _12427_ (
    .A(large_1[17]),
    .ZN(_00653_)
  );
  INV_X1 _12428_ (
    .A(large_1[16]),
    .ZN(_00654_)
  );
  INV_X1 _12429_ (
    .A(large_1[15]),
    .ZN(_00655_)
  );
  INV_X1 _12430_ (
    .A(large_1[14]),
    .ZN(_00656_)
  );
  INV_X1 _12431_ (
    .A(large_1[13]),
    .ZN(_00657_)
  );
  INV_X1 _12432_ (
    .A(large_1[12]),
    .ZN(_00658_)
  );
  INV_X1 _12433_ (
    .A(large_1[11]),
    .ZN(_00659_)
  );
  INV_X1 _12434_ (
    .A(large_1[10]),
    .ZN(_00660_)
  );
  INV_X1 _12435_ (
    .A(large_1[9]),
    .ZN(_00661_)
  );
  INV_X1 _12436_ (
    .A(large_1[8]),
    .ZN(_00662_)
  );
  INV_X1 _12437_ (
    .A(large_1[7]),
    .ZN(_00663_)
  );
  INV_X1 _12438_ (
    .A(large_1[6]),
    .ZN(_00664_)
  );
  INV_X1 _12439_ (
    .A(large_1[5]),
    .ZN(_00665_)
  );
  INV_X1 _12440_ (
    .A(large_1[4]),
    .ZN(_00666_)
  );
  INV_X1 _12441_ (
    .A(large_1[3]),
    .ZN(_00667_)
  );
  INV_X1 _12442_ (
    .A(large_1[2]),
    .ZN(_00668_)
  );
  INV_X1 _12443_ (
    .A(large_1[1]),
    .ZN(_00669_)
  );
  INV_X1 _12444_ (
    .A(reg_pmp_7_cfg_l),
    .ZN(_00670_)
  );
  INV_X1 _12445_ (
    .A(reg_pmp_7_cfg_a[1]),
    .ZN(_00671_)
  );
  INV_X1 _12446_ (
    .A(reg_pmp_7_cfg_a[0]),
    .ZN(_00672_)
  );
  INV_X1 _12447_ (
    .A(reg_mtvec[31]),
    .ZN(_00673_)
  );
  INV_X1 _12448_ (
    .A(reg_mtvec[30]),
    .ZN(_00674_)
  );
  INV_X1 _12449_ (
    .A(reg_mtvec[29]),
    .ZN(_00675_)
  );
  INV_X1 _12450_ (
    .A(reg_mtvec[28]),
    .ZN(_00676_)
  );
  INV_X1 _12451_ (
    .A(reg_mtvec[27]),
    .ZN(_00677_)
  );
  INV_X1 _12452_ (
    .A(reg_mtvec[26]),
    .ZN(_00678_)
  );
  INV_X1 _12453_ (
    .A(reg_mtvec[25]),
    .ZN(_00679_)
  );
  INV_X1 _12454_ (
    .A(reg_mtvec[24]),
    .ZN(_00680_)
  );
  INV_X1 _12455_ (
    .A(reg_mtvec[23]),
    .ZN(_00681_)
  );
  INV_X1 _12456_ (
    .A(reg_mtvec[22]),
    .ZN(_00682_)
  );
  INV_X1 _12457_ (
    .A(reg_mtvec[21]),
    .ZN(_00683_)
  );
  INV_X1 _12458_ (
    .A(reg_mtvec[20]),
    .ZN(_00684_)
  );
  INV_X1 _12459_ (
    .A(reg_mtvec[19]),
    .ZN(_00685_)
  );
  INV_X1 _12460_ (
    .A(reg_mtvec[18]),
    .ZN(_00686_)
  );
  INV_X1 _12461_ (
    .A(reg_mtvec[17]),
    .ZN(_00687_)
  );
  INV_X1 _12462_ (
    .A(reg_mtvec[16]),
    .ZN(_00688_)
  );
  INV_X1 _12463_ (
    .A(reg_mtvec[15]),
    .ZN(_00689_)
  );
  INV_X1 _12464_ (
    .A(reg_mtvec[14]),
    .ZN(_00690_)
  );
  INV_X1 _12465_ (
    .A(reg_mtvec[13]),
    .ZN(_00691_)
  );
  INV_X1 _12466_ (
    .A(reg_mtvec[12]),
    .ZN(_00692_)
  );
  INV_X1 _12467_ (
    .A(reg_mtvec[11]),
    .ZN(_00693_)
  );
  INV_X1 _12468_ (
    .A(reg_mtvec[10]),
    .ZN(_00694_)
  );
  INV_X1 _12469_ (
    .A(reg_mtvec[9]),
    .ZN(_00695_)
  );
  INV_X1 _12470_ (
    .A(reg_mtvec[8]),
    .ZN(_00696_)
  );
  INV_X1 _12471_ (
    .A(reg_mtvec[7]),
    .ZN(_00697_)
  );
  INV_X1 _12472_ (
    .A(reg_mtvec[6]),
    .ZN(_00698_)
  );
  INV_X1 _12473_ (
    .A(reg_mtvec[5]),
    .ZN(_00699_)
  );
  INV_X1 _12474_ (
    .A(reg_mtvec[4]),
    .ZN(_00700_)
  );
  INV_X1 _12475_ (
    .A(reg_mtvec[3]),
    .ZN(_00701_)
  );
  INV_X1 _12476_ (
    .A(reg_mtvec[2]),
    .ZN(_00702_)
  );
  INV_X1 _12477_ (
    .A(reg_mtvec[0]),
    .ZN(_00703_)
  );
  INV_X1 _12478_ (
    .A(small_[5]),
    .ZN(_00704_)
  );
  INV_X1 _12479_ (
    .A(small_[4]),
    .ZN(_00705_)
  );
  INV_X1 _12480_ (
    .A(small_[3]),
    .ZN(_00706_)
  );
  INV_X1 _12481_ (
    .A(small_[2]),
    .ZN(_00707_)
  );
  INV_X1 _12482_ (
    .A(small_[1]),
    .ZN(_00708_)
  );
  INV_X1 _12483_ (
    .A(small_[0]),
    .ZN(_00709_)
  );
  INV_X1 _12484_ (
    .A(large_[57]),
    .ZN(_00710_)
  );
  INV_X1 _12485_ (
    .A(large_[56]),
    .ZN(_00711_)
  );
  INV_X1 _12486_ (
    .A(large_[55]),
    .ZN(_00712_)
  );
  INV_X1 _12487_ (
    .A(large_[54]),
    .ZN(_00713_)
  );
  INV_X1 _12488_ (
    .A(large_[53]),
    .ZN(_00714_)
  );
  INV_X1 _12489_ (
    .A(large_[52]),
    .ZN(_00715_)
  );
  INV_X1 _12490_ (
    .A(large_[51]),
    .ZN(_00716_)
  );
  INV_X1 _12491_ (
    .A(large_[50]),
    .ZN(_00717_)
  );
  INV_X1 _12492_ (
    .A(large_[49]),
    .ZN(_00718_)
  );
  INV_X1 _12493_ (
    .A(large_[48]),
    .ZN(_00719_)
  );
  INV_X1 _12494_ (
    .A(large_[47]),
    .ZN(_00720_)
  );
  INV_X1 _12495_ (
    .A(large_[46]),
    .ZN(_00721_)
  );
  INV_X1 _12496_ (
    .A(large_[45]),
    .ZN(_00722_)
  );
  INV_X1 _12497_ (
    .A(large_[44]),
    .ZN(_00723_)
  );
  INV_X1 _12498_ (
    .A(large_[43]),
    .ZN(_00724_)
  );
  INV_X1 _12499_ (
    .A(large_[42]),
    .ZN(_00725_)
  );
  INV_X1 _12500_ (
    .A(large_[41]),
    .ZN(_00726_)
  );
  INV_X1 _12501_ (
    .A(large_[40]),
    .ZN(_00727_)
  );
  INV_X1 _12502_ (
    .A(large_[39]),
    .ZN(_00728_)
  );
  INV_X1 _12503_ (
    .A(large_[38]),
    .ZN(_00729_)
  );
  INV_X1 _12504_ (
    .A(large_[37]),
    .ZN(_00730_)
  );
  INV_X1 _12505_ (
    .A(large_[36]),
    .ZN(_00731_)
  );
  INV_X1 _12506_ (
    .A(large_[35]),
    .ZN(_00732_)
  );
  INV_X1 _12507_ (
    .A(large_[34]),
    .ZN(_00733_)
  );
  INV_X1 _12508_ (
    .A(large_[33]),
    .ZN(_00734_)
  );
  INV_X1 _12509_ (
    .A(large_[32]),
    .ZN(_00735_)
  );
  INV_X1 _12510_ (
    .A(large_[31]),
    .ZN(_00736_)
  );
  INV_X1 _12511_ (
    .A(large_[30]),
    .ZN(_00737_)
  );
  INV_X1 _12512_ (
    .A(large_[29]),
    .ZN(_00738_)
  );
  INV_X1 _12513_ (
    .A(large_[28]),
    .ZN(_00739_)
  );
  INV_X1 _12514_ (
    .A(large_[27]),
    .ZN(_00740_)
  );
  INV_X1 _12515_ (
    .A(large_[26]),
    .ZN(_00741_)
  );
  INV_X1 _12516_ (
    .A(reg_misa[2]),
    .ZN(_00742_)
  );
  INV_X1 _12517_ (
    .A(reg_misa[0]),
    .ZN(_00743_)
  );
  INV_X1 _12518_ (
    .A(small_1[5]),
    .ZN(_00744_)
  );
  INV_X1 _12519_ (
    .A(small_1[4]),
    .ZN(_00745_)
  );
  INV_X1 _12520_ (
    .A(small_1[3]),
    .ZN(_00746_)
  );
  INV_X1 _12521_ (
    .A(small_1[2]),
    .ZN(_00747_)
  );
  INV_X1 _12522_ (
    .A(small_1[1]),
    .ZN(_00748_)
  );
  INV_X1 _12523_ (
    .A(small_1[0]),
    .ZN(_00749_)
  );
  INV_X1 _12524_ (
    .A(large_1[57]),
    .ZN(_00750_)
  );
  INV_X1 _12525_ (
    .A(large_1[56]),
    .ZN(_00751_)
  );
  INV_X1 _12526_ (
    .A(large_1[55]),
    .ZN(_00752_)
  );
  INV_X1 _12527_ (
    .A(large_1[54]),
    .ZN(_00753_)
  );
  INV_X1 _12528_ (
    .A(large_1[53]),
    .ZN(_00754_)
  );
  INV_X1 _12529_ (
    .A(large_1[52]),
    .ZN(_00755_)
  );
  INV_X1 _12530_ (
    .A(large_1[51]),
    .ZN(_00756_)
  );
  INV_X1 _12531_ (
    .A(large_1[50]),
    .ZN(_00757_)
  );
  INV_X1 _12532_ (
    .A(large_1[49]),
    .ZN(_00758_)
  );
  INV_X1 _12533_ (
    .A(large_1[48]),
    .ZN(_00759_)
  );
  INV_X1 _12534_ (
    .A(large_1[47]),
    .ZN(_00760_)
  );
  INV_X1 _12535_ (
    .A(large_1[46]),
    .ZN(_00761_)
  );
  INV_X1 _12536_ (
    .A(large_1[45]),
    .ZN(_00762_)
  );
  INV_X1 _12537_ (
    .A(large_1[44]),
    .ZN(_00763_)
  );
  INV_X1 _12538_ (
    .A(large_1[43]),
    .ZN(_00764_)
  );
  INV_X1 _12539_ (
    .A(large_1[42]),
    .ZN(_00765_)
  );
  INV_X1 _12540_ (
    .A(large_1[41]),
    .ZN(_00766_)
  );
  INV_X1 _12541_ (
    .A(large_1[40]),
    .ZN(_00767_)
  );
  INV_X1 _12542_ (
    .A(large_1[39]),
    .ZN(_00768_)
  );
  INV_X1 _12543_ (
    .A(large_1[38]),
    .ZN(_00769_)
  );
  INV_X1 _12544_ (
    .A(large_1[37]),
    .ZN(_00770_)
  );
  INV_X1 _12545_ (
    .A(large_1[36]),
    .ZN(_00771_)
  );
  INV_X1 _12546_ (
    .A(large_1[35]),
    .ZN(_00772_)
  );
  INV_X1 _12547_ (
    .A(large_1[34]),
    .ZN(_00773_)
  );
  INV_X1 _12548_ (
    .A(large_1[33]),
    .ZN(_00774_)
  );
  INV_X1 _12549_ (
    .A(large_1[32]),
    .ZN(_00775_)
  );
  INV_X1 _12550_ (
    .A(large_1[31]),
    .ZN(_00776_)
  );
  INV_X1 _12551_ (
    .A(large_1[30]),
    .ZN(_00777_)
  );
  INV_X1 _12552_ (
    .A(large_1[29]),
    .ZN(_00778_)
  );
  INV_X1 _12553_ (
    .A(large_1[28]),
    .ZN(_00779_)
  );
  INV_X1 _12554_ (
    .A(large_1[27]),
    .ZN(_00780_)
  );
  INV_X1 _12555_ (
    .A(large_1[26]),
    .ZN(_00781_)
  );
  INV_X1 _12556_ (
    .A(reg_mcountinhibit[2]),
    .ZN(_00782_)
  );
  INV_X1 _12557_ (
    .A(reg_mcountinhibit[0]),
    .ZN(_00783_)
  );
  INV_X1 _12558_ (
    .A(reg_dcsr_ebreakm),
    .ZN(_00784_)
  );
  INV_X1 _12559_ (
    .A(reg_singleStepped),
    .ZN(_00785_)
  );
  INV_X1 _12560_ (
    .A(reg_dcsr_step),
    .ZN(_00786_)
  );
  INV_X1 _12561_ (
    .A(reg_bp_0_control_x),
    .ZN(_00787_)
  );
  INV_X1 _12562_ (
    .A(reg_bp_0_control_w),
    .ZN(_00788_)
  );
  INV_X1 _12563_ (
    .A(reg_bp_0_control_r),
    .ZN(_00789_)
  );
  INV_X1 _12564_ (
    .A(reg_pmp_0_cfg_l),
    .ZN(_00790_)
  );
  INV_X1 _12565_ (
    .A(reg_pmp_0_cfg_a[1]),
    .ZN(_00791_)
  );
  INV_X1 _12566_ (
    .A(reg_pmp_0_cfg_a[0]),
    .ZN(_00792_)
  );
  INV_X1 _12567_ (
    .A(reg_pmp_1_cfg_l),
    .ZN(_00793_)
  );
  INV_X1 _12568_ (
    .A(reg_pmp_1_cfg_a[1]),
    .ZN(_00794_)
  );
  INV_X1 _12569_ (
    .A(reg_pmp_1_cfg_a[0]),
    .ZN(_00795_)
  );
  INV_X1 _12570_ (
    .A(reg_pmp_2_cfg_l),
    .ZN(_00796_)
  );
  INV_X1 _12571_ (
    .A(reg_pmp_2_cfg_a[1]),
    .ZN(_00797_)
  );
  INV_X1 _12572_ (
    .A(reg_pmp_2_cfg_a[0]),
    .ZN(_00798_)
  );
  INV_X1 _12573_ (
    .A(reg_pmp_3_cfg_l),
    .ZN(_00799_)
  );
  INV_X1 _12574_ (
    .A(reg_pmp_3_cfg_a[1]),
    .ZN(_00800_)
  );
  INV_X1 _12575_ (
    .A(reg_pmp_3_cfg_a[0]),
    .ZN(_00801_)
  );
  INV_X1 _12576_ (
    .A(reg_pmp_4_cfg_l),
    .ZN(_00802_)
  );
  INV_X1 _12577_ (
    .A(reg_pmp_4_cfg_a[1]),
    .ZN(_00803_)
  );
  INV_X1 _12578_ (
    .A(reg_pmp_4_cfg_a[0]),
    .ZN(_00804_)
  );
  INV_X1 _12579_ (
    .A(reg_pmp_5_cfg_l),
    .ZN(_00805_)
  );
  INV_X1 _12580_ (
    .A(reg_pmp_5_cfg_a[1]),
    .ZN(_00806_)
  );
  INV_X1 _12581_ (
    .A(reg_pmp_5_cfg_a[0]),
    .ZN(_00807_)
  );
  INV_X1 _12582_ (
    .A(reg_pmp_6_cfg_l),
    .ZN(_00808_)
  );
  INV_X1 _12583_ (
    .A(reg_pmp_6_cfg_a[1]),
    .ZN(_00809_)
  );
  INV_X1 _12584_ (
    .A(reg_pmp_6_cfg_a[0]),
    .ZN(_00810_)
  );
  INV_X1 _12585_ (
    .A(reset),
    .ZN(_00811_)
  );
  INV_X1 _12586_ (
    .A(io_rw_cmd[1]),
    .ZN(_00812_)
  );
  INV_X1 _12587_ (
    .A(io_rw_cmd[0]),
    .ZN(_00813_)
  );
  INV_X1 _12588_ (
    .A(io_decode_0_inst[22]),
    .ZN(_00814_)
  );
  INV_X1 _12589_ (
    .A(io_decode_0_inst[26]),
    .ZN(_00815_)
  );
  INV_X1 _12590_ (
    .A(io_decode_0_inst[31]),
    .ZN(_00816_)
  );
  INV_X1 _12591_ (
    .A(io_decode_0_inst[21]),
    .ZN(_00817_)
  );
  INV_X1 _12592_ (
    .A(io_decode_0_inst[20]),
    .ZN(_00818_)
  );
  INV_X1 _12593_ (
    .A(io_decode_0_inst[23]),
    .ZN(_00819_)
  );
  INV_X1 _12594_ (
    .A(io_decode_0_inst[25]),
    .ZN(_00820_)
  );
  INV_X1 _12595_ (
    .A(io_decode_0_inst[24]),
    .ZN(_00821_)
  );
  INV_X1 _12596_ (
    .A(io_decode_0_inst[27]),
    .ZN(_00822_)
  );
  INV_X1 _12597_ (
    .A(io_decode_0_inst[30]),
    .ZN(_00823_)
  );
  INV_X1 _12598_ (
    .A(io_rw_addr[6]),
    .ZN(_00824_)
  );
  INV_X1 _12599_ (
    .A(io_rw_addr[5]),
    .ZN(_00825_)
  );
  INV_X1 _12600_ (
    .A(io_rw_addr[4]),
    .ZN(_00826_)
  );
  INV_X1 _12601_ (
    .A(io_rw_addr[1]),
    .ZN(_00827_)
  );
  INV_X1 _12602_ (
    .A(io_rw_addr[10]),
    .ZN(_00828_)
  );
  INV_X1 _12603_ (
    .A(io_rw_addr[7]),
    .ZN(_00829_)
  );
  INV_X1 _12604_ (
    .A(io_rw_addr[11]),
    .ZN(_00830_)
  );
  INV_X1 _12605_ (
    .A(io_rw_addr[0]),
    .ZN(_00831_)
  );
  INV_X1 _12606_ (
    .A(io_rw_addr[8]),
    .ZN(_00832_)
  );
  INV_X1 _12607_ (
    .A(io_rw_addr[9]),
    .ZN(_00833_)
  );
  INV_X1 _12608_ (
    .A(io_rw_addr[2]),
    .ZN(_00834_)
  );
  INV_X1 _12609_ (
    .A(io_interrupts_debug),
    .ZN(_00835_)
  );
  INV_X1 _12610_ (
    .A(io_rw_wdata[0]),
    .ZN(_00836_)
  );
  INV_X1 _12611_ (
    .A(io_rw_wdata[1]),
    .ZN(_00837_)
  );
  INV_X1 _12612_ (
    .A(io_rw_wdata[2]),
    .ZN(_00838_)
  );
  INV_X1 _12613_ (
    .A(io_rw_wdata[3]),
    .ZN(_00839_)
  );
  INV_X1 _12614_ (
    .A(io_rw_wdata[4]),
    .ZN(_00840_)
  );
  INV_X1 _12615_ (
    .A(io_rw_wdata[5]),
    .ZN(_00841_)
  );
  INV_X1 _12616_ (
    .A(io_rw_wdata[6]),
    .ZN(_00842_)
  );
  INV_X1 _12617_ (
    .A(io_rw_wdata[7]),
    .ZN(_00843_)
  );
  INV_X1 _12618_ (
    .A(io_rw_wdata[8]),
    .ZN(_00844_)
  );
  INV_X1 _12619_ (
    .A(io_rw_wdata[9]),
    .ZN(_00845_)
  );
  INV_X1 _12620_ (
    .A(io_rw_wdata[10]),
    .ZN(_00846_)
  );
  INV_X1 _12621_ (
    .A(io_rw_wdata[11]),
    .ZN(_00847_)
  );
  INV_X1 _12622_ (
    .A(io_rw_wdata[13]),
    .ZN(_00848_)
  );
  INV_X1 _12623_ (
    .A(io_rw_wdata[14]),
    .ZN(_00849_)
  );
  INV_X1 _12624_ (
    .A(io_rw_wdata[15]),
    .ZN(_00850_)
  );
  INV_X1 _12625_ (
    .A(io_rw_wdata[16]),
    .ZN(_00851_)
  );
  INV_X1 _12626_ (
    .A(io_rw_wdata[17]),
    .ZN(_00852_)
  );
  INV_X1 _12627_ (
    .A(io_rw_wdata[18]),
    .ZN(_00853_)
  );
  INV_X1 _12628_ (
    .A(io_rw_wdata[19]),
    .ZN(_00854_)
  );
  INV_X1 _12629_ (
    .A(io_rw_wdata[20]),
    .ZN(_00855_)
  );
  INV_X1 _12630_ (
    .A(io_rw_wdata[21]),
    .ZN(_00856_)
  );
  INV_X1 _12631_ (
    .A(io_rw_wdata[22]),
    .ZN(_00857_)
  );
  INV_X1 _12632_ (
    .A(io_rw_wdata[23]),
    .ZN(_00858_)
  );
  INV_X1 _12633_ (
    .A(io_rw_wdata[24]),
    .ZN(_00859_)
  );
  INV_X1 _12634_ (
    .A(io_rw_wdata[25]),
    .ZN(_00860_)
  );
  INV_X1 _12635_ (
    .A(io_rw_wdata[26]),
    .ZN(_00861_)
  );
  INV_X1 _12636_ (
    .A(io_rw_wdata[27]),
    .ZN(_00862_)
  );
  INV_X1 _12637_ (
    .A(io_rw_wdata[28]),
    .ZN(_00863_)
  );
  INV_X1 _12638_ (
    .A(io_rw_wdata[29]),
    .ZN(_00864_)
  );
  INV_X1 _12639_ (
    .A(io_rw_wdata[30]),
    .ZN(_00865_)
  );
  INV_X1 _12640_ (
    .A(io_rw_wdata[31]),
    .ZN(_00866_)
  );
  INV_X1 _12641_ (
    .A(io_cause[0]),
    .ZN(_00867_)
  );
  INV_X1 _12642_ (
    .A(io_cause[1]),
    .ZN(_00868_)
  );
  INV_X1 _12643_ (
    .A(io_cause[4]),
    .ZN(_00869_)
  );
  INV_X1 _12644_ (
    .A(reg_debug),
    .ZN(_00870_)
  );
  INV_X1 _12645_ (
    .A(reg_mcause[1]),
    .ZN(_00871_)
  );
  INV_X1 _12646_ (
    .A(reg_mcause[3]),
    .ZN(_00872_)
  );
  INV_X1 _12647_ (
    .A(io_rw_addr[3]),
    .ZN(_00873_)
  );
  INV_X1 _12648_ (
    .A(_T_18[1]),
    .ZN(_00874_)
  );
  INV_X1 _12649_ (
    .A(_GEN_586[1]),
    .ZN(_00875_)
  );
  INV_X1 _12650_ (
    .A(_T_24[1]),
    .ZN(_00876_)
  );
  INV_X1 _12651_ (
    .A(reg_wfi),
    .ZN(_00877_)
  );
  INV_X1 _12652_ (
    .A(io_retire),
    .ZN(_00878_)
  );
  INV_X1 _12653_ (
    .A(io_status_cease_r),
    .ZN(_00879_)
  );
  INV_X1 _12654_ (
    .A(io_exception),
    .ZN(_00880_)
  );
  INV_X1 _12655_ (
    .A(_00005_),
    .ZN(_00881_)
  );
  AND2_X1 _12656_ (
    .A1(_00834_),
    .A2(_00873_),
    .ZN(_00882_)
  );
  AND2_X1 _12657_ (
    .A1(_00827_),
    .A2(_00882_),
    .ZN(_00883_)
  );
  AND2_X1 _12658_ (
    .A1(io_rw_addr[0]),
    .A2(_00883_),
    .ZN(_00884_)
  );
  AND2_X1 _12659_ (
    .A1(_00828_),
    .A2(_00830_),
    .ZN(_00885_)
  );
  AND2_X1 _12660_ (
    .A1(io_rw_addr[8]),
    .A2(io_rw_addr[9]),
    .ZN(_00886_)
  );
  AND2_X1 _12661_ (
    .A1(io_rw_addr[8]),
    .A2(_00885_),
    .ZN(_00887_)
  );
  AND2_X1 _12662_ (
    .A1(_00885_),
    .A2(_00886_),
    .ZN(_00888_)
  );
  AND2_X1 _12663_ (
    .A1(_00824_),
    .A2(io_rw_addr[7]),
    .ZN(_00889_)
  );
  AND2_X1 _12664_ (
    .A1(io_rw_addr[5]),
    .A2(_00826_),
    .ZN(_00890_)
  );
  AND2_X1 _12665_ (
    .A1(_00889_),
    .A2(_00890_),
    .ZN(_00891_)
  );
  AND2_X1 _12666_ (
    .A1(_00888_),
    .A2(_00890_),
    .ZN(_00892_)
  );
  AND2_X1 _12667_ (
    .A1(_00888_),
    .A2(_00891_),
    .ZN(_00893_)
  );
  AND2_X1 _12668_ (
    .A1(_00884_),
    .A2(_00893_),
    .ZN(_00894_)
  );
  AND2_X1 _12669_ (
    .A1(_00812_),
    .A2(_00813_),
    .ZN(_00895_)
  );
  INV_X1 _12670_ (
    .A(_00895_),
    .ZN(_00896_)
  );
  AND2_X1 _12671_ (
    .A1(io_rw_cmd[2]),
    .A2(_00896_),
    .ZN(_00897_)
  );
  INV_X1 _12672_ (
    .A(_00897_),
    .ZN(_00898_)
  );
  AND2_X1 _12673_ (
    .A1(_00017_),
    .A2(_00894_),
    .ZN(_00899_)
  );
  AND2_X1 _12674_ (
    .A1(_00897_),
    .A2(_00899_),
    .ZN(_00900_)
  );
  INV_X1 _12675_ (
    .A(_00900_),
    .ZN(_00901_)
  );
  AND2_X1 _12676_ (
    .A1(io_rw_cmd[1]),
    .A2(io_rw_cmd[0]),
    .ZN(_00902_)
  );
  INV_X1 _12677_ (
    .A(_00902_),
    .ZN(_00903_)
  );
  AND2_X1 _12678_ (
    .A1(io_rw_wdata[16]),
    .A2(_00903_),
    .ZN(_00904_)
  );
  INV_X1 _12679_ (
    .A(_00904_),
    .ZN(_00905_)
  );
  AND2_X1 _12680_ (
    .A1(io_rw_addr[5]),
    .A2(io_rw_addr[4]),
    .ZN(_00906_)
  );
  AND2_X1 _12681_ (
    .A1(_00889_),
    .A2(_00906_),
    .ZN(_00907_)
  );
  AND2_X1 _12682_ (
    .A1(io_rw_addr[10]),
    .A2(_00830_),
    .ZN(_00908_)
  );
  INV_X1 _12683_ (
    .A(_00908_),
    .ZN(_00909_)
  );
  AND2_X1 _12684_ (
    .A1(_00886_),
    .A2(_00908_),
    .ZN(_00910_)
  );
  AND2_X1 _12685_ (
    .A1(_00907_),
    .A2(_00910_),
    .ZN(_00911_)
  );
  AND2_X1 _12686_ (
    .A1(_00884_),
    .A2(_00911_),
    .ZN(_00912_)
  );
  AND2_X1 _12687_ (
    .A1(reg_dpc[16]),
    .A2(_00912_),
    .ZN(_00913_)
  );
  INV_X1 _12688_ (
    .A(_00913_),
    .ZN(_00914_)
  );
  AND2_X1 _12689_ (
    .A1(_00831_),
    .A2(_00883_),
    .ZN(_00915_)
  );
  AND2_X1 _12690_ (
    .A1(_00893_),
    .A2(_00915_),
    .ZN(_00916_)
  );
  AND2_X1 _12691_ (
    .A1(reg_pmp_2_cfg_r),
    .A2(_00916_),
    .ZN(_00917_)
  );
  INV_X1 _12692_ (
    .A(_00917_),
    .ZN(_00918_)
  );
  AND2_X1 _12693_ (
    .A1(_00914_),
    .A2(_00918_),
    .ZN(_00919_)
  );
  AND2_X1 _12694_ (
    .A1(_00825_),
    .A2(_00826_),
    .ZN(_00920_)
  );
  AND2_X1 _12695_ (
    .A1(io_rw_addr[6]),
    .A2(_00829_),
    .ZN(_00921_)
  );
  AND2_X1 _12696_ (
    .A1(_00920_),
    .A2(_00921_),
    .ZN(_00922_)
  );
  AND2_X1 _12697_ (
    .A1(_00888_),
    .A2(_00922_),
    .ZN(_00923_)
  );
  AND2_X1 _12698_ (
    .A1(io_rw_addr[1]),
    .A2(_00882_),
    .ZN(_00924_)
  );
  AND2_X1 _12699_ (
    .A1(io_rw_addr[0]),
    .A2(_00924_),
    .ZN(_00925_)
  );
  AND2_X1 _12700_ (
    .A1(_00923_),
    .A2(_00925_),
    .ZN(_00926_)
  );
  AND2_X1 _12701_ (
    .A1(reg_mtval[16]),
    .A2(_00926_),
    .ZN(_00927_)
  );
  INV_X1 _12702_ (
    .A(_00927_),
    .ZN(_00928_)
  );
  AND2_X1 _12703_ (
    .A1(_00915_),
    .A2(_00923_),
    .ZN(_00929_)
  );
  AND2_X1 _12704_ (
    .A1(reg_mscratch[16]),
    .A2(_00929_),
    .ZN(_00930_)
  );
  INV_X1 _12705_ (
    .A(_00930_),
    .ZN(_00931_)
  );
  AND2_X1 _12706_ (
    .A1(_00928_),
    .A2(_00931_),
    .ZN(_00932_)
  );
  AND2_X1 _12707_ (
    .A1(_00919_),
    .A2(_00932_),
    .ZN(_00933_)
  );
  AND2_X1 _12708_ (
    .A1(_00824_),
    .A2(_00829_),
    .ZN(_00934_)
  );
  AND2_X1 _12709_ (
    .A1(_00920_),
    .A2(_00934_),
    .ZN(_00935_)
  );
  AND2_X1 _12710_ (
    .A1(_00888_),
    .A2(_00935_),
    .ZN(_00936_)
  );
  AND2_X1 _12711_ (
    .A1(io_rw_addr[2]),
    .A2(_00873_),
    .ZN(_00937_)
  );
  AND2_X1 _12712_ (
    .A1(io_rw_addr[0]),
    .A2(_00937_),
    .ZN(_00938_)
  );
  AND2_X1 _12713_ (
    .A1(_00827_),
    .A2(_00938_),
    .ZN(_00939_)
  );
  AND2_X1 _12714_ (
    .A1(_00936_),
    .A2(_00939_),
    .ZN(_00940_)
  );
  AND2_X1 _12715_ (
    .A1(reg_mtvec[16]),
    .A2(_00940_),
    .ZN(_00941_)
  );
  INV_X1 _12716_ (
    .A(_00941_),
    .ZN(_00942_)
  );
  AND2_X1 _12717_ (
    .A1(_00884_),
    .A2(_00923_),
    .ZN(_00943_)
  );
  AND2_X1 _12718_ (
    .A1(reg_mepc[16]),
    .A2(_00943_),
    .ZN(_00944_)
  );
  INV_X1 _12719_ (
    .A(_00944_),
    .ZN(_00945_)
  );
  AND2_X1 _12720_ (
    .A1(_00942_),
    .A2(_00945_),
    .ZN(_00946_)
  );
  AND2_X1 _12721_ (
    .A1(_00888_),
    .A2(_00907_),
    .ZN(_00947_)
  );
  AND2_X1 _12722_ (
    .A1(_00939_),
    .A2(_00947_),
    .ZN(_00948_)
  );
  AND2_X1 _12723_ (
    .A1(reg_pmp_5_addr[16]),
    .A2(_00948_),
    .ZN(_00949_)
  );
  INV_X1 _12724_ (
    .A(_00949_),
    .ZN(_00950_)
  );
  AND2_X1 _12725_ (
    .A1(_00831_),
    .A2(_00924_),
    .ZN(_00951_)
  );
  INV_X1 _12726_ (
    .A(_00951_),
    .ZN(_00952_)
  );
  AND2_X1 _12727_ (
    .A1(_00947_),
    .A2(_00951_),
    .ZN(_00953_)
  );
  AND2_X1 _12728_ (
    .A1(reg_pmp_2_addr[16]),
    .A2(_00953_),
    .ZN(_00954_)
  );
  INV_X1 _12729_ (
    .A(_00954_),
    .ZN(_00955_)
  );
  AND2_X1 _12730_ (
    .A1(_00950_),
    .A2(_00955_),
    .ZN(_00956_)
  );
  AND2_X1 _12731_ (
    .A1(_00946_),
    .A2(_00956_),
    .ZN(_00957_)
  );
  AND2_X1 _12732_ (
    .A1(_00911_),
    .A2(_00924_),
    .ZN(_00958_)
  );
  AND2_X1 _12733_ (
    .A1(reg_dscratch0[16]),
    .A2(_00958_),
    .ZN(_00959_)
  );
  INV_X1 _12734_ (
    .A(_00959_),
    .ZN(_00960_)
  );
  AND2_X1 _12735_ (
    .A1(_00891_),
    .A2(_00910_),
    .ZN(_00961_)
  );
  AND2_X1 _12736_ (
    .A1(_00951_),
    .A2(_00961_),
    .ZN(_00962_)
  );
  AND2_X1 _12737_ (
    .A1(reg_bp_0_address[16]),
    .A2(_00962_),
    .ZN(_00963_)
  );
  INV_X1 _12738_ (
    .A(_00963_),
    .ZN(_00964_)
  );
  AND2_X1 _12739_ (
    .A1(_00960_),
    .A2(_00964_),
    .ZN(_00965_)
  );
  AND2_X1 _12740_ (
    .A1(_00831_),
    .A2(_00937_),
    .ZN(_00966_)
  );
  AND2_X1 _12741_ (
    .A1(_00827_),
    .A2(_00966_),
    .ZN(_00967_)
  );
  AND2_X1 _12742_ (
    .A1(_00947_),
    .A2(_00967_),
    .ZN(_00968_)
  );
  AND2_X1 _12743_ (
    .A1(reg_pmp_4_addr[16]),
    .A2(_00968_),
    .ZN(_00969_)
  );
  INV_X1 _12744_ (
    .A(_00969_),
    .ZN(_00970_)
  );
  AND2_X1 _12745_ (
    .A1(reg_pmp_6_cfg_r),
    .A2(_00894_),
    .ZN(_00971_)
  );
  INV_X1 _12746_ (
    .A(_00971_),
    .ZN(_00972_)
  );
  AND2_X1 _12747_ (
    .A1(_00970_),
    .A2(_00972_),
    .ZN(_00973_)
  );
  AND2_X1 _12748_ (
    .A1(_00965_),
    .A2(_00973_),
    .ZN(_00974_)
  );
  AND2_X1 _12749_ (
    .A1(_00957_),
    .A2(_00974_),
    .ZN(_00975_)
  );
  AND2_X1 _12750_ (
    .A1(_00933_),
    .A2(_00975_),
    .ZN(_00976_)
  );
  AND2_X1 _12751_ (
    .A1(io_rw_addr[1]),
    .A2(_00947_),
    .ZN(_00977_)
  );
  AND2_X1 _12752_ (
    .A1(_00966_),
    .A2(_00977_),
    .ZN(_00978_)
  );
  AND2_X1 _12753_ (
    .A1(reg_pmp_6_addr[16]),
    .A2(_00978_),
    .ZN(_00979_)
  );
  INV_X1 _12754_ (
    .A(_00979_),
    .ZN(_00980_)
  );
  AND2_X1 _12755_ (
    .A1(io_rw_addr[11]),
    .A2(_00886_),
    .ZN(_00981_)
  );
  AND2_X1 _12756_ (
    .A1(_00828_),
    .A2(_00920_),
    .ZN(_00982_)
  );
  AND2_X1 _12757_ (
    .A1(_00981_),
    .A2(_00982_),
    .ZN(_00983_)
  );
  AND2_X1 _12758_ (
    .A1(_00934_),
    .A2(_00983_),
    .ZN(_00984_)
  );
  AND2_X1 _12759_ (
    .A1(_00951_),
    .A2(_00984_),
    .ZN(_00985_)
  );
  AND2_X1 _12760_ (
    .A1(large_[10]),
    .A2(_00985_),
    .ZN(_00986_)
  );
  INV_X1 _12761_ (
    .A(_00986_),
    .ZN(_00987_)
  );
  AND2_X1 _12762_ (
    .A1(_00980_),
    .A2(_00987_),
    .ZN(_00988_)
  );
  AND2_X1 _12763_ (
    .A1(_00828_),
    .A2(_00981_),
    .ZN(_00989_)
  );
  AND2_X1 _12764_ (
    .A1(_00889_),
    .A2(_00983_),
    .ZN(_00990_)
  );
  AND2_X1 _12765_ (
    .A1(_00951_),
    .A2(_00990_),
    .ZN(_00991_)
  );
  INV_X1 _12766_ (
    .A(_00991_),
    .ZN(_00992_)
  );
  AND2_X1 _12767_ (
    .A1(large_[42]),
    .A2(_00991_),
    .ZN(_00993_)
  );
  INV_X1 _12768_ (
    .A(_00993_),
    .ZN(_00994_)
  );
  AND2_X1 _12769_ (
    .A1(_00883_),
    .A2(_00984_),
    .ZN(_00995_)
  );
  INV_X1 _12770_ (
    .A(_00995_),
    .ZN(_00996_)
  );
  AND2_X1 _12771_ (
    .A1(large_1[10]),
    .A2(_00995_),
    .ZN(_00997_)
  );
  INV_X1 _12772_ (
    .A(_00997_),
    .ZN(_00998_)
  );
  AND2_X1 _12773_ (
    .A1(_00994_),
    .A2(_00998_),
    .ZN(_00999_)
  );
  AND2_X1 _12774_ (
    .A1(_00988_),
    .A2(_00999_),
    .ZN(_01000_)
  );
  AND2_X1 _12775_ (
    .A1(_00923_),
    .A2(_00951_),
    .ZN(_01001_)
  );
  AND2_X1 _12776_ (
    .A1(reg_mcause[16]),
    .A2(_01001_),
    .ZN(_01002_)
  );
  INV_X1 _12777_ (
    .A(_01002_),
    .ZN(_01003_)
  );
  AND2_X1 _12778_ (
    .A1(_00915_),
    .A2(_00947_),
    .ZN(_01004_)
  );
  AND2_X1 _12779_ (
    .A1(reg_pmp_0_addr[16]),
    .A2(_01004_),
    .ZN(_01005_)
  );
  INV_X1 _12780_ (
    .A(_01005_),
    .ZN(_01006_)
  );
  AND2_X1 _12781_ (
    .A1(_01003_),
    .A2(_01006_),
    .ZN(_01007_)
  );
  AND2_X1 _12782_ (
    .A1(_00884_),
    .A2(_00947_),
    .ZN(_01008_)
  );
  AND2_X1 _12783_ (
    .A1(reg_pmp_1_addr[16]),
    .A2(_01008_),
    .ZN(_01009_)
  );
  INV_X1 _12784_ (
    .A(_01009_),
    .ZN(_01010_)
  );
  AND2_X1 _12785_ (
    .A1(_00925_),
    .A2(_00947_),
    .ZN(_01011_)
  );
  AND2_X1 _12786_ (
    .A1(reg_pmp_3_addr[16]),
    .A2(_01011_),
    .ZN(_01012_)
  );
  INV_X1 _12787_ (
    .A(_01012_),
    .ZN(_01013_)
  );
  AND2_X1 _12788_ (
    .A1(_01010_),
    .A2(_01013_),
    .ZN(_01014_)
  );
  AND2_X1 _12789_ (
    .A1(_01007_),
    .A2(_01014_),
    .ZN(_01015_)
  );
  AND2_X1 _12790_ (
    .A1(_00938_),
    .A2(_00977_),
    .ZN(_01016_)
  );
  AND2_X1 _12791_ (
    .A1(reg_pmp_7_addr[16]),
    .A2(_01016_),
    .ZN(_01017_)
  );
  INV_X1 _12792_ (
    .A(_01017_),
    .ZN(_01018_)
  );
  AND2_X1 _12793_ (
    .A1(_00883_),
    .A2(_00990_),
    .ZN(_01019_)
  );
  INV_X1 _12794_ (
    .A(_01019_),
    .ZN(_01020_)
  );
  AND2_X1 _12795_ (
    .A1(large_1[42]),
    .A2(_01019_),
    .ZN(_01021_)
  );
  INV_X1 _12796_ (
    .A(_01021_),
    .ZN(_01022_)
  );
  AND2_X1 _12797_ (
    .A1(_01018_),
    .A2(_01022_),
    .ZN(_01023_)
  );
  AND2_X1 _12798_ (
    .A1(_01015_),
    .A2(_01023_),
    .ZN(_01024_)
  );
  AND2_X1 _12799_ (
    .A1(_01000_),
    .A2(_01024_),
    .ZN(_01025_)
  );
  AND2_X1 _12800_ (
    .A1(_00935_),
    .A2(_00989_),
    .ZN(_01026_)
  );
  AND2_X1 _12801_ (
    .A1(_00951_),
    .A2(_01026_),
    .ZN(_01027_)
  );
  INV_X1 _12802_ (
    .A(_01027_),
    .ZN(_01028_)
  );
  AND2_X1 _12803_ (
    .A1(_00883_),
    .A2(_01026_),
    .ZN(_01029_)
  );
  AND2_X1 _12804_ (
    .A1(_00976_),
    .A2(_01025_),
    .ZN(_01030_)
  );
  INV_X1 _12805_ (
    .A(_01030_),
    .ZN(io_rw_rdata[16])
  );
  AND2_X1 _12806_ (
    .A1(io_rw_cmd[1]),
    .A2(_00851_),
    .ZN(_01031_)
  );
  AND2_X1 _12807_ (
    .A1(io_rw_rdata[16]),
    .A2(_01031_),
    .ZN(_01032_)
  );
  INV_X1 _12808_ (
    .A(_01032_),
    .ZN(_01033_)
  );
  AND2_X1 _12809_ (
    .A1(_00905_),
    .A2(_01033_),
    .ZN(_01034_)
  );
  INV_X1 _12810_ (
    .A(_01034_),
    .ZN(_01035_)
  );
  MUX2_X1 _12811_ (
    .A(reg_pmp_6_cfg_r),
    .B(_01035_),
    .S(_00900_),
    .Z(_00019_)
  );
  AND2_X1 _12812_ (
    .A1(io_rw_wdata[18]),
    .A2(_00903_),
    .ZN(_01036_)
  );
  INV_X1 _12813_ (
    .A(_01036_),
    .ZN(_01037_)
  );
  AND2_X1 _12814_ (
    .A1(reg_pmp_2_cfg_x),
    .A2(_00916_),
    .ZN(_01038_)
  );
  INV_X1 _12815_ (
    .A(_01038_),
    .ZN(_01039_)
  );
  AND2_X1 _12816_ (
    .A1(reg_pmp_3_addr[18]),
    .A2(_01011_),
    .ZN(_01040_)
  );
  INV_X1 _12817_ (
    .A(_01040_),
    .ZN(_01041_)
  );
  AND2_X1 _12818_ (
    .A1(_01039_),
    .A2(_01041_),
    .ZN(_01042_)
  );
  AND2_X1 _12819_ (
    .A1(reg_mepc[18]),
    .A2(_00943_),
    .ZN(_01043_)
  );
  INV_X1 _12820_ (
    .A(_01043_),
    .ZN(_01044_)
  );
  AND2_X1 _12821_ (
    .A1(reg_mtval[18]),
    .A2(_00926_),
    .ZN(_01045_)
  );
  INV_X1 _12822_ (
    .A(_01045_),
    .ZN(_01046_)
  );
  AND2_X1 _12823_ (
    .A1(_01044_),
    .A2(_01046_),
    .ZN(_01047_)
  );
  AND2_X1 _12824_ (
    .A1(_01042_),
    .A2(_01047_),
    .ZN(_01048_)
  );
  AND2_X1 _12825_ (
    .A1(reg_mcause[18]),
    .A2(_01001_),
    .ZN(_01049_)
  );
  INV_X1 _12826_ (
    .A(_01049_),
    .ZN(_01050_)
  );
  AND2_X1 _12827_ (
    .A1(reg_pmp_0_addr[18]),
    .A2(_01004_),
    .ZN(_01051_)
  );
  INV_X1 _12828_ (
    .A(_01051_),
    .ZN(_01052_)
  );
  AND2_X1 _12829_ (
    .A1(_01050_),
    .A2(_01052_),
    .ZN(_01053_)
  );
  AND2_X1 _12830_ (
    .A1(reg_dpc[18]),
    .A2(_00912_),
    .ZN(_01054_)
  );
  INV_X1 _12831_ (
    .A(_01054_),
    .ZN(_01055_)
  );
  AND2_X1 _12832_ (
    .A1(reg_pmp_2_addr[18]),
    .A2(_00953_),
    .ZN(_01056_)
  );
  INV_X1 _12833_ (
    .A(_01056_),
    .ZN(_01057_)
  );
  AND2_X1 _12834_ (
    .A1(_01055_),
    .A2(_01057_),
    .ZN(_01058_)
  );
  AND2_X1 _12835_ (
    .A1(_01053_),
    .A2(_01058_),
    .ZN(_01059_)
  );
  AND2_X1 _12836_ (
    .A1(reg_pmp_4_addr[18]),
    .A2(_00968_),
    .ZN(_01060_)
  );
  INV_X1 _12837_ (
    .A(_01060_),
    .ZN(_01061_)
  );
  AND2_X1 _12838_ (
    .A1(reg_mtvec[18]),
    .A2(_00940_),
    .ZN(_01062_)
  );
  INV_X1 _12839_ (
    .A(_01062_),
    .ZN(_01063_)
  );
  AND2_X1 _12840_ (
    .A1(_01061_),
    .A2(_01063_),
    .ZN(_01064_)
  );
  AND2_X1 _12841_ (
    .A1(reg_mscratch[18]),
    .A2(_00929_),
    .ZN(_01065_)
  );
  INV_X1 _12842_ (
    .A(_01065_),
    .ZN(_01066_)
  );
  AND2_X1 _12843_ (
    .A1(reg_pmp_6_cfg_x),
    .A2(_00894_),
    .ZN(_01067_)
  );
  INV_X1 _12844_ (
    .A(_01067_),
    .ZN(_01068_)
  );
  AND2_X1 _12845_ (
    .A1(_01066_),
    .A2(_01068_),
    .ZN(_01069_)
  );
  AND2_X1 _12846_ (
    .A1(_01064_),
    .A2(_01069_),
    .ZN(_01070_)
  );
  AND2_X1 _12847_ (
    .A1(_01059_),
    .A2(_01070_),
    .ZN(_01071_)
  );
  AND2_X1 _12848_ (
    .A1(_01048_),
    .A2(_01071_),
    .ZN(_01072_)
  );
  AND2_X1 _12849_ (
    .A1(large_1[44]),
    .A2(_01019_),
    .ZN(_01073_)
  );
  INV_X1 _12850_ (
    .A(_01073_),
    .ZN(_01074_)
  );
  AND2_X1 _12851_ (
    .A1(large_1[12]),
    .A2(_00995_),
    .ZN(_01075_)
  );
  INV_X1 _12852_ (
    .A(_01075_),
    .ZN(_01076_)
  );
  AND2_X1 _12853_ (
    .A1(_01074_),
    .A2(_01076_),
    .ZN(_01077_)
  );
  AND2_X1 _12854_ (
    .A1(large_[44]),
    .A2(_00991_),
    .ZN(_01078_)
  );
  INV_X1 _12855_ (
    .A(_01078_),
    .ZN(_01079_)
  );
  AND2_X1 _12856_ (
    .A1(large_[12]),
    .A2(_00985_),
    .ZN(_01080_)
  );
  INV_X1 _12857_ (
    .A(_01080_),
    .ZN(_01081_)
  );
  AND2_X1 _12858_ (
    .A1(_01079_),
    .A2(_01081_),
    .ZN(_01082_)
  );
  AND2_X1 _12859_ (
    .A1(_01077_),
    .A2(_01082_),
    .ZN(_01083_)
  );
  AND2_X1 _12860_ (
    .A1(reg_pmp_5_addr[18]),
    .A2(_00948_),
    .ZN(_01084_)
  );
  INV_X1 _12861_ (
    .A(_01084_),
    .ZN(_01085_)
  );
  AND2_X1 _12862_ (
    .A1(reg_bp_0_address[18]),
    .A2(_00962_),
    .ZN(_01086_)
  );
  INV_X1 _12863_ (
    .A(_01086_),
    .ZN(_01087_)
  );
  AND2_X1 _12864_ (
    .A1(_01085_),
    .A2(_01087_),
    .ZN(_01088_)
  );
  AND2_X1 _12865_ (
    .A1(reg_dscratch0[18]),
    .A2(_00958_),
    .ZN(_01089_)
  );
  INV_X1 _12866_ (
    .A(_01089_),
    .ZN(_01090_)
  );
  AND2_X1 _12867_ (
    .A1(reg_pmp_1_addr[18]),
    .A2(_01008_),
    .ZN(_01091_)
  );
  INV_X1 _12868_ (
    .A(_01091_),
    .ZN(_01092_)
  );
  AND2_X1 _12869_ (
    .A1(_01090_),
    .A2(_01092_),
    .ZN(_01093_)
  );
  AND2_X1 _12870_ (
    .A1(_01088_),
    .A2(_01093_),
    .ZN(_01094_)
  );
  AND2_X1 _12871_ (
    .A1(reg_pmp_6_addr[18]),
    .A2(_00978_),
    .ZN(_01095_)
  );
  INV_X1 _12872_ (
    .A(_01095_),
    .ZN(_01096_)
  );
  AND2_X1 _12873_ (
    .A1(reg_pmp_7_addr[18]),
    .A2(_01016_),
    .ZN(_01097_)
  );
  INV_X1 _12874_ (
    .A(_01097_),
    .ZN(_01098_)
  );
  AND2_X1 _12875_ (
    .A1(_01096_),
    .A2(_01098_),
    .ZN(_01099_)
  );
  AND2_X1 _12876_ (
    .A1(_01094_),
    .A2(_01099_),
    .ZN(_01100_)
  );
  AND2_X1 _12877_ (
    .A1(_01083_),
    .A2(_01100_),
    .ZN(_01101_)
  );
  AND2_X1 _12878_ (
    .A1(_01072_),
    .A2(_01101_),
    .ZN(_01102_)
  );
  INV_X1 _12879_ (
    .A(_01102_),
    .ZN(io_rw_rdata[18])
  );
  AND2_X1 _12880_ (
    .A1(io_rw_cmd[1]),
    .A2(_00853_),
    .ZN(_01103_)
  );
  AND2_X1 _12881_ (
    .A1(io_rw_rdata[18]),
    .A2(_01103_),
    .ZN(_01104_)
  );
  INV_X1 _12882_ (
    .A(_01104_),
    .ZN(_01105_)
  );
  AND2_X1 _12883_ (
    .A1(_01037_),
    .A2(_01105_),
    .ZN(_01106_)
  );
  INV_X1 _12884_ (
    .A(_01106_),
    .ZN(_01107_)
  );
  MUX2_X1 _12885_ (
    .A(reg_pmp_6_cfg_x),
    .B(_01107_),
    .S(_00900_),
    .Z(_00020_)
  );
  AND2_X1 _12886_ (
    .A1(io_rw_cmd[2]),
    .A2(_00895_),
    .ZN(_01108_)
  );
  AND2_X1 _12887_ (
    .A1(_00937_),
    .A2(_01108_),
    .ZN(_01109_)
  );
  AND2_X1 _12888_ (
    .A1(_00936_),
    .A2(_01109_),
    .ZN(_01110_)
  );
  INV_X1 _12889_ (
    .A(_01110_),
    .ZN(_01111_)
  );
  AND2_X1 _12890_ (
    .A1(_00879_),
    .A2(_01111_),
    .ZN(_01112_)
  );
  INV_X1 _12891_ (
    .A(_01112_),
    .ZN(_01113_)
  );
  AND2_X1 _12892_ (
    .A1(_00811_),
    .A2(_01113_),
    .ZN(_00021_)
  );
  AND2_X1 _12893_ (
    .A1(_00810_),
    .A2(_00901_),
    .ZN(_01114_)
  );
  INV_X1 _12894_ (
    .A(_01114_),
    .ZN(_01115_)
  );
  AND2_X1 _12895_ (
    .A1(_00811_),
    .A2(_01115_),
    .ZN(_01116_)
  );
  AND2_X1 _12896_ (
    .A1(io_rw_wdata[19]),
    .A2(_00903_),
    .ZN(_01117_)
  );
  INV_X1 _12897_ (
    .A(_01117_),
    .ZN(_01118_)
  );
  AND2_X1 _12898_ (
    .A1(io_rw_cmd[1]),
    .A2(_00854_),
    .ZN(_01119_)
  );
  AND2_X1 _12899_ (
    .A1(reg_bp_0_address[19]),
    .A2(_00962_),
    .ZN(_01120_)
  );
  INV_X1 _12900_ (
    .A(_01120_),
    .ZN(_01121_)
  );
  AND2_X1 _12901_ (
    .A1(reg_pmp_5_addr[19]),
    .A2(_00948_),
    .ZN(_01122_)
  );
  INV_X1 _12902_ (
    .A(_01122_),
    .ZN(_01123_)
  );
  AND2_X1 _12903_ (
    .A1(_01121_),
    .A2(_01123_),
    .ZN(_01124_)
  );
  AND2_X1 _12904_ (
    .A1(reg_pmp_2_cfg_a[0]),
    .A2(_00916_),
    .ZN(_01125_)
  );
  INV_X1 _12905_ (
    .A(_01125_),
    .ZN(_01126_)
  );
  AND2_X1 _12906_ (
    .A1(_00825_),
    .A2(io_rw_addr[4]),
    .ZN(_01127_)
  );
  AND2_X1 _12907_ (
    .A1(io_rw_addr[10]),
    .A2(_01127_),
    .ZN(_01128_)
  );
  AND2_X1 _12908_ (
    .A1(_00934_),
    .A2(_01128_),
    .ZN(_01129_)
  );
  AND2_X1 _12909_ (
    .A1(_00981_),
    .A2(_01129_),
    .ZN(_01130_)
  );
  AND2_X1 _12910_ (
    .A1(_00925_),
    .A2(_01130_),
    .ZN(_01131_)
  );
  INV_X1 _12911_ (
    .A(_01131_),
    .ZN(_01132_)
  );
  AND2_X1 _12912_ (
    .A1(_01126_),
    .A2(_01132_),
    .ZN(_01133_)
  );
  AND2_X1 _12913_ (
    .A1(_01124_),
    .A2(_01133_),
    .ZN(_01134_)
  );
  AND2_X1 _12914_ (
    .A1(reg_mtvec[19]),
    .A2(_00940_),
    .ZN(_01135_)
  );
  INV_X1 _12915_ (
    .A(_01135_),
    .ZN(_01136_)
  );
  AND2_X1 _12916_ (
    .A1(reg_dpc[19]),
    .A2(_00912_),
    .ZN(_01137_)
  );
  INV_X1 _12917_ (
    .A(_01137_),
    .ZN(_01138_)
  );
  AND2_X1 _12918_ (
    .A1(_01136_),
    .A2(_01138_),
    .ZN(_01139_)
  );
  AND2_X1 _12919_ (
    .A1(reg_mepc[19]),
    .A2(_00943_),
    .ZN(_01140_)
  );
  INV_X1 _12920_ (
    .A(_01140_),
    .ZN(_01141_)
  );
  AND2_X1 _12921_ (
    .A1(reg_mcause[19]),
    .A2(_01001_),
    .ZN(_01142_)
  );
  INV_X1 _12922_ (
    .A(_01142_),
    .ZN(_01143_)
  );
  AND2_X1 _12923_ (
    .A1(_01141_),
    .A2(_01143_),
    .ZN(_01144_)
  );
  AND2_X1 _12924_ (
    .A1(_01139_),
    .A2(_01144_),
    .ZN(_01145_)
  );
  AND2_X1 _12925_ (
    .A1(_01134_),
    .A2(_01145_),
    .ZN(_01146_)
  );
  AND2_X1 _12926_ (
    .A1(reg_pmp_2_addr[19]),
    .A2(_00953_),
    .ZN(_01147_)
  );
  INV_X1 _12927_ (
    .A(_01147_),
    .ZN(_01148_)
  );
  AND2_X1 _12928_ (
    .A1(reg_pmp_6_cfg_a[0]),
    .A2(_00894_),
    .ZN(_01149_)
  );
  INV_X1 _12929_ (
    .A(_01149_),
    .ZN(_01150_)
  );
  AND2_X1 _12930_ (
    .A1(reg_pmp_4_addr[19]),
    .A2(_00968_),
    .ZN(_01151_)
  );
  INV_X1 _12931_ (
    .A(_01151_),
    .ZN(_01152_)
  );
  AND2_X1 _12932_ (
    .A1(_01150_),
    .A2(_01152_),
    .ZN(_01153_)
  );
  AND2_X1 _12933_ (
    .A1(_01148_),
    .A2(_01153_),
    .ZN(_01154_)
  );
  AND2_X1 _12934_ (
    .A1(reg_dscratch0[19]),
    .A2(_00958_),
    .ZN(_01155_)
  );
  INV_X1 _12935_ (
    .A(_01155_),
    .ZN(_01156_)
  );
  AND2_X1 _12936_ (
    .A1(reg_pmp_1_addr[19]),
    .A2(_01008_),
    .ZN(_01157_)
  );
  INV_X1 _12937_ (
    .A(_01157_),
    .ZN(_01158_)
  );
  AND2_X1 _12938_ (
    .A1(_01156_),
    .A2(_01158_),
    .ZN(_01159_)
  );
  AND2_X1 _12939_ (
    .A1(reg_mtval[19]),
    .A2(_00926_),
    .ZN(_01160_)
  );
  INV_X1 _12940_ (
    .A(_01160_),
    .ZN(_01161_)
  );
  AND2_X1 _12941_ (
    .A1(reg_pmp_3_addr[19]),
    .A2(_01011_),
    .ZN(_01162_)
  );
  INV_X1 _12942_ (
    .A(_01162_),
    .ZN(_01163_)
  );
  AND2_X1 _12943_ (
    .A1(_01161_),
    .A2(_01163_),
    .ZN(_01164_)
  );
  AND2_X1 _12944_ (
    .A1(_01159_),
    .A2(_01164_),
    .ZN(_01165_)
  );
  AND2_X1 _12945_ (
    .A1(_01154_),
    .A2(_01165_),
    .ZN(_01166_)
  );
  AND2_X1 _12946_ (
    .A1(_01146_),
    .A2(_01166_),
    .ZN(_01167_)
  );
  AND2_X1 _12947_ (
    .A1(large_1[45]),
    .A2(_01019_),
    .ZN(_01168_)
  );
  INV_X1 _12948_ (
    .A(_01168_),
    .ZN(_01169_)
  );
  AND2_X1 _12949_ (
    .A1(reg_pmp_7_addr[19]),
    .A2(_01016_),
    .ZN(_01170_)
  );
  INV_X1 _12950_ (
    .A(_01170_),
    .ZN(_01171_)
  );
  AND2_X1 _12951_ (
    .A1(large_[13]),
    .A2(_00985_),
    .ZN(_01172_)
  );
  INV_X1 _12952_ (
    .A(_01172_),
    .ZN(_01173_)
  );
  AND2_X1 _12953_ (
    .A1(_01171_),
    .A2(_01173_),
    .ZN(_01174_)
  );
  AND2_X1 _12954_ (
    .A1(_01169_),
    .A2(_01174_),
    .ZN(_01175_)
  );
  AND2_X1 _12955_ (
    .A1(large_[45]),
    .A2(_00991_),
    .ZN(_01176_)
  );
  INV_X1 _12956_ (
    .A(_01176_),
    .ZN(_01177_)
  );
  AND2_X1 _12957_ (
    .A1(reg_pmp_0_addr[19]),
    .A2(_01004_),
    .ZN(_01178_)
  );
  INV_X1 _12958_ (
    .A(_01178_),
    .ZN(_01179_)
  );
  AND2_X1 _12959_ (
    .A1(reg_mscratch[19]),
    .A2(_00929_),
    .ZN(_01180_)
  );
  INV_X1 _12960_ (
    .A(_01180_),
    .ZN(_01181_)
  );
  AND2_X1 _12961_ (
    .A1(_01179_),
    .A2(_01181_),
    .ZN(_01182_)
  );
  AND2_X1 _12962_ (
    .A1(_01177_),
    .A2(_01182_),
    .ZN(_01183_)
  );
  AND2_X1 _12963_ (
    .A1(reg_pmp_6_addr[19]),
    .A2(_00978_),
    .ZN(_01184_)
  );
  INV_X1 _12964_ (
    .A(_01184_),
    .ZN(_01185_)
  );
  AND2_X1 _12965_ (
    .A1(large_1[13]),
    .A2(_00995_),
    .ZN(_01186_)
  );
  INV_X1 _12966_ (
    .A(_01186_),
    .ZN(_01187_)
  );
  AND2_X1 _12967_ (
    .A1(_01185_),
    .A2(_01187_),
    .ZN(_01188_)
  );
  AND2_X1 _12968_ (
    .A1(_01183_),
    .A2(_01188_),
    .ZN(_01189_)
  );
  AND2_X1 _12969_ (
    .A1(_01175_),
    .A2(_01189_),
    .ZN(_01190_)
  );
  AND2_X1 _12970_ (
    .A1(_01167_),
    .A2(_01190_),
    .ZN(_01191_)
  );
  INV_X1 _12971_ (
    .A(_01191_),
    .ZN(io_rw_rdata[19])
  );
  AND2_X1 _12972_ (
    .A1(_01119_),
    .A2(io_rw_rdata[19]),
    .ZN(_01192_)
  );
  INV_X1 _12973_ (
    .A(_01192_),
    .ZN(_01193_)
  );
  AND2_X1 _12974_ (
    .A1(io_rw_addr[4]),
    .A2(io_rw_addr[10]),
    .ZN(_01194_)
  );
  AND2_X1 _12975_ (
    .A1(_00825_),
    .A2(_00934_),
    .ZN(_01195_)
  );
  AND2_X1 _12976_ (
    .A1(_00981_),
    .A2(_01195_),
    .ZN(_01196_)
  );
  AND2_X1 _12977_ (
    .A1(_01194_),
    .A2(_01196_),
    .ZN(_01197_)
  );
  AND2_X1 _12978_ (
    .A1(_01118_),
    .A2(_01193_),
    .ZN(_01198_)
  );
  INV_X1 _12979_ (
    .A(_01198_),
    .ZN(_01199_)
  );
  AND2_X1 _12980_ (
    .A1(_00900_),
    .A2(_01198_),
    .ZN(_01200_)
  );
  INV_X1 _12981_ (
    .A(_01200_),
    .ZN(_01201_)
  );
  AND2_X1 _12982_ (
    .A1(_01116_),
    .A2(_01201_),
    .ZN(_00022_)
  );
  AND2_X1 _12983_ (
    .A1(_00809_),
    .A2(_00901_),
    .ZN(_01202_)
  );
  INV_X1 _12984_ (
    .A(_01202_),
    .ZN(_01203_)
  );
  AND2_X1 _12985_ (
    .A1(_00811_),
    .A2(_01203_),
    .ZN(_01204_)
  );
  AND2_X1 _12986_ (
    .A1(io_rw_wdata[20]),
    .A2(_00903_),
    .ZN(_01205_)
  );
  INV_X1 _12987_ (
    .A(_01205_),
    .ZN(_01206_)
  );
  AND2_X1 _12988_ (
    .A1(reg_pmp_4_addr[20]),
    .A2(_00968_),
    .ZN(_01207_)
  );
  INV_X1 _12989_ (
    .A(_01207_),
    .ZN(_01208_)
  );
  AND2_X1 _12990_ (
    .A1(reg_bp_0_address[20]),
    .A2(_00962_),
    .ZN(_01209_)
  );
  INV_X1 _12991_ (
    .A(_01209_),
    .ZN(_01210_)
  );
  AND2_X1 _12992_ (
    .A1(_01208_),
    .A2(_01210_),
    .ZN(_01211_)
  );
  AND2_X1 _12993_ (
    .A1(reg_pmp_2_addr[20]),
    .A2(_00953_),
    .ZN(_01212_)
  );
  INV_X1 _12994_ (
    .A(_01212_),
    .ZN(_01213_)
  );
  AND2_X1 _12995_ (
    .A1(reg_dpc[20]),
    .A2(_00912_),
    .ZN(_01214_)
  );
  INV_X1 _12996_ (
    .A(_01214_),
    .ZN(_01215_)
  );
  AND2_X1 _12997_ (
    .A1(_01213_),
    .A2(_01215_),
    .ZN(_01216_)
  );
  AND2_X1 _12998_ (
    .A1(_01211_),
    .A2(_01216_),
    .ZN(_01217_)
  );
  AND2_X1 _12999_ (
    .A1(reg_pmp_2_cfg_a[1]),
    .A2(_00916_),
    .ZN(_01218_)
  );
  INV_X1 _13000_ (
    .A(_01218_),
    .ZN(_01219_)
  );
  AND2_X1 _13001_ (
    .A1(reg_pmp_5_addr[20]),
    .A2(_00948_),
    .ZN(_01220_)
  );
  INV_X1 _13002_ (
    .A(_01220_),
    .ZN(_01221_)
  );
  AND2_X1 _13003_ (
    .A1(_01219_),
    .A2(_01221_),
    .ZN(_01222_)
  );
  AND2_X1 _13004_ (
    .A1(reg_mepc[20]),
    .A2(_00943_),
    .ZN(_01223_)
  );
  INV_X1 _13005_ (
    .A(_01223_),
    .ZN(_01224_)
  );
  AND2_X1 _13006_ (
    .A1(reg_mscratch[20]),
    .A2(_00929_),
    .ZN(_01225_)
  );
  INV_X1 _13007_ (
    .A(_01225_),
    .ZN(_01226_)
  );
  AND2_X1 _13008_ (
    .A1(_01224_),
    .A2(_01226_),
    .ZN(_01227_)
  );
  AND2_X1 _13009_ (
    .A1(_01222_),
    .A2(_01227_),
    .ZN(_01228_)
  );
  AND2_X1 _13010_ (
    .A1(_01217_),
    .A2(_01228_),
    .ZN(_01229_)
  );
  AND2_X1 _13011_ (
    .A1(reg_pmp_0_addr[20]),
    .A2(_01004_),
    .ZN(_01230_)
  );
  INV_X1 _13012_ (
    .A(_01230_),
    .ZN(_01231_)
  );
  AND2_X1 _13013_ (
    .A1(reg_pmp_3_addr[20]),
    .A2(_01011_),
    .ZN(_01232_)
  );
  INV_X1 _13014_ (
    .A(_01232_),
    .ZN(_01233_)
  );
  AND2_X1 _13015_ (
    .A1(reg_pmp_1_addr[20]),
    .A2(_01008_),
    .ZN(_01234_)
  );
  INV_X1 _13016_ (
    .A(_01234_),
    .ZN(_01235_)
  );
  AND2_X1 _13017_ (
    .A1(_01233_),
    .A2(_01235_),
    .ZN(_01236_)
  );
  AND2_X1 _13018_ (
    .A1(_01231_),
    .A2(_01236_),
    .ZN(_01237_)
  );
  AND2_X1 _13019_ (
    .A1(reg_mtvec[20]),
    .A2(_00940_),
    .ZN(_01238_)
  );
  INV_X1 _13020_ (
    .A(_01238_),
    .ZN(_01239_)
  );
  AND2_X1 _13021_ (
    .A1(reg_mcause[20]),
    .A2(_01001_),
    .ZN(_01240_)
  );
  INV_X1 _13022_ (
    .A(_01240_),
    .ZN(_01241_)
  );
  AND2_X1 _13023_ (
    .A1(_01239_),
    .A2(_01241_),
    .ZN(_01242_)
  );
  AND2_X1 _13024_ (
    .A1(reg_mtval[20]),
    .A2(_00926_),
    .ZN(_01243_)
  );
  INV_X1 _13025_ (
    .A(_01243_),
    .ZN(_01244_)
  );
  AND2_X1 _13026_ (
    .A1(reg_dscratch0[20]),
    .A2(_00958_),
    .ZN(_01245_)
  );
  INV_X1 _13027_ (
    .A(_01245_),
    .ZN(_01246_)
  );
  AND2_X1 _13028_ (
    .A1(_01244_),
    .A2(_01246_),
    .ZN(_01247_)
  );
  AND2_X1 _13029_ (
    .A1(_01242_),
    .A2(_01247_),
    .ZN(_01248_)
  );
  AND2_X1 _13030_ (
    .A1(_01237_),
    .A2(_01248_),
    .ZN(_01249_)
  );
  AND2_X1 _13031_ (
    .A1(_01229_),
    .A2(_01249_),
    .ZN(_01250_)
  );
  AND2_X1 _13032_ (
    .A1(large_1[14]),
    .A2(_00995_),
    .ZN(_01251_)
  );
  INV_X1 _13033_ (
    .A(_01251_),
    .ZN(_01252_)
  );
  AND2_X1 _13034_ (
    .A1(reg_pmp_6_addr[20]),
    .A2(_00978_),
    .ZN(_01253_)
  );
  INV_X1 _13035_ (
    .A(_01253_),
    .ZN(_01254_)
  );
  AND2_X1 _13036_ (
    .A1(large_1[46]),
    .A2(_01019_),
    .ZN(_01255_)
  );
  INV_X1 _13037_ (
    .A(_01255_),
    .ZN(_01256_)
  );
  AND2_X1 _13038_ (
    .A1(_01254_),
    .A2(_01256_),
    .ZN(_01257_)
  );
  AND2_X1 _13039_ (
    .A1(_01252_),
    .A2(_01257_),
    .ZN(_01258_)
  );
  AND2_X1 _13040_ (
    .A1(large_[46]),
    .A2(_00991_),
    .ZN(_01259_)
  );
  INV_X1 _13041_ (
    .A(_01259_),
    .ZN(_01260_)
  );
  AND2_X1 _13042_ (
    .A1(reg_pmp_6_cfg_a[1]),
    .A2(_00894_),
    .ZN(_01261_)
  );
  INV_X1 _13043_ (
    .A(_01261_),
    .ZN(_01262_)
  );
  AND2_X1 _13044_ (
    .A1(_01132_),
    .A2(_01262_),
    .ZN(_01263_)
  );
  AND2_X1 _13045_ (
    .A1(_01260_),
    .A2(_01263_),
    .ZN(_01264_)
  );
  AND2_X1 _13046_ (
    .A1(reg_pmp_7_addr[20]),
    .A2(_01016_),
    .ZN(_01265_)
  );
  INV_X1 _13047_ (
    .A(_01265_),
    .ZN(_01266_)
  );
  AND2_X1 _13048_ (
    .A1(large_[14]),
    .A2(_00985_),
    .ZN(_01267_)
  );
  INV_X1 _13049_ (
    .A(_01267_),
    .ZN(_01268_)
  );
  AND2_X1 _13050_ (
    .A1(_01266_),
    .A2(_01268_),
    .ZN(_01269_)
  );
  AND2_X1 _13051_ (
    .A1(_01264_),
    .A2(_01269_),
    .ZN(_01270_)
  );
  AND2_X1 _13052_ (
    .A1(_01258_),
    .A2(_01270_),
    .ZN(_01271_)
  );
  AND2_X1 _13053_ (
    .A1(_01250_),
    .A2(_01271_),
    .ZN(_01272_)
  );
  INV_X1 _13054_ (
    .A(_01272_),
    .ZN(io_rw_rdata[20])
  );
  AND2_X1 _13055_ (
    .A1(io_rw_cmd[1]),
    .A2(_00855_),
    .ZN(_01273_)
  );
  AND2_X1 _13056_ (
    .A1(io_rw_rdata[20]),
    .A2(_01273_),
    .ZN(_01274_)
  );
  INV_X1 _13057_ (
    .A(_01274_),
    .ZN(_01275_)
  );
  AND2_X1 _13058_ (
    .A1(_01206_),
    .A2(_01275_),
    .ZN(_01276_)
  );
  INV_X1 _13059_ (
    .A(_01276_),
    .ZN(_01277_)
  );
  AND2_X1 _13060_ (
    .A1(_00900_),
    .A2(_01276_),
    .ZN(_01278_)
  );
  INV_X1 _13061_ (
    .A(_01278_),
    .ZN(_01279_)
  );
  AND2_X1 _13062_ (
    .A1(_01204_),
    .A2(_01279_),
    .ZN(_00023_)
  );
  AND2_X1 _13063_ (
    .A1(_00808_),
    .A2(_00901_),
    .ZN(_01280_)
  );
  INV_X1 _13064_ (
    .A(_01280_),
    .ZN(_01281_)
  );
  AND2_X1 _13065_ (
    .A1(_00811_),
    .A2(_01281_),
    .ZN(_01282_)
  );
  AND2_X1 _13066_ (
    .A1(io_rw_wdata[23]),
    .A2(_00903_),
    .ZN(_01283_)
  );
  INV_X1 _13067_ (
    .A(_01283_),
    .ZN(_01284_)
  );
  AND2_X1 _13068_ (
    .A1(reg_pmp_5_addr[23]),
    .A2(_00948_),
    .ZN(_01285_)
  );
  INV_X1 _13069_ (
    .A(_01285_),
    .ZN(_01286_)
  );
  AND2_X1 _13070_ (
    .A1(reg_bp_0_address[23]),
    .A2(_00962_),
    .ZN(_01287_)
  );
  INV_X1 _13071_ (
    .A(_01287_),
    .ZN(_01288_)
  );
  AND2_X1 _13072_ (
    .A1(_01286_),
    .A2(_01288_),
    .ZN(_01289_)
  );
  AND2_X1 _13073_ (
    .A1(reg_pmp_2_addr[23]),
    .A2(_00953_),
    .ZN(_01290_)
  );
  INV_X1 _13074_ (
    .A(_01290_),
    .ZN(_01291_)
  );
  AND2_X1 _13075_ (
    .A1(reg_pmp_0_addr[23]),
    .A2(_01004_),
    .ZN(_01292_)
  );
  INV_X1 _13076_ (
    .A(_01292_),
    .ZN(_01293_)
  );
  AND2_X1 _13077_ (
    .A1(_01291_),
    .A2(_01293_),
    .ZN(_01294_)
  );
  AND2_X1 _13078_ (
    .A1(_01289_),
    .A2(_01294_),
    .ZN(_01295_)
  );
  AND2_X1 _13079_ (
    .A1(reg_pmp_4_addr[23]),
    .A2(_00968_),
    .ZN(_01296_)
  );
  INV_X1 _13080_ (
    .A(_01296_),
    .ZN(_01297_)
  );
  AND2_X1 _13081_ (
    .A1(reg_mtvec[23]),
    .A2(_00940_),
    .ZN(_01298_)
  );
  INV_X1 _13082_ (
    .A(_01298_),
    .ZN(_01299_)
  );
  AND2_X1 _13083_ (
    .A1(_01297_),
    .A2(_01299_),
    .ZN(_01300_)
  );
  AND2_X1 _13084_ (
    .A1(reg_dpc[23]),
    .A2(_00912_),
    .ZN(_01301_)
  );
  INV_X1 _13085_ (
    .A(_01301_),
    .ZN(_01302_)
  );
  AND2_X1 _13086_ (
    .A1(reg_pmp_1_addr[23]),
    .A2(_01008_),
    .ZN(_01303_)
  );
  INV_X1 _13087_ (
    .A(_01303_),
    .ZN(_01304_)
  );
  AND2_X1 _13088_ (
    .A1(_01302_),
    .A2(_01304_),
    .ZN(_01305_)
  );
  AND2_X1 _13089_ (
    .A1(_01300_),
    .A2(_01305_),
    .ZN(_01306_)
  );
  AND2_X1 _13090_ (
    .A1(_01295_),
    .A2(_01306_),
    .ZN(_01307_)
  );
  AND2_X1 _13091_ (
    .A1(reg_mcause[23]),
    .A2(_01001_),
    .ZN(_01308_)
  );
  INV_X1 _13092_ (
    .A(_01308_),
    .ZN(_01309_)
  );
  AND2_X1 _13093_ (
    .A1(reg_mtval[23]),
    .A2(_00926_),
    .ZN(_01310_)
  );
  INV_X1 _13094_ (
    .A(_01310_),
    .ZN(_01311_)
  );
  AND2_X1 _13095_ (
    .A1(reg_mscratch[23]),
    .A2(_00929_),
    .ZN(_01312_)
  );
  INV_X1 _13096_ (
    .A(_01312_),
    .ZN(_01313_)
  );
  AND2_X1 _13097_ (
    .A1(_01311_),
    .A2(_01313_),
    .ZN(_01314_)
  );
  AND2_X1 _13098_ (
    .A1(_01309_),
    .A2(_01314_),
    .ZN(_01315_)
  );
  AND2_X1 _13099_ (
    .A1(reg_pmp_2_cfg_l),
    .A2(_00916_),
    .ZN(_01316_)
  );
  INV_X1 _13100_ (
    .A(_01316_),
    .ZN(_01317_)
  );
  AND2_X1 _13101_ (
    .A1(reg_pmp_6_cfg_l),
    .A2(_00894_),
    .ZN(_01318_)
  );
  INV_X1 _13102_ (
    .A(_01318_),
    .ZN(_01319_)
  );
  AND2_X1 _13103_ (
    .A1(_01317_),
    .A2(_01319_),
    .ZN(_01320_)
  );
  AND2_X1 _13104_ (
    .A1(reg_dscratch0[23]),
    .A2(_00958_),
    .ZN(_01321_)
  );
  INV_X1 _13105_ (
    .A(_01321_),
    .ZN(_01322_)
  );
  AND2_X1 _13106_ (
    .A1(reg_pmp_3_addr[23]),
    .A2(_01011_),
    .ZN(_01323_)
  );
  INV_X1 _13107_ (
    .A(_01323_),
    .ZN(_01324_)
  );
  AND2_X1 _13108_ (
    .A1(_01322_),
    .A2(_01324_),
    .ZN(_01325_)
  );
  AND2_X1 _13109_ (
    .A1(_01320_),
    .A2(_01325_),
    .ZN(_01326_)
  );
  AND2_X1 _13110_ (
    .A1(_01315_),
    .A2(_01326_),
    .ZN(_01327_)
  );
  AND2_X1 _13111_ (
    .A1(_01307_),
    .A2(_01327_),
    .ZN(_01328_)
  );
  AND2_X1 _13112_ (
    .A1(large_1[17]),
    .A2(_00995_),
    .ZN(_01329_)
  );
  INV_X1 _13113_ (
    .A(_01329_),
    .ZN(_01330_)
  );
  AND2_X1 _13114_ (
    .A1(large_1[49]),
    .A2(_01019_),
    .ZN(_01331_)
  );
  INV_X1 _13115_ (
    .A(_01331_),
    .ZN(_01332_)
  );
  AND2_X1 _13116_ (
    .A1(reg_pmp_6_addr[23]),
    .A2(_00978_),
    .ZN(_01333_)
  );
  INV_X1 _13117_ (
    .A(_01333_),
    .ZN(_01334_)
  );
  AND2_X1 _13118_ (
    .A1(_01332_),
    .A2(_01334_),
    .ZN(_01335_)
  );
  AND2_X1 _13119_ (
    .A1(_01330_),
    .A2(_01335_),
    .ZN(_01336_)
  );
  AND2_X1 _13120_ (
    .A1(reg_pmp_7_addr[23]),
    .A2(_01016_),
    .ZN(_01337_)
  );
  INV_X1 _13121_ (
    .A(_01337_),
    .ZN(_01338_)
  );
  AND2_X1 _13122_ (
    .A1(_00884_),
    .A2(_00936_),
    .ZN(_01339_)
  );
  INV_X1 _13123_ (
    .A(_01339_),
    .ZN(_01340_)
  );
  AND2_X1 _13124_ (
    .A1(_00884_),
    .A2(_00961_),
    .ZN(_01341_)
  );
  INV_X1 _13125_ (
    .A(_01341_),
    .ZN(_01342_)
  );
  AND2_X1 _13126_ (
    .A1(_01340_),
    .A2(_01342_),
    .ZN(_01343_)
  );
  AND2_X1 _13127_ (
    .A1(reg_mepc[23]),
    .A2(_00943_),
    .ZN(_01344_)
  );
  INV_X1 _13128_ (
    .A(_01344_),
    .ZN(_01345_)
  );
  AND2_X1 _13129_ (
    .A1(_01343_),
    .A2(_01345_),
    .ZN(_01346_)
  );
  AND2_X1 _13130_ (
    .A1(_01338_),
    .A2(_01346_),
    .ZN(_01347_)
  );
  AND2_X1 _13131_ (
    .A1(large_[49]),
    .A2(_00991_),
    .ZN(_01348_)
  );
  INV_X1 _13132_ (
    .A(_01348_),
    .ZN(_01349_)
  );
  AND2_X1 _13133_ (
    .A1(large_[17]),
    .A2(_00985_),
    .ZN(_01350_)
  );
  INV_X1 _13134_ (
    .A(_01350_),
    .ZN(_01351_)
  );
  AND2_X1 _13135_ (
    .A1(_01349_),
    .A2(_01351_),
    .ZN(_01352_)
  );
  AND2_X1 _13136_ (
    .A1(_01347_),
    .A2(_01352_),
    .ZN(_01353_)
  );
  AND2_X1 _13137_ (
    .A1(_01336_),
    .A2(_01353_),
    .ZN(_01354_)
  );
  AND2_X1 _13138_ (
    .A1(_01328_),
    .A2(_01354_),
    .ZN(_01355_)
  );
  INV_X1 _13139_ (
    .A(_01355_),
    .ZN(io_rw_rdata[23])
  );
  AND2_X1 _13140_ (
    .A1(io_rw_cmd[1]),
    .A2(_00858_),
    .ZN(_01356_)
  );
  AND2_X1 _13141_ (
    .A1(io_rw_rdata[23]),
    .A2(_01356_),
    .ZN(_01357_)
  );
  INV_X1 _13142_ (
    .A(_01357_),
    .ZN(_01358_)
  );
  AND2_X1 _13143_ (
    .A1(_01284_),
    .A2(_01358_),
    .ZN(_01359_)
  );
  INV_X1 _13144_ (
    .A(_01359_),
    .ZN(_01360_)
  );
  AND2_X1 _13145_ (
    .A1(_00900_),
    .A2(_01359_),
    .ZN(_01361_)
  );
  INV_X1 _13146_ (
    .A(_01361_),
    .ZN(_01362_)
  );
  AND2_X1 _13147_ (
    .A1(_01282_),
    .A2(_01362_),
    .ZN(_00024_)
  );
  AND2_X1 _13148_ (
    .A1(_00015_),
    .A2(_00894_),
    .ZN(_01363_)
  );
  AND2_X1 _13149_ (
    .A1(_00897_),
    .A2(_01363_),
    .ZN(_01364_)
  );
  INV_X1 _13150_ (
    .A(_01364_),
    .ZN(_01365_)
  );
  AND2_X1 _13151_ (
    .A1(io_rw_wdata[8]),
    .A2(_00903_),
    .ZN(_01366_)
  );
  INV_X1 _13152_ (
    .A(_01366_),
    .ZN(_01367_)
  );
  AND2_X1 _13153_ (
    .A1(reg_pmp_0_addr[8]),
    .A2(_01004_),
    .ZN(_01368_)
  );
  INV_X1 _13154_ (
    .A(_01368_),
    .ZN(_01369_)
  );
  AND2_X1 _13155_ (
    .A1(reg_mtvec[8]),
    .A2(_00940_),
    .ZN(_01370_)
  );
  INV_X1 _13156_ (
    .A(_01370_),
    .ZN(_01371_)
  );
  AND2_X1 _13157_ (
    .A1(_01369_),
    .A2(_01371_),
    .ZN(_01372_)
  );
  AND2_X1 _13158_ (
    .A1(reg_mtval[8]),
    .A2(_00926_),
    .ZN(_01373_)
  );
  INV_X1 _13159_ (
    .A(_01373_),
    .ZN(_01374_)
  );
  AND2_X1 _13160_ (
    .A1(reg_dpc[8]),
    .A2(_00912_),
    .ZN(_01375_)
  );
  INV_X1 _13161_ (
    .A(_01375_),
    .ZN(_01376_)
  );
  AND2_X1 _13162_ (
    .A1(_01374_),
    .A2(_01376_),
    .ZN(_01377_)
  );
  AND2_X1 _13163_ (
    .A1(_01372_),
    .A2(_01377_),
    .ZN(_01378_)
  );
  AND2_X1 _13164_ (
    .A1(reg_bp_0_control_tmatch[1]),
    .A2(_01341_),
    .ZN(_01379_)
  );
  INV_X1 _13165_ (
    .A(_01379_),
    .ZN(_01380_)
  );
  AND2_X1 _13166_ (
    .A1(_00911_),
    .A2(_00915_),
    .ZN(_01381_)
  );
  INV_X1 _13167_ (
    .A(_01381_),
    .ZN(_01382_)
  );
  AND2_X1 _13168_ (
    .A1(reg_dcsr_cause[2]),
    .A2(_01381_),
    .ZN(_01383_)
  );
  INV_X1 _13169_ (
    .A(_01383_),
    .ZN(_01384_)
  );
  AND2_X1 _13170_ (
    .A1(_01380_),
    .A2(_01384_),
    .ZN(_01385_)
  );
  AND2_X1 _13171_ (
    .A1(reg_bp_0_address[8]),
    .A2(_00962_),
    .ZN(_01386_)
  );
  INV_X1 _13172_ (
    .A(_01386_),
    .ZN(_01387_)
  );
  AND2_X1 _13173_ (
    .A1(reg_dscratch0[8]),
    .A2(_00958_),
    .ZN(_01388_)
  );
  INV_X1 _13174_ (
    .A(_01388_),
    .ZN(_01389_)
  );
  AND2_X1 _13175_ (
    .A1(_01387_),
    .A2(_01389_),
    .ZN(_01390_)
  );
  AND2_X1 _13176_ (
    .A1(_01385_),
    .A2(_01390_),
    .ZN(_01391_)
  );
  AND2_X1 _13177_ (
    .A1(_01378_),
    .A2(_01391_),
    .ZN(_01392_)
  );
  AND2_X1 _13178_ (
    .A1(reg_pmp_4_addr[8]),
    .A2(_00968_),
    .ZN(_01393_)
  );
  INV_X1 _13179_ (
    .A(_01393_),
    .ZN(_01394_)
  );
  AND2_X1 _13180_ (
    .A1(reg_mscratch[8]),
    .A2(_00929_),
    .ZN(_01395_)
  );
  INV_X1 _13181_ (
    .A(_01395_),
    .ZN(_01396_)
  );
  AND2_X1 _13182_ (
    .A1(reg_mepc[8]),
    .A2(_00943_),
    .ZN(_01397_)
  );
  INV_X1 _13183_ (
    .A(_01397_),
    .ZN(_01398_)
  );
  AND2_X1 _13184_ (
    .A1(_01396_),
    .A2(_01398_),
    .ZN(_01399_)
  );
  AND2_X1 _13185_ (
    .A1(_01394_),
    .A2(_01399_),
    .ZN(_01400_)
  );
  AND2_X1 _13186_ (
    .A1(reg_pmp_2_addr[8]),
    .A2(_00953_),
    .ZN(_01401_)
  );
  INV_X1 _13187_ (
    .A(_01401_),
    .ZN(_01402_)
  );
  AND2_X1 _13188_ (
    .A1(reg_pmp_5_cfg_r),
    .A2(_00894_),
    .ZN(_01403_)
  );
  INV_X1 _13189_ (
    .A(_01403_),
    .ZN(_01404_)
  );
  AND2_X1 _13190_ (
    .A1(_01402_),
    .A2(_01404_),
    .ZN(_01405_)
  );
  AND2_X1 _13191_ (
    .A1(reg_pmp_1_cfg_r),
    .A2(_00916_),
    .ZN(_01406_)
  );
  INV_X1 _13192_ (
    .A(_01406_),
    .ZN(_01407_)
  );
  AND2_X1 _13193_ (
    .A1(reg_mcause[8]),
    .A2(_01001_),
    .ZN(_01408_)
  );
  INV_X1 _13194_ (
    .A(_01408_),
    .ZN(_01409_)
  );
  AND2_X1 _13195_ (
    .A1(_01407_),
    .A2(_01409_),
    .ZN(_01410_)
  );
  AND2_X1 _13196_ (
    .A1(_01405_),
    .A2(_01410_),
    .ZN(_01411_)
  );
  AND2_X1 _13197_ (
    .A1(_01400_),
    .A2(_01411_),
    .ZN(_01412_)
  );
  AND2_X1 _13198_ (
    .A1(_01392_),
    .A2(_01412_),
    .ZN(_01413_)
  );
  AND2_X1 _13199_ (
    .A1(reg_pmp_7_addr[8]),
    .A2(_01016_),
    .ZN(_01414_)
  );
  INV_X1 _13200_ (
    .A(_01414_),
    .ZN(_01415_)
  );
  AND2_X1 _13201_ (
    .A1(reg_pmp_6_addr[8]),
    .A2(_00978_),
    .ZN(_01416_)
  );
  INV_X1 _13202_ (
    .A(_01416_),
    .ZN(_01417_)
  );
  AND2_X1 _13203_ (
    .A1(_01415_),
    .A2(_01417_),
    .ZN(_01418_)
  );
  AND2_X1 _13204_ (
    .A1(large_[34]),
    .A2(_00991_),
    .ZN(_01419_)
  );
  INV_X1 _13205_ (
    .A(_01419_),
    .ZN(_01420_)
  );
  AND2_X1 _13206_ (
    .A1(large_[2]),
    .A2(_00985_),
    .ZN(_01421_)
  );
  INV_X1 _13207_ (
    .A(_01421_),
    .ZN(_01422_)
  );
  AND2_X1 _13208_ (
    .A1(_01420_),
    .A2(_01422_),
    .ZN(_01423_)
  );
  AND2_X1 _13209_ (
    .A1(_01418_),
    .A2(_01423_),
    .ZN(_01424_)
  );
  AND2_X1 _13210_ (
    .A1(reg_pmp_3_addr[8]),
    .A2(_01011_),
    .ZN(_01425_)
  );
  INV_X1 _13211_ (
    .A(_01425_),
    .ZN(_01426_)
  );
  AND2_X1 _13212_ (
    .A1(_01340_),
    .A2(_01426_),
    .ZN(_01427_)
  );
  AND2_X1 _13213_ (
    .A1(reg_pmp_5_addr[8]),
    .A2(_00948_),
    .ZN(_01428_)
  );
  INV_X1 _13214_ (
    .A(_01428_),
    .ZN(_01429_)
  );
  AND2_X1 _13215_ (
    .A1(reg_pmp_1_addr[8]),
    .A2(_01008_),
    .ZN(_01430_)
  );
  INV_X1 _13216_ (
    .A(_01430_),
    .ZN(_01431_)
  );
  AND2_X1 _13217_ (
    .A1(_01429_),
    .A2(_01431_),
    .ZN(_01432_)
  );
  AND2_X1 _13218_ (
    .A1(_01427_),
    .A2(_01432_),
    .ZN(_01433_)
  );
  AND2_X1 _13219_ (
    .A1(large_1[34]),
    .A2(_01019_),
    .ZN(_01434_)
  );
  INV_X1 _13220_ (
    .A(_01434_),
    .ZN(_01435_)
  );
  AND2_X1 _13221_ (
    .A1(large_1[2]),
    .A2(_00995_),
    .ZN(_01436_)
  );
  INV_X1 _13222_ (
    .A(_01436_),
    .ZN(_01437_)
  );
  AND2_X1 _13223_ (
    .A1(_01435_),
    .A2(_01437_),
    .ZN(_01438_)
  );
  AND2_X1 _13224_ (
    .A1(_01433_),
    .A2(_01438_),
    .ZN(_01439_)
  );
  AND2_X1 _13225_ (
    .A1(_01424_),
    .A2(_01439_),
    .ZN(_01440_)
  );
  AND2_X1 _13226_ (
    .A1(_01413_),
    .A2(_01440_),
    .ZN(_01441_)
  );
  INV_X1 _13227_ (
    .A(_01441_),
    .ZN(io_rw_rdata[8])
  );
  AND2_X1 _13228_ (
    .A1(io_rw_cmd[1]),
    .A2(_00844_),
    .ZN(_01442_)
  );
  AND2_X1 _13229_ (
    .A1(io_rw_rdata[8]),
    .A2(_01442_),
    .ZN(_01443_)
  );
  INV_X1 _13230_ (
    .A(_01443_),
    .ZN(_01444_)
  );
  AND2_X1 _13231_ (
    .A1(_01367_),
    .A2(_01444_),
    .ZN(_01445_)
  );
  INV_X1 _13232_ (
    .A(_01445_),
    .ZN(_01446_)
  );
  MUX2_X1 _13233_ (
    .A(reg_pmp_5_cfg_r),
    .B(_01446_),
    .S(_01364_),
    .Z(_00025_)
  );
  AND2_X1 _13234_ (
    .A1(io_rw_wdata[9]),
    .A2(_00903_),
    .ZN(_01447_)
  );
  INV_X1 _13235_ (
    .A(_01447_),
    .ZN(_01448_)
  );
  AND2_X1 _13236_ (
    .A1(reg_mscratch[9]),
    .A2(_00929_),
    .ZN(_01449_)
  );
  INV_X1 _13237_ (
    .A(_01449_),
    .ZN(_01450_)
  );
  AND2_X1 _13238_ (
    .A1(reg_mtvec[9]),
    .A2(_00940_),
    .ZN(_01451_)
  );
  INV_X1 _13239_ (
    .A(_01451_),
    .ZN(_01452_)
  );
  AND2_X1 _13240_ (
    .A1(_01450_),
    .A2(_01452_),
    .ZN(_01453_)
  );
  AND2_X1 _13241_ (
    .A1(reg_pmp_1_addr[9]),
    .A2(_01008_),
    .ZN(_01454_)
  );
  INV_X1 _13242_ (
    .A(_01454_),
    .ZN(_01455_)
  );
  AND2_X1 _13243_ (
    .A1(reg_pmp_2_addr[9]),
    .A2(_00953_),
    .ZN(_01456_)
  );
  INV_X1 _13244_ (
    .A(_01456_),
    .ZN(_01457_)
  );
  AND2_X1 _13245_ (
    .A1(_01455_),
    .A2(_01457_),
    .ZN(_01458_)
  );
  AND2_X1 _13246_ (
    .A1(_01453_),
    .A2(_01458_),
    .ZN(_01459_)
  );
  AND2_X1 _13247_ (
    .A1(reg_mtval[9]),
    .A2(_00926_),
    .ZN(_01460_)
  );
  INV_X1 _13248_ (
    .A(_01460_),
    .ZN(_01461_)
  );
  AND2_X1 _13249_ (
    .A1(reg_mcause[9]),
    .A2(_01001_),
    .ZN(_01462_)
  );
  INV_X1 _13250_ (
    .A(_01462_),
    .ZN(_01463_)
  );
  AND2_X1 _13251_ (
    .A1(_01461_),
    .A2(_01463_),
    .ZN(_01464_)
  );
  AND2_X1 _13252_ (
    .A1(reg_pmp_0_addr[9]),
    .A2(_01004_),
    .ZN(_01465_)
  );
  INV_X1 _13253_ (
    .A(_01465_),
    .ZN(_01466_)
  );
  AND2_X1 _13254_ (
    .A1(reg_pmp_5_addr[9]),
    .A2(_00948_),
    .ZN(_01467_)
  );
  INV_X1 _13255_ (
    .A(_01467_),
    .ZN(_01468_)
  );
  AND2_X1 _13256_ (
    .A1(_01466_),
    .A2(_01468_),
    .ZN(_01469_)
  );
  AND2_X1 _13257_ (
    .A1(_01464_),
    .A2(_01469_),
    .ZN(_01470_)
  );
  AND2_X1 _13258_ (
    .A1(reg_dscratch0[9]),
    .A2(_00958_),
    .ZN(_01471_)
  );
  INV_X1 _13259_ (
    .A(_01471_),
    .ZN(_01472_)
  );
  AND2_X1 _13260_ (
    .A1(reg_bp_0_address[9]),
    .A2(_00962_),
    .ZN(_01473_)
  );
  INV_X1 _13261_ (
    .A(_01473_),
    .ZN(_01474_)
  );
  AND2_X1 _13262_ (
    .A1(_01472_),
    .A2(_01474_),
    .ZN(_01475_)
  );
  AND2_X1 _13263_ (
    .A1(reg_dpc[9]),
    .A2(_00912_),
    .ZN(_01476_)
  );
  INV_X1 _13264_ (
    .A(_01476_),
    .ZN(_01477_)
  );
  AND2_X1 _13265_ (
    .A1(reg_pmp_4_addr[9]),
    .A2(_00968_),
    .ZN(_01478_)
  );
  INV_X1 _13266_ (
    .A(_01478_),
    .ZN(_01479_)
  );
  AND2_X1 _13267_ (
    .A1(_01477_),
    .A2(_01479_),
    .ZN(_01480_)
  );
  AND2_X1 _13268_ (
    .A1(_01475_),
    .A2(_01480_),
    .ZN(_01481_)
  );
  AND2_X1 _13269_ (
    .A1(_01470_),
    .A2(_01481_),
    .ZN(_01482_)
  );
  AND2_X1 _13270_ (
    .A1(_01459_),
    .A2(_01482_),
    .ZN(_01483_)
  );
  AND2_X1 _13271_ (
    .A1(reg_pmp_7_addr[9]),
    .A2(_01016_),
    .ZN(_01484_)
  );
  INV_X1 _13272_ (
    .A(_01484_),
    .ZN(_01485_)
  );
  AND2_X1 _13273_ (
    .A1(large_1[35]),
    .A2(_01019_),
    .ZN(_01486_)
  );
  INV_X1 _13274_ (
    .A(_01486_),
    .ZN(_01487_)
  );
  AND2_X1 _13275_ (
    .A1(_01485_),
    .A2(_01487_),
    .ZN(_01488_)
  );
  AND2_X1 _13276_ (
    .A1(reg_pmp_6_addr[9]),
    .A2(_00978_),
    .ZN(_01489_)
  );
  INV_X1 _13277_ (
    .A(_01489_),
    .ZN(_01490_)
  );
  AND2_X1 _13278_ (
    .A1(large_1[3]),
    .A2(_00995_),
    .ZN(_01491_)
  );
  INV_X1 _13279_ (
    .A(_01491_),
    .ZN(_01492_)
  );
  AND2_X1 _13280_ (
    .A1(_01490_),
    .A2(_01492_),
    .ZN(_01493_)
  );
  AND2_X1 _13281_ (
    .A1(_01488_),
    .A2(_01493_),
    .ZN(_01494_)
  );
  AND2_X1 _13282_ (
    .A1(reg_pmp_5_cfg_w),
    .A2(_00894_),
    .ZN(_01495_)
  );
  INV_X1 _13283_ (
    .A(_01495_),
    .ZN(_01496_)
  );
  AND2_X1 _13284_ (
    .A1(reg_mepc[9]),
    .A2(_00943_),
    .ZN(_01497_)
  );
  INV_X1 _13285_ (
    .A(_01497_),
    .ZN(_01498_)
  );
  AND2_X1 _13286_ (
    .A1(_01496_),
    .A2(_01498_),
    .ZN(_01499_)
  );
  AND2_X1 _13287_ (
    .A1(reg_pmp_1_cfg_w),
    .A2(_00916_),
    .ZN(_01500_)
  );
  INV_X1 _13288_ (
    .A(_01500_),
    .ZN(_01501_)
  );
  AND2_X1 _13289_ (
    .A1(reg_pmp_3_addr[9]),
    .A2(_01011_),
    .ZN(_01502_)
  );
  INV_X1 _13290_ (
    .A(_01502_),
    .ZN(_01503_)
  );
  AND2_X1 _13291_ (
    .A1(_01501_),
    .A2(_01503_),
    .ZN(_01504_)
  );
  AND2_X1 _13292_ (
    .A1(_01499_),
    .A2(_01504_),
    .ZN(_01505_)
  );
  AND2_X1 _13293_ (
    .A1(large_[35]),
    .A2(_00991_),
    .ZN(_01506_)
  );
  INV_X1 _13294_ (
    .A(_01506_),
    .ZN(_01507_)
  );
  AND2_X1 _13295_ (
    .A1(large_[3]),
    .A2(_00985_),
    .ZN(_01508_)
  );
  INV_X1 _13296_ (
    .A(_01508_),
    .ZN(_01509_)
  );
  AND2_X1 _13297_ (
    .A1(_01507_),
    .A2(_01509_),
    .ZN(_01510_)
  );
  AND2_X1 _13298_ (
    .A1(_01505_),
    .A2(_01510_),
    .ZN(_01511_)
  );
  AND2_X1 _13299_ (
    .A1(_01494_),
    .A2(_01511_),
    .ZN(_01512_)
  );
  AND2_X1 _13300_ (
    .A1(_01483_),
    .A2(_01512_),
    .ZN(_01513_)
  );
  INV_X1 _13301_ (
    .A(_01513_),
    .ZN(io_rw_rdata[9])
  );
  AND2_X1 _13302_ (
    .A1(io_rw_cmd[1]),
    .A2(_00845_),
    .ZN(_01514_)
  );
  AND2_X1 _13303_ (
    .A1(io_rw_rdata[9]),
    .A2(_01514_),
    .ZN(_01515_)
  );
  INV_X1 _13304_ (
    .A(_01515_),
    .ZN(_01516_)
  );
  AND2_X1 _13305_ (
    .A1(_01448_),
    .A2(_01516_),
    .ZN(_01517_)
  );
  INV_X1 _13306_ (
    .A(_01517_),
    .ZN(_01518_)
  );
  AND2_X1 _13307_ (
    .A1(_01446_),
    .A2(_01518_),
    .ZN(_01519_)
  );
  MUX2_X1 _13308_ (
    .A(reg_pmp_5_cfg_w),
    .B(_01519_),
    .S(_01364_),
    .Z(_00026_)
  );
  AND2_X1 _13309_ (
    .A1(reg_pmp_6_cfg_l),
    .A2(reg_pmp_6_cfg_a[0]),
    .ZN(_01520_)
  );
  AND2_X1 _13310_ (
    .A1(_00018_),
    .A2(_01520_),
    .ZN(_01521_)
  );
  INV_X1 _13311_ (
    .A(_01521_),
    .ZN(_01522_)
  );
  AND2_X1 _13312_ (
    .A1(_00805_),
    .A2(_01522_),
    .ZN(_01523_)
  );
  AND2_X1 _13313_ (
    .A1(_00897_),
    .A2(_01523_),
    .ZN(_01524_)
  );
  AND2_X1 _13314_ (
    .A1(_00948_),
    .A2(_01524_),
    .ZN(_01525_)
  );
  AND2_X1 _13315_ (
    .A1(io_rw_wdata[0]),
    .A2(_00903_),
    .ZN(_01526_)
  );
  INV_X1 _13316_ (
    .A(_01526_),
    .ZN(_01527_)
  );
  AND2_X1 _13317_ (
    .A1(reg_misa[0]),
    .A2(_01339_),
    .ZN(_01528_)
  );
  INV_X1 _13318_ (
    .A(_01528_),
    .ZN(_01529_)
  );
  AND2_X1 _13319_ (
    .A1(reg_pmp_5_addr[0]),
    .A2(_00948_),
    .ZN(_01530_)
  );
  INV_X1 _13320_ (
    .A(_01530_),
    .ZN(_01531_)
  );
  AND2_X1 _13321_ (
    .A1(reg_mscratch[0]),
    .A2(_00929_),
    .ZN(_01532_)
  );
  INV_X1 _13322_ (
    .A(_01532_),
    .ZN(_01533_)
  );
  AND2_X1 _13323_ (
    .A1(io_hartid),
    .A2(_00937_),
    .ZN(_01534_)
  );
  INV_X1 _13324_ (
    .A(_01534_),
    .ZN(_01535_)
  );
  AND2_X1 _13325_ (
    .A1(_00952_),
    .A2(_01535_),
    .ZN(_01536_)
  );
  INV_X1 _13326_ (
    .A(_01536_),
    .ZN(_01537_)
  );
  AND2_X1 _13327_ (
    .A1(reg_pmp_2_addr[0]),
    .A2(_00953_),
    .ZN(_01538_)
  );
  INV_X1 _13328_ (
    .A(_01538_),
    .ZN(_01539_)
  );
  AND2_X1 _13329_ (
    .A1(reg_pmp_3_addr[0]),
    .A2(_01011_),
    .ZN(_01540_)
  );
  INV_X1 _13330_ (
    .A(_01540_),
    .ZN(_01541_)
  );
  AND2_X1 _13331_ (
    .A1(reg_dscratch0[0]),
    .A2(_00958_),
    .ZN(_01542_)
  );
  INV_X1 _13332_ (
    .A(_01542_),
    .ZN(_01543_)
  );
  AND2_X1 _13333_ (
    .A1(reg_pmp_1_addr[0]),
    .A2(_01008_),
    .ZN(_01544_)
  );
  INV_X1 _13334_ (
    .A(_01544_),
    .ZN(_01545_)
  );
  AND2_X1 _13335_ (
    .A1(reg_mtvec[0]),
    .A2(_00940_),
    .ZN(_01546_)
  );
  INV_X1 _13336_ (
    .A(_01546_),
    .ZN(_01547_)
  );
  AND2_X1 _13337_ (
    .A1(reg_mcause[0]),
    .A2(_01001_),
    .ZN(_01548_)
  );
  INV_X1 _13338_ (
    .A(_01548_),
    .ZN(_01549_)
  );
  AND2_X1 _13339_ (
    .A1(_00890_),
    .A2(_00934_),
    .ZN(_01550_)
  );
  AND2_X1 _13340_ (
    .A1(_00883_),
    .A2(_01550_),
    .ZN(_01551_)
  );
  AND2_X1 _13341_ (
    .A1(_00888_),
    .A2(_01551_),
    .ZN(_01552_)
  );
  AND2_X1 _13342_ (
    .A1(reg_mcountinhibit[0]),
    .A2(_01552_),
    .ZN(_01553_)
  );
  INV_X1 _13343_ (
    .A(_01553_),
    .ZN(_01554_)
  );
  AND2_X1 _13344_ (
    .A1(_01549_),
    .A2(_01554_),
    .ZN(_01555_)
  );
  AND2_X1 _13345_ (
    .A1(reg_pmp_0_cfg_r),
    .A2(_00916_),
    .ZN(_01556_)
  );
  INV_X1 _13346_ (
    .A(_01556_),
    .ZN(_01557_)
  );
  AND2_X1 _13347_ (
    .A1(reg_pmp_4_cfg_r),
    .A2(_00894_),
    .ZN(_01558_)
  );
  INV_X1 _13348_ (
    .A(_01558_),
    .ZN(_01559_)
  );
  AND2_X1 _13349_ (
    .A1(_01557_),
    .A2(_01559_),
    .ZN(_01560_)
  );
  AND2_X1 _13350_ (
    .A1(reg_mtval[0]),
    .A2(_00926_),
    .ZN(_01561_)
  );
  INV_X1 _13351_ (
    .A(_01561_),
    .ZN(_01562_)
  );
  AND2_X1 _13352_ (
    .A1(reg_pmp_4_addr[0]),
    .A2(_00968_),
    .ZN(_01563_)
  );
  INV_X1 _13353_ (
    .A(_01563_),
    .ZN(_01564_)
  );
  AND2_X1 _13354_ (
    .A1(reg_pmp_7_addr[0]),
    .A2(_01016_),
    .ZN(_01565_)
  );
  INV_X1 _13355_ (
    .A(_01565_),
    .ZN(_01566_)
  );
  AND2_X1 _13356_ (
    .A1(reg_pmp_6_addr[0]),
    .A2(_00978_),
    .ZN(_01567_)
  );
  INV_X1 _13357_ (
    .A(_01567_),
    .ZN(_01568_)
  );
  AND2_X1 _13358_ (
    .A1(reg_bp_0_address[0]),
    .A2(_00962_),
    .ZN(_01569_)
  );
  INV_X1 _13359_ (
    .A(_01569_),
    .ZN(_01570_)
  );
  AND2_X1 _13360_ (
    .A1(reg_pmp_0_addr[0]),
    .A2(_01004_),
    .ZN(_01571_)
  );
  INV_X1 _13361_ (
    .A(_01571_),
    .ZN(_01572_)
  );
  AND2_X1 _13362_ (
    .A1(reg_bp_0_control_r),
    .A2(_01341_),
    .ZN(_01573_)
  );
  INV_X1 _13363_ (
    .A(_01573_),
    .ZN(_01574_)
  );
  AND2_X1 _13364_ (
    .A1(large_[26]),
    .A2(_00991_),
    .ZN(_01575_)
  );
  INV_X1 _13365_ (
    .A(_01575_),
    .ZN(_01576_)
  );
  AND2_X1 _13366_ (
    .A1(large_1[26]),
    .A2(_01019_),
    .ZN(_01577_)
  );
  INV_X1 _13367_ (
    .A(_01577_),
    .ZN(_01578_)
  );
  AND2_X1 _13368_ (
    .A1(_01529_),
    .A2(_01543_),
    .ZN(_01579_)
  );
  AND2_X1 _13369_ (
    .A1(_01382_),
    .A2(_01579_),
    .ZN(_01580_)
  );
  AND2_X1 _13370_ (
    .A1(_01539_),
    .A2(_01545_),
    .ZN(_01581_)
  );
  AND2_X1 _13371_ (
    .A1(_01578_),
    .A2(_01581_),
    .ZN(_01582_)
  );
  AND2_X1 _13372_ (
    .A1(small_[0]),
    .A2(_01027_),
    .ZN(_01583_)
  );
  INV_X1 _13373_ (
    .A(_01583_),
    .ZN(_01584_)
  );
  AND2_X1 _13374_ (
    .A1(_01572_),
    .A2(_01584_),
    .ZN(_01585_)
  );
  AND2_X1 _13375_ (
    .A1(_01582_),
    .A2(_01585_),
    .ZN(_01586_)
  );
  AND2_X1 _13376_ (
    .A1(_01541_),
    .A2(_01564_),
    .ZN(_01587_)
  );
  AND2_X1 _13377_ (
    .A1(_01531_),
    .A2(_01587_),
    .ZN(_01588_)
  );
  AND2_X1 _13378_ (
    .A1(small_1[0]),
    .A2(_01029_),
    .ZN(_01589_)
  );
  INV_X1 _13379_ (
    .A(_01589_),
    .ZN(_01590_)
  );
  AND2_X1 _13380_ (
    .A1(_01547_),
    .A2(_01590_),
    .ZN(_01591_)
  );
  AND2_X1 _13381_ (
    .A1(_01533_),
    .A2(_01591_),
    .ZN(_01592_)
  );
  AND2_X1 _13382_ (
    .A1(_01588_),
    .A2(_01592_),
    .ZN(_01593_)
  );
  AND2_X1 _13383_ (
    .A1(_01586_),
    .A2(_01593_),
    .ZN(_01594_)
  );
  AND2_X1 _13384_ (
    .A1(_01560_),
    .A2(_01566_),
    .ZN(_01595_)
  );
  AND2_X1 _13385_ (
    .A1(_01568_),
    .A2(_01595_),
    .ZN(_01596_)
  );
  AND2_X1 _13386_ (
    .A1(_01197_),
    .A2(_01537_),
    .ZN(_01597_)
  );
  INV_X1 _13387_ (
    .A(_01597_),
    .ZN(_01598_)
  );
  AND2_X1 _13388_ (
    .A1(_01570_),
    .A2(_01574_),
    .ZN(_01599_)
  );
  AND2_X1 _13389_ (
    .A1(_01598_),
    .A2(_01599_),
    .ZN(_01600_)
  );
  AND2_X1 _13390_ (
    .A1(_01555_),
    .A2(_01562_),
    .ZN(_01601_)
  );
  AND2_X1 _13391_ (
    .A1(_01576_),
    .A2(_01601_),
    .ZN(_01602_)
  );
  AND2_X1 _13392_ (
    .A1(_01600_),
    .A2(_01602_),
    .ZN(_01603_)
  );
  AND2_X1 _13393_ (
    .A1(_01596_),
    .A2(_01603_),
    .ZN(_01604_)
  );
  AND2_X1 _13394_ (
    .A1(_01594_),
    .A2(_01604_),
    .ZN(_01605_)
  );
  AND2_X1 _13395_ (
    .A1(_00883_),
    .A2(_00892_),
    .ZN(_01606_)
  );
  AND2_X1 _13396_ (
    .A1(_00934_),
    .A2(_01606_),
    .ZN(_01607_)
  );
  AND2_X1 _13397_ (
    .A1(_01580_),
    .A2(_01605_),
    .ZN(_01608_)
  );
  INV_X1 _13398_ (
    .A(_01608_),
    .ZN(io_rw_rdata[0])
  );
  AND2_X1 _13399_ (
    .A1(io_rw_cmd[1]),
    .A2(_00836_),
    .ZN(_01609_)
  );
  AND2_X1 _13400_ (
    .A1(io_rw_rdata[0]),
    .A2(_01609_),
    .ZN(_01610_)
  );
  INV_X1 _13401_ (
    .A(_01610_),
    .ZN(_01611_)
  );
  AND2_X1 _13402_ (
    .A1(_01527_),
    .A2(_01611_),
    .ZN(_01612_)
  );
  INV_X1 _13403_ (
    .A(_01612_),
    .ZN(_01613_)
  );
  MUX2_X1 _13404_ (
    .A(reg_pmp_5_addr[0]),
    .B(_01613_),
    .S(_01525_),
    .Z(_00027_)
  );
  AND2_X1 _13405_ (
    .A1(io_rw_wdata[1]),
    .A2(_00903_),
    .ZN(_01614_)
  );
  INV_X1 _13406_ (
    .A(_01614_),
    .ZN(_01615_)
  );
  AND2_X1 _13407_ (
    .A1(io_rw_cmd[1]),
    .A2(_00837_),
    .ZN(_01616_)
  );
  AND2_X1 _13408_ (
    .A1(reg_pmp_1_addr[1]),
    .A2(_01008_),
    .ZN(_01617_)
  );
  INV_X1 _13409_ (
    .A(_01617_),
    .ZN(_01618_)
  );
  AND2_X1 _13410_ (
    .A1(reg_pmp_4_addr[1]),
    .A2(_00968_),
    .ZN(_01619_)
  );
  INV_X1 _13411_ (
    .A(_01619_),
    .ZN(_01620_)
  );
  AND2_X1 _13412_ (
    .A1(_01618_),
    .A2(_01620_),
    .ZN(_01621_)
  );
  AND2_X1 _13413_ (
    .A1(reg_pmp_0_addr[1]),
    .A2(_01004_),
    .ZN(_01622_)
  );
  INV_X1 _13414_ (
    .A(_01622_),
    .ZN(_01623_)
  );
  AND2_X1 _13415_ (
    .A1(reg_bp_0_address[1]),
    .A2(_00962_),
    .ZN(_01624_)
  );
  INV_X1 _13416_ (
    .A(_01624_),
    .ZN(_01625_)
  );
  AND2_X1 _13417_ (
    .A1(_01623_),
    .A2(_01625_),
    .ZN(_01626_)
  );
  AND2_X1 _13418_ (
    .A1(_01621_),
    .A2(_01626_),
    .ZN(_01627_)
  );
  AND2_X1 _13419_ (
    .A1(reg_dscratch0[1]),
    .A2(_00958_),
    .ZN(_01628_)
  );
  INV_X1 _13420_ (
    .A(_01628_),
    .ZN(_01629_)
  );
  AND2_X1 _13421_ (
    .A1(_00875_),
    .A2(_00876_),
    .ZN(_01630_)
  );
  AND2_X1 _13422_ (
    .A1(_00912_),
    .A2(_01630_),
    .ZN(_01631_)
  );
  INV_X1 _13423_ (
    .A(_01631_),
    .ZN(_01632_)
  );
  AND2_X1 _13424_ (
    .A1(_01629_),
    .A2(_01632_),
    .ZN(_01633_)
  );
  AND2_X1 _13425_ (
    .A1(reg_pmp_2_addr[1]),
    .A2(_00953_),
    .ZN(_01634_)
  );
  INV_X1 _13426_ (
    .A(_01634_),
    .ZN(_01635_)
  );
  AND2_X1 _13427_ (
    .A1(reg_bp_0_control_w),
    .A2(_01341_),
    .ZN(_01636_)
  );
  INV_X1 _13428_ (
    .A(_01636_),
    .ZN(_01637_)
  );
  AND2_X1 _13429_ (
    .A1(_01635_),
    .A2(_01637_),
    .ZN(_01638_)
  );
  AND2_X1 _13430_ (
    .A1(_01633_),
    .A2(_01638_),
    .ZN(_01639_)
  );
  AND2_X1 _13431_ (
    .A1(_01627_),
    .A2(_01639_),
    .ZN(_01640_)
  );
  AND2_X1 _13432_ (
    .A1(_00874_),
    .A2(_00875_),
    .ZN(_01641_)
  );
  AND2_X1 _13433_ (
    .A1(_00943_),
    .A2(_01641_),
    .ZN(_01642_)
  );
  INV_X1 _13434_ (
    .A(_01642_),
    .ZN(_01643_)
  );
  AND2_X1 _13435_ (
    .A1(reg_mcause[1]),
    .A2(_01001_),
    .ZN(_01644_)
  );
  INV_X1 _13436_ (
    .A(_01644_),
    .ZN(_01645_)
  );
  AND2_X1 _13437_ (
    .A1(reg_mscratch[1]),
    .A2(_00929_),
    .ZN(_01646_)
  );
  INV_X1 _13438_ (
    .A(_01646_),
    .ZN(_01647_)
  );
  AND2_X1 _13439_ (
    .A1(_01645_),
    .A2(_01647_),
    .ZN(_01648_)
  );
  AND2_X1 _13440_ (
    .A1(_01643_),
    .A2(_01648_),
    .ZN(_01649_)
  );
  AND2_X1 _13441_ (
    .A1(reg_pmp_5_addr[1]),
    .A2(_00948_),
    .ZN(_01650_)
  );
  INV_X1 _13442_ (
    .A(_01650_),
    .ZN(_01651_)
  );
  AND2_X1 _13443_ (
    .A1(reg_pmp_4_cfg_w),
    .A2(_00894_),
    .ZN(_01652_)
  );
  INV_X1 _13444_ (
    .A(_01652_),
    .ZN(_01653_)
  );
  AND2_X1 _13445_ (
    .A1(_01651_),
    .A2(_01653_),
    .ZN(_01654_)
  );
  AND2_X1 _13446_ (
    .A1(reg_mtval[1]),
    .A2(_00926_),
    .ZN(_01655_)
  );
  INV_X1 _13447_ (
    .A(_01655_),
    .ZN(_01656_)
  );
  AND2_X1 _13448_ (
    .A1(reg_pmp_3_addr[1]),
    .A2(_01011_),
    .ZN(_01657_)
  );
  INV_X1 _13449_ (
    .A(_01657_),
    .ZN(_01658_)
  );
  AND2_X1 _13450_ (
    .A1(_01656_),
    .A2(_01658_),
    .ZN(_01659_)
  );
  AND2_X1 _13451_ (
    .A1(_01654_),
    .A2(_01659_),
    .ZN(_01660_)
  );
  AND2_X1 _13452_ (
    .A1(_01649_),
    .A2(_01660_),
    .ZN(_01661_)
  );
  AND2_X1 _13453_ (
    .A1(_01640_),
    .A2(_01661_),
    .ZN(_01662_)
  );
  AND2_X1 _13454_ (
    .A1(large_1[27]),
    .A2(_01019_),
    .ZN(_01663_)
  );
  INV_X1 _13455_ (
    .A(_01663_),
    .ZN(_01664_)
  );
  AND2_X1 _13456_ (
    .A1(small_1[1]),
    .A2(_00995_),
    .ZN(_01665_)
  );
  INV_X1 _13457_ (
    .A(_01665_),
    .ZN(_01666_)
  );
  AND2_X1 _13458_ (
    .A1(small_[1]),
    .A2(_00985_),
    .ZN(_01667_)
  );
  INV_X1 _13459_ (
    .A(_01667_),
    .ZN(_01668_)
  );
  AND2_X1 _13460_ (
    .A1(_01666_),
    .A2(_01668_),
    .ZN(_01669_)
  );
  AND2_X1 _13461_ (
    .A1(_01664_),
    .A2(_01669_),
    .ZN(_01670_)
  );
  AND2_X1 _13462_ (
    .A1(reg_pmp_6_addr[1]),
    .A2(_00978_),
    .ZN(_01671_)
  );
  INV_X1 _13463_ (
    .A(_01671_),
    .ZN(_01672_)
  );
  AND2_X1 _13464_ (
    .A1(reg_pmp_0_cfg_w),
    .A2(_00916_),
    .ZN(_01673_)
  );
  INV_X1 _13465_ (
    .A(_01673_),
    .ZN(_01674_)
  );
  AND2_X1 _13466_ (
    .A1(_01382_),
    .A2(_01674_),
    .ZN(_01675_)
  );
  AND2_X1 _13467_ (
    .A1(_01672_),
    .A2(_01675_),
    .ZN(_01676_)
  );
  AND2_X1 _13468_ (
    .A1(large_[27]),
    .A2(_00991_),
    .ZN(_01677_)
  );
  INV_X1 _13469_ (
    .A(_01677_),
    .ZN(_01678_)
  );
  AND2_X1 _13470_ (
    .A1(reg_pmp_7_addr[1]),
    .A2(_01016_),
    .ZN(_01679_)
  );
  INV_X1 _13471_ (
    .A(_01679_),
    .ZN(_01680_)
  );
  AND2_X1 _13472_ (
    .A1(_01678_),
    .A2(_01680_),
    .ZN(_01681_)
  );
  AND2_X1 _13473_ (
    .A1(_01676_),
    .A2(_01681_),
    .ZN(_01682_)
  );
  AND2_X1 _13474_ (
    .A1(_01670_),
    .A2(_01682_),
    .ZN(_01683_)
  );
  AND2_X1 _13475_ (
    .A1(_01662_),
    .A2(_01683_),
    .ZN(_01684_)
  );
  INV_X1 _13476_ (
    .A(_01684_),
    .ZN(io_rw_rdata[1])
  );
  AND2_X1 _13477_ (
    .A1(_01616_),
    .A2(io_rw_rdata[1]),
    .ZN(_01685_)
  );
  INV_X1 _13478_ (
    .A(_01685_),
    .ZN(_01686_)
  );
  AND2_X1 _13479_ (
    .A1(_01615_),
    .A2(_01686_),
    .ZN(_01687_)
  );
  INV_X1 _13480_ (
    .A(_01687_),
    .ZN(_01688_)
  );
  MUX2_X1 _13481_ (
    .A(reg_pmp_5_addr[1]),
    .B(_01688_),
    .S(_01525_),
    .Z(_00028_)
  );
  AND2_X1 _13482_ (
    .A1(io_rw_wdata[2]),
    .A2(_00903_),
    .ZN(_01689_)
  );
  INV_X1 _13483_ (
    .A(_01689_),
    .ZN(_01690_)
  );
  AND2_X1 _13484_ (
    .A1(reg_mepc[2]),
    .A2(_00943_),
    .ZN(_01691_)
  );
  INV_X1 _13485_ (
    .A(_01691_),
    .ZN(_01692_)
  );
  AND2_X1 _13486_ (
    .A1(reg_mscratch[2]),
    .A2(_00929_),
    .ZN(_01693_)
  );
  INV_X1 _13487_ (
    .A(_01693_),
    .ZN(_01694_)
  );
  AND2_X1 _13488_ (
    .A1(reg_dscratch0[2]),
    .A2(_00958_),
    .ZN(_01695_)
  );
  INV_X1 _13489_ (
    .A(_01695_),
    .ZN(_01696_)
  );
  AND2_X1 _13490_ (
    .A1(_01694_),
    .A2(_01696_),
    .ZN(_01697_)
  );
  AND2_X1 _13491_ (
    .A1(_01692_),
    .A2(_01697_),
    .ZN(_01698_)
  );
  AND2_X1 _13492_ (
    .A1(reg_pmp_0_addr[2]),
    .A2(_01004_),
    .ZN(_01699_)
  );
  INV_X1 _13493_ (
    .A(_01699_),
    .ZN(_01700_)
  );
  AND2_X1 _13494_ (
    .A1(reg_mcause[2]),
    .A2(_01001_),
    .ZN(_01701_)
  );
  INV_X1 _13495_ (
    .A(_01701_),
    .ZN(_01702_)
  );
  AND2_X1 _13496_ (
    .A1(_01700_),
    .A2(_01702_),
    .ZN(_01703_)
  );
  AND2_X1 _13497_ (
    .A1(reg_misa[2]),
    .A2(_01339_),
    .ZN(_01704_)
  );
  INV_X1 _13498_ (
    .A(_01704_),
    .ZN(_01705_)
  );
  AND2_X1 _13499_ (
    .A1(reg_mcountinhibit[2]),
    .A2(_01552_),
    .ZN(_01706_)
  );
  INV_X1 _13500_ (
    .A(_01706_),
    .ZN(_01707_)
  );
  AND2_X1 _13501_ (
    .A1(_01705_),
    .A2(_01707_),
    .ZN(_01708_)
  );
  AND2_X1 _13502_ (
    .A1(_01703_),
    .A2(_01708_),
    .ZN(_01709_)
  );
  AND2_X1 _13503_ (
    .A1(reg_bp_0_address[2]),
    .A2(_00962_),
    .ZN(_01710_)
  );
  INV_X1 _13504_ (
    .A(_01710_),
    .ZN(_01711_)
  );
  AND2_X1 _13505_ (
    .A1(reg_dcsr_step),
    .A2(_01381_),
    .ZN(_01712_)
  );
  INV_X1 _13506_ (
    .A(_01712_),
    .ZN(_01713_)
  );
  AND2_X1 _13507_ (
    .A1(_01711_),
    .A2(_01713_),
    .ZN(_01714_)
  );
  AND2_X1 _13508_ (
    .A1(reg_bp_0_control_x),
    .A2(_01341_),
    .ZN(_01715_)
  );
  INV_X1 _13509_ (
    .A(_01715_),
    .ZN(_01716_)
  );
  AND2_X1 _13510_ (
    .A1(reg_mtvec[2]),
    .A2(_read_mtvec_T_4[6]),
    .ZN(_01717_)
  );
  AND2_X1 _13511_ (
    .A1(_00940_),
    .A2(_01717_),
    .ZN(_01718_)
  );
  INV_X1 _13512_ (
    .A(_01718_),
    .ZN(_01719_)
  );
  AND2_X1 _13513_ (
    .A1(_01716_),
    .A2(_01719_),
    .ZN(_01720_)
  );
  AND2_X1 _13514_ (
    .A1(_01714_),
    .A2(_01720_),
    .ZN(_01721_)
  );
  AND2_X1 _13515_ (
    .A1(_01709_),
    .A2(_01721_),
    .ZN(_01722_)
  );
  AND2_X1 _13516_ (
    .A1(_01698_),
    .A2(_01722_),
    .ZN(_01723_)
  );
  AND2_X1 _13517_ (
    .A1(reg_pmp_6_addr[2]),
    .A2(_00978_),
    .ZN(_01724_)
  );
  INV_X1 _13518_ (
    .A(_01724_),
    .ZN(_01725_)
  );
  AND2_X1 _13519_ (
    .A1(reg_pmp_7_addr[2]),
    .A2(_01016_),
    .ZN(_01726_)
  );
  INV_X1 _13520_ (
    .A(_01726_),
    .ZN(_01727_)
  );
  AND2_X1 _13521_ (
    .A1(small_1[2]),
    .A2(_00995_),
    .ZN(_01728_)
  );
  INV_X1 _13522_ (
    .A(_01728_),
    .ZN(_01729_)
  );
  AND2_X1 _13523_ (
    .A1(_01727_),
    .A2(_01729_),
    .ZN(_01730_)
  );
  AND2_X1 _13524_ (
    .A1(_01725_),
    .A2(_01730_),
    .ZN(_01731_)
  );
  AND2_X1 _13525_ (
    .A1(small_[2]),
    .A2(_00985_),
    .ZN(_01732_)
  );
  INV_X1 _13526_ (
    .A(_01732_),
    .ZN(_01733_)
  );
  AND2_X1 _13527_ (
    .A1(reg_pmp_5_addr[2]),
    .A2(_00948_),
    .ZN(_01734_)
  );
  INV_X1 _13528_ (
    .A(_01734_),
    .ZN(_01735_)
  );
  AND2_X1 _13529_ (
    .A1(_01132_),
    .A2(_01735_),
    .ZN(_01736_)
  );
  AND2_X1 _13530_ (
    .A1(_01733_),
    .A2(_01736_),
    .ZN(_01737_)
  );
  AND2_X1 _13531_ (
    .A1(large_[28]),
    .A2(_00991_),
    .ZN(_01738_)
  );
  INV_X1 _13532_ (
    .A(_01738_),
    .ZN(_01739_)
  );
  AND2_X1 _13533_ (
    .A1(large_1[28]),
    .A2(_01019_),
    .ZN(_01740_)
  );
  INV_X1 _13534_ (
    .A(_01740_),
    .ZN(_01741_)
  );
  AND2_X1 _13535_ (
    .A1(_01739_),
    .A2(_01741_),
    .ZN(_01742_)
  );
  AND2_X1 _13536_ (
    .A1(_01737_),
    .A2(_01742_),
    .ZN(_01743_)
  );
  AND2_X1 _13537_ (
    .A1(reg_pmp_3_addr[2]),
    .A2(_01011_),
    .ZN(_01744_)
  );
  INV_X1 _13538_ (
    .A(_01744_),
    .ZN(_01745_)
  );
  AND2_X1 _13539_ (
    .A1(reg_pmp_4_addr[2]),
    .A2(_00968_),
    .ZN(_01746_)
  );
  INV_X1 _13540_ (
    .A(_01746_),
    .ZN(_01747_)
  );
  AND2_X1 _13541_ (
    .A1(_01745_),
    .A2(_01747_),
    .ZN(_01748_)
  );
  AND2_X1 _13542_ (
    .A1(reg_pmp_1_addr[2]),
    .A2(_01008_),
    .ZN(_01749_)
  );
  INV_X1 _13543_ (
    .A(_01749_),
    .ZN(_01750_)
  );
  AND2_X1 _13544_ (
    .A1(reg_mtval[2]),
    .A2(_00926_),
    .ZN(_01751_)
  );
  INV_X1 _13545_ (
    .A(_01751_),
    .ZN(_01752_)
  );
  AND2_X1 _13546_ (
    .A1(_01750_),
    .A2(_01752_),
    .ZN(_01753_)
  );
  AND2_X1 _13547_ (
    .A1(_01748_),
    .A2(_01753_),
    .ZN(_01754_)
  );
  AND2_X1 _13548_ (
    .A1(reg_pmp_4_cfg_x),
    .A2(_00894_),
    .ZN(_01755_)
  );
  INV_X1 _13549_ (
    .A(_01755_),
    .ZN(_01756_)
  );
  AND2_X1 _13550_ (
    .A1(reg_pmp_0_cfg_x),
    .A2(_00916_),
    .ZN(_01757_)
  );
  INV_X1 _13551_ (
    .A(_01757_),
    .ZN(_01758_)
  );
  AND2_X1 _13552_ (
    .A1(_01756_),
    .A2(_01758_),
    .ZN(_01759_)
  );
  AND2_X1 _13553_ (
    .A1(reg_pmp_2_addr[2]),
    .A2(_00953_),
    .ZN(_01760_)
  );
  INV_X1 _13554_ (
    .A(_01760_),
    .ZN(_01761_)
  );
  AND2_X1 _13555_ (
    .A1(reg_dpc[2]),
    .A2(_00912_),
    .ZN(_01762_)
  );
  INV_X1 _13556_ (
    .A(_01762_),
    .ZN(_01763_)
  );
  AND2_X1 _13557_ (
    .A1(_01761_),
    .A2(_01763_),
    .ZN(_01764_)
  );
  AND2_X1 _13558_ (
    .A1(_01759_),
    .A2(_01764_),
    .ZN(_01765_)
  );
  AND2_X1 _13559_ (
    .A1(_01754_),
    .A2(_01765_),
    .ZN(_01766_)
  );
  AND2_X1 _13560_ (
    .A1(_01743_),
    .A2(_01766_),
    .ZN(_01767_)
  );
  AND2_X1 _13561_ (
    .A1(_01731_),
    .A2(_01767_),
    .ZN(_01768_)
  );
  AND2_X1 _13562_ (
    .A1(_01723_),
    .A2(_01768_),
    .ZN(_01769_)
  );
  INV_X1 _13563_ (
    .A(_01769_),
    .ZN(io_rw_rdata[2])
  );
  AND2_X1 _13564_ (
    .A1(io_rw_cmd[1]),
    .A2(_00838_),
    .ZN(_01770_)
  );
  AND2_X1 _13565_ (
    .A1(io_rw_rdata[2]),
    .A2(_01770_),
    .ZN(_01771_)
  );
  INV_X1 _13566_ (
    .A(_01771_),
    .ZN(_01772_)
  );
  AND2_X1 _13567_ (
    .A1(_01690_),
    .A2(_01772_),
    .ZN(_01773_)
  );
  INV_X1 _13568_ (
    .A(_01773_),
    .ZN(_01774_)
  );
  MUX2_X1 _13569_ (
    .A(reg_pmp_5_addr[2]),
    .B(_01774_),
    .S(_01525_),
    .Z(_00029_)
  );
  AND2_X1 _13570_ (
    .A1(io_rw_wdata[3]),
    .A2(_00903_),
    .ZN(_01775_)
  );
  INV_X1 _13571_ (
    .A(_01775_),
    .ZN(_01776_)
  );
  AND2_X1 _13572_ (
    .A1(reg_pmp_4_cfg_a[0]),
    .A2(_00894_),
    .ZN(_01777_)
  );
  INV_X1 _13573_ (
    .A(_01777_),
    .ZN(_01778_)
  );
  AND2_X1 _13574_ (
    .A1(reg_pmp_2_addr[3]),
    .A2(_00953_),
    .ZN(_01779_)
  );
  INV_X1 _13575_ (
    .A(_01779_),
    .ZN(_01780_)
  );
  AND2_X1 _13576_ (
    .A1(_01778_),
    .A2(_01780_),
    .ZN(_01781_)
  );
  AND2_X1 _13577_ (
    .A1(_00936_),
    .A2(_00967_),
    .ZN(_01782_)
  );
  AND2_X1 _13578_ (
    .A1(reg_mie[3]),
    .A2(_01782_),
    .ZN(_01783_)
  );
  INV_X1 _13579_ (
    .A(_01783_),
    .ZN(_01784_)
  );
  AND2_X1 _13580_ (
    .A1(reg_pmp_0_addr[3]),
    .A2(_01004_),
    .ZN(_01785_)
  );
  INV_X1 _13581_ (
    .A(_01785_),
    .ZN(_01786_)
  );
  AND2_X1 _13582_ (
    .A1(_01784_),
    .A2(_01786_),
    .ZN(_01787_)
  );
  AND2_X1 _13583_ (
    .A1(_01781_),
    .A2(_01787_),
    .ZN(_01788_)
  );
  AND2_X1 _13584_ (
    .A1(reg_pmp_4_addr[3]),
    .A2(_00968_),
    .ZN(_01789_)
  );
  INV_X1 _13585_ (
    .A(_01789_),
    .ZN(_01790_)
  );
  AND2_X1 _13586_ (
    .A1(reg_dscratch0[3]),
    .A2(_00958_),
    .ZN(_01791_)
  );
  INV_X1 _13587_ (
    .A(_01791_),
    .ZN(_01792_)
  );
  AND2_X1 _13588_ (
    .A1(_01790_),
    .A2(_01792_),
    .ZN(_01793_)
  );
  AND2_X1 _13589_ (
    .A1(reg_bp_0_address[3]),
    .A2(_00962_),
    .ZN(_01794_)
  );
  INV_X1 _13590_ (
    .A(_01794_),
    .ZN(_01795_)
  );
  AND2_X1 _13591_ (
    .A1(reg_pmp_0_cfg_a[0]),
    .A2(_00916_),
    .ZN(_01796_)
  );
  INV_X1 _13592_ (
    .A(_01796_),
    .ZN(_01797_)
  );
  AND2_X1 _13593_ (
    .A1(_01795_),
    .A2(_01797_),
    .ZN(_01798_)
  );
  AND2_X1 _13594_ (
    .A1(_01793_),
    .A2(_01798_),
    .ZN(_01799_)
  );
  AND2_X1 _13595_ (
    .A1(_01788_),
    .A2(_01799_),
    .ZN(_01800_)
  );
  AND2_X1 _13596_ (
    .A1(reg_mepc[3]),
    .A2(_00943_),
    .ZN(_01801_)
  );
  INV_X1 _13597_ (
    .A(_01801_),
    .ZN(_01802_)
  );
  AND2_X1 _13598_ (
    .A1(_00923_),
    .A2(_00937_),
    .ZN(_01803_)
  );
  AND2_X1 _13599_ (
    .A1(io_interrupts_msip),
    .A2(_01803_),
    .ZN(_01804_)
  );
  INV_X1 _13600_ (
    .A(_01804_),
    .ZN(_01805_)
  );
  AND2_X1 _13601_ (
    .A1(_01802_),
    .A2(_01805_),
    .ZN(_01806_)
  );
  AND2_X1 _13602_ (
    .A1(reg_mscratch[3]),
    .A2(_00929_),
    .ZN(_01807_)
  );
  INV_X1 _13603_ (
    .A(_01807_),
    .ZN(_01808_)
  );
  AND2_X1 _13604_ (
    .A1(reg_mtval[3]),
    .A2(_00926_),
    .ZN(_01809_)
  );
  INV_X1 _13605_ (
    .A(_01809_),
    .ZN(_01810_)
  );
  AND2_X1 _13606_ (
    .A1(_01808_),
    .A2(_01810_),
    .ZN(_01811_)
  );
  AND2_X1 _13607_ (
    .A1(_01806_),
    .A2(_01811_),
    .ZN(_01812_)
  );
  AND2_X1 _13608_ (
    .A1(_00915_),
    .A2(_00936_),
    .ZN(_01813_)
  );
  INV_X1 _13609_ (
    .A(_01813_),
    .ZN(_01814_)
  );
  AND2_X1 _13610_ (
    .A1(reg_mstatus_mie),
    .A2(_01813_),
    .ZN(_01815_)
  );
  INV_X1 _13611_ (
    .A(_01815_),
    .ZN(_01816_)
  );
  AND2_X1 _13612_ (
    .A1(reg_pmp_3_addr[3]),
    .A2(_01011_),
    .ZN(_01817_)
  );
  INV_X1 _13613_ (
    .A(_01817_),
    .ZN(_01818_)
  );
  AND2_X1 _13614_ (
    .A1(_01816_),
    .A2(_01818_),
    .ZN(_01819_)
  );
  AND2_X1 _13615_ (
    .A1(reg_pmp_5_addr[3]),
    .A2(_00948_),
    .ZN(_01820_)
  );
  INV_X1 _13616_ (
    .A(_01820_),
    .ZN(_01821_)
  );
  AND2_X1 _13617_ (
    .A1(reg_mcause[3]),
    .A2(_01001_),
    .ZN(_01822_)
  );
  INV_X1 _13618_ (
    .A(_01822_),
    .ZN(_01823_)
  );
  AND2_X1 _13619_ (
    .A1(_01821_),
    .A2(_01823_),
    .ZN(_01824_)
  );
  AND2_X1 _13620_ (
    .A1(_01819_),
    .A2(_01824_),
    .ZN(_01825_)
  );
  AND2_X1 _13621_ (
    .A1(_01812_),
    .A2(_01825_),
    .ZN(_01826_)
  );
  AND2_X1 _13622_ (
    .A1(_01800_),
    .A2(_01826_),
    .ZN(_01827_)
  );
  AND2_X1 _13623_ (
    .A1(reg_pmp_7_addr[3]),
    .A2(_01016_),
    .ZN(_01828_)
  );
  INV_X1 _13624_ (
    .A(_01828_),
    .ZN(_01829_)
  );
  AND2_X1 _13625_ (
    .A1(reg_pmp_6_addr[3]),
    .A2(_00978_),
    .ZN(_01830_)
  );
  INV_X1 _13626_ (
    .A(_01830_),
    .ZN(_01831_)
  );
  AND2_X1 _13627_ (
    .A1(_01829_),
    .A2(_01831_),
    .ZN(_01832_)
  );
  AND2_X1 _13628_ (
    .A1(large_1[29]),
    .A2(_01019_),
    .ZN(_01833_)
  );
  INV_X1 _13629_ (
    .A(_01833_),
    .ZN(_01834_)
  );
  AND2_X1 _13630_ (
    .A1(small_1[3]),
    .A2(_00995_),
    .ZN(_01835_)
  );
  INV_X1 _13631_ (
    .A(_01835_),
    .ZN(_01836_)
  );
  AND2_X1 _13632_ (
    .A1(_01834_),
    .A2(_01836_),
    .ZN(_01837_)
  );
  AND2_X1 _13633_ (
    .A1(_01832_),
    .A2(_01837_),
    .ZN(_01838_)
  );
  AND2_X1 _13634_ (
    .A1(reg_pmp_1_addr[3]),
    .A2(_01008_),
    .ZN(_01839_)
  );
  INV_X1 _13635_ (
    .A(_01839_),
    .ZN(_01840_)
  );
  AND2_X1 _13636_ (
    .A1(io_rw_addr[6]),
    .A2(io_rw_addr[7]),
    .ZN(_01841_)
  );
  AND2_X1 _13637_ (
    .A1(_00910_),
    .A2(_01841_),
    .ZN(_01842_)
  );
  AND2_X1 _13638_ (
    .A1(reg_custom_0[3]),
    .A2(_01842_),
    .ZN(_01843_)
  );
  INV_X1 _13639_ (
    .A(_01843_),
    .ZN(_01844_)
  );
  AND2_X1 _13640_ (
    .A1(_01840_),
    .A2(_01844_),
    .ZN(_01845_)
  );
  AND2_X1 _13641_ (
    .A1(reg_mtvec[3]),
    .A2(_read_mtvec_T_4[6]),
    .ZN(_01846_)
  );
  AND2_X1 _13642_ (
    .A1(_00940_),
    .A2(_01846_),
    .ZN(_01847_)
  );
  INV_X1 _13643_ (
    .A(_01847_),
    .ZN(_01848_)
  );
  AND2_X1 _13644_ (
    .A1(reg_dpc[3]),
    .A2(_00912_),
    .ZN(_01849_)
  );
  INV_X1 _13645_ (
    .A(_01849_),
    .ZN(_01850_)
  );
  AND2_X1 _13646_ (
    .A1(_01848_),
    .A2(_01850_),
    .ZN(_01851_)
  );
  AND2_X1 _13647_ (
    .A1(_01845_),
    .A2(_01851_),
    .ZN(_01852_)
  );
  AND2_X1 _13648_ (
    .A1(large_[29]),
    .A2(_00991_),
    .ZN(_01853_)
  );
  INV_X1 _13649_ (
    .A(_01853_),
    .ZN(_01854_)
  );
  AND2_X1 _13650_ (
    .A1(small_[3]),
    .A2(_00985_),
    .ZN(_01855_)
  );
  INV_X1 _13651_ (
    .A(_01855_),
    .ZN(_01856_)
  );
  AND2_X1 _13652_ (
    .A1(_01854_),
    .A2(_01856_),
    .ZN(_01857_)
  );
  AND2_X1 _13653_ (
    .A1(_01852_),
    .A2(_01857_),
    .ZN(_01858_)
  );
  AND2_X1 _13654_ (
    .A1(_01838_),
    .A2(_01858_),
    .ZN(_01859_)
  );
  AND2_X1 _13655_ (
    .A1(_01827_),
    .A2(_01859_),
    .ZN(_01860_)
  );
  INV_X1 _13656_ (
    .A(_01860_),
    .ZN(io_rw_rdata[3])
  );
  AND2_X1 _13657_ (
    .A1(io_rw_cmd[1]),
    .A2(_00839_),
    .ZN(_01861_)
  );
  AND2_X1 _13658_ (
    .A1(io_rw_rdata[3]),
    .A2(_01861_),
    .ZN(_01862_)
  );
  INV_X1 _13659_ (
    .A(_01862_),
    .ZN(_01863_)
  );
  AND2_X1 _13660_ (
    .A1(_01776_),
    .A2(_01863_),
    .ZN(_01864_)
  );
  INV_X1 _13661_ (
    .A(_01864_),
    .ZN(_01865_)
  );
  MUX2_X1 _13662_ (
    .A(reg_pmp_5_addr[3]),
    .B(_01865_),
    .S(_01525_),
    .Z(_00030_)
  );
  AND2_X1 _13663_ (
    .A1(io_rw_wdata[4]),
    .A2(_00903_),
    .ZN(_01866_)
  );
  INV_X1 _13664_ (
    .A(_01866_),
    .ZN(_01867_)
  );
  AND2_X1 _13665_ (
    .A1(reg_mscratch[4]),
    .A2(_00929_),
    .ZN(_01868_)
  );
  INV_X1 _13666_ (
    .A(_01868_),
    .ZN(_01869_)
  );
  AND2_X1 _13667_ (
    .A1(reg_mepc[4]),
    .A2(_00943_),
    .ZN(_01870_)
  );
  INV_X1 _13668_ (
    .A(_01870_),
    .ZN(_01871_)
  );
  AND2_X1 _13669_ (
    .A1(_01869_),
    .A2(_01871_),
    .ZN(_01872_)
  );
  AND2_X1 _13670_ (
    .A1(reg_pmp_0_addr[4]),
    .A2(_01004_),
    .ZN(_01873_)
  );
  INV_X1 _13671_ (
    .A(_01873_),
    .ZN(_01874_)
  );
  AND2_X1 _13672_ (
    .A1(reg_pmp_1_addr[4]),
    .A2(_01008_),
    .ZN(_01875_)
  );
  INV_X1 _13673_ (
    .A(_01875_),
    .ZN(_01876_)
  );
  AND2_X1 _13674_ (
    .A1(_01874_),
    .A2(_01876_),
    .ZN(_01877_)
  );
  AND2_X1 _13675_ (
    .A1(_01872_),
    .A2(_01877_),
    .ZN(_01878_)
  );
  AND2_X1 _13676_ (
    .A1(reg_mtvec[4]),
    .A2(_read_mtvec_T_4[6]),
    .ZN(_01879_)
  );
  AND2_X1 _13677_ (
    .A1(_00940_),
    .A2(_01879_),
    .ZN(_01880_)
  );
  INV_X1 _13678_ (
    .A(_01880_),
    .ZN(_01881_)
  );
  AND2_X1 _13679_ (
    .A1(reg_mtval[4]),
    .A2(_00926_),
    .ZN(_01882_)
  );
  INV_X1 _13680_ (
    .A(_01882_),
    .ZN(_01883_)
  );
  AND2_X1 _13681_ (
    .A1(_01881_),
    .A2(_01883_),
    .ZN(_01884_)
  );
  AND2_X1 _13682_ (
    .A1(reg_pmp_5_addr[4]),
    .A2(_00948_),
    .ZN(_01885_)
  );
  INV_X1 _13683_ (
    .A(_01885_),
    .ZN(_01886_)
  );
  AND2_X1 _13684_ (
    .A1(reg_mcause[4]),
    .A2(_01001_),
    .ZN(_01887_)
  );
  INV_X1 _13685_ (
    .A(_01887_),
    .ZN(_01888_)
  );
  AND2_X1 _13686_ (
    .A1(_01886_),
    .A2(_01888_),
    .ZN(_01889_)
  );
  AND2_X1 _13687_ (
    .A1(_01884_),
    .A2(_01889_),
    .ZN(_01890_)
  );
  AND2_X1 _13688_ (
    .A1(reg_pmp_4_addr[4]),
    .A2(_00968_),
    .ZN(_01891_)
  );
  INV_X1 _13689_ (
    .A(_01891_),
    .ZN(_01892_)
  );
  AND2_X1 _13690_ (
    .A1(reg_pmp_0_cfg_a[1]),
    .A2(_00916_),
    .ZN(_01893_)
  );
  INV_X1 _13691_ (
    .A(_01893_),
    .ZN(_01894_)
  );
  AND2_X1 _13692_ (
    .A1(_01892_),
    .A2(_01894_),
    .ZN(_01895_)
  );
  AND2_X1 _13693_ (
    .A1(reg_bp_0_address[4]),
    .A2(_00962_),
    .ZN(_01896_)
  );
  INV_X1 _13694_ (
    .A(_01896_),
    .ZN(_01897_)
  );
  AND2_X1 _13695_ (
    .A1(reg_pmp_4_cfg_a[1]),
    .A2(_00894_),
    .ZN(_01898_)
  );
  INV_X1 _13696_ (
    .A(_01898_),
    .ZN(_01899_)
  );
  AND2_X1 _13697_ (
    .A1(_01897_),
    .A2(_01899_),
    .ZN(_01900_)
  );
  AND2_X1 _13698_ (
    .A1(_01895_),
    .A2(_01900_),
    .ZN(_01901_)
  );
  AND2_X1 _13699_ (
    .A1(_01890_),
    .A2(_01901_),
    .ZN(_01902_)
  );
  AND2_X1 _13700_ (
    .A1(_01878_),
    .A2(_01902_),
    .ZN(_01903_)
  );
  AND2_X1 _13701_ (
    .A1(reg_pmp_6_addr[4]),
    .A2(_00978_),
    .ZN(_01904_)
  );
  INV_X1 _13702_ (
    .A(_01904_),
    .ZN(_01905_)
  );
  AND2_X1 _13703_ (
    .A1(large_1[30]),
    .A2(_01019_),
    .ZN(_01906_)
  );
  INV_X1 _13704_ (
    .A(_01906_),
    .ZN(_01907_)
  );
  AND2_X1 _13705_ (
    .A1(_01905_),
    .A2(_01907_),
    .ZN(_01908_)
  );
  AND2_X1 _13706_ (
    .A1(reg_pmp_7_addr[4]),
    .A2(_01016_),
    .ZN(_01909_)
  );
  INV_X1 _13707_ (
    .A(_01909_),
    .ZN(_01910_)
  );
  AND2_X1 _13708_ (
    .A1(small_1[4]),
    .A2(_00995_),
    .ZN(_01911_)
  );
  INV_X1 _13709_ (
    .A(_01911_),
    .ZN(_01912_)
  );
  AND2_X1 _13710_ (
    .A1(_01910_),
    .A2(_01912_),
    .ZN(_01913_)
  );
  AND2_X1 _13711_ (
    .A1(_01908_),
    .A2(_01913_),
    .ZN(_01914_)
  );
  AND2_X1 _13712_ (
    .A1(reg_pmp_3_addr[4]),
    .A2(_01011_),
    .ZN(_01915_)
  );
  INV_X1 _13713_ (
    .A(_01915_),
    .ZN(_01916_)
  );
  AND2_X1 _13714_ (
    .A1(reg_pmp_2_addr[4]),
    .A2(_00953_),
    .ZN(_01917_)
  );
  INV_X1 _13715_ (
    .A(_01917_),
    .ZN(_01918_)
  );
  AND2_X1 _13716_ (
    .A1(_01916_),
    .A2(_01918_),
    .ZN(_01919_)
  );
  AND2_X1 _13717_ (
    .A1(reg_dpc[4]),
    .A2(_00912_),
    .ZN(_01920_)
  );
  INV_X1 _13718_ (
    .A(_01920_),
    .ZN(_01921_)
  );
  AND2_X1 _13719_ (
    .A1(reg_dscratch0[4]),
    .A2(_00958_),
    .ZN(_01922_)
  );
  INV_X1 _13720_ (
    .A(_01922_),
    .ZN(_01923_)
  );
  AND2_X1 _13721_ (
    .A1(_01921_),
    .A2(_01923_),
    .ZN(_01924_)
  );
  AND2_X1 _13722_ (
    .A1(_01919_),
    .A2(_01924_),
    .ZN(_01925_)
  );
  AND2_X1 _13723_ (
    .A1(large_[30]),
    .A2(_00991_),
    .ZN(_01926_)
  );
  INV_X1 _13724_ (
    .A(_01926_),
    .ZN(_01927_)
  );
  AND2_X1 _13725_ (
    .A1(small_[4]),
    .A2(_00985_),
    .ZN(_01928_)
  );
  INV_X1 _13726_ (
    .A(_01928_),
    .ZN(_01929_)
  );
  AND2_X1 _13727_ (
    .A1(_01927_),
    .A2(_01929_),
    .ZN(_01930_)
  );
  AND2_X1 _13728_ (
    .A1(_01925_),
    .A2(_01930_),
    .ZN(_01931_)
  );
  AND2_X1 _13729_ (
    .A1(_01914_),
    .A2(_01931_),
    .ZN(_01932_)
  );
  AND2_X1 _13730_ (
    .A1(_01903_),
    .A2(_01932_),
    .ZN(_01933_)
  );
  INV_X1 _13731_ (
    .A(_01933_),
    .ZN(io_rw_rdata[4])
  );
  AND2_X1 _13732_ (
    .A1(io_rw_cmd[1]),
    .A2(_00840_),
    .ZN(_01934_)
  );
  AND2_X1 _13733_ (
    .A1(io_rw_rdata[4]),
    .A2(_01934_),
    .ZN(_01935_)
  );
  INV_X1 _13734_ (
    .A(_01935_),
    .ZN(_01936_)
  );
  AND2_X1 _13735_ (
    .A1(_01867_),
    .A2(_01936_),
    .ZN(_01937_)
  );
  INV_X1 _13736_ (
    .A(_01937_),
    .ZN(_01938_)
  );
  MUX2_X1 _13737_ (
    .A(reg_pmp_5_addr[4]),
    .B(_01938_),
    .S(_01525_),
    .Z(_00031_)
  );
  AND2_X1 _13738_ (
    .A1(io_rw_wdata[5]),
    .A2(_00903_),
    .ZN(_01939_)
  );
  INV_X1 _13739_ (
    .A(_01939_),
    .ZN(_01940_)
  );
  AND2_X1 _13740_ (
    .A1(reg_pmp_1_addr[5]),
    .A2(_01008_),
    .ZN(_01941_)
  );
  INV_X1 _13741_ (
    .A(_01941_),
    .ZN(_01942_)
  );
  AND2_X1 _13742_ (
    .A1(reg_pmp_4_addr[5]),
    .A2(_00968_),
    .ZN(_01943_)
  );
  INV_X1 _13743_ (
    .A(_01943_),
    .ZN(_01944_)
  );
  AND2_X1 _13744_ (
    .A1(reg_pmp_2_addr[5]),
    .A2(_00953_),
    .ZN(_01945_)
  );
  INV_X1 _13745_ (
    .A(_01945_),
    .ZN(_01946_)
  );
  AND2_X1 _13746_ (
    .A1(reg_dpc[5]),
    .A2(_00912_),
    .ZN(_01947_)
  );
  INV_X1 _13747_ (
    .A(_01947_),
    .ZN(_01948_)
  );
  AND2_X1 _13748_ (
    .A1(reg_pmp_0_addr[5]),
    .A2(_01004_),
    .ZN(_01949_)
  );
  INV_X1 _13749_ (
    .A(_01949_),
    .ZN(_01950_)
  );
  AND2_X1 _13750_ (
    .A1(reg_bp_0_address[5]),
    .A2(_00962_),
    .ZN(_01951_)
  );
  INV_X1 _13751_ (
    .A(_01951_),
    .ZN(_01952_)
  );
  AND2_X1 _13752_ (
    .A1(reg_mepc[5]),
    .A2(_00943_),
    .ZN(_01953_)
  );
  INV_X1 _13753_ (
    .A(_01953_),
    .ZN(_01954_)
  );
  AND2_X1 _13754_ (
    .A1(reg_mtvec[5]),
    .A2(_read_mtvec_T_4[6]),
    .ZN(_01955_)
  );
  AND2_X1 _13755_ (
    .A1(_00940_),
    .A2(_01955_),
    .ZN(_01956_)
  );
  INV_X1 _13756_ (
    .A(_01956_),
    .ZN(_01957_)
  );
  AND2_X1 _13757_ (
    .A1(reg_pmp_5_addr[5]),
    .A2(_00948_),
    .ZN(_01958_)
  );
  INV_X1 _13758_ (
    .A(_01958_),
    .ZN(_01959_)
  );
  AND2_X1 _13759_ (
    .A1(reg_dscratch0[5]),
    .A2(_00958_),
    .ZN(_01960_)
  );
  INV_X1 _13760_ (
    .A(_01960_),
    .ZN(_01961_)
  );
  AND2_X1 _13761_ (
    .A1(reg_mscratch[5]),
    .A2(_00929_),
    .ZN(_01962_)
  );
  INV_X1 _13762_ (
    .A(_01962_),
    .ZN(_01963_)
  );
  AND2_X1 _13763_ (
    .A1(reg_pmp_3_addr[5]),
    .A2(_01011_),
    .ZN(_01964_)
  );
  INV_X1 _13764_ (
    .A(_01964_),
    .ZN(_01965_)
  );
  AND2_X1 _13765_ (
    .A1(reg_pmp_6_addr[5]),
    .A2(_00978_),
    .ZN(_01966_)
  );
  INV_X1 _13766_ (
    .A(_01966_),
    .ZN(_01967_)
  );
  AND2_X1 _13767_ (
    .A1(reg_pmp_7_addr[5]),
    .A2(_01016_),
    .ZN(_01968_)
  );
  INV_X1 _13768_ (
    .A(_01968_),
    .ZN(_01969_)
  );
  AND2_X1 _13769_ (
    .A1(large_1[31]),
    .A2(_01019_),
    .ZN(_01970_)
  );
  INV_X1 _13770_ (
    .A(_01970_),
    .ZN(_01971_)
  );
  AND2_X1 _13771_ (
    .A1(reg_mtval[5]),
    .A2(_00926_),
    .ZN(_01972_)
  );
  INV_X1 _13772_ (
    .A(_01972_),
    .ZN(_01973_)
  );
  AND2_X1 _13773_ (
    .A1(reg_mcause[5]),
    .A2(_01001_),
    .ZN(_01974_)
  );
  INV_X1 _13774_ (
    .A(_01974_),
    .ZN(_01975_)
  );
  AND2_X1 _13775_ (
    .A1(large_[31]),
    .A2(_00991_),
    .ZN(_01976_)
  );
  INV_X1 _13776_ (
    .A(_01976_),
    .ZN(_01977_)
  );
  AND2_X1 _13777_ (
    .A1(_01942_),
    .A2(_01950_),
    .ZN(_01978_)
  );
  AND2_X1 _13778_ (
    .A1(small_[5]),
    .A2(_01027_),
    .ZN(_01979_)
  );
  INV_X1 _13779_ (
    .A(_01979_),
    .ZN(_01980_)
  );
  AND2_X1 _13780_ (
    .A1(small_1[5]),
    .A2(_01029_),
    .ZN(_01981_)
  );
  INV_X1 _13781_ (
    .A(_01981_),
    .ZN(_01982_)
  );
  AND2_X1 _13782_ (
    .A1(_01946_),
    .A2(_01969_),
    .ZN(_01983_)
  );
  AND2_X1 _13783_ (
    .A1(_01954_),
    .A2(_01975_),
    .ZN(_01984_)
  );
  AND2_X1 _13784_ (
    .A1(_01973_),
    .A2(_01984_),
    .ZN(_01985_)
  );
  AND2_X1 _13785_ (
    .A1(_01983_),
    .A2(_01985_),
    .ZN(_01986_)
  );
  AND2_X1 _13786_ (
    .A1(_01959_),
    .A2(_01978_),
    .ZN(_01987_)
  );
  AND2_X1 _13787_ (
    .A1(_01971_),
    .A2(_01977_),
    .ZN(_01988_)
  );
  AND2_X1 _13788_ (
    .A1(_01987_),
    .A2(_01988_),
    .ZN(_01989_)
  );
  AND2_X1 _13789_ (
    .A1(_01986_),
    .A2(_01989_),
    .ZN(_01990_)
  );
  AND2_X1 _13790_ (
    .A1(_01944_),
    .A2(_01957_),
    .ZN(_01991_)
  );
  AND2_X1 _13791_ (
    .A1(_01967_),
    .A2(_01991_),
    .ZN(_01992_)
  );
  AND2_X1 _13792_ (
    .A1(_01952_),
    .A2(_01963_),
    .ZN(_01993_)
  );
  AND2_X1 _13793_ (
    .A1(_01992_),
    .A2(_01993_),
    .ZN(_01994_)
  );
  AND2_X1 _13794_ (
    .A1(_01948_),
    .A2(_01965_),
    .ZN(_01995_)
  );
  AND2_X1 _13795_ (
    .A1(_01961_),
    .A2(_01980_),
    .ZN(_01996_)
  );
  AND2_X1 _13796_ (
    .A1(_01982_),
    .A2(_01996_),
    .ZN(_01997_)
  );
  AND2_X1 _13797_ (
    .A1(_01995_),
    .A2(_01997_),
    .ZN(_01998_)
  );
  AND2_X1 _13798_ (
    .A1(_01994_),
    .A2(_01998_),
    .ZN(_01999_)
  );
  AND2_X1 _13799_ (
    .A1(_01990_),
    .A2(_01999_),
    .ZN(_02000_)
  );
  INV_X1 _13800_ (
    .A(_02000_),
    .ZN(io_rw_rdata[5])
  );
  AND2_X1 _13801_ (
    .A1(io_rw_cmd[1]),
    .A2(_00841_),
    .ZN(_02001_)
  );
  AND2_X1 _13802_ (
    .A1(io_rw_rdata[5]),
    .A2(_02001_),
    .ZN(_02002_)
  );
  INV_X1 _13803_ (
    .A(_02002_),
    .ZN(_02003_)
  );
  AND2_X1 _13804_ (
    .A1(_01940_),
    .A2(_02003_),
    .ZN(_02004_)
  );
  INV_X1 _13805_ (
    .A(_02004_),
    .ZN(_02005_)
  );
  MUX2_X1 _13806_ (
    .A(reg_pmp_5_addr[5]),
    .B(_02005_),
    .S(_01525_),
    .Z(_00032_)
  );
  AND2_X1 _13807_ (
    .A1(io_rw_wdata[6]),
    .A2(_00903_),
    .ZN(_02006_)
  );
  INV_X1 _13808_ (
    .A(_02006_),
    .ZN(_02007_)
  );
  AND2_X1 _13809_ (
    .A1(reg_pmp_3_addr[6]),
    .A2(_01011_),
    .ZN(_02008_)
  );
  INV_X1 _13810_ (
    .A(_02008_),
    .ZN(_02009_)
  );
  AND2_X1 _13811_ (
    .A1(reg_pmp_2_addr[6]),
    .A2(_00953_),
    .ZN(_02010_)
  );
  INV_X1 _13812_ (
    .A(_02010_),
    .ZN(_02011_)
  );
  AND2_X1 _13813_ (
    .A1(reg_dcsr_cause[0]),
    .A2(_01381_),
    .ZN(_02012_)
  );
  INV_X1 _13814_ (
    .A(_02012_),
    .ZN(_02013_)
  );
  AND2_X1 _13815_ (
    .A1(reg_mepc[6]),
    .A2(_00943_),
    .ZN(_02014_)
  );
  INV_X1 _13816_ (
    .A(_02014_),
    .ZN(_02015_)
  );
  AND2_X1 _13817_ (
    .A1(reg_pmp_5_addr[6]),
    .A2(_00948_),
    .ZN(_02016_)
  );
  INV_X1 _13818_ (
    .A(_02016_),
    .ZN(_02017_)
  );
  AND2_X1 _13819_ (
    .A1(reg_dpc[6]),
    .A2(_00912_),
    .ZN(_02018_)
  );
  INV_X1 _13820_ (
    .A(_02018_),
    .ZN(_02019_)
  );
  AND2_X1 _13821_ (
    .A1(reg_pmp_1_addr[6]),
    .A2(_01008_),
    .ZN(_02020_)
  );
  INV_X1 _13822_ (
    .A(_02020_),
    .ZN(_02021_)
  );
  AND2_X1 _13823_ (
    .A1(reg_pmp_0_addr[6]),
    .A2(_01004_),
    .ZN(_02022_)
  );
  INV_X1 _13824_ (
    .A(_02022_),
    .ZN(_02023_)
  );
  AND2_X1 _13825_ (
    .A1(reg_pmp_4_addr[6]),
    .A2(_00968_),
    .ZN(_02024_)
  );
  INV_X1 _13826_ (
    .A(_02024_),
    .ZN(_02025_)
  );
  AND2_X1 _13827_ (
    .A1(reg_mcause[6]),
    .A2(_01001_),
    .ZN(_02026_)
  );
  INV_X1 _13828_ (
    .A(_02026_),
    .ZN(_02027_)
  );
  AND2_X1 _13829_ (
    .A1(reg_mtval[6]),
    .A2(_00926_),
    .ZN(_02028_)
  );
  INV_X1 _13830_ (
    .A(_02028_),
    .ZN(_02029_)
  );
  AND2_X1 _13831_ (
    .A1(reg_mscratch[6]),
    .A2(_00929_),
    .ZN(_02030_)
  );
  INV_X1 _13832_ (
    .A(_02030_),
    .ZN(_02031_)
  );
  AND2_X1 _13833_ (
    .A1(large_[32]),
    .A2(_00991_),
    .ZN(_02032_)
  );
  INV_X1 _13834_ (
    .A(_02032_),
    .ZN(_02033_)
  );
  AND2_X1 _13835_ (
    .A1(large_1[32]),
    .A2(_01019_),
    .ZN(_02034_)
  );
  INV_X1 _13836_ (
    .A(_02034_),
    .ZN(_02035_)
  );
  AND2_X1 _13837_ (
    .A1(reg_dscratch0[6]),
    .A2(_00958_),
    .ZN(_02036_)
  );
  INV_X1 _13838_ (
    .A(_02036_),
    .ZN(_02037_)
  );
  AND2_X1 _13839_ (
    .A1(reg_bp_0_address[6]),
    .A2(_00962_),
    .ZN(_02038_)
  );
  INV_X1 _13840_ (
    .A(_02038_),
    .ZN(_02039_)
  );
  AND2_X1 _13841_ (
    .A1(reg_mtvec[6]),
    .A2(_read_mtvec_T_4[6]),
    .ZN(_02040_)
  );
  AND2_X1 _13842_ (
    .A1(_00940_),
    .A2(_02040_),
    .ZN(_02041_)
  );
  INV_X1 _13843_ (
    .A(_02041_),
    .ZN(_02042_)
  );
  AND2_X1 _13844_ (
    .A1(reg_pmp_6_addr[6]),
    .A2(_00978_),
    .ZN(_02043_)
  );
  INV_X1 _13845_ (
    .A(_02043_),
    .ZN(_02044_)
  );
  AND2_X1 _13846_ (
    .A1(reg_pmp_7_addr[6]),
    .A2(_01016_),
    .ZN(_02045_)
  );
  INV_X1 _13847_ (
    .A(_02045_),
    .ZN(_02046_)
  );
  AND2_X1 _13848_ (
    .A1(_02011_),
    .A2(_02023_),
    .ZN(_02047_)
  );
  AND2_X1 _13849_ (
    .A1(large_[0]),
    .A2(_01027_),
    .ZN(_02048_)
  );
  INV_X1 _13850_ (
    .A(_02048_),
    .ZN(_02049_)
  );
  AND2_X1 _13851_ (
    .A1(large_1[0]),
    .A2(_01029_),
    .ZN(_02050_)
  );
  INV_X1 _13852_ (
    .A(_02050_),
    .ZN(_02051_)
  );
  AND2_X1 _13853_ (
    .A1(_02017_),
    .A2(_02025_),
    .ZN(_02052_)
  );
  AND2_X1 _13854_ (
    .A1(_02013_),
    .A2(_02052_),
    .ZN(_02053_)
  );
  AND2_X1 _13855_ (
    .A1(_02019_),
    .A2(_02037_),
    .ZN(_02054_)
  );
  AND2_X1 _13856_ (
    .A1(_02015_),
    .A2(_02029_),
    .ZN(_02055_)
  );
  AND2_X1 _13857_ (
    .A1(_02054_),
    .A2(_02055_),
    .ZN(_02056_)
  );
  AND2_X1 _13858_ (
    .A1(_02053_),
    .A2(_02056_),
    .ZN(_02057_)
  );
  AND2_X1 _13859_ (
    .A1(_02027_),
    .A2(_02044_),
    .ZN(_02058_)
  );
  AND2_X1 _13860_ (
    .A1(_02021_),
    .A2(_02058_),
    .ZN(_02059_)
  );
  AND2_X1 _13861_ (
    .A1(_02057_),
    .A2(_02059_),
    .ZN(_02060_)
  );
  AND2_X1 _13862_ (
    .A1(_01342_),
    .A2(_02039_),
    .ZN(_02061_)
  );
  AND2_X1 _13863_ (
    .A1(_02046_),
    .A2(_02061_),
    .ZN(_02062_)
  );
  AND2_X1 _13864_ (
    .A1(_02031_),
    .A2(_02033_),
    .ZN(_02063_)
  );
  AND2_X1 _13865_ (
    .A1(_02062_),
    .A2(_02063_),
    .ZN(_02064_)
  );
  AND2_X1 _13866_ (
    .A1(_02049_),
    .A2(_02051_),
    .ZN(_02065_)
  );
  AND2_X1 _13867_ (
    .A1(_02009_),
    .A2(_02042_),
    .ZN(_02066_)
  );
  AND2_X1 _13868_ (
    .A1(_02065_),
    .A2(_02066_),
    .ZN(_02067_)
  );
  AND2_X1 _13869_ (
    .A1(_02035_),
    .A2(_02047_),
    .ZN(_02068_)
  );
  AND2_X1 _13870_ (
    .A1(_02067_),
    .A2(_02068_),
    .ZN(_02069_)
  );
  AND2_X1 _13871_ (
    .A1(_02064_),
    .A2(_02069_),
    .ZN(_02070_)
  );
  AND2_X1 _13872_ (
    .A1(_02060_),
    .A2(_02070_),
    .ZN(_02071_)
  );
  INV_X1 _13873_ (
    .A(_02071_),
    .ZN(io_rw_rdata[6])
  );
  AND2_X1 _13874_ (
    .A1(io_rw_cmd[1]),
    .A2(_00842_),
    .ZN(_02072_)
  );
  AND2_X1 _13875_ (
    .A1(io_rw_rdata[6]),
    .A2(_02072_),
    .ZN(_02073_)
  );
  INV_X1 _13876_ (
    .A(_02073_),
    .ZN(_02074_)
  );
  AND2_X1 _13877_ (
    .A1(_02007_),
    .A2(_02074_),
    .ZN(_02075_)
  );
  INV_X1 _13878_ (
    .A(_02075_),
    .ZN(_02076_)
  );
  MUX2_X1 _13879_ (
    .A(reg_pmp_5_addr[6]),
    .B(_02076_),
    .S(_01525_),
    .Z(_00033_)
  );
  AND2_X1 _13880_ (
    .A1(io_rw_wdata[7]),
    .A2(_00903_),
    .ZN(_02077_)
  );
  INV_X1 _13881_ (
    .A(_02077_),
    .ZN(_02078_)
  );
  AND2_X1 _13882_ (
    .A1(reg_pmp_0_cfg_l),
    .A2(_00916_),
    .ZN(_02079_)
  );
  INV_X1 _13883_ (
    .A(_02079_),
    .ZN(_02080_)
  );
  AND2_X1 _13884_ (
    .A1(reg_mscratch[7]),
    .A2(_00929_),
    .ZN(_02081_)
  );
  INV_X1 _13885_ (
    .A(_02081_),
    .ZN(_02082_)
  );
  AND2_X1 _13886_ (
    .A1(reg_pmp_4_cfg_l),
    .A2(_00894_),
    .ZN(_02083_)
  );
  INV_X1 _13887_ (
    .A(_02083_),
    .ZN(_02084_)
  );
  AND2_X1 _13888_ (
    .A1(reg_mie[7]),
    .A2(_01782_),
    .ZN(_02085_)
  );
  INV_X1 _13889_ (
    .A(_02085_),
    .ZN(_02086_)
  );
  AND2_X1 _13890_ (
    .A1(reg_dpc[7]),
    .A2(_00912_),
    .ZN(_02087_)
  );
  INV_X1 _13891_ (
    .A(_02087_),
    .ZN(_02088_)
  );
  AND2_X1 _13892_ (
    .A1(reg_bp_0_control_tmatch[0]),
    .A2(_01341_),
    .ZN(_02089_)
  );
  INV_X1 _13893_ (
    .A(_02089_),
    .ZN(_02090_)
  );
  AND2_X1 _13894_ (
    .A1(reg_mtvec[7]),
    .A2(_00940_),
    .ZN(_02091_)
  );
  INV_X1 _13895_ (
    .A(_02091_),
    .ZN(_02092_)
  );
  AND2_X1 _13896_ (
    .A1(reg_pmp_5_addr[7]),
    .A2(_00948_),
    .ZN(_02093_)
  );
  INV_X1 _13897_ (
    .A(_02093_),
    .ZN(_02094_)
  );
  AND2_X1 _13898_ (
    .A1(reg_mtval[7]),
    .A2(_00926_),
    .ZN(_02095_)
  );
  INV_X1 _13899_ (
    .A(_02095_),
    .ZN(_02096_)
  );
  AND2_X1 _13900_ (
    .A1(reg_dscratch0[7]),
    .A2(_00958_),
    .ZN(_02097_)
  );
  INV_X1 _13901_ (
    .A(_02097_),
    .ZN(_02098_)
  );
  AND2_X1 _13902_ (
    .A1(reg_pmp_2_addr[7]),
    .A2(_00953_),
    .ZN(_02099_)
  );
  INV_X1 _13903_ (
    .A(_02099_),
    .ZN(_02100_)
  );
  AND2_X1 _13904_ (
    .A1(reg_pmp_7_addr[7]),
    .A2(_01016_),
    .ZN(_02101_)
  );
  INV_X1 _13905_ (
    .A(_02101_),
    .ZN(_02102_)
  );
  AND2_X1 _13906_ (
    .A1(large_1[33]),
    .A2(_01019_),
    .ZN(_02103_)
  );
  INV_X1 _13907_ (
    .A(_02103_),
    .ZN(_02104_)
  );
  AND2_X1 _13908_ (
    .A1(large_[33]),
    .A2(_00991_),
    .ZN(_02105_)
  );
  INV_X1 _13909_ (
    .A(_02105_),
    .ZN(_02106_)
  );
  AND2_X1 _13910_ (
    .A1(reg_pmp_4_addr[7]),
    .A2(_00968_),
    .ZN(_02107_)
  );
  INV_X1 _13911_ (
    .A(_02107_),
    .ZN(_02108_)
  );
  AND2_X1 _13912_ (
    .A1(reg_pmp_1_addr[7]),
    .A2(_01008_),
    .ZN(_02109_)
  );
  INV_X1 _13913_ (
    .A(_02109_),
    .ZN(_02110_)
  );
  AND2_X1 _13914_ (
    .A1(reg_pmp_6_addr[7]),
    .A2(_00978_),
    .ZN(_02111_)
  );
  INV_X1 _13915_ (
    .A(_02111_),
    .ZN(_02112_)
  );
  AND2_X1 _13916_ (
    .A1(io_interrupts_mtip),
    .A2(_01803_),
    .ZN(_02113_)
  );
  INV_X1 _13917_ (
    .A(_02113_),
    .ZN(_02114_)
  );
  AND2_X1 _13918_ (
    .A1(reg_mcause[7]),
    .A2(_01001_),
    .ZN(_02115_)
  );
  INV_X1 _13919_ (
    .A(_02115_),
    .ZN(_02116_)
  );
  AND2_X1 _13920_ (
    .A1(reg_mstatus_mpie),
    .A2(_01813_),
    .ZN(_02117_)
  );
  INV_X1 _13921_ (
    .A(_02117_),
    .ZN(_02118_)
  );
  AND2_X1 _13922_ (
    .A1(reg_pmp_0_addr[7]),
    .A2(_01004_),
    .ZN(_02119_)
  );
  INV_X1 _13923_ (
    .A(_02119_),
    .ZN(_02120_)
  );
  AND2_X1 _13924_ (
    .A1(reg_dcsr_cause[1]),
    .A2(_01381_),
    .ZN(_02121_)
  );
  INV_X1 _13925_ (
    .A(_02121_),
    .ZN(_02122_)
  );
  AND2_X1 _13926_ (
    .A1(reg_mepc[7]),
    .A2(_00943_),
    .ZN(_02123_)
  );
  INV_X1 _13927_ (
    .A(_02123_),
    .ZN(_02124_)
  );
  AND2_X1 _13928_ (
    .A1(reg_pmp_3_addr[7]),
    .A2(_01011_),
    .ZN(_02125_)
  );
  INV_X1 _13929_ (
    .A(_02125_),
    .ZN(_02126_)
  );
  AND2_X1 _13930_ (
    .A1(reg_bp_0_address[7]),
    .A2(_00962_),
    .ZN(_02127_)
  );
  INV_X1 _13931_ (
    .A(_02127_),
    .ZN(_02128_)
  );
  AND2_X1 _13932_ (
    .A1(_02082_),
    .A2(_02092_),
    .ZN(_02129_)
  );
  AND2_X1 _13933_ (
    .A1(large_1[1]),
    .A2(_01029_),
    .ZN(_02130_)
  );
  INV_X1 _13934_ (
    .A(_02130_),
    .ZN(_02131_)
  );
  AND2_X1 _13935_ (
    .A1(_02096_),
    .A2(_02131_),
    .ZN(_02132_)
  );
  AND2_X1 _13936_ (
    .A1(_02129_),
    .A2(_02132_),
    .ZN(_02133_)
  );
  AND2_X1 _13937_ (
    .A1(large_[1]),
    .A2(_01027_),
    .ZN(_02134_)
  );
  INV_X1 _13938_ (
    .A(_02134_),
    .ZN(_02135_)
  );
  AND2_X1 _13939_ (
    .A1(_02100_),
    .A2(_02110_),
    .ZN(_02136_)
  );
  AND2_X1 _13940_ (
    .A1(_02106_),
    .A2(_02136_),
    .ZN(_02137_)
  );
  AND2_X1 _13941_ (
    .A1(_02086_),
    .A2(_02118_),
    .ZN(_02138_)
  );
  AND2_X1 _13942_ (
    .A1(_02080_),
    .A2(_02084_),
    .ZN(_02139_)
  );
  AND2_X1 _13943_ (
    .A1(_02112_),
    .A2(_02139_),
    .ZN(_02140_)
  );
  AND2_X1 _13944_ (
    .A1(_02108_),
    .A2(_02126_),
    .ZN(_02141_)
  );
  AND2_X1 _13945_ (
    .A1(_02090_),
    .A2(_02141_),
    .ZN(_02142_)
  );
  AND2_X1 _13946_ (
    .A1(_02114_),
    .A2(_02138_),
    .ZN(_02143_)
  );
  AND2_X1 _13947_ (
    .A1(_02094_),
    .A2(_02120_),
    .ZN(_02144_)
  );
  AND2_X1 _13948_ (
    .A1(_02104_),
    .A2(_02144_),
    .ZN(_02145_)
  );
  AND2_X1 _13949_ (
    .A1(_02143_),
    .A2(_02145_),
    .ZN(_02146_)
  );
  AND2_X1 _13950_ (
    .A1(_02142_),
    .A2(_02146_),
    .ZN(_02147_)
  );
  AND2_X1 _13951_ (
    .A1(_02116_),
    .A2(_02122_),
    .ZN(_02148_)
  );
  AND2_X1 _13952_ (
    .A1(_02135_),
    .A2(_02148_),
    .ZN(_02149_)
  );
  AND2_X1 _13953_ (
    .A1(_02098_),
    .A2(_02128_),
    .ZN(_02150_)
  );
  AND2_X1 _13954_ (
    .A1(_02149_),
    .A2(_02150_),
    .ZN(_02151_)
  );
  AND2_X1 _13955_ (
    .A1(_02088_),
    .A2(_02124_),
    .ZN(_02152_)
  );
  AND2_X1 _13956_ (
    .A1(_02133_),
    .A2(_02152_),
    .ZN(_02153_)
  );
  AND2_X1 _13957_ (
    .A1(_02151_),
    .A2(_02153_),
    .ZN(_02154_)
  );
  AND2_X1 _13958_ (
    .A1(_02102_),
    .A2(_02137_),
    .ZN(_02155_)
  );
  AND2_X1 _13959_ (
    .A1(_02140_),
    .A2(_02155_),
    .ZN(_02156_)
  );
  AND2_X1 _13960_ (
    .A1(_02154_),
    .A2(_02156_),
    .ZN(_02157_)
  );
  AND2_X1 _13961_ (
    .A1(_02147_),
    .A2(_02157_),
    .ZN(_02158_)
  );
  INV_X1 _13962_ (
    .A(_02158_),
    .ZN(io_rw_rdata[7])
  );
  AND2_X1 _13963_ (
    .A1(io_rw_cmd[1]),
    .A2(_00843_),
    .ZN(_02159_)
  );
  AND2_X1 _13964_ (
    .A1(io_rw_rdata[7]),
    .A2(_02159_),
    .ZN(_02160_)
  );
  INV_X1 _13965_ (
    .A(_02160_),
    .ZN(_02161_)
  );
  AND2_X1 _13966_ (
    .A1(_02078_),
    .A2(_02161_),
    .ZN(_02162_)
  );
  INV_X1 _13967_ (
    .A(_02162_),
    .ZN(_02163_)
  );
  MUX2_X1 _13968_ (
    .A(reg_pmp_5_addr[7]),
    .B(_02163_),
    .S(_01525_),
    .Z(_00034_)
  );
  MUX2_X1 _13969_ (
    .A(reg_pmp_5_addr[8]),
    .B(_01446_),
    .S(_01525_),
    .Z(_00035_)
  );
  MUX2_X1 _13970_ (
    .A(reg_pmp_5_addr[9]),
    .B(_01518_),
    .S(_01525_),
    .Z(_00036_)
  );
  AND2_X1 _13971_ (
    .A1(io_rw_wdata[10]),
    .A2(_00903_),
    .ZN(_02164_)
  );
  INV_X1 _13972_ (
    .A(_02164_),
    .ZN(_02165_)
  );
  AND2_X1 _13973_ (
    .A1(reg_dscratch0[10]),
    .A2(_00958_),
    .ZN(_02166_)
  );
  INV_X1 _13974_ (
    .A(_02166_),
    .ZN(_02167_)
  );
  AND2_X1 _13975_ (
    .A1(reg_pmp_1_addr[10]),
    .A2(_01008_),
    .ZN(_02168_)
  );
  INV_X1 _13976_ (
    .A(_02168_),
    .ZN(_02169_)
  );
  AND2_X1 _13977_ (
    .A1(_02167_),
    .A2(_02169_),
    .ZN(_02170_)
  );
  AND2_X1 _13978_ (
    .A1(reg_bp_0_address[10]),
    .A2(_00962_),
    .ZN(_02171_)
  );
  INV_X1 _13979_ (
    .A(_02171_),
    .ZN(_02172_)
  );
  AND2_X1 _13980_ (
    .A1(reg_pmp_5_addr[10]),
    .A2(_00948_),
    .ZN(_02173_)
  );
  INV_X1 _13981_ (
    .A(_02173_),
    .ZN(_02174_)
  );
  AND2_X1 _13982_ (
    .A1(_02172_),
    .A2(_02174_),
    .ZN(_02175_)
  );
  AND2_X1 _13983_ (
    .A1(_02170_),
    .A2(_02175_),
    .ZN(_02176_)
  );
  AND2_X1 _13984_ (
    .A1(reg_mepc[10]),
    .A2(_00943_),
    .ZN(_02177_)
  );
  INV_X1 _13985_ (
    .A(_02177_),
    .ZN(_02178_)
  );
  AND2_X1 _13986_ (
    .A1(reg_pmp_0_addr[10]),
    .A2(_01004_),
    .ZN(_02179_)
  );
  INV_X1 _13987_ (
    .A(_02179_),
    .ZN(_02180_)
  );
  AND2_X1 _13988_ (
    .A1(_02178_),
    .A2(_02180_),
    .ZN(_02181_)
  );
  AND2_X1 _13989_ (
    .A1(reg_pmp_1_cfg_x),
    .A2(_00916_),
    .ZN(_02182_)
  );
  INV_X1 _13990_ (
    .A(_02182_),
    .ZN(_02183_)
  );
  AND2_X1 _13991_ (
    .A1(reg_pmp_3_addr[10]),
    .A2(_01011_),
    .ZN(_02184_)
  );
  INV_X1 _13992_ (
    .A(_02184_),
    .ZN(_02185_)
  );
  AND2_X1 _13993_ (
    .A1(_02183_),
    .A2(_02185_),
    .ZN(_02186_)
  );
  AND2_X1 _13994_ (
    .A1(_02181_),
    .A2(_02186_),
    .ZN(_02187_)
  );
  AND2_X1 _13995_ (
    .A1(reg_mtvec[10]),
    .A2(_00940_),
    .ZN(_02188_)
  );
  INV_X1 _13996_ (
    .A(_02188_),
    .ZN(_02189_)
  );
  AND2_X1 _13997_ (
    .A1(reg_mtval[10]),
    .A2(_00926_),
    .ZN(_02190_)
  );
  INV_X1 _13998_ (
    .A(_02190_),
    .ZN(_02191_)
  );
  AND2_X1 _13999_ (
    .A1(_02189_),
    .A2(_02191_),
    .ZN(_02192_)
  );
  AND2_X1 _14000_ (
    .A1(reg_pmp_5_cfg_x),
    .A2(_00894_),
    .ZN(_02193_)
  );
  INV_X1 _14001_ (
    .A(_02193_),
    .ZN(_02194_)
  );
  AND2_X1 _14002_ (
    .A1(reg_mcause[10]),
    .A2(_01001_),
    .ZN(_02195_)
  );
  INV_X1 _14003_ (
    .A(_02195_),
    .ZN(_02196_)
  );
  AND2_X1 _14004_ (
    .A1(_02194_),
    .A2(_02196_),
    .ZN(_02197_)
  );
  AND2_X1 _14005_ (
    .A1(_02192_),
    .A2(_02197_),
    .ZN(_02198_)
  );
  AND2_X1 _14006_ (
    .A1(_02187_),
    .A2(_02198_),
    .ZN(_02199_)
  );
  AND2_X1 _14007_ (
    .A1(_02176_),
    .A2(_02199_),
    .ZN(_02200_)
  );
  AND2_X1 _14008_ (
    .A1(reg_pmp_7_addr[10]),
    .A2(_01016_),
    .ZN(_02201_)
  );
  INV_X1 _14009_ (
    .A(_02201_),
    .ZN(_02202_)
  );
  AND2_X1 _14010_ (
    .A1(large_[36]),
    .A2(_00991_),
    .ZN(_02203_)
  );
  INV_X1 _14011_ (
    .A(_02203_),
    .ZN(_02204_)
  );
  AND2_X1 _14012_ (
    .A1(_02202_),
    .A2(_02204_),
    .ZN(_02205_)
  );
  AND2_X1 _14013_ (
    .A1(large_1[36]),
    .A2(_01019_),
    .ZN(_02206_)
  );
  INV_X1 _14014_ (
    .A(_02206_),
    .ZN(_02207_)
  );
  AND2_X1 _14015_ (
    .A1(large_[4]),
    .A2(_00985_),
    .ZN(_02208_)
  );
  INV_X1 _14016_ (
    .A(_02208_),
    .ZN(_02209_)
  );
  AND2_X1 _14017_ (
    .A1(_02207_),
    .A2(_02209_),
    .ZN(_02210_)
  );
  AND2_X1 _14018_ (
    .A1(_02205_),
    .A2(_02210_),
    .ZN(_02211_)
  );
  AND2_X1 _14019_ (
    .A1(reg_dpc[10]),
    .A2(_00912_),
    .ZN(_02212_)
  );
  INV_X1 _14020_ (
    .A(_02212_),
    .ZN(_02213_)
  );
  AND2_X1 _14021_ (
    .A1(reg_mscratch[10]),
    .A2(_00929_),
    .ZN(_02214_)
  );
  INV_X1 _14022_ (
    .A(_02214_),
    .ZN(_02215_)
  );
  AND2_X1 _14023_ (
    .A1(_02213_),
    .A2(_02215_),
    .ZN(_02216_)
  );
  AND2_X1 _14024_ (
    .A1(reg_pmp_4_addr[10]),
    .A2(_00968_),
    .ZN(_02217_)
  );
  INV_X1 _14025_ (
    .A(_02217_),
    .ZN(_02218_)
  );
  AND2_X1 _14026_ (
    .A1(reg_pmp_2_addr[10]),
    .A2(_00953_),
    .ZN(_02219_)
  );
  INV_X1 _14027_ (
    .A(_02219_),
    .ZN(_02220_)
  );
  AND2_X1 _14028_ (
    .A1(_02218_),
    .A2(_02220_),
    .ZN(_02221_)
  );
  AND2_X1 _14029_ (
    .A1(_02216_),
    .A2(_02221_),
    .ZN(_02222_)
  );
  AND2_X1 _14030_ (
    .A1(reg_pmp_6_addr[10]),
    .A2(_00978_),
    .ZN(_02223_)
  );
  INV_X1 _14031_ (
    .A(_02223_),
    .ZN(_02224_)
  );
  AND2_X1 _14032_ (
    .A1(large_1[4]),
    .A2(_00995_),
    .ZN(_02225_)
  );
  INV_X1 _14033_ (
    .A(_02225_),
    .ZN(_02226_)
  );
  AND2_X1 _14034_ (
    .A1(_02224_),
    .A2(_02226_),
    .ZN(_02227_)
  );
  AND2_X1 _14035_ (
    .A1(_02222_),
    .A2(_02227_),
    .ZN(_02228_)
  );
  AND2_X1 _14036_ (
    .A1(_02211_),
    .A2(_02228_),
    .ZN(_02229_)
  );
  AND2_X1 _14037_ (
    .A1(_02200_),
    .A2(_02229_),
    .ZN(_02230_)
  );
  INV_X1 _14038_ (
    .A(_02230_),
    .ZN(io_rw_rdata[10])
  );
  AND2_X1 _14039_ (
    .A1(io_rw_cmd[1]),
    .A2(_00846_),
    .ZN(_02231_)
  );
  AND2_X1 _14040_ (
    .A1(io_rw_rdata[10]),
    .A2(_02231_),
    .ZN(_02232_)
  );
  INV_X1 _14041_ (
    .A(_02232_),
    .ZN(_02233_)
  );
  DFF_X1 \io_status_cease_r$_SDFF_PP0_  (
    .CK(clock),
    .D(_00021_),
    .Q(io_status_cease_r),
    .QN(_07071_)
  );
  DFF_X1 \large_1[0]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00569_),
    .Q(large_1[0]),
    .QN(_large_r_T_3[0])
  );
  DFF_X1 \large_1[10]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00579_),
    .Q(large_1[10]),
    .QN(_06534_)
  );
  DFF_X1 \large_1[11]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00580_),
    .Q(large_1[11]),
    .QN(_06533_)
  );
  DFF_X1 \large_1[12]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00581_),
    .Q(large_1[12]),
    .QN(_06532_)
  );
  DFF_X1 \large_1[13]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00582_),
    .Q(large_1[13]),
    .QN(_06531_)
  );
  DFF_X1 \large_1[14]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00583_),
    .Q(large_1[14]),
    .QN(_06530_)
  );
  DFF_X1 \large_1[15]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00584_),
    .Q(large_1[15]),
    .QN(_06529_)
  );
  DFF_X1 \large_1[16]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00585_),
    .Q(large_1[16]),
    .QN(_06528_)
  );
  DFF_X1 \large_1[17]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00586_),
    .Q(large_1[17]),
    .QN(_06527_)
  );
  DFF_X1 \large_1[18]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00587_),
    .Q(large_1[18]),
    .QN(_06526_)
  );
  DFF_X1 \large_1[19]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00588_),
    .Q(large_1[19]),
    .QN(_06525_)
  );
  DFF_X1 \large_1[1]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00570_),
    .Q(large_1[1]),
    .QN(_06543_)
  );
  DFF_X1 \large_1[20]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00589_),
    .Q(large_1[20]),
    .QN(_06524_)
  );
  DFF_X1 \large_1[21]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00590_),
    .Q(large_1[21]),
    .QN(_06523_)
  );
  DFF_X1 \large_1[22]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00591_),
    .Q(large_1[22]),
    .QN(_06522_)
  );
  DFF_X1 \large_1[23]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00592_),
    .Q(large_1[23]),
    .QN(_06521_)
  );
  DFF_X1 \large_1[24]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00593_),
    .Q(large_1[24]),
    .QN(_06520_)
  );
  DFF_X1 \large_1[25]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00594_),
    .Q(large_1[25]),
    .QN(_06519_)
  );
  DFF_X1 \large_1[26]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00294_),
    .Q(large_1[26]),
    .QN(_06814_)
  );
  DFF_X1 \large_1[27]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00295_),
    .Q(large_1[27]),
    .QN(_06813_)
  );
  DFF_X1 \large_1[28]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00296_),
    .Q(large_1[28]),
    .QN(_06812_)
  );
  DFF_X1 \large_1[29]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00297_),
    .Q(large_1[29]),
    .QN(_06811_)
  );
  DFF_X1 \large_1[2]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00571_),
    .Q(large_1[2]),
    .QN(_06542_)
  );
  DFF_X1 \large_1[30]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00298_),
    .Q(large_1[30]),
    .QN(_06810_)
  );
  DFF_X1 \large_1[31]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00299_),
    .Q(large_1[31]),
    .QN(_06809_)
  );
  DFF_X1 \large_1[32]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00300_),
    .Q(large_1[32]),
    .QN(_06808_)
  );
  DFF_X1 \large_1[33]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00301_),
    .Q(large_1[33]),
    .QN(_06807_)
  );
  DFF_X1 \large_1[34]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00302_),
    .Q(large_1[34]),
    .QN(_06806_)
  );
  DFF_X1 \large_1[35]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00303_),
    .Q(large_1[35]),
    .QN(_06805_)
  );
  DFF_X1 \large_1[36]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00304_),
    .Q(large_1[36]),
    .QN(_06804_)
  );
  DFF_X1 \large_1[37]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00305_),
    .Q(large_1[37]),
    .QN(_06803_)
  );
  DFF_X1 \large_1[38]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00306_),
    .Q(large_1[38]),
    .QN(_06802_)
  );
  DFF_X1 \large_1[39]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00307_),
    .Q(large_1[39]),
    .QN(_06801_)
  );
  DFF_X1 \large_1[3]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00572_),
    .Q(large_1[3]),
    .QN(_06541_)
  );
  DFF_X1 \large_1[40]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00308_),
    .Q(large_1[40]),
    .QN(_06800_)
  );
  DFF_X1 \large_1[41]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00309_),
    .Q(large_1[41]),
    .QN(_06799_)
  );
  DFF_X1 \large_1[42]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00310_),
    .Q(large_1[42]),
    .QN(_06798_)
  );
  DFF_X1 \large_1[43]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00311_),
    .Q(large_1[43]),
    .QN(_06797_)
  );
  DFF_X1 \large_1[44]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00312_),
    .Q(large_1[44]),
    .QN(_06796_)
  );
  DFF_X1 \large_1[45]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00313_),
    .Q(large_1[45]),
    .QN(_06795_)
  );
  DFF_X1 \large_1[46]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00314_),
    .Q(large_1[46]),
    .QN(_06794_)
  );
  DFF_X1 \large_1[47]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00315_),
    .Q(large_1[47]),
    .QN(_06793_)
  );
  DFF_X1 \large_1[48]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00316_),
    .Q(large_1[48]),
    .QN(_06792_)
  );
  DFF_X1 \large_1[49]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00317_),
    .Q(large_1[49]),
    .QN(_06791_)
  );
  DFF_X1 \large_1[4]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00573_),
    .Q(large_1[4]),
    .QN(_06540_)
  );
  DFF_X1 \large_1[50]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00318_),
    .Q(large_1[50]),
    .QN(_06790_)
  );
  DFF_X1 \large_1[51]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00319_),
    .Q(large_1[51]),
    .QN(_06789_)
  );
  DFF_X1 \large_1[52]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00320_),
    .Q(large_1[52]),
    .QN(_06788_)
  );
  DFF_X1 \large_1[53]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00321_),
    .Q(large_1[53]),
    .QN(_06787_)
  );
  DFF_X1 \large_1[54]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00322_),
    .Q(large_1[54]),
    .QN(_06786_)
  );
  DFF_X1 \large_1[55]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00323_),
    .Q(large_1[55]),
    .QN(_06785_)
  );
  DFF_X1 \large_1[56]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00324_),
    .Q(large_1[56]),
    .QN(_06784_)
  );
  DFF_X1 \large_1[57]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00325_),
    .Q(large_1[57]),
    .QN(_06783_)
  );
  DFF_X1 \large_1[5]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00574_),
    .Q(large_1[5]),
    .QN(_06539_)
  );
  DFF_X1 \large_1[6]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00575_),
    .Q(large_1[6]),
    .QN(_06538_)
  );
  DFF_X1 \large_1[7]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00576_),
    .Q(large_1[7]),
    .QN(_06537_)
  );
  DFF_X1 \large_1[8]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00577_),
    .Q(large_1[8]),
    .QN(_06536_)
  );
  DFF_X1 \large_1[9]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00578_),
    .Q(large_1[9]),
    .QN(_06535_)
  );
  DFF_X1 \large_[0]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00595_),
    .Q(large_[0]),
    .QN(_large_r_T_1[0])
  );
  DFF_X1 \large_[10]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00605_),
    .Q(large_[10]),
    .QN(_06509_)
  );
  DFF_X1 \large_[11]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00606_),
    .Q(large_[11]),
    .QN(_06508_)
  );
  DFF_X1 \large_[12]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00607_),
    .Q(large_[12]),
    .QN(_06507_)
  );
  DFF_X1 \large_[13]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00608_),
    .Q(large_[13]),
    .QN(_06506_)
  );
  DFF_X1 \large_[14]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00609_),
    .Q(large_[14]),
    .QN(_06505_)
  );
  DFF_X1 \large_[15]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00610_),
    .Q(large_[15]),
    .QN(_06504_)
  );
  DFF_X1 \large_[16]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00611_),
    .Q(large_[16]),
    .QN(_06503_)
  );
  DFF_X1 \large_[17]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00612_),
    .Q(large_[17]),
    .QN(_06502_)
  );
  DFF_X1 \large_[18]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00613_),
    .Q(large_[18]),
    .QN(_06501_)
  );
  DFF_X1 \large_[19]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00614_),
    .Q(large_[19]),
    .QN(_06500_)
  );
  DFF_X1 \large_[1]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00596_),
    .Q(large_[1]),
    .QN(_06518_)
  );
  DFF_X1 \large_[20]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00615_),
    .Q(large_[20]),
    .QN(_06499_)
  );
  DFF_X1 \large_[21]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00616_),
    .Q(large_[21]),
    .QN(_06498_)
  );
  DFF_X1 \large_[22]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00617_),
    .Q(large_[22]),
    .QN(_06497_)
  );
  DFF_X1 \large_[23]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00618_),
    .Q(large_[23]),
    .QN(_06496_)
  );
  DFF_X1 \large_[24]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00619_),
    .Q(large_[24]),
    .QN(_06495_)
  );
  DFF_X1 \large_[25]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00620_),
    .Q(large_[25]),
    .QN(_06494_)
  );
  DFF_X1 \large_[26]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00429_),
    .Q(large_[26]),
    .QN(_06680_)
  );
  DFF_X1 \large_[27]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00430_),
    .Q(large_[27]),
    .QN(_06679_)
  );
  DFF_X1 \large_[28]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00431_),
    .Q(large_[28]),
    .QN(_06678_)
  );
  DFF_X1 \large_[29]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00432_),
    .Q(large_[29]),
    .QN(_06677_)
  );
  DFF_X1 \large_[2]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00597_),
    .Q(large_[2]),
    .QN(_06517_)
  );
  DFF_X1 \large_[30]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00433_),
    .Q(large_[30]),
    .QN(_06676_)
  );
  DFF_X1 \large_[31]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00434_),
    .Q(large_[31]),
    .QN(_06675_)
  );
  DFF_X1 \large_[32]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00435_),
    .Q(large_[32]),
    .QN(_06674_)
  );
  DFF_X1 \large_[33]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00436_),
    .Q(large_[33]),
    .QN(_06673_)
  );
  DFF_X1 \large_[34]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00437_),
    .Q(large_[34]),
    .QN(_06672_)
  );
  DFF_X1 \large_[35]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00438_),
    .Q(large_[35]),
    .QN(_06671_)
  );
  DFF_X1 \large_[36]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00439_),
    .Q(large_[36]),
    .QN(_06670_)
  );
  DFF_X1 \large_[37]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00440_),
    .Q(large_[37]),
    .QN(_06669_)
  );
  DFF_X1 \large_[38]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00441_),
    .Q(large_[38]),
    .QN(_06668_)
  );
  DFF_X1 \large_[39]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00442_),
    .Q(large_[39]),
    .QN(_06667_)
  );
  DFF_X1 \large_[3]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00598_),
    .Q(large_[3]),
    .QN(_06516_)
  );
  DFF_X1 \large_[40]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00443_),
    .Q(large_[40]),
    .QN(_06666_)
  );
  DFF_X1 \large_[41]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00444_),
    .Q(large_[41]),
    .QN(_06665_)
  );
  DFF_X1 \large_[42]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00445_),
    .Q(large_[42]),
    .QN(_06664_)
  );
  DFF_X1 \large_[43]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00446_),
    .Q(large_[43]),
    .QN(_06663_)
  );
  DFF_X1 \large_[44]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00447_),
    .Q(large_[44]),
    .QN(_06662_)
  );
  DFF_X1 \large_[45]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00448_),
    .Q(large_[45]),
    .QN(_06661_)
  );
  DFF_X1 \large_[46]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00449_),
    .Q(large_[46]),
    .QN(_06660_)
  );
  DFF_X1 \large_[47]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00450_),
    .Q(large_[47]),
    .QN(_06659_)
  );
  DFF_X1 \large_[48]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00451_),
    .Q(large_[48]),
    .QN(_06658_)
  );
  DFF_X1 \large_[49]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00452_),
    .Q(large_[49]),
    .QN(_06657_)
  );
  DFF_X1 \large_[4]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00599_),
    .Q(large_[4]),
    .QN(_06515_)
  );
  DFF_X1 \large_[50]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00453_),
    .Q(large_[50]),
    .QN(_06656_)
  );
  DFF_X1 \large_[51]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00454_),
    .Q(large_[51]),
    .QN(_06655_)
  );
  DFF_X1 \large_[52]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00455_),
    .Q(large_[52]),
    .QN(_06654_)
  );
  DFF_X1 \large_[53]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00456_),
    .Q(large_[53]),
    .QN(_06653_)
  );
  DFF_X1 \large_[54]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00457_),
    .Q(large_[54]),
    .QN(_06652_)
  );
  DFF_X1 \large_[55]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00458_),
    .Q(large_[55]),
    .QN(_06651_)
  );
  DFF_X1 \large_[56]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00459_),
    .Q(large_[56]),
    .QN(_06650_)
  );
  DFF_X1 \large_[57]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00460_),
    .Q(large_[57]),
    .QN(_06649_)
  );
  DFF_X1 \large_[5]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00600_),
    .Q(large_[5]),
    .QN(_06514_)
  );
  DFF_X1 \large_[6]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00601_),
    .Q(large_[6]),
    .QN(_06513_)
  );
  DFF_X1 \large_[7]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00602_),
    .Q(large_[7]),
    .QN(_06512_)
  );
  DFF_X1 \large_[8]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00603_),
    .Q(large_[8]),
    .QN(_06511_)
  );
  DFF_X1 \large_[9]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00604_),
    .Q(large_[9]),
    .QN(_06510_)
  );
  DFF_X1 \reg_bp_0_address[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00207_),
    .Q(reg_bp_0_address[0]),
    .QN(_06897_)
  );
  DFF_X1 \reg_bp_0_address[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00217_),
    .Q(reg_bp_0_address[10]),
    .QN(_06887_)
  );
  DFF_X1 \reg_bp_0_address[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00218_),
    .Q(reg_bp_0_address[11]),
    .QN(_06886_)
  );
  DFF_X1 \reg_bp_0_address[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00219_),
    .Q(reg_bp_0_address[12]),
    .QN(_06885_)
  );
  DFF_X1 \reg_bp_0_address[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00220_),
    .Q(reg_bp_0_address[13]),
    .QN(_06884_)
  );
  DFF_X1 \reg_bp_0_address[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00221_),
    .Q(reg_bp_0_address[14]),
    .QN(_06883_)
  );
  DFF_X1 \reg_bp_0_address[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00222_),
    .Q(reg_bp_0_address[15]),
    .QN(_06882_)
  );
  DFF_X1 \reg_bp_0_address[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00223_),
    .Q(reg_bp_0_address[16]),
    .QN(_06881_)
  );
  DFF_X1 \reg_bp_0_address[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00224_),
    .Q(reg_bp_0_address[17]),
    .QN(_06880_)
  );
  DFF_X1 \reg_bp_0_address[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00225_),
    .Q(reg_bp_0_address[18]),
    .QN(_06879_)
  );
  DFF_X1 \reg_bp_0_address[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00226_),
    .Q(reg_bp_0_address[19]),
    .QN(_06878_)
  );
  DFF_X1 \reg_bp_0_address[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00208_),
    .Q(reg_bp_0_address[1]),
    .QN(_06896_)
  );
  DFF_X1 \reg_bp_0_address[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00227_),
    .Q(reg_bp_0_address[20]),
    .QN(_06877_)
  );
  DFF_X1 \reg_bp_0_address[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00228_),
    .Q(reg_bp_0_address[21]),
    .QN(_06876_)
  );
  DFF_X1 \reg_bp_0_address[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00229_),
    .Q(reg_bp_0_address[22]),
    .QN(_06875_)
  );
  DFF_X1 \reg_bp_0_address[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00230_),
    .Q(reg_bp_0_address[23]),
    .QN(_06874_)
  );
  DFF_X1 \reg_bp_0_address[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00231_),
    .Q(reg_bp_0_address[24]),
    .QN(_06873_)
  );
  DFF_X1 \reg_bp_0_address[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00232_),
    .Q(reg_bp_0_address[25]),
    .QN(_06872_)
  );
  DFF_X1 \reg_bp_0_address[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00233_),
    .Q(reg_bp_0_address[26]),
    .QN(_06871_)
  );
  DFF_X1 \reg_bp_0_address[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00234_),
    .Q(reg_bp_0_address[27]),
    .QN(_06870_)
  );
  DFF_X1 \reg_bp_0_address[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00235_),
    .Q(reg_bp_0_address[28]),
    .QN(_06869_)
  );
  DFF_X1 \reg_bp_0_address[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00236_),
    .Q(reg_bp_0_address[29]),
    .QN(_06868_)
  );
  DFF_X1 \reg_bp_0_address[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00209_),
    .Q(reg_bp_0_address[2]),
    .QN(_06895_)
  );
  DFF_X1 \reg_bp_0_address[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00237_),
    .Q(reg_bp_0_address[30]),
    .QN(_06867_)
  );
  DFF_X1 \reg_bp_0_address[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00238_),
    .Q(reg_bp_0_address[31]),
    .QN(_06866_)
  );
  DFF_X1 \reg_bp_0_address[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00210_),
    .Q(reg_bp_0_address[3]),
    .QN(_06894_)
  );
  DFF_X1 \reg_bp_0_address[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00211_),
    .Q(reg_bp_0_address[4]),
    .QN(_06893_)
  );
  DFF_X1 \reg_bp_0_address[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00212_),
    .Q(reg_bp_0_address[5]),
    .QN(_06892_)
  );
  DFF_X1 \reg_bp_0_address[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00213_),
    .Q(reg_bp_0_address[6]),
    .QN(_06891_)
  );
  DFF_X1 \reg_bp_0_address[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00214_),
    .Q(reg_bp_0_address[7]),
    .QN(_06890_)
  );
  DFF_X1 \reg_bp_0_address[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00215_),
    .Q(reg_bp_0_address[8]),
    .QN(_06889_)
  );
  DFF_X1 \reg_bp_0_address[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00216_),
    .Q(reg_bp_0_address[9]),
    .QN(_06888_)
  );
  DFF_X1 \reg_bp_0_control_action$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00248_),
    .Q(reg_bp_0_control_action),
    .QN(_06857_)
  );
  DFF_X1 \reg_bp_0_control_dmode$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00249_),
    .Q(reg_bp_0_control_dmode),
    .QN(_00005_)
  );
  DFF_X1 \reg_bp_0_control_r$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00244_),
    .Q(reg_bp_0_control_r),
    .QN(_06861_)
  );
  DFF_X1 \reg_bp_0_control_tmatch[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00242_),
    .Q(reg_bp_0_control_tmatch[0]),
    .QN(_06863_)
  );
  DFF_X1 \reg_bp_0_control_tmatch[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00243_),
    .Q(reg_bp_0_control_tmatch[1]),
    .QN(_06862_)
  );
  DFF_X1 \reg_bp_0_control_w$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00245_),
    .Q(reg_bp_0_control_w),
    .QN(_06860_)
  );
  DFF_X1 \reg_bp_0_control_x$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00246_),
    .Q(reg_bp_0_control_x),
    .QN(_06859_)
  );
  DFF_X1 \reg_custom_0[3]$_SDFFE_PP1P_  (
    .CK(clock),
    .D(_00425_),
    .Q(reg_custom_0[3]),
    .QN(_06683_)
  );
  DFF_X1 \reg_dcsr_cause[0]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00285_),
    .Q(reg_dcsr_cause[0]),
    .QN(_06821_)
  );
  DFF_X1 \reg_dcsr_cause[1]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00286_),
    .Q(reg_dcsr_cause[1]),
    .QN(_06820_)
  );
  DFF_X1 \reg_dcsr_cause[2]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00287_),
    .Q(reg_dcsr_cause[2]),
    .QN(_06819_)
  );
  DFF_X1 \reg_dcsr_ebreakm$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00288_),
    .Q(reg_dcsr_ebreakm),
    .QN(_06818_)
  );
  DFF_X1 \reg_dcsr_step$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00284_),
    .Q(reg_dcsr_step),
    .QN(_06822_)
  );
  DFF_X1 \reg_debug$_SDFF_PP0_  (
    .CK(clock),
    .D(_00282_),
    .Q(reg_debug),
    .QN(_io_decode_0_read_illegal_T_15)
  );
  DFF_X1 \reg_dpc[10]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[10]),
    .Q(reg_dpc[10]),
    .QN(_07082_)
  );
  DFF_X1 \reg_dpc[11]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[11]),
    .Q(reg_dpc[11]),
    .QN(_07083_)
  );
  DFF_X1 \reg_dpc[12]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[12]),
    .Q(reg_dpc[12]),
    .QN(_07084_)
  );
  DFF_X1 \reg_dpc[13]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[13]),
    .Q(reg_dpc[13]),
    .QN(_07085_)
  );
  DFF_X1 \reg_dpc[14]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[14]),
    .Q(reg_dpc[14]),
    .QN(_07086_)
  );
  DFF_X1 \reg_dpc[15]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[15]),
    .Q(reg_dpc[15]),
    .QN(_07087_)
  );
  DFF_X1 \reg_dpc[16]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[16]),
    .Q(reg_dpc[16]),
    .QN(_07088_)
  );
  DFF_X1 \reg_dpc[17]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[17]),
    .Q(reg_dpc[17]),
    .QN(_07089_)
  );
  DFF_X1 \reg_dpc[18]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[18]),
    .Q(reg_dpc[18]),
    .QN(_07090_)
  );
  DFF_X1 \reg_dpc[19]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[19]),
    .Q(reg_dpc[19]),
    .QN(_07091_)
  );
  DFF_X1 \reg_dpc[1]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[1]),
    .Q(reg_dpc[1]),
    .QN(_T_24[1])
  );
  DFF_X1 \reg_dpc[20]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[20]),
    .Q(reg_dpc[20]),
    .QN(_07092_)
  );
  DFF_X1 \reg_dpc[21]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[21]),
    .Q(reg_dpc[21]),
    .QN(_07093_)
  );
  DFF_X1 \reg_dpc[22]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[22]),
    .Q(reg_dpc[22]),
    .QN(_07094_)
  );
  DFF_X1 \reg_dpc[23]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[23]),
    .Q(reg_dpc[23]),
    .QN(_07095_)
  );
  DFF_X1 \reg_dpc[24]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[24]),
    .Q(reg_dpc[24]),
    .QN(_07096_)
  );
  DFF_X1 \reg_dpc[25]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[25]),
    .Q(reg_dpc[25]),
    .QN(_07097_)
  );
  DFF_X1 \reg_dpc[26]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[26]),
    .Q(reg_dpc[26]),
    .QN(_07098_)
  );
  DFF_X1 \reg_dpc[27]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[27]),
    .Q(reg_dpc[27]),
    .QN(_07099_)
  );
  DFF_X1 \reg_dpc[28]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[28]),
    .Q(reg_dpc[28]),
    .QN(_07100_)
  );
  DFF_X1 \reg_dpc[29]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[29]),
    .Q(reg_dpc[29]),
    .QN(_07101_)
  );
  DFF_X1 \reg_dpc[2]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[2]),
    .Q(reg_dpc[2]),
    .QN(_07074_)
  );
  DFF_X1 \reg_dpc[30]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[30]),
    .Q(reg_dpc[30]),
    .QN(_07102_)
  );
  DFF_X1 \reg_dpc[31]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[31]),
    .Q(reg_dpc[31]),
    .QN(_06824_)
  );
  DFF_X1 \reg_dpc[3]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[3]),
    .Q(reg_dpc[3]),
    .QN(_07075_)
  );
  DFF_X1 \reg_dpc[4]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[4]),
    .Q(reg_dpc[4]),
    .QN(_07076_)
  );
  DFF_X1 \reg_dpc[5]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[5]),
    .Q(reg_dpc[5]),
    .QN(_07077_)
  );
  DFF_X1 \reg_dpc[6]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[6]),
    .Q(reg_dpc[6]),
    .QN(_07078_)
  );
  DFF_X1 \reg_dpc[7]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[7]),
    .Q(reg_dpc[7]),
    .QN(_07079_)
  );
  DFF_X1 \reg_dpc[8]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[8]),
    .Q(reg_dpc[8]),
    .QN(_07080_)
  );
  DFF_X1 \reg_dpc[9]$_DFF_P_  (
    .CK(clock),
    .D(_00000_[9]),
    .Q(reg_dpc[9]),
    .QN(_07081_)
  );
  DFF_X1 \reg_dscratch0[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00250_),
    .Q(reg_dscratch0[0]),
    .QN(_06856_)
  );
  DFF_X1 \reg_dscratch0[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00260_),
    .Q(reg_dscratch0[10]),
    .QN(_06846_)
  );
  DFF_X1 \reg_dscratch0[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00261_),
    .Q(reg_dscratch0[11]),
    .QN(_06845_)
  );
  DFF_X1 \reg_dscratch0[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00262_),
    .Q(reg_dscratch0[12]),
    .QN(_06844_)
  );
  DFF_X1 \reg_dscratch0[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00263_),
    .Q(reg_dscratch0[13]),
    .QN(_06843_)
  );
  DFF_X1 \reg_dscratch0[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00264_),
    .Q(reg_dscratch0[14]),
    .QN(_06842_)
  );
  DFF_X1 \reg_dscratch0[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00265_),
    .Q(reg_dscratch0[15]),
    .QN(_06841_)
  );
  DFF_X1 \reg_dscratch0[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00266_),
    .Q(reg_dscratch0[16]),
    .QN(_06840_)
  );
  DFF_X1 \reg_dscratch0[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00267_),
    .Q(reg_dscratch0[17]),
    .QN(_06839_)
  );
  DFF_X1 \reg_dscratch0[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00268_),
    .Q(reg_dscratch0[18]),
    .QN(_06838_)
  );
  DFF_X1 \reg_dscratch0[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00269_),
    .Q(reg_dscratch0[19]),
    .QN(_06837_)
  );
  DFF_X1 \reg_dscratch0[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00251_),
    .Q(reg_dscratch0[1]),
    .QN(_06855_)
  );
  DFF_X1 \reg_dscratch0[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00270_),
    .Q(reg_dscratch0[20]),
    .QN(_06836_)
  );
  DFF_X1 \reg_dscratch0[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00271_),
    .Q(reg_dscratch0[21]),
    .QN(_06835_)
  );
  DFF_X1 \reg_dscratch0[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00272_),
    .Q(reg_dscratch0[22]),
    .QN(_06834_)
  );
  DFF_X1 \reg_dscratch0[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00273_),
    .Q(reg_dscratch0[23]),
    .QN(_06833_)
  );
  DFF_X1 \reg_dscratch0[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00274_),
    .Q(reg_dscratch0[24]),
    .QN(_06832_)
  );
  DFF_X1 \reg_dscratch0[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00275_),
    .Q(reg_dscratch0[25]),
    .QN(_06831_)
  );
  DFF_X1 \reg_dscratch0[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00276_),
    .Q(reg_dscratch0[26]),
    .QN(_06830_)
  );
  DFF_X1 \reg_dscratch0[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00277_),
    .Q(reg_dscratch0[27]),
    .QN(_06829_)
  );
  DFF_X1 \reg_dscratch0[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00278_),
    .Q(reg_dscratch0[28]),
    .QN(_06828_)
  );
  DFF_X1 \reg_dscratch0[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00279_),
    .Q(reg_dscratch0[29]),
    .QN(_06827_)
  );
  DFF_X1 \reg_dscratch0[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00252_),
    .Q(reg_dscratch0[2]),
    .QN(_06854_)
  );
  DFF_X1 \reg_dscratch0[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00280_),
    .Q(reg_dscratch0[30]),
    .QN(_06826_)
  );
  DFF_X1 \reg_dscratch0[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00281_),
    .Q(reg_dscratch0[31]),
    .QN(_06825_)
  );
  DFF_X1 \reg_dscratch0[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00253_),
    .Q(reg_dscratch0[3]),
    .QN(_06853_)
  );
  DFF_X1 \reg_dscratch0[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00254_),
    .Q(reg_dscratch0[4]),
    .QN(_06852_)
  );
  DFF_X1 \reg_dscratch0[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00255_),
    .Q(reg_dscratch0[5]),
    .QN(_06851_)
  );
  DFF_X1 \reg_dscratch0[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00256_),
    .Q(reg_dscratch0[6]),
    .QN(_06850_)
  );
  DFF_X1 \reg_dscratch0[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00257_),
    .Q(reg_dscratch0[7]),
    .QN(_06849_)
  );
  DFF_X1 \reg_dscratch0[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00258_),
    .Q(reg_dscratch0[8]),
    .QN(_06848_)
  );
  DFF_X1 \reg_dscratch0[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00259_),
    .Q(reg_dscratch0[9]),
    .QN(_06847_)
  );
  DFF_X1 \reg_mcause[0]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00498_),
    .Q(reg_mcause[0]),
    .QN(_06612_)
  );
  DFF_X1 \reg_mcause[10]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00508_),
    .Q(reg_mcause[10]),
    .QN(_06602_)
  );
  DFF_X1 \reg_mcause[11]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00509_),
    .Q(reg_mcause[11]),
    .QN(_06601_)
  );
  DFF_X1 \reg_mcause[12]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00510_),
    .Q(reg_mcause[12]),
    .QN(_06600_)
  );
  DFF_X1 \reg_mcause[13]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00511_),
    .Q(reg_mcause[13]),
    .QN(_06599_)
  );
  DFF_X1 \reg_mcause[14]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00512_),
    .Q(reg_mcause[14]),
    .QN(_06598_)
  );
  DFF_X1 \reg_mcause[15]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00513_),
    .Q(reg_mcause[15]),
    .QN(_06597_)
  );
  DFF_X1 \reg_mcause[16]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00514_),
    .Q(reg_mcause[16]),
    .QN(_06596_)
  );
  DFF_X1 \reg_mcause[17]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00515_),
    .Q(reg_mcause[17]),
    .QN(_06595_)
  );
  DFF_X1 \reg_mcause[18]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00516_),
    .Q(reg_mcause[18]),
    .QN(_06594_)
  );
  DFF_X1 \reg_mcause[19]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00517_),
    .Q(reg_mcause[19]),
    .QN(_06593_)
  );
  DFF_X1 \reg_mcause[1]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00499_),
    .Q(reg_mcause[1]),
    .QN(_06611_)
  );
  DFF_X1 \reg_mcause[20]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00518_),
    .Q(reg_mcause[20]),
    .QN(_06592_)
  );
  DFF_X1 \reg_mcause[21]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00519_),
    .Q(reg_mcause[21]),
    .QN(_06591_)
  );
  DFF_X1 \reg_mcause[22]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00520_),
    .Q(reg_mcause[22]),
    .QN(_06590_)
  );
  DFF_X1 \reg_mcause[23]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00521_),
    .Q(reg_mcause[23]),
    .QN(_06589_)
  );
  DFF_X1 \reg_mcause[24]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00522_),
    .Q(reg_mcause[24]),
    .QN(_06588_)
  );
  DFF_X1 \reg_mcause[25]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00523_),
    .Q(reg_mcause[25]),
    .QN(_06587_)
  );
  DFF_X1 \reg_mcause[26]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00524_),
    .Q(reg_mcause[26]),
    .QN(_06586_)
  );
  DFF_X1 \reg_mcause[27]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00525_),
    .Q(reg_mcause[27]),
    .QN(_06585_)
  );
  DFF_X1 \reg_mcause[28]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00526_),
    .Q(reg_mcause[28]),
    .QN(_06584_)
  );
  DFF_X1 \reg_mcause[29]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00527_),
    .Q(reg_mcause[29]),
    .QN(_06583_)
  );
  DFF_X1 \reg_mcause[2]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00500_),
    .Q(reg_mcause[2]),
    .QN(_06610_)
  );
  DFF_X1 \reg_mcause[30]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00528_),
    .Q(reg_mcause[30]),
    .QN(_06582_)
  );
  DFF_X1 \reg_mcause[31]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00529_),
    .Q(reg_mcause[31]),
    .QN(_07103_)
  );
  DFF_X1 \reg_mcause[3]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00501_),
    .Q(reg_mcause[3]),
    .QN(_06609_)
  );
  DFF_X1 \reg_mcause[4]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00502_),
    .Q(reg_mcause[4]),
    .QN(_06608_)
  );
  DFF_X1 \reg_mcause[5]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00503_),
    .Q(reg_mcause[5]),
    .QN(_06607_)
  );
  DFF_X1 \reg_mcause[6]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00504_),
    .Q(reg_mcause[6]),
    .QN(_06606_)
  );
  DFF_X1 \reg_mcause[7]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00505_),
    .Q(reg_mcause[7]),
    .QN(_06605_)
  );
  DFF_X1 \reg_mcause[8]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00506_),
    .Q(reg_mcause[8]),
    .QN(_06604_)
  );
  DFF_X1 \reg_mcause[9]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00507_),
    .Q(reg_mcause[9]),
    .QN(_06603_)
  );
  DFF_X1 \reg_mcountinhibit[0]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00290_),
    .Q(reg_mcountinhibit[0]),
    .QN(_T_15)
  );
  DFF_X1 \reg_mcountinhibit[2]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00291_),
    .Q(reg_mcountinhibit[2]),
    .QN(_T_14)
  );
  DFF_X1 \reg_mepc[10]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[10]),
    .Q(reg_mepc[10]),
    .QN(_07144_)
  );
  DFF_X1 \reg_mepc[11]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[11]),
    .Q(reg_mepc[11]),
    .QN(_07145_)
  );
  DFF_X1 \reg_mepc[12]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[12]),
    .Q(reg_mepc[12]),
    .QN(_07146_)
  );
  DFF_X1 \reg_mepc[13]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[13]),
    .Q(reg_mepc[13]),
    .QN(_07147_)
  );
  DFF_X1 \reg_mepc[14]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[14]),
    .Q(reg_mepc[14]),
    .QN(_07148_)
  );
  DFF_X1 \reg_mepc[15]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[15]),
    .Q(reg_mepc[15]),
    .QN(_07149_)
  );
  DFF_X1 \reg_mepc[16]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[16]),
    .Q(reg_mepc[16]),
    .QN(_07150_)
  );
  DFF_X1 \reg_mepc[17]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[17]),
    .Q(reg_mepc[17]),
    .QN(_07151_)
  );
  DFF_X1 \reg_mepc[18]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[18]),
    .Q(reg_mepc[18]),
    .QN(_07152_)
  );
  DFF_X1 \reg_mepc[19]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[19]),
    .Q(reg_mepc[19]),
    .QN(_07153_)
  );
  DFF_X1 \reg_mepc[1]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[1]),
    .Q(reg_mepc[1]),
    .QN(_T_18[1])
  );
  DFF_X1 \reg_mepc[20]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[20]),
    .Q(reg_mepc[20]),
    .QN(_07154_)
  );
  DFF_X1 \reg_mepc[21]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[21]),
    .Q(reg_mepc[21]),
    .QN(_07155_)
  );
  DFF_X1 \reg_mepc[22]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[22]),
    .Q(reg_mepc[22]),
    .QN(_07156_)
  );
  DFF_X1 \reg_mepc[23]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[23]),
    .Q(reg_mepc[23]),
    .QN(_07157_)
  );
  DFF_X1 \reg_mepc[24]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[24]),
    .Q(reg_mepc[24]),
    .QN(_07158_)
  );
  DFF_X1 \reg_mepc[25]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[25]),
    .Q(reg_mepc[25]),
    .QN(_07159_)
  );
  DFF_X1 \reg_mepc[26]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[26]),
    .Q(reg_mepc[26]),
    .QN(_07160_)
  );
  DFF_X1 \reg_mepc[27]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[27]),
    .Q(reg_mepc[27]),
    .QN(_07161_)
  );
  DFF_X1 \reg_mepc[28]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[28]),
    .Q(reg_mepc[28]),
    .QN(_07162_)
  );
  DFF_X1 \reg_mepc[29]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[29]),
    .Q(reg_mepc[29]),
    .QN(_07163_)
  );
  DFF_X1 \reg_mepc[2]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[2]),
    .Q(reg_mepc[2]),
    .QN(_07136_)
  );
  DFF_X1 \reg_mepc[30]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[30]),
    .Q(reg_mepc[30]),
    .QN(_07164_)
  );
  DFF_X1 \reg_mepc[31]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[31]),
    .Q(reg_mepc[31]),
    .QN(_06581_)
  );
  DFF_X1 \reg_mepc[3]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[3]),
    .Q(reg_mepc[3]),
    .QN(_07137_)
  );
  DFF_X1 \reg_mepc[4]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[4]),
    .Q(reg_mepc[4]),
    .QN(_07138_)
  );
  DFF_X1 \reg_mepc[5]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[5]),
    .Q(reg_mepc[5]),
    .QN(_07139_)
  );
  DFF_X1 \reg_mepc[6]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[6]),
    .Q(reg_mepc[6]),
    .QN(_07140_)
  );
  DFF_X1 \reg_mepc[7]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[7]),
    .Q(reg_mepc[7]),
    .QN(_07141_)
  );
  DFF_X1 \reg_mepc[8]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[8]),
    .Q(reg_mepc[8]),
    .QN(_07142_)
  );
  DFF_X1 \reg_mepc[9]$_DFF_P_  (
    .CK(clock),
    .D(_00001_[9]),
    .Q(reg_mepc[9]),
    .QN(_07143_)
  );
  DFF_X1 \reg_mie[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00532_),
    .Q(reg_mie[11]),
    .QN(_06578_)
  );
  DFF_X1 \reg_mie[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00530_),
    .Q(reg_mie[3]),
    .QN(_06580_)
  );
  DFF_X1 \reg_mie[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00531_),
    .Q(reg_mie[7]),
    .QN(_06579_)
  );
  DFF_X1 \reg_misa[0]$_SDFFE_PP1P_  (
    .CK(clock),
    .D(_00426_),
    .Q(reg_misa[0]),
    .QN(_06682_)
  );
  DFF_X1 \reg_misa[12]$_SDFFE_PP1P_  (
    .CK(clock),
    .D(_00428_),
    .Q(reg_misa[12]),
    .QN(_06681_)
  );
  DFF_X1 \reg_misa[2]$_SDFFE_PP1P_  (
    .CK(clock),
    .D(_00427_),
    .Q(reg_misa[2]),
    .QN(_GEN_586[1])
  );
  DFF_X1 \reg_mscratch[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00332_),
    .Q(reg_mscratch[0]),
    .QN(_06776_)
  );
  DFF_X1 \reg_mscratch[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00342_),
    .Q(reg_mscratch[10]),
    .QN(_06766_)
  );
  DFF_X1 \reg_mscratch[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00343_),
    .Q(reg_mscratch[11]),
    .QN(_06765_)
  );
  DFF_X1 \reg_mscratch[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00344_),
    .Q(reg_mscratch[12]),
    .QN(_06764_)
  );
  DFF_X1 \reg_mscratch[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00345_),
    .Q(reg_mscratch[13]),
    .QN(_06763_)
  );
  DFF_X1 \reg_mscratch[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00346_),
    .Q(reg_mscratch[14]),
    .QN(_06762_)
  );
  DFF_X1 \reg_mscratch[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00347_),
    .Q(reg_mscratch[15]),
    .QN(_06761_)
  );
  DFF_X1 \reg_mscratch[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00348_),
    .Q(reg_mscratch[16]),
    .QN(_06760_)
  );
  DFF_X1 \reg_mscratch[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00349_),
    .Q(reg_mscratch[17]),
    .QN(_06759_)
  );
  DFF_X1 \reg_mscratch[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00350_),
    .Q(reg_mscratch[18]),
    .QN(_06758_)
  );
  DFF_X1 \reg_mscratch[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00351_),
    .Q(reg_mscratch[19]),
    .QN(_06757_)
  );
  DFF_X1 \reg_mscratch[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00333_),
    .Q(reg_mscratch[1]),
    .QN(_06775_)
  );
  DFF_X1 \reg_mscratch[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00352_),
    .Q(reg_mscratch[20]),
    .QN(_06756_)
  );
  DFF_X1 \reg_mscratch[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00353_),
    .Q(reg_mscratch[21]),
    .QN(_06755_)
  );
  DFF_X1 \reg_mscratch[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00354_),
    .Q(reg_mscratch[22]),
    .QN(_06754_)
  );
  DFF_X1 \reg_mscratch[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00355_),
    .Q(reg_mscratch[23]),
    .QN(_06753_)
  );
  DFF_X1 \reg_mscratch[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00356_),
    .Q(reg_mscratch[24]),
    .QN(_06752_)
  );
  DFF_X1 \reg_mscratch[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00357_),
    .Q(reg_mscratch[25]),
    .QN(_06751_)
  );
  DFF_X1 \reg_mscratch[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00358_),
    .Q(reg_mscratch[26]),
    .QN(_06750_)
  );
  DFF_X1 \reg_mscratch[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00359_),
    .Q(reg_mscratch[27]),
    .QN(_06749_)
  );
  DFF_X1 \reg_mscratch[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00360_),
    .Q(reg_mscratch[28]),
    .QN(_06748_)
  );
  DFF_X1 \reg_mscratch[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00361_),
    .Q(reg_mscratch[29]),
    .QN(_06747_)
  );
  DFF_X1 \reg_mscratch[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00334_),
    .Q(reg_mscratch[2]),
    .QN(_06774_)
  );
  DFF_X1 \reg_mscratch[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00362_),
    .Q(reg_mscratch[30]),
    .QN(_06746_)
  );
  DFF_X1 \reg_mscratch[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00363_),
    .Q(reg_mscratch[31]),
    .QN(_06745_)
  );
  DFF_X1 \reg_mscratch[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00335_),
    .Q(reg_mscratch[3]),
    .QN(_06773_)
  );
  DFF_X1 \reg_mscratch[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00336_),
    .Q(reg_mscratch[4]),
    .QN(_06772_)
  );
  DFF_X1 \reg_mscratch[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00337_),
    .Q(reg_mscratch[5]),
    .QN(_06771_)
  );
  DFF_X1 \reg_mscratch[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00338_),
    .Q(reg_mscratch[6]),
    .QN(_06770_)
  );
  DFF_X1 \reg_mscratch[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00339_),
    .Q(reg_mscratch[7]),
    .QN(_06769_)
  );
  DFF_X1 \reg_mscratch[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00340_),
    .Q(reg_mscratch[8]),
    .QN(_06768_)
  );
  DFF_X1 \reg_mscratch[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00341_),
    .Q(reg_mscratch[9]),
    .QN(_06767_)
  );
  DFF_X1 \reg_mstatus_gva$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00293_),
    .Q(reg_mstatus_gva),
    .QN(_06815_)
  );
  DFF_X1 \reg_mstatus_mie$_SDFF_PP0_  (
    .CK(clock),
    .D(_00283_),
    .Q(reg_mstatus_mie),
    .QN(_06823_)
  );
  DFF_X1 \reg_mstatus_mpie$_SDFF_PP0_  (
    .CK(clock),
    .D(_00289_),
    .Q(reg_mstatus_mpie),
    .QN(_06817_)
  );
  DFF_X1 \reg_mtval[0]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[0]),
    .Q(reg_mtval[0]),
    .QN(_07104_)
  );
  DFF_X1 \reg_mtval[10]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[10]),
    .Q(reg_mtval[10]),
    .QN(_07114_)
  );
  DFF_X1 \reg_mtval[11]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[11]),
    .Q(reg_mtval[11]),
    .QN(_07115_)
  );
  DFF_X1 \reg_mtval[12]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[12]),
    .Q(reg_mtval[12]),
    .QN(_07116_)
  );
  DFF_X1 \reg_mtval[13]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[13]),
    .Q(reg_mtval[13]),
    .QN(_07117_)
  );
  DFF_X1 \reg_mtval[14]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[14]),
    .Q(reg_mtval[14]),
    .QN(_07118_)
  );
  DFF_X1 \reg_mtval[15]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[15]),
    .Q(reg_mtval[15]),
    .QN(_07119_)
  );
  DFF_X1 \reg_mtval[16]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[16]),
    .Q(reg_mtval[16]),
    .QN(_07120_)
  );
  DFF_X1 \reg_mtval[17]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[17]),
    .Q(reg_mtval[17]),
    .QN(_07121_)
  );
  DFF_X1 \reg_mtval[18]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[18]),
    .Q(reg_mtval[18]),
    .QN(_07122_)
  );
  DFF_X1 \reg_mtval[19]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[19]),
    .Q(reg_mtval[19]),
    .QN(_07123_)
  );
  DFF_X1 \reg_mtval[1]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[1]),
    .Q(reg_mtval[1]),
    .QN(_07105_)
  );
  DFF_X1 \reg_mtval[20]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[20]),
    .Q(reg_mtval[20]),
    .QN(_07124_)
  );
  DFF_X1 \reg_mtval[21]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[21]),
    .Q(reg_mtval[21]),
    .QN(_07125_)
  );
  DFF_X1 \reg_mtval[22]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[22]),
    .Q(reg_mtval[22]),
    .QN(_07126_)
  );
  DFF_X1 \reg_mtval[23]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[23]),
    .Q(reg_mtval[23]),
    .QN(_07127_)
  );
  DFF_X1 \reg_mtval[24]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[24]),
    .Q(reg_mtval[24]),
    .QN(_07128_)
  );
  DFF_X1 \reg_mtval[25]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[25]),
    .Q(reg_mtval[25]),
    .QN(_07129_)
  );
  DFF_X1 \reg_mtval[26]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[26]),
    .Q(reg_mtval[26]),
    .QN(_07130_)
  );
  DFF_X1 \reg_mtval[27]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[27]),
    .Q(reg_mtval[27]),
    .QN(_07131_)
  );
  DFF_X1 \reg_mtval[28]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[28]),
    .Q(reg_mtval[28]),
    .QN(_07132_)
  );
  DFF_X1 \reg_mtval[29]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[29]),
    .Q(reg_mtval[29]),
    .QN(_07133_)
  );
  DFF_X1 \reg_mtval[2]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[2]),
    .Q(reg_mtval[2]),
    .QN(_07106_)
  );
  DFF_X1 \reg_mtval[30]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[30]),
    .Q(reg_mtval[30]),
    .QN(_07134_)
  );
  DFF_X1 \reg_mtval[31]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[31]),
    .Q(reg_mtval[31]),
    .QN(_07135_)
  );
  DFF_X1 \reg_mtval[3]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[3]),
    .Q(reg_mtval[3]),
    .QN(_07107_)
  );
  DFF_X1 \reg_mtval[4]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[4]),
    .Q(reg_mtval[4]),
    .QN(_07108_)
  );
  DFF_X1 \reg_mtval[5]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[5]),
    .Q(reg_mtval[5]),
    .QN(_07109_)
  );
  DFF_X1 \reg_mtval[6]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[6]),
    .Q(reg_mtval[6]),
    .QN(_07110_)
  );
  DFF_X1 \reg_mtval[7]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[7]),
    .Q(reg_mtval[7]),
    .QN(_07111_)
  );
  DFF_X1 \reg_mtval[8]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[8]),
    .Q(reg_mtval[8]),
    .QN(_07112_)
  );
  DFF_X1 \reg_mtval[9]$_DFF_P_  (
    .CK(clock),
    .D(_00002_[9]),
    .Q(reg_mtval[9]),
    .QN(_07113_)
  );
  DFF_X1 \reg_mtvec[0]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00467_),
    .Q(reg_mtvec[0]),
    .QN(_read_mtvec_T_4[6])
  );
  DFF_X1 \reg_mtvec[10]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00476_),
    .Q(reg_mtvec[10]),
    .QN(_06634_)
  );
  DFF_X1 \reg_mtvec[11]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00477_),
    .Q(reg_mtvec[11]),
    .QN(_06633_)
  );
  DFF_X1 \reg_mtvec[12]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00478_),
    .Q(reg_mtvec[12]),
    .QN(_06632_)
  );
  DFF_X1 \reg_mtvec[13]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00479_),
    .Q(reg_mtvec[13]),
    .QN(_06631_)
  );
  DFF_X1 \reg_mtvec[14]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00480_),
    .Q(reg_mtvec[14]),
    .QN(_06630_)
  );
  DFF_X1 \reg_mtvec[15]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00481_),
    .Q(reg_mtvec[15]),
    .QN(_06629_)
  );
  DFF_X1 \reg_mtvec[16]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00482_),
    .Q(reg_mtvec[16]),
    .QN(_06628_)
  );
  DFF_X1 \reg_mtvec[17]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00483_),
    .Q(reg_mtvec[17]),
    .QN(_06627_)
  );
  DFF_X1 \reg_mtvec[18]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00484_),
    .Q(reg_mtvec[18]),
    .QN(_06626_)
  );
  DFF_X1 \reg_mtvec[19]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00485_),
    .Q(reg_mtvec[19]),
    .QN(_06625_)
  );
  DFF_X1 \reg_mtvec[20]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00486_),
    .Q(reg_mtvec[20]),
    .QN(_06624_)
  );
  DFF_X1 \reg_mtvec[21]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00487_),
    .Q(reg_mtvec[21]),
    .QN(_06623_)
  );
  DFF_X1 \reg_mtvec[22]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00488_),
    .Q(reg_mtvec[22]),
    .QN(_06622_)
  );
  DFF_X1 \reg_mtvec[23]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00489_),
    .Q(reg_mtvec[23]),
    .QN(_06621_)
  );
  DFF_X1 \reg_mtvec[24]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00490_),
    .Q(reg_mtvec[24]),
    .QN(_06620_)
  );
  DFF_X1 \reg_mtvec[25]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00491_),
    .Q(reg_mtvec[25]),
    .QN(_06619_)
  );
  DFF_X1 \reg_mtvec[26]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00492_),
    .Q(reg_mtvec[26]),
    .QN(_06618_)
  );
  DFF_X1 \reg_mtvec[27]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00493_),
    .Q(reg_mtvec[27]),
    .QN(_06617_)
  );
  DFF_X1 \reg_mtvec[28]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00494_),
    .Q(reg_mtvec[28]),
    .QN(_06616_)
  );
  DFF_X1 \reg_mtvec[29]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00495_),
    .Q(reg_mtvec[29]),
    .QN(_06615_)
  );
  DFF_X1 \reg_mtvec[2]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00468_),
    .Q(reg_mtvec[2]),
    .QN(_06642_)
  );
  DFF_X1 \reg_mtvec[30]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00496_),
    .Q(reg_mtvec[30]),
    .QN(_06614_)
  );
  DFF_X1 \reg_mtvec[31]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00497_),
    .Q(reg_mtvec[31]),
    .QN(_06613_)
  );
  DFF_X1 \reg_mtvec[3]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00469_),
    .Q(reg_mtvec[3]),
    .QN(_06641_)
  );
  DFF_X1 \reg_mtvec[4]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00470_),
    .Q(reg_mtvec[4]),
    .QN(_06640_)
  );
  DFF_X1 \reg_mtvec[5]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00471_),
    .Q(reg_mtvec[5]),
    .QN(_06639_)
  );
  DFF_X1 \reg_mtvec[6]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00472_),
    .Q(reg_mtvec[6]),
    .QN(_06638_)
  );
  DFF_X1 \reg_mtvec[7]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00473_),
    .Q(reg_mtvec[7]),
    .QN(_06637_)
  );
  DFF_X1 \reg_mtvec[8]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00474_),
    .Q(reg_mtvec[8]),
    .QN(_06636_)
  );
  DFF_X1 \reg_mtvec[9]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00475_),
    .Q(reg_mtvec[9]),
    .QN(_06635_)
  );
  DFF_X1 \reg_pmp_0_addr[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00176_),
    .Q(reg_pmp_0_addr[0]),
    .QN(_06928_)
  );
  DFF_X1 \reg_pmp_0_addr[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00186_),
    .Q(reg_pmp_0_addr[10]),
    .QN(_06918_)
  );
  DFF_X1 \reg_pmp_0_addr[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00187_),
    .Q(reg_pmp_0_addr[11]),
    .QN(_06917_)
  );
  DFF_X1 \reg_pmp_0_addr[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00188_),
    .Q(reg_pmp_0_addr[12]),
    .QN(_06916_)
  );
  DFF_X1 \reg_pmp_0_addr[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00189_),
    .Q(reg_pmp_0_addr[13]),
    .QN(_06915_)
  );
  DFF_X1 \reg_pmp_0_addr[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00190_),
    .Q(reg_pmp_0_addr[14]),
    .QN(_06914_)
  );
  DFF_X1 \reg_pmp_0_addr[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00191_),
    .Q(reg_pmp_0_addr[15]),
    .QN(_06913_)
  );
  DFF_X1 \reg_pmp_0_addr[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00192_),
    .Q(reg_pmp_0_addr[16]),
    .QN(_06912_)
  );
  DFF_X1 \reg_pmp_0_addr[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00193_),
    .Q(reg_pmp_0_addr[17]),
    .QN(_06911_)
  );
  DFF_X1 \reg_pmp_0_addr[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00194_),
    .Q(reg_pmp_0_addr[18]),
    .QN(_06910_)
  );
  DFF_X1 \reg_pmp_0_addr[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00195_),
    .Q(reg_pmp_0_addr[19]),
    .QN(_06909_)
  );
  DFF_X1 \reg_pmp_0_addr[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00177_),
    .Q(reg_pmp_0_addr[1]),
    .QN(_06927_)
  );
  DFF_X1 \reg_pmp_0_addr[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00196_),
    .Q(reg_pmp_0_addr[20]),
    .QN(_06908_)
  );
  DFF_X1 \reg_pmp_0_addr[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00197_),
    .Q(reg_pmp_0_addr[21]),
    .QN(_06907_)
  );
  DFF_X1 \reg_pmp_0_addr[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00198_),
    .Q(reg_pmp_0_addr[22]),
    .QN(_06906_)
  );
  DFF_X1 \reg_pmp_0_addr[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00199_),
    .Q(reg_pmp_0_addr[23]),
    .QN(_06905_)
  );
  DFF_X1 \reg_pmp_0_addr[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00200_),
    .Q(reg_pmp_0_addr[24]),
    .QN(_06904_)
  );
  DFF_X1 \reg_pmp_0_addr[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00201_),
    .Q(reg_pmp_0_addr[25]),
    .QN(_06903_)
  );
  DFF_X1 \reg_pmp_0_addr[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00202_),
    .Q(reg_pmp_0_addr[26]),
    .QN(_06902_)
  );
  DFF_X1 \reg_pmp_0_addr[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00203_),
    .Q(reg_pmp_0_addr[27]),
    .QN(_06901_)
  );
  DFF_X1 \reg_pmp_0_addr[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00204_),
    .Q(reg_pmp_0_addr[28]),
    .QN(_06900_)
  );
  DFF_X1 \reg_pmp_0_addr[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00205_),
    .Q(reg_pmp_0_addr[29]),
    .QN(_06899_)
  );
  DFF_X1 \reg_pmp_0_addr[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00178_),
    .Q(reg_pmp_0_addr[2]),
    .QN(_06926_)
  );
  DFF_X1 \reg_pmp_0_addr[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00179_),
    .Q(reg_pmp_0_addr[3]),
    .QN(_06925_)
  );
  DFF_X1 \reg_pmp_0_addr[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00180_),
    .Q(reg_pmp_0_addr[4]),
    .QN(_06924_)
  );
  DFF_X1 \reg_pmp_0_addr[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00181_),
    .Q(reg_pmp_0_addr[5]),
    .QN(_06923_)
  );
  DFF_X1 \reg_pmp_0_addr[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00182_),
    .Q(reg_pmp_0_addr[6]),
    .QN(_06922_)
  );
  DFF_X1 \reg_pmp_0_addr[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00183_),
    .Q(reg_pmp_0_addr[7]),
    .QN(_06921_)
  );
  DFF_X1 \reg_pmp_0_addr[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00184_),
    .Q(reg_pmp_0_addr[8]),
    .QN(_06920_)
  );
  DFF_X1 \reg_pmp_0_addr[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00185_),
    .Q(reg_pmp_0_addr[9]),
    .QN(_06919_)
  );
  DFF_X1 \reg_pmp_0_cfg_a[0]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00239_),
    .Q(reg_pmp_0_cfg_a[0]),
    .QN(_06865_)
  );
  DFF_X1 \reg_pmp_0_cfg_a[1]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00240_),
    .Q(reg_pmp_0_cfg_a[1]),
    .QN(_06864_)
  );
  DFF_X1 \reg_pmp_0_cfg_l$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00241_),
    .Q(reg_pmp_0_cfg_l),
    .QN(_00006_)
  );
  DFF_X1 \reg_pmp_0_cfg_r$_DFFE_PP_  (
    .CK(clock),
    .D(_00175_),
    .Q(reg_pmp_0_cfg_r),
    .QN(_06929_)
  );
  DFF_X1 \reg_pmp_0_cfg_w$_DFFE_PP_  (
    .CK(clock),
    .D(_00057_),
    .Q(reg_pmp_0_cfg_w),
    .QN(_07037_)
  );
  DFF_X1 \reg_pmp_0_cfg_x$_DFFE_PP_  (
    .CK(clock),
    .D(_00206_),
    .Q(reg_pmp_0_cfg_x),
    .QN(_06898_)
  );
  DFF_X1 \reg_pmp_1_addr[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00365_),
    .Q(reg_pmp_1_addr[0]),
    .QN(_06743_)
  );
  DFF_X1 \reg_pmp_1_addr[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00375_),
    .Q(reg_pmp_1_addr[10]),
    .QN(_06733_)
  );
  DFF_X1 \reg_pmp_1_addr[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00376_),
    .Q(reg_pmp_1_addr[11]),
    .QN(_06732_)
  );
  DFF_X1 \reg_pmp_1_addr[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00377_),
    .Q(reg_pmp_1_addr[12]),
    .QN(_06731_)
  );
  DFF_X1 \reg_pmp_1_addr[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00378_),
    .Q(reg_pmp_1_addr[13]),
    .QN(_06730_)
  );
  DFF_X1 \reg_pmp_1_addr[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00379_),
    .Q(reg_pmp_1_addr[14]),
    .QN(_06729_)
  );
  DFF_X1 \reg_pmp_1_addr[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00380_),
    .Q(reg_pmp_1_addr[15]),
    .QN(_06728_)
  );
  DFF_X1 \reg_pmp_1_addr[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00381_),
    .Q(reg_pmp_1_addr[16]),
    .QN(_06727_)
  );
  DFF_X1 \reg_pmp_1_addr[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00382_),
    .Q(reg_pmp_1_addr[17]),
    .QN(_06726_)
  );
  DFF_X1 \reg_pmp_1_addr[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00383_),
    .Q(reg_pmp_1_addr[18]),
    .QN(_06725_)
  );
  DFF_X1 \reg_pmp_1_addr[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00384_),
    .Q(reg_pmp_1_addr[19]),
    .QN(_06724_)
  );
  DFF_X1 \reg_pmp_1_addr[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00366_),
    .Q(reg_pmp_1_addr[1]),
    .QN(_06742_)
  );
  DFF_X1 \reg_pmp_1_addr[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00385_),
    .Q(reg_pmp_1_addr[20]),
    .QN(_06723_)
  );
  DFF_X1 \reg_pmp_1_addr[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00386_),
    .Q(reg_pmp_1_addr[21]),
    .QN(_06722_)
  );
  DFF_X1 \reg_pmp_1_addr[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00387_),
    .Q(reg_pmp_1_addr[22]),
    .QN(_06721_)
  );
  DFF_X1 \reg_pmp_1_addr[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00388_),
    .Q(reg_pmp_1_addr[23]),
    .QN(_06720_)
  );
  DFF_X1 \reg_pmp_1_addr[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00389_),
    .Q(reg_pmp_1_addr[24]),
    .QN(_06719_)
  );
  DFF_X1 \reg_pmp_1_addr[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00390_),
    .Q(reg_pmp_1_addr[25]),
    .QN(_06718_)
  );
  DFF_X1 \reg_pmp_1_addr[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00391_),
    .Q(reg_pmp_1_addr[26]),
    .QN(_06717_)
  );
  DFF_X1 \reg_pmp_1_addr[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00392_),
    .Q(reg_pmp_1_addr[27]),
    .QN(_06716_)
  );
  DFF_X1 \reg_pmp_1_addr[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00393_),
    .Q(reg_pmp_1_addr[28]),
    .QN(_06715_)
  );
  DFF_X1 \reg_pmp_1_addr[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00394_),
    .Q(reg_pmp_1_addr[29]),
    .QN(_06714_)
  );
  DFF_X1 \reg_pmp_1_addr[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00367_),
    .Q(reg_pmp_1_addr[2]),
    .QN(_06741_)
  );
  DFF_X1 \reg_pmp_1_addr[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00368_),
    .Q(reg_pmp_1_addr[3]),
    .QN(_06740_)
  );
  DFF_X1 \reg_pmp_1_addr[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00369_),
    .Q(reg_pmp_1_addr[4]),
    .QN(_06739_)
  );
  DFF_X1 \reg_pmp_1_addr[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00370_),
    .Q(reg_pmp_1_addr[5]),
    .QN(_06738_)
  );
  DFF_X1 \reg_pmp_1_addr[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00371_),
    .Q(reg_pmp_1_addr[6]),
    .QN(_06737_)
  );
  DFF_X1 \reg_pmp_1_addr[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00372_),
    .Q(reg_pmp_1_addr[7]),
    .QN(_06736_)
  );
  DFF_X1 \reg_pmp_1_addr[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00373_),
    .Q(reg_pmp_1_addr[8]),
    .QN(_06735_)
  );
  DFF_X1 \reg_pmp_1_addr[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00374_),
    .Q(reg_pmp_1_addr[9]),
    .QN(_06734_)
  );
  DFF_X1 \reg_pmp_1_cfg_a[0]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00172_),
    .Q(reg_pmp_1_cfg_a[0]),
    .QN(_06930_)
  );
  DFF_X1 \reg_pmp_1_cfg_a[1]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00173_),
    .Q(reg_pmp_1_cfg_a[1]),
    .QN(_00008_)
  );
  DFF_X1 \reg_pmp_1_cfg_l$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00174_),
    .Q(reg_pmp_1_cfg_l),
    .QN(_00007_)
  );
  DFF_X1 \reg_pmp_1_cfg_r$_DFFE_PP_  (
    .CK(clock),
    .D(_00168_),
    .Q(reg_pmp_1_cfg_r),
    .QN(_06934_)
  );
  DFF_X1 \reg_pmp_1_cfg_w$_DFFE_PP_  (
    .CK(clock),
    .D(_00133_),
    .Q(reg_pmp_1_cfg_w),
    .QN(_06967_)
  );
  DFF_X1 \reg_pmp_1_cfg_x$_DFFE_PP_  (
    .CK(clock),
    .D(_00170_),
    .Q(reg_pmp_1_cfg_x),
    .QN(_06932_)
  );
  DFF_X1 \reg_pmp_2_addr[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00103_),
    .Q(reg_pmp_2_addr[0]),
    .QN(_06997_)
  );
  DFF_X1 \reg_pmp_2_addr[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00113_),
    .Q(reg_pmp_2_addr[10]),
    .QN(_06987_)
  );
  DFF_X1 \reg_pmp_2_addr[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00114_),
    .Q(reg_pmp_2_addr[11]),
    .QN(_06986_)
  );
  DFF_X1 \reg_pmp_2_addr[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00115_),
    .Q(reg_pmp_2_addr[12]),
    .QN(_06985_)
  );
  DFF_X1 \reg_pmp_2_addr[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00116_),
    .Q(reg_pmp_2_addr[13]),
    .QN(_06984_)
  );
  DFF_X1 \reg_pmp_2_addr[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00117_),
    .Q(reg_pmp_2_addr[14]),
    .QN(_06983_)
  );
  DFF_X1 \reg_pmp_2_addr[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00118_),
    .Q(reg_pmp_2_addr[15]),
    .QN(_06982_)
  );
  DFF_X1 \reg_pmp_2_addr[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00119_),
    .Q(reg_pmp_2_addr[16]),
    .QN(_06981_)
  );
  DFF_X1 \reg_pmp_2_addr[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00120_),
    .Q(reg_pmp_2_addr[17]),
    .QN(_06980_)
  );
  DFF_X1 \reg_pmp_2_addr[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00121_),
    .Q(reg_pmp_2_addr[18]),
    .QN(_06979_)
  );
  DFF_X1 \reg_pmp_2_addr[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00122_),
    .Q(reg_pmp_2_addr[19]),
    .QN(_06978_)
  );
  DFF_X1 \reg_pmp_2_addr[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00104_),
    .Q(reg_pmp_2_addr[1]),
    .QN(_06996_)
  );
  DFF_X1 \reg_pmp_2_addr[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00123_),
    .Q(reg_pmp_2_addr[20]),
    .QN(_06977_)
  );
  DFF_X1 \reg_pmp_2_addr[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00124_),
    .Q(reg_pmp_2_addr[21]),
    .QN(_06976_)
  );
  DFF_X1 \reg_pmp_2_addr[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00125_),
    .Q(reg_pmp_2_addr[22]),
    .QN(_06975_)
  );
  DFF_X1 \reg_pmp_2_addr[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00126_),
    .Q(reg_pmp_2_addr[23]),
    .QN(_06974_)
  );
  DFF_X1 \reg_pmp_2_addr[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00127_),
    .Q(reg_pmp_2_addr[24]),
    .QN(_06973_)
  );
  DFF_X1 \reg_pmp_2_addr[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00128_),
    .Q(reg_pmp_2_addr[25]),
    .QN(_06972_)
  );
  DFF_X1 \reg_pmp_2_addr[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00129_),
    .Q(reg_pmp_2_addr[26]),
    .QN(_06971_)
  );
  DFF_X1 \reg_pmp_2_addr[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00130_),
    .Q(reg_pmp_2_addr[27]),
    .QN(_06970_)
  );
  DFF_X1 \reg_pmp_2_addr[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00131_),
    .Q(reg_pmp_2_addr[28]),
    .QN(_06969_)
  );
  DFF_X1 \reg_pmp_2_addr[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00132_),
    .Q(reg_pmp_2_addr[29]),
    .QN(_06968_)
  );
  DFF_X1 \reg_pmp_2_addr[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00105_),
    .Q(reg_pmp_2_addr[2]),
    .QN(_06995_)
  );
  DFF_X1 \reg_pmp_2_addr[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00106_),
    .Q(reg_pmp_2_addr[3]),
    .QN(_06994_)
  );
  DFF_X1 \reg_pmp_2_addr[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00107_),
    .Q(reg_pmp_2_addr[4]),
    .QN(_06993_)
  );
  DFF_X1 \reg_pmp_2_addr[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00108_),
    .Q(reg_pmp_2_addr[5]),
    .QN(_06992_)
  );
  DFF_X1 \reg_pmp_2_addr[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00109_),
    .Q(reg_pmp_2_addr[6]),
    .QN(_06991_)
  );
  DFF_X1 \reg_pmp_2_addr[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00110_),
    .Q(reg_pmp_2_addr[7]),
    .QN(_06990_)
  );
  DFF_X1 \reg_pmp_2_addr[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00111_),
    .Q(reg_pmp_2_addr[8]),
    .QN(_06989_)
  );
  DFF_X1 \reg_pmp_2_addr[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00112_),
    .Q(reg_pmp_2_addr[9]),
    .QN(_06988_)
  );
  DFF_X1 \reg_pmp_2_cfg_a[0]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00165_),
    .Q(reg_pmp_2_cfg_a[0]),
    .QN(_06935_)
  );
  DFF_X1 \reg_pmp_2_cfg_a[1]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00166_),
    .Q(reg_pmp_2_cfg_a[1]),
    .QN(_00010_)
  );
  DFF_X1 \reg_pmp_2_cfg_l$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00167_),
    .Q(reg_pmp_2_cfg_l),
    .QN(_00009_)
  );
  DFF_X1 \reg_pmp_2_cfg_r$_DFFE_PP_  (
    .CK(clock),
    .D(_00134_),
    .Q(reg_pmp_2_cfg_r),
    .QN(_06966_)
  );
  DFF_X1 \reg_pmp_2_cfg_w$_DFFE_PP_  (
    .CK(clock),
    .D(_00099_),
    .Q(reg_pmp_2_cfg_w),
    .QN(_06999_)
  );
  DFF_X1 \reg_pmp_2_cfg_x$_DFFE_PP_  (
    .CK(clock),
    .D(_00171_),
    .Q(reg_pmp_2_cfg_x),
    .QN(_06931_)
  );
  DFF_X1 \reg_pmp_3_addr[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00135_),
    .Q(reg_pmp_3_addr[0]),
    .QN(_06965_)
  );
  DFF_X1 \reg_pmp_3_addr[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00145_),
    .Q(reg_pmp_3_addr[10]),
    .QN(_06955_)
  );
  DFF_X1 \reg_pmp_3_addr[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00146_),
    .Q(reg_pmp_3_addr[11]),
    .QN(_06954_)
  );
  DFF_X1 \reg_pmp_3_addr[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00147_),
    .Q(reg_pmp_3_addr[12]),
    .QN(_06953_)
  );
  DFF_X1 \reg_pmp_3_addr[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00148_),
    .Q(reg_pmp_3_addr[13]),
    .QN(_06952_)
  );
  DFF_X1 \reg_pmp_3_addr[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00149_),
    .Q(reg_pmp_3_addr[14]),
    .QN(_06951_)
  );
  DFF_X1 \reg_pmp_3_addr[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00150_),
    .Q(reg_pmp_3_addr[15]),
    .QN(_06950_)
  );
  DFF_X1 \reg_pmp_3_addr[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00151_),
    .Q(reg_pmp_3_addr[16]),
    .QN(_06949_)
  );
  DFF_X1 \reg_pmp_3_addr[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00152_),
    .Q(reg_pmp_3_addr[17]),
    .QN(_06948_)
  );
  DFF_X1 \reg_pmp_3_addr[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00153_),
    .Q(reg_pmp_3_addr[18]),
    .QN(_06947_)
  );
  DFF_X1 \reg_pmp_3_addr[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00154_),
    .Q(reg_pmp_3_addr[19]),
    .QN(_06946_)
  );
  DFF_X1 \reg_pmp_3_addr[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00136_),
    .Q(reg_pmp_3_addr[1]),
    .QN(_06964_)
  );
  DFF_X1 \reg_pmp_3_addr[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00155_),
    .Q(reg_pmp_3_addr[20]),
    .QN(_06945_)
  );
  DFF_X1 \reg_pmp_3_addr[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00156_),
    .Q(reg_pmp_3_addr[21]),
    .QN(_06944_)
  );
  DFF_X1 \reg_pmp_3_addr[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00157_),
    .Q(reg_pmp_3_addr[22]),
    .QN(_06943_)
  );
  DFF_X1 \reg_pmp_3_addr[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00158_),
    .Q(reg_pmp_3_addr[23]),
    .QN(_06942_)
  );
  DFF_X1 \reg_pmp_3_addr[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00159_),
    .Q(reg_pmp_3_addr[24]),
    .QN(_06941_)
  );
  DFF_X1 \reg_pmp_3_addr[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00160_),
    .Q(reg_pmp_3_addr[25]),
    .QN(_06940_)
  );
  DFF_X1 \reg_pmp_3_addr[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00161_),
    .Q(reg_pmp_3_addr[26]),
    .QN(_06939_)
  );
  DFF_X1 \reg_pmp_3_addr[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00162_),
    .Q(reg_pmp_3_addr[27]),
    .QN(_06938_)
  );
  DFF_X1 \reg_pmp_3_addr[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00163_),
    .Q(reg_pmp_3_addr[28]),
    .QN(_06937_)
  );
  DFF_X1 \reg_pmp_3_addr[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00164_),
    .Q(reg_pmp_3_addr[29]),
    .QN(_06936_)
  );
  DFF_X1 \reg_pmp_3_addr[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00137_),
    .Q(reg_pmp_3_addr[2]),
    .QN(_06963_)
  );
  DFF_X1 \reg_pmp_3_addr[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00138_),
    .Q(reg_pmp_3_addr[3]),
    .QN(_06962_)
  );
  DFF_X1 \reg_pmp_3_addr[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00139_),
    .Q(reg_pmp_3_addr[4]),
    .QN(_06961_)
  );
  DFF_X1 \reg_pmp_3_addr[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00140_),
    .Q(reg_pmp_3_addr[5]),
    .QN(_06960_)
  );
  DFF_X1 \reg_pmp_3_addr[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00141_),
    .Q(reg_pmp_3_addr[6]),
    .QN(_06959_)
  );
  DFF_X1 \reg_pmp_3_addr[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00142_),
    .Q(reg_pmp_3_addr[7]),
    .QN(_06958_)
  );
  DFF_X1 \reg_pmp_3_addr[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00143_),
    .Q(reg_pmp_3_addr[8]),
    .QN(_06957_)
  );
  DFF_X1 \reg_pmp_3_addr[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00144_),
    .Q(reg_pmp_3_addr[9]),
    .QN(_06956_)
  );
  DFF_X1 \reg_pmp_3_cfg_a[0]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00100_),
    .Q(reg_pmp_3_cfg_a[0]),
    .QN(_06998_)
  );
  DFF_X1 \reg_pmp_3_cfg_a[1]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00101_),
    .Q(reg_pmp_3_cfg_a[1]),
    .QN(_00012_)
  );
  DFF_X1 \reg_pmp_3_cfg_l$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00102_),
    .Q(reg_pmp_3_cfg_l),
    .QN(_00011_)
  );
  DFF_X1 \reg_pmp_3_cfg_r$_DFFE_PP_  (
    .CK(clock),
    .D(_00098_),
    .Q(reg_pmp_3_cfg_r),
    .QN(_07000_)
  );
  DFF_X1 \reg_pmp_3_cfg_w$_DFFE_PP_  (
    .CK(clock),
    .D(_00096_),
    .Q(reg_pmp_3_cfg_w),
    .QN(_07002_)
  );
  DFF_X1 \reg_pmp_3_cfg_x$_DFFE_PP_  (
    .CK(clock),
    .D(_00097_),
    .Q(reg_pmp_3_cfg_x),
    .QN(_07001_)
  );
  DFF_X1 \reg_pmp_4_addr[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00061_),
    .Q(reg_pmp_4_addr[0]),
    .QN(_07035_)
  );
  DFF_X1 \reg_pmp_4_addr[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00071_),
    .Q(reg_pmp_4_addr[10]),
    .QN(_07025_)
  );
  DFF_X1 \reg_pmp_4_addr[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00072_),
    .Q(reg_pmp_4_addr[11]),
    .QN(_07024_)
  );
  DFF_X1 \reg_pmp_4_addr[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00073_),
    .Q(reg_pmp_4_addr[12]),
    .QN(_07023_)
  );
  DFF_X1 \reg_pmp_4_addr[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00074_),
    .Q(reg_pmp_4_addr[13]),
    .QN(_07022_)
  );
  DFF_X1 \reg_pmp_4_addr[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00075_),
    .Q(reg_pmp_4_addr[14]),
    .QN(_07021_)
  );
  DFF_X1 \reg_pmp_4_addr[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00076_),
    .Q(reg_pmp_4_addr[15]),
    .QN(_07020_)
  );
  DFF_X1 \reg_pmp_4_addr[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00077_),
    .Q(reg_pmp_4_addr[16]),
    .QN(_07019_)
  );
  DFF_X1 \reg_pmp_4_addr[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00078_),
    .Q(reg_pmp_4_addr[17]),
    .QN(_07018_)
  );
  DFF_X1 \reg_pmp_4_addr[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00079_),
    .Q(reg_pmp_4_addr[18]),
    .QN(_07017_)
  );
  DFF_X1 \reg_pmp_4_addr[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00080_),
    .Q(reg_pmp_4_addr[19]),
    .QN(_07016_)
  );
  DFF_X1 \reg_pmp_4_addr[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00062_),
    .Q(reg_pmp_4_addr[1]),
    .QN(_07034_)
  );
  DFF_X1 \reg_pmp_4_addr[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00081_),
    .Q(reg_pmp_4_addr[20]),
    .QN(_07015_)
  );
  DFF_X1 \reg_pmp_4_addr[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00082_),
    .Q(reg_pmp_4_addr[21]),
    .QN(_07014_)
  );
  DFF_X1 \reg_pmp_4_addr[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00083_),
    .Q(reg_pmp_4_addr[22]),
    .QN(_07013_)
  );
  DFF_X1 \reg_pmp_4_addr[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00084_),
    .Q(reg_pmp_4_addr[23]),
    .QN(_07012_)
  );
  DFF_X1 \reg_pmp_4_addr[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00085_),
    .Q(reg_pmp_4_addr[24]),
    .QN(_07011_)
  );
  DFF_X1 \reg_pmp_4_addr[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00086_),
    .Q(reg_pmp_4_addr[25]),
    .QN(_07010_)
  );
  DFF_X1 \reg_pmp_4_addr[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00087_),
    .Q(reg_pmp_4_addr[26]),
    .QN(_07009_)
  );
  DFF_X1 \reg_pmp_4_addr[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00088_),
    .Q(reg_pmp_4_addr[27]),
    .QN(_07008_)
  );
  DFF_X1 \reg_pmp_4_addr[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00089_),
    .Q(reg_pmp_4_addr[28]),
    .QN(_07007_)
  );
  DFF_X1 \reg_pmp_4_addr[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00090_),
    .Q(reg_pmp_4_addr[29]),
    .QN(_07006_)
  );
  DFF_X1 \reg_pmp_4_addr[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00063_),
    .Q(reg_pmp_4_addr[2]),
    .QN(_07033_)
  );
  DFF_X1 \reg_pmp_4_addr[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00064_),
    .Q(reg_pmp_4_addr[3]),
    .QN(_07032_)
  );
  DFF_X1 \reg_pmp_4_addr[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00065_),
    .Q(reg_pmp_4_addr[4]),
    .QN(_07031_)
  );
  DFF_X1 \reg_pmp_4_addr[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00066_),
    .Q(reg_pmp_4_addr[5]),
    .QN(_07030_)
  );
  DFF_X1 \reg_pmp_4_addr[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00067_),
    .Q(reg_pmp_4_addr[6]),
    .QN(_07029_)
  );
  DFF_X1 \reg_pmp_4_addr[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00068_),
    .Q(reg_pmp_4_addr[7]),
    .QN(_07028_)
  );
  DFF_X1 \reg_pmp_4_addr[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00069_),
    .Q(reg_pmp_4_addr[8]),
    .QN(_07027_)
  );
  DFF_X1 \reg_pmp_4_addr[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00070_),
    .Q(reg_pmp_4_addr[9]),
    .QN(_07026_)
  );
  DFF_X1 \reg_pmp_4_cfg_a[0]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00093_),
    .Q(reg_pmp_4_cfg_a[0]),
    .QN(_07003_)
  );
  DFF_X1 \reg_pmp_4_cfg_a[1]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00094_),
    .Q(reg_pmp_4_cfg_a[1]),
    .QN(_00014_)
  );
  DFF_X1 \reg_pmp_4_cfg_l$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00095_),
    .Q(reg_pmp_4_cfg_l),
    .QN(_00013_)
  );
  DFF_X1 \reg_pmp_4_cfg_r$_DFFE_PP_  (
    .CK(clock),
    .D(_00169_),
    .Q(reg_pmp_4_cfg_r),
    .QN(_06933_)
  );
  DFF_X1 \reg_pmp_4_cfg_w$_DFFE_PP_  (
    .CK(clock),
    .D(_00091_),
    .Q(reg_pmp_4_cfg_w),
    .QN(_07005_)
  );
  DFF_X1 \reg_pmp_4_cfg_x$_DFFE_PP_  (
    .CK(clock),
    .D(_00092_),
    .Q(reg_pmp_4_cfg_x),
    .QN(_07004_)
  );
  DFF_X1 \reg_pmp_5_addr[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00027_),
    .Q(reg_pmp_5_addr[0]),
    .QN(_07067_)
  );
  DFF_X1 \reg_pmp_5_addr[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00037_),
    .Q(reg_pmp_5_addr[10]),
    .QN(_07057_)
  );
  DFF_X1 \reg_pmp_5_addr[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00038_),
    .Q(reg_pmp_5_addr[11]),
    .QN(_07056_)
  );
  DFF_X1 \reg_pmp_5_addr[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00039_),
    .Q(reg_pmp_5_addr[12]),
    .QN(_07055_)
  );
  DFF_X1 \reg_pmp_5_addr[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00040_),
    .Q(reg_pmp_5_addr[13]),
    .QN(_07054_)
  );
  DFF_X1 \reg_pmp_5_addr[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00041_),
    .Q(reg_pmp_5_addr[14]),
    .QN(_07053_)
  );
  DFF_X1 \reg_pmp_5_addr[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00042_),
    .Q(reg_pmp_5_addr[15]),
    .QN(_07052_)
  );
  DFF_X1 \reg_pmp_5_addr[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00043_),
    .Q(reg_pmp_5_addr[16]),
    .QN(_07051_)
  );
  DFF_X1 \reg_pmp_5_addr[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00044_),
    .Q(reg_pmp_5_addr[17]),
    .QN(_07050_)
  );
  DFF_X1 \reg_pmp_5_addr[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00045_),
    .Q(reg_pmp_5_addr[18]),
    .QN(_07049_)
  );
  DFF_X1 \reg_pmp_5_addr[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00046_),
    .Q(reg_pmp_5_addr[19]),
    .QN(_07048_)
  );
  DFF_X1 \reg_pmp_5_addr[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00028_),
    .Q(reg_pmp_5_addr[1]),
    .QN(_07066_)
  );
  DFF_X1 \reg_pmp_5_addr[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00047_),
    .Q(reg_pmp_5_addr[20]),
    .QN(_07047_)
  );
  DFF_X1 \reg_pmp_5_addr[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00048_),
    .Q(reg_pmp_5_addr[21]),
    .QN(_07046_)
  );
  DFF_X1 \reg_pmp_5_addr[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00049_),
    .Q(reg_pmp_5_addr[22]),
    .QN(_07045_)
  );
  DFF_X1 \reg_pmp_5_addr[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00050_),
    .Q(reg_pmp_5_addr[23]),
    .QN(_07044_)
  );
  DFF_X1 \reg_pmp_5_addr[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00051_),
    .Q(reg_pmp_5_addr[24]),
    .QN(_07043_)
  );
  DFF_X1 \reg_pmp_5_addr[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00052_),
    .Q(reg_pmp_5_addr[25]),
    .QN(_07042_)
  );
  DFF_X1 \reg_pmp_5_addr[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00053_),
    .Q(reg_pmp_5_addr[26]),
    .QN(_07041_)
  );
  DFF_X1 \reg_pmp_5_addr[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00054_),
    .Q(reg_pmp_5_addr[27]),
    .QN(_07040_)
  );
  DFF_X1 \reg_pmp_5_addr[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00055_),
    .Q(reg_pmp_5_addr[28]),
    .QN(_07039_)
  );
  DFF_X1 \reg_pmp_5_addr[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00056_),
    .Q(reg_pmp_5_addr[29]),
    .QN(_07038_)
  );
  DFF_X1 \reg_pmp_5_addr[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00029_),
    .Q(reg_pmp_5_addr[2]),
    .QN(_07065_)
  );
  DFF_X1 \reg_pmp_5_addr[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00030_),
    .Q(reg_pmp_5_addr[3]),
    .QN(_07064_)
  );
  DFF_X1 \reg_pmp_5_addr[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00031_),
    .Q(reg_pmp_5_addr[4]),
    .QN(_07063_)
  );
  DFF_X1 \reg_pmp_5_addr[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00032_),
    .Q(reg_pmp_5_addr[5]),
    .QN(_07062_)
  );
  DFF_X1 \reg_pmp_5_addr[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00033_),
    .Q(reg_pmp_5_addr[6]),
    .QN(_07061_)
  );
  DFF_X1 \reg_pmp_5_addr[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00034_),
    .Q(reg_pmp_5_addr[7]),
    .QN(_07060_)
  );
  DFF_X1 \reg_pmp_5_addr[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00035_),
    .Q(reg_pmp_5_addr[8]),
    .QN(_07059_)
  );
  DFF_X1 \reg_pmp_5_addr[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00036_),
    .Q(reg_pmp_5_addr[9]),
    .QN(_07058_)
  );
  DFF_X1 \reg_pmp_5_cfg_a[0]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00058_),
    .Q(reg_pmp_5_cfg_a[0]),
    .QN(_07036_)
  );
  DFF_X1 \reg_pmp_5_cfg_a[1]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00059_),
    .Q(reg_pmp_5_cfg_a[1]),
    .QN(_00016_)
  );
  DFF_X1 \reg_pmp_5_cfg_l$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00060_),
    .Q(reg_pmp_5_cfg_l),
    .QN(_00015_)
  );
  DFF_X1 \reg_pmp_5_cfg_r$_DFFE_PP_  (
    .CK(clock),
    .D(_00025_),
    .Q(reg_pmp_5_cfg_r),
    .QN(_07069_)
  );
  DFF_X1 \reg_pmp_5_cfg_w$_DFFE_PP_  (
    .CK(clock),
    .D(_00026_),
    .Q(reg_pmp_5_cfg_w),
    .QN(_07068_)
  );
  DFF_X1 \reg_pmp_5_cfg_x$_DFFE_PP_  (
    .CK(clock),
    .D(_00364_),
    .Q(reg_pmp_5_cfg_x),
    .QN(_06744_)
  );
  DFF_X1 \reg_pmp_6_addr[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00395_),
    .Q(reg_pmp_6_addr[0]),
    .QN(_06713_)
  );
  DFF_X1 \reg_pmp_6_addr[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00405_),
    .Q(reg_pmp_6_addr[10]),
    .QN(_06703_)
  );
  DFF_X1 \reg_pmp_6_addr[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00406_),
    .Q(reg_pmp_6_addr[11]),
    .QN(_06702_)
  );
  DFF_X1 \reg_pmp_6_addr[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00407_),
    .Q(reg_pmp_6_addr[12]),
    .QN(_06701_)
  );
  DFF_X1 \reg_pmp_6_addr[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00408_),
    .Q(reg_pmp_6_addr[13]),
    .QN(_06700_)
  );
  DFF_X1 \reg_pmp_6_addr[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00409_),
    .Q(reg_pmp_6_addr[14]),
    .QN(_06699_)
  );
  DFF_X1 \reg_pmp_6_addr[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00410_),
    .Q(reg_pmp_6_addr[15]),
    .QN(_06698_)
  );
  DFF_X1 \reg_pmp_6_addr[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00411_),
    .Q(reg_pmp_6_addr[16]),
    .QN(_06697_)
  );
  DFF_X1 \reg_pmp_6_addr[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00412_),
    .Q(reg_pmp_6_addr[17]),
    .QN(_06696_)
  );
  DFF_X1 \reg_pmp_6_addr[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00413_),
    .Q(reg_pmp_6_addr[18]),
    .QN(_06695_)
  );
  DFF_X1 \reg_pmp_6_addr[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00414_),
    .Q(reg_pmp_6_addr[19]),
    .QN(_06694_)
  );
  DFF_X1 \reg_pmp_6_addr[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00396_),
    .Q(reg_pmp_6_addr[1]),
    .QN(_06712_)
  );
  DFF_X1 \reg_pmp_6_addr[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00415_),
    .Q(reg_pmp_6_addr[20]),
    .QN(_06693_)
  );
  DFF_X1 \reg_pmp_6_addr[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00416_),
    .Q(reg_pmp_6_addr[21]),
    .QN(_06692_)
  );
  DFF_X1 \reg_pmp_6_addr[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00417_),
    .Q(reg_pmp_6_addr[22]),
    .QN(_06691_)
  );
  DFF_X1 \reg_pmp_6_addr[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00418_),
    .Q(reg_pmp_6_addr[23]),
    .QN(_06690_)
  );
  DFF_X1 \reg_pmp_6_addr[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00419_),
    .Q(reg_pmp_6_addr[24]),
    .QN(_06689_)
  );
  DFF_X1 \reg_pmp_6_addr[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00420_),
    .Q(reg_pmp_6_addr[25]),
    .QN(_06688_)
  );
  DFF_X1 \reg_pmp_6_addr[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00421_),
    .Q(reg_pmp_6_addr[26]),
    .QN(_06687_)
  );
  DFF_X1 \reg_pmp_6_addr[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00422_),
    .Q(reg_pmp_6_addr[27]),
    .QN(_06686_)
  );
  DFF_X1 \reg_pmp_6_addr[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00423_),
    .Q(reg_pmp_6_addr[28]),
    .QN(_06685_)
  );
  DFF_X1 \reg_pmp_6_addr[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00424_),
    .Q(reg_pmp_6_addr[29]),
    .QN(_06684_)
  );
  DFF_X1 \reg_pmp_6_addr[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00397_),
    .Q(reg_pmp_6_addr[2]),
    .QN(_06711_)
  );
  DFF_X1 \reg_pmp_6_addr[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00398_),
    .Q(reg_pmp_6_addr[3]),
    .QN(_06710_)
  );
  DFF_X1 \reg_pmp_6_addr[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00399_),
    .Q(reg_pmp_6_addr[4]),
    .QN(_06709_)
  );
  DFF_X1 \reg_pmp_6_addr[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00400_),
    .Q(reg_pmp_6_addr[5]),
    .QN(_06708_)
  );
  DFF_X1 \reg_pmp_6_addr[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00401_),
    .Q(reg_pmp_6_addr[6]),
    .QN(_06707_)
  );
  DFF_X1 \reg_pmp_6_addr[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00402_),
    .Q(reg_pmp_6_addr[7]),
    .QN(_06706_)
  );
  DFF_X1 \reg_pmp_6_addr[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00403_),
    .Q(reg_pmp_6_addr[8]),
    .QN(_06705_)
  );
  DFF_X1 \reg_pmp_6_addr[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00404_),
    .Q(reg_pmp_6_addr[9]),
    .QN(_06704_)
  );
  DFF_X1 \reg_pmp_6_cfg_a[0]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00022_),
    .Q(reg_pmp_6_cfg_a[0]),
    .QN(_07070_)
  );
  DFF_X1 \reg_pmp_6_cfg_a[1]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00023_),
    .Q(reg_pmp_6_cfg_a[1]),
    .QN(_00018_)
  );
  DFF_X1 \reg_pmp_6_cfg_l$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00024_),
    .Q(reg_pmp_6_cfg_l),
    .QN(_00017_)
  );
  DFF_X1 \reg_pmp_6_cfg_r$_DFFE_PP_  (
    .CK(clock),
    .D(_00019_),
    .Q(reg_pmp_6_cfg_r),
    .QN(_07073_)
  );
  DFF_X1 \reg_pmp_6_cfg_w$_DFFE_PP_  (
    .CK(clock),
    .D(_00621_),
    .Q(reg_pmp_6_cfg_w),
    .QN(_06493_)
  );
  DFF_X1 \reg_pmp_6_cfg_x$_DFFE_PP_  (
    .CK(clock),
    .D(_00020_),
    .Q(reg_pmp_6_cfg_x),
    .QN(_07072_)
  );
  DFF_X1 \reg_pmp_7_addr[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00536_),
    .Q(reg_pmp_7_addr[0]),
    .QN(_06574_)
  );
  DFF_X1 \reg_pmp_7_addr[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00546_),
    .Q(reg_pmp_7_addr[10]),
    .QN(_06564_)
  );
  DFF_X1 \reg_pmp_7_addr[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00547_),
    .Q(reg_pmp_7_addr[11]),
    .QN(_06563_)
  );
  DFF_X1 \reg_pmp_7_addr[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00548_),
    .Q(reg_pmp_7_addr[12]),
    .QN(_06562_)
  );
  DFF_X1 \reg_pmp_7_addr[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00549_),
    .Q(reg_pmp_7_addr[13]),
    .QN(_06561_)
  );
  DFF_X1 \reg_pmp_7_addr[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00550_),
    .Q(reg_pmp_7_addr[14]),
    .QN(_06560_)
  );
  DFF_X1 \reg_pmp_7_addr[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00551_),
    .Q(reg_pmp_7_addr[15]),
    .QN(_06559_)
  );
  DFF_X1 \reg_pmp_7_addr[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00552_),
    .Q(reg_pmp_7_addr[16]),
    .QN(_06558_)
  );
  DFF_X1 \reg_pmp_7_addr[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00553_),
    .Q(reg_pmp_7_addr[17]),
    .QN(_06557_)
  );
  DFF_X1 \reg_pmp_7_addr[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00554_),
    .Q(reg_pmp_7_addr[18]),
    .QN(_06556_)
  );
  DFF_X1 \reg_pmp_7_addr[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00555_),
    .Q(reg_pmp_7_addr[19]),
    .QN(_06555_)
  );
  DFF_X1 \reg_pmp_7_addr[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00537_),
    .Q(reg_pmp_7_addr[1]),
    .QN(_06573_)
  );
  DFF_X1 \reg_pmp_7_addr[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00556_),
    .Q(reg_pmp_7_addr[20]),
    .QN(_06554_)
  );
  DFF_X1 \reg_pmp_7_addr[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00557_),
    .Q(reg_pmp_7_addr[21]),
    .QN(_06553_)
  );
  DFF_X1 \reg_pmp_7_addr[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00558_),
    .Q(reg_pmp_7_addr[22]),
    .QN(_06552_)
  );
  DFF_X1 \reg_pmp_7_addr[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00559_),
    .Q(reg_pmp_7_addr[23]),
    .QN(_06551_)
  );
  DFF_X1 \reg_pmp_7_addr[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00560_),
    .Q(reg_pmp_7_addr[24]),
    .QN(_06550_)
  );
  DFF_X1 \reg_pmp_7_addr[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00561_),
    .Q(reg_pmp_7_addr[25]),
    .QN(_06549_)
  );
  DFF_X1 \reg_pmp_7_addr[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00562_),
    .Q(reg_pmp_7_addr[26]),
    .QN(_06548_)
  );
  DFF_X1 \reg_pmp_7_addr[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00563_),
    .Q(reg_pmp_7_addr[27]),
    .QN(_06547_)
  );
  DFF_X1 \reg_pmp_7_addr[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00564_),
    .Q(reg_pmp_7_addr[28]),
    .QN(_06546_)
  );
  DFF_X1 \reg_pmp_7_addr[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00565_),
    .Q(reg_pmp_7_addr[29]),
    .QN(_06545_)
  );
  DFF_X1 \reg_pmp_7_addr[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00538_),
    .Q(reg_pmp_7_addr[2]),
    .QN(_06572_)
  );
  DFF_X1 \reg_pmp_7_addr[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00539_),
    .Q(reg_pmp_7_addr[3]),
    .QN(_06571_)
  );
  DFF_X1 \reg_pmp_7_addr[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00540_),
    .Q(reg_pmp_7_addr[4]),
    .QN(_06570_)
  );
  DFF_X1 \reg_pmp_7_addr[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00541_),
    .Q(reg_pmp_7_addr[5]),
    .QN(_06569_)
  );
  DFF_X1 \reg_pmp_7_addr[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00542_),
    .Q(reg_pmp_7_addr[6]),
    .QN(_06568_)
  );
  DFF_X1 \reg_pmp_7_addr[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00543_),
    .Q(reg_pmp_7_addr[7]),
    .QN(_06567_)
  );
  DFF_X1 \reg_pmp_7_addr[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00544_),
    .Q(reg_pmp_7_addr[8]),
    .QN(_06566_)
  );
  DFF_X1 \reg_pmp_7_addr[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00545_),
    .Q(reg_pmp_7_addr[9]),
    .QN(_06565_)
  );
  DFF_X1 \reg_pmp_7_cfg_a[0]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00566_),
    .Q(reg_pmp_7_cfg_a[0]),
    .QN(_06544_)
  );
  DFF_X1 \reg_pmp_7_cfg_a[1]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00567_),
    .Q(reg_pmp_7_cfg_a[1]),
    .QN(_00004_)
  );
  DFF_X1 \reg_pmp_7_cfg_l$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00568_),
    .Q(reg_pmp_7_cfg_l),
    .QN(_00003_)
  );
  DFF_X1 \reg_pmp_7_cfg_r$_DFFE_PP_  (
    .CK(clock),
    .D(_00533_),
    .Q(reg_pmp_7_cfg_r),
    .QN(_06577_)
  );
  DFF_X1 \reg_pmp_7_cfg_w$_DFFE_PP_  (
    .CK(clock),
    .D(_00534_),
    .Q(reg_pmp_7_cfg_w),
    .QN(_06576_)
  );
  DFF_X1 \reg_pmp_7_cfg_x$_DFFE_PP_  (
    .CK(clock),
    .D(_00535_),
    .Q(reg_pmp_7_cfg_x),
    .QN(_06575_)
  );
  DFF_X1 \reg_singleStepped$_SDFF_PN0_  (
    .CK(clock),
    .D(_00247_),
    .Q(reg_singleStepped),
    .QN(_06858_)
  );
  DFF_X1 \reg_wfi$_SDFF_PP0_  (
    .CK(io_ungated_clock),
    .D(_00292_),
    .Q(reg_wfi),
    .QN(_06816_)
  );
  DFF_X1 \small_1[0]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00326_),
    .Q(small_1[0]),
    .QN(_06782_)
  );
  DFF_X1 \small_1[1]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00327_),
    .Q(small_1[1]),
    .QN(_06781_)
  );
  DFF_X1 \small_1[2]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00328_),
    .Q(small_1[2]),
    .QN(_06780_)
  );
  DFF_X1 \small_1[3]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00329_),
    .Q(small_1[3]),
    .QN(_06779_)
  );
  DFF_X1 \small_1[4]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00330_),
    .Q(small_1[4]),
    .QN(_06778_)
  );
  DFF_X1 \small_1[5]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_00331_),
    .Q(small_1[5]),
    .QN(_06777_)
  );
  DFF_X1 \small_[0]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00461_),
    .Q(small_[0]),
    .QN(_06648_)
  );
  DFF_X1 \small_[1]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00462_),
    .Q(small_[1]),
    .QN(_06647_)
  );
  DFF_X1 \small_[2]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00463_),
    .Q(small_[2]),
    .QN(_06646_)
  );
  DFF_X1 \small_[3]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00464_),
    .Q(small_[3]),
    .QN(_06645_)
  );
  DFF_X1 \small_[4]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00465_),
    .Q(small_[4]),
    .QN(_06644_)
  );
  DFF_X1 \small_[5]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00466_),
    .Q(small_[5]),
    .QN(_06643_)
  );
  assign _GEN_170 = 2'h0;
  assign _GEN_207 = 2'h0;
  assign _GEN_239[0] = 1'h0;
  assign _GEN_34 = { 5'h00, io_retire };
  assign _GEN_35[5:1] = 5'h00;
  assign _GEN_40 = { 20'h00000, io_interrupts_meip, 3'h0, io_interrupts_mtip, 3'h0, io_interrupts_msip, 3'h0 };
  assign _GEN_41 = { 28'h0000000, io_interrupt_cause[3:0] };
  assign _GEN_51 = 1'h1;
  assign { _GEN_586[31:2], _GEN_586[0] } = 31'h00000001;
  assign { _GEN_592[31:12], _GEN_592[10:8], _GEN_592[6:4], _GEN_592[2:0] } = 29'h00000000;
  assign _GEN_593[31:1] = 31'h00000000;
  assign { _GEN_594[31:3], _GEN_594[1] } = 30'h00000000;
  assign _GEN_595[63:32] = 32'd0;
  assign _GEN_596[63:32] = 32'd0;
  assign _GEN_597[63:32] = 32'd0;
  assign { _GEN_598[63:32], _GEN_598[30:29], _GEN_598[22:21], _GEN_598[14:13], _GEN_598[6:5] } = 40'h0000000000;
  assign { _GEN_599[63:32], _GEN_599[30:29], _GEN_599[22:21], _GEN_599[14:13], _GEN_599[6:5] } = 40'h0000000000;
  assign _GEN_600[63:30] = 34'h000000000;
  assign _GEN_601[63:30] = 34'h000000000;
  assign _GEN_602[63:30] = 34'h000000000;
  assign _GEN_603[63:30] = 34'h000000000;
  assign _GEN_604[63:30] = 34'h000000000;
  assign _GEN_605[63:30] = 34'h000000000;
  assign _GEN_606[63:30] = 34'h000000000;
  assign _GEN_607[63:30] = 34'h000000000;
  assign { _GEN_608[63:4], _GEN_608[2:0] } = 63'h0000000000000000;
  assign _GEN_609[63:1] = 63'h0000000000000000;
  assign { _GEN_610[63:30], _GEN_610[28:0] } = { 42'h00000000000, _GEN_610[29], _GEN_610[29], 6'h00, _GEN_610[29], 9'h000, _GEN_610[29], 2'h0 };
  assign { _GEN_611[31:4], _GEN_611[2:0] } = 31'h00000000;
  assign _GEN_73 = 2'h0;
  assign _T_16 = { 4'h2, reg_bp_0_control_dmode, 14'h0400, reg_bp_0_control_action, 3'h0, reg_bp_0_control_tmatch, 4'h8, reg_bp_0_control_x, reg_bp_0_control_w, reg_bp_0_control_r };
  assign _T_20 = { _GEN_586[1], 1'h1 };
  assign _T_2000[63:32] = large_1[57:26];
  assign _T_2003 = { _T_2000[31:0], large_1[25:0], small_1 };
  assign _T_2005 = { large_[57:26], _T_2000[31:0] };
  assign _T_2008 = { _T_2000[31:0], large_[25:0], small_ };
  assign { _T_21[31:2], _T_21[0] } = { _T_18[31:2], 1'h1 };
  assign _T_213 = { io_rw_addr, 20'h00000 };
  assign { _T_22[31:2], _T_22[0] } = { reg_mepc[31:2], 1'h0 };
  assign _T_23 = { 16'h4000, reg_dcsr_ebreakm, 6'h00, reg_dcsr_cause, 3'h0, reg_dcsr_step, 2'h3 };
  assign { _T_27[31:2], _T_27[0] } = { _T_24[31:2], 1'h1 };
  assign { _T_28[31:2], _T_28[0] } = { reg_dpc[31:2], 1'h0 };
  assign _T_60 = { reg_pmp_0_cfg_l, 2'h0, reg_pmp_0_cfg_a, reg_pmp_0_cfg_x, reg_pmp_0_cfg_w, reg_pmp_0_cfg_r };
  assign _T_62 = { reg_pmp_2_cfg_l, 2'h0, reg_pmp_2_cfg_a, reg_pmp_2_cfg_x, reg_pmp_2_cfg_w, reg_pmp_2_cfg_r };
  assign _T_64 = { reg_pmp_3_cfg_l, 2'h0, reg_pmp_3_cfg_a, reg_pmp_3_cfg_x, reg_pmp_3_cfg_w, reg_pmp_3_cfg_r, reg_pmp_2_cfg_l, 2'h0, reg_pmp_2_cfg_a, reg_pmp_2_cfg_x, reg_pmp_2_cfg_w, reg_pmp_2_cfg_r, reg_pmp_1_cfg_l, 2'h0, reg_pmp_1_cfg_a, reg_pmp_1_cfg_x, reg_pmp_1_cfg_w, reg_pmp_1_cfg_r, reg_pmp_0_cfg_l, 2'h0, reg_pmp_0_cfg_a, reg_pmp_0_cfg_x, reg_pmp_0_cfg_w, reg_pmp_0_cfg_r };
  assign _T_65 = { reg_pmp_4_cfg_l, 2'h0, reg_pmp_4_cfg_a, reg_pmp_4_cfg_x, reg_pmp_4_cfg_w, reg_pmp_4_cfg_r };
  assign _T_67 = { reg_pmp_6_cfg_l, 2'h0, reg_pmp_6_cfg_a, reg_pmp_6_cfg_x, reg_pmp_6_cfg_w, reg_pmp_6_cfg_r };
  assign _T_69 = { reg_pmp_7_cfg_l, 2'h0, reg_pmp_7_cfg_a, reg_pmp_7_cfg_x, reg_pmp_7_cfg_w, reg_pmp_7_cfg_r, reg_pmp_6_cfg_l, 2'h0, reg_pmp_6_cfg_a, reg_pmp_6_cfg_x, reg_pmp_6_cfg_w, reg_pmp_6_cfg_r, reg_pmp_5_cfg_l, 2'h0, reg_pmp_5_cfg_a, reg_pmp_5_cfg_x, reg_pmp_5_cfg_w, reg_pmp_5_cfg_r, reg_pmp_4_cfg_l, 2'h0, reg_pmp_4_cfg_a, reg_pmp_4_cfg_x, reg_pmp_4_cfg_w, reg_pmp_4_cfg_r };
  assign _any_T_78 = io_interrupts_debug;
  assign _causeIsDebugBreak_T_3 = { reg_dcsr_ebreakm, 3'h0 };
  assign _causeIsDebugBreak_T_4 = { 3'h0, reg_dcsr_ebreakm };
  assign { _debugTVec_T[11:4], _debugTVec_T[2:0] } = 11'h400;
  assign _decoded_T_10[1] = io_rw_addr[10];
  assign _decoded_T_14[11] = io_decode_0_inst[20];
  assign _decoded_T_16[3] = io_decode_0_inst[28];
  assign _decoded_T_18[3:2] = { io_decode_0_inst[28], io_decode_0_inst[29] };
  assign _decoded_T_2[11] = io_rw_addr[0];
  assign { _decoded_T_20[9], _decoded_T_20[3:2] } = { io_decode_0_inst[22], io_decode_0_inst[28], io_decode_0_inst[29] };
  assign _decoded_T_22[1] = io_decode_0_inst[30];
  assign _decoded_T_4[3] = io_rw_addr[8];
  assign _decoded_T_6[3:2] = { io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_T_8[9], _decoded_T_8[3:2] } = { io_rw_addr[2], io_rw_addr[8], io_rw_addr[9] };
  assign _decoded_decoded_T[3:2] = { io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_10[10], _decoded_decoded_T_10[6], _decoded_decoded_T_10[3:2] } = { io_rw_addr[1], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_100[11:9], _decoded_decoded_T_100[7:6], _decoded_decoded_T_100[4:2] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[2], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_102[8:6], _decoded_decoded_T_102[4:2] } = { io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_104[11], _decoded_decoded_T_104[8:6], _decoded_decoded_T_104[4:2] } = { io_rw_addr[0], io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_106[10], _decoded_decoded_T_106[8:6], _decoded_decoded_T_106[4:2] } = { io_rw_addr[1], io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_108[11:10], _decoded_decoded_T_108[8:6], _decoded_decoded_T_108[4:2] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_110[9:6], _decoded_decoded_T_110[4:2] } = { io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_112[11], _decoded_decoded_T_112[9:6], _decoded_decoded_T_112[4:2] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_114[10:6], _decoded_decoded_T_114[4:2] } = { io_rw_addr[1], io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_116[11:6], _decoded_decoded_T_116[4:2] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_118[6], _decoded_decoded_T_118[4:1] } = { io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[10] };
  assign { _decoded_decoded_T_12[9], _decoded_decoded_T_12[6], _decoded_decoded_T_12[3:2] } = { io_rw_addr[2], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_120[11], _decoded_decoded_T_120[6], _decoded_decoded_T_120[4:1] } = { io_rw_addr[0], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[10] };
  assign { _decoded_decoded_T_122[10], _decoded_decoded_T_122[6], _decoded_decoded_T_122[4:1] } = { io_rw_addr[1], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[10] };
  assign { _decoded_decoded_T_124[11:10], _decoded_decoded_T_124[6], _decoded_decoded_T_124[4:1] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[10] };
  assign { _decoded_decoded_T_126[7:6], _decoded_decoded_T_126[4:1] } = { io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[10] };
  assign { _decoded_decoded_T_128[11], _decoded_decoded_T_128[7:6], _decoded_decoded_T_128[4:1] } = { io_rw_addr[0], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[10] };
  assign { _decoded_decoded_T_130[10], _decoded_decoded_T_130[7:6], _decoded_decoded_T_130[4:1] } = { io_rw_addr[1], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[10] };
  assign _decoded_decoded_T_132[5:1] = { io_rw_addr[6], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[10] };
  assign { _decoded_decoded_T_134[3:2], _decoded_decoded_T_134[0] } = { io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_136[10], _decoded_decoded_T_136[3:2], _decoded_decoded_T_136[0] } = { io_rw_addr[1], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_138[11:10], _decoded_decoded_T_138[3:2], _decoded_decoded_T_138[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_14[11], _decoded_decoded_T_14[9], _decoded_decoded_T_14[6], _decoded_decoded_T_14[3:2] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_140[9], _decoded_decoded_T_140[3:2], _decoded_decoded_T_140[0] } = { io_rw_addr[2], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_142[11], _decoded_decoded_T_142[9], _decoded_decoded_T_142[3:2], _decoded_decoded_T_142[0] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_144[10:9], _decoded_decoded_T_144[3:2], _decoded_decoded_T_144[0] } = { io_rw_addr[1], io_rw_addr[2], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_146[11:9], _decoded_decoded_T_146[3:2], _decoded_decoded_T_146[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[2], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_148[8], _decoded_decoded_T_148[3:2], _decoded_decoded_T_148[0] } = { io_rw_addr[3], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_150[11], _decoded_decoded_T_150[8], _decoded_decoded_T_150[3:2], _decoded_decoded_T_150[0] } = { io_rw_addr[0], io_rw_addr[3], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_152[10], _decoded_decoded_T_152[8], _decoded_decoded_T_152[3:2], _decoded_decoded_T_152[0] } = { io_rw_addr[1], io_rw_addr[3], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_154[11:10], _decoded_decoded_T_154[8], _decoded_decoded_T_154[3:2], _decoded_decoded_T_154[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[3], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_156[9:8], _decoded_decoded_T_156[3:2], _decoded_decoded_T_156[0] } = { io_rw_addr[2], io_rw_addr[3], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_158[11], _decoded_decoded_T_158[9:8], _decoded_decoded_T_158[3:2], _decoded_decoded_T_158[0] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[3], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_16[10:9], _decoded_decoded_T_16[6], _decoded_decoded_T_16[3:2] } = { io_rw_addr[1], io_rw_addr[2], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_160[10:8], _decoded_decoded_T_160[3:2], _decoded_decoded_T_160[0] } = { io_rw_addr[1], io_rw_addr[2], io_rw_addr[3], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_162[11:8], _decoded_decoded_T_162[3:2], _decoded_decoded_T_162[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[2], io_rw_addr[3], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_164[7], _decoded_decoded_T_164[3:2], _decoded_decoded_T_164[0] } = { io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_166[11], _decoded_decoded_T_166[7], _decoded_decoded_T_166[3:2], _decoded_decoded_T_166[0] } = { io_rw_addr[0], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_168[10], _decoded_decoded_T_168[7], _decoded_decoded_T_168[3:2], _decoded_decoded_T_168[0] } = { io_rw_addr[1], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_170[11:10], _decoded_decoded_T_170[7], _decoded_decoded_T_170[3:2], _decoded_decoded_T_170[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_172[9], _decoded_decoded_T_172[7], _decoded_decoded_T_172[3:2], _decoded_decoded_T_172[0] } = { io_rw_addr[2], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_174[11], _decoded_decoded_T_174[9], _decoded_decoded_T_174[7], _decoded_decoded_T_174[3:2], _decoded_decoded_T_174[0] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_176[10:9], _decoded_decoded_T_176[7], _decoded_decoded_T_176[3:2], _decoded_decoded_T_176[0] } = { io_rw_addr[1], io_rw_addr[2], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_178[11:9], _decoded_decoded_T_178[7], _decoded_decoded_T_178[3:2], _decoded_decoded_T_178[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[2], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_18[11:9], _decoded_decoded_T_18[6], _decoded_decoded_T_18[3:2] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[2], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_180[8:7], _decoded_decoded_T_180[3:2], _decoded_decoded_T_180[0] } = { io_rw_addr[3], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_182[11], _decoded_decoded_T_182[8:7], _decoded_decoded_T_182[3:2], _decoded_decoded_T_182[0] } = { io_rw_addr[0], io_rw_addr[3], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_184[10], _decoded_decoded_T_184[8:7], _decoded_decoded_T_184[3:2], _decoded_decoded_T_184[0] } = { io_rw_addr[1], io_rw_addr[3], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_186[11:10], _decoded_decoded_T_186[8:7], _decoded_decoded_T_186[3:2], _decoded_decoded_T_186[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[3], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_188[9:7], _decoded_decoded_T_188[3:2], _decoded_decoded_T_188[0] } = { io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_190[11], _decoded_decoded_T_190[9:7], _decoded_decoded_T_190[3:2], _decoded_decoded_T_190[0] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_192[10:7], _decoded_decoded_T_192[3:2], _decoded_decoded_T_192[0] } = { io_rw_addr[1], io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_194[11:7], _decoded_decoded_T_194[3:2], _decoded_decoded_T_194[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_196[4:2], _decoded_decoded_T_196[0] } = { io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_198[10], _decoded_decoded_T_198[4:2], _decoded_decoded_T_198[0] } = { io_rw_addr[1], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_2[11], _decoded_decoded_T_2[3:2] } = { io_rw_addr[0], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_20[8], _decoded_decoded_T_20[6], _decoded_decoded_T_20[3:2] } = { io_rw_addr[3], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_200[11:10], _decoded_decoded_T_200[4:2], _decoded_decoded_T_200[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_202[9], _decoded_decoded_T_202[4:2], _decoded_decoded_T_202[0] } = { io_rw_addr[2], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_204[11], _decoded_decoded_T_204[9], _decoded_decoded_T_204[4:2], _decoded_decoded_T_204[0] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_206[10:9], _decoded_decoded_T_206[4:2], _decoded_decoded_T_206[0] } = { io_rw_addr[1], io_rw_addr[2], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_208[11:9], _decoded_decoded_T_208[4:2], _decoded_decoded_T_208[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[2], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_210[8], _decoded_decoded_T_210[4:2], _decoded_decoded_T_210[0] } = { io_rw_addr[3], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_212[11], _decoded_decoded_T_212[8], _decoded_decoded_T_212[4:2], _decoded_decoded_T_212[0] } = { io_rw_addr[0], io_rw_addr[3], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_214[10], _decoded_decoded_T_214[8], _decoded_decoded_T_214[4:2], _decoded_decoded_T_214[0] } = { io_rw_addr[1], io_rw_addr[3], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_216[11:10], _decoded_decoded_T_216[8], _decoded_decoded_T_216[4:2], _decoded_decoded_T_216[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[3], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_218[9:8], _decoded_decoded_T_218[4:2], _decoded_decoded_T_218[0] } = { io_rw_addr[2], io_rw_addr[3], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_22[11], _decoded_decoded_T_22[8], _decoded_decoded_T_22[6], _decoded_decoded_T_22[3:2] } = { io_rw_addr[0], io_rw_addr[3], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_220[11], _decoded_decoded_T_220[9:8], _decoded_decoded_T_220[4:2], _decoded_decoded_T_220[0] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[3], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_222[10:8], _decoded_decoded_T_222[4:2], _decoded_decoded_T_222[0] } = { io_rw_addr[1], io_rw_addr[2], io_rw_addr[3], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_224[11:8], _decoded_decoded_T_224[4:2], _decoded_decoded_T_224[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[2], io_rw_addr[3], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_226[7], _decoded_decoded_T_226[4:2], _decoded_decoded_T_226[0] } = { io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_228[11], _decoded_decoded_T_228[7], _decoded_decoded_T_228[4:2], _decoded_decoded_T_228[0] } = { io_rw_addr[0], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_230[10], _decoded_decoded_T_230[7], _decoded_decoded_T_230[4:2], _decoded_decoded_T_230[0] } = { io_rw_addr[1], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_232[11:10], _decoded_decoded_T_232[7], _decoded_decoded_T_232[4:2], _decoded_decoded_T_232[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_234[9], _decoded_decoded_T_234[7], _decoded_decoded_T_234[4:2], _decoded_decoded_T_234[0] } = { io_rw_addr[2], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_236[11], _decoded_decoded_T_236[9], _decoded_decoded_T_236[7], _decoded_decoded_T_236[4:2], _decoded_decoded_T_236[0] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_238[10:9], _decoded_decoded_T_238[7], _decoded_decoded_T_238[4:2], _decoded_decoded_T_238[0] } = { io_rw_addr[1], io_rw_addr[2], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_24[10], _decoded_decoded_T_24[8], _decoded_decoded_T_24[6], _decoded_decoded_T_24[3:2] } = { io_rw_addr[1], io_rw_addr[3], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_240[11:9], _decoded_decoded_T_240[7], _decoded_decoded_T_240[4:2], _decoded_decoded_T_240[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[2], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_242[8:7], _decoded_decoded_T_242[4:2], _decoded_decoded_T_242[0] } = { io_rw_addr[3], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_244[11], _decoded_decoded_T_244[8:7], _decoded_decoded_T_244[4:2], _decoded_decoded_T_244[0] } = { io_rw_addr[0], io_rw_addr[3], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_246[10], _decoded_decoded_T_246[8:7], _decoded_decoded_T_246[4:2], _decoded_decoded_T_246[0] } = { io_rw_addr[1], io_rw_addr[3], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_248[11:10], _decoded_decoded_T_248[8:7], _decoded_decoded_T_248[4:2], _decoded_decoded_T_248[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[3], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_250[9:7], _decoded_decoded_T_250[4:2], _decoded_decoded_T_250[0] } = { io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_252[11], _decoded_decoded_T_252[9:7], _decoded_decoded_T_252[4:2], _decoded_decoded_T_252[0] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_254[10:7], _decoded_decoded_T_254[4:2], _decoded_decoded_T_254[0] } = { io_rw_addr[1], io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_256[11:7], _decoded_decoded_T_256[4:2], _decoded_decoded_T_256[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_258[7], _decoded_decoded_T_258[3:0] } = { io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[10], io_rw_addr[11] };
  assign { _decoded_decoded_T_26[11:10], _decoded_decoded_T_26[8], _decoded_decoded_T_26[6], _decoded_decoded_T_26[3:2] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[3], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_260[10], _decoded_decoded_T_260[7], _decoded_decoded_T_260[3:0] } = { io_rw_addr[1], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[10], io_rw_addr[11] };
  assign _decoded_decoded_T_261 = _GEN_609[0];
  assign { _decoded_decoded_T_262[11:10], _decoded_decoded_T_262[7], _decoded_decoded_T_262[3:0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[10], io_rw_addr[11] };
  assign _decoded_decoded_T_263 = _GEN_610[29];
  assign { _decoded_decoded_T_264[9], _decoded_decoded_T_264[7], _decoded_decoded_T_264[3:0] } = { io_rw_addr[2], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[10], io_rw_addr[11] };
  assign { _decoded_decoded_T_28[9:8], _decoded_decoded_T_28[6], _decoded_decoded_T_28[3:2] } = { io_rw_addr[2], io_rw_addr[3], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_30[11], _decoded_decoded_T_30[9:8], _decoded_decoded_T_30[6], _decoded_decoded_T_30[3:2] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[3], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_32[10:8], _decoded_decoded_T_32[6], _decoded_decoded_T_32[3:2] } = { io_rw_addr[1], io_rw_addr[2], io_rw_addr[3], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_34[11:8], _decoded_decoded_T_34[6], _decoded_decoded_T_34[3:2] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[2], io_rw_addr[3], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_36[7:6], _decoded_decoded_T_36[3:2] } = { io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_38[11], _decoded_decoded_T_38[7:6], _decoded_decoded_T_38[3:2] } = { io_rw_addr[0], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_4[9], _decoded_decoded_T_4[3:2] } = { io_rw_addr[2], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_40[10], _decoded_decoded_T_40[7:6], _decoded_decoded_T_40[3:2] } = { io_rw_addr[1], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_42[11:10], _decoded_decoded_T_42[7:6], _decoded_decoded_T_42[3:2] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_44[9], _decoded_decoded_T_44[7:6], _decoded_decoded_T_44[3:2] } = { io_rw_addr[2], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_46[11], _decoded_decoded_T_46[9], _decoded_decoded_T_46[7:6], _decoded_decoded_T_46[3:2] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_48[10:9], _decoded_decoded_T_48[7:6], _decoded_decoded_T_48[3:2] } = { io_rw_addr[1], io_rw_addr[2], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_50[11:9], _decoded_decoded_T_50[7:6], _decoded_decoded_T_50[3:2] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[2], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_52[8:6], _decoded_decoded_T_52[3:2] } = { io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_54[11], _decoded_decoded_T_54[8:6], _decoded_decoded_T_54[3:2] } = { io_rw_addr[0], io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_56[10], _decoded_decoded_T_56[8:6], _decoded_decoded_T_56[3:2] } = { io_rw_addr[1], io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_58[11:10], _decoded_decoded_T_58[8:6], _decoded_decoded_T_58[3:2] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_6[11], _decoded_decoded_T_6[9], _decoded_decoded_T_6[3:2] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_60[9:6], _decoded_decoded_T_60[3:2] } = { io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_62[11], _decoded_decoded_T_62[9:6], _decoded_decoded_T_62[3:2] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_64[10:6], _decoded_decoded_T_64[3:2] } = { io_rw_addr[1], io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_66[11:6], _decoded_decoded_T_66[3:2] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_68[5], _decoded_decoded_T_68[3:2] } = { io_rw_addr[6], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_70[11], _decoded_decoded_T_70[5], _decoded_decoded_T_70[3:2] } = { io_rw_addr[0], io_rw_addr[6], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_72[10], _decoded_decoded_T_72[5], _decoded_decoded_T_72[3:2] } = { io_rw_addr[1], io_rw_addr[6], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_74[11:10], _decoded_decoded_T_74[5], _decoded_decoded_T_74[3:2] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[6], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_76[9], _decoded_decoded_T_76[5], _decoded_decoded_T_76[3:2] } = { io_rw_addr[2], io_rw_addr[6], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_78[6], _decoded_decoded_T_78[4:2] } = { io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_8[6], _decoded_decoded_T_8[3:2] } = { io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_80[11], _decoded_decoded_T_80[6], _decoded_decoded_T_80[4:2] } = { io_rw_addr[0], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_82[10], _decoded_decoded_T_82[6], _decoded_decoded_T_82[4:2] } = { io_rw_addr[1], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_84[11:10], _decoded_decoded_T_84[6], _decoded_decoded_T_84[4:2] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_86[7:6], _decoded_decoded_T_86[4:2] } = { io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_88[11], _decoded_decoded_T_88[7:6], _decoded_decoded_T_88[4:2] } = { io_rw_addr[0], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_90[10], _decoded_decoded_T_90[7:6], _decoded_decoded_T_90[4:2] } = { io_rw_addr[1], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_92[11:10], _decoded_decoded_T_92[7:6], _decoded_decoded_T_92[4:2] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_94[9], _decoded_decoded_T_94[7:6], _decoded_decoded_T_94[4:2] } = { io_rw_addr[2], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_96[11], _decoded_decoded_T_96[9], _decoded_decoded_T_96[7:6], _decoded_decoded_T_96[4:2] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_98[10:9], _decoded_decoded_T_98[7:6], _decoded_decoded_T_98[4:2] } = { io_rw_addr[1], io_rw_addr[2], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign _decoded_decoded_orMatrixOutputs_T = _GEN_610[29];
  assign _decoded_decoded_orMatrixOutputs_T_2 = _GEN_609[0];
  assign _epc_T_1[0] = 1'h1;
  assign { _io_decode_0_read_illegal_T_12[7:6], _io_decode_0_read_illegal_T_12[4:1] } = { io_decode_0_inst[24], io_decode_0_inst[25], io_decode_0_inst[27], io_decode_0_inst[28], io_decode_0_inst[29], io_decode_0_inst[30] };
  assign _io_decode_0_read_illegal_T_17 = io_decode_0_read_illegal;
  assign _io_decode_0_read_illegal_T_21 = 1'h0;
  assign { _io_rw_rdata_T_1[31:30], _io_rw_rdata_T_1[28], _io_rw_rdata_T_1[26:24], _io_rw_rdata_T_1[22:13], _io_rw_rdata_T_1[11:9], _io_rw_rdata_T_1[5:3] } = 22'h000000;
  assign _io_rw_rdata_T_10[0] = 1'h0;
  assign _io_rw_rdata_T_107 = _GEN_596[31:0];
  assign _io_rw_rdata_T_108 = _GEN_597[31:0];
  assign _io_rw_rdata_T_109 = { _GEN_598[31], 2'h0, _GEN_598[28:23], 2'h0, _GEN_598[20:15], 2'h0, _GEN_598[12:7], 2'h0, _GEN_598[4:0] };
  assign _io_rw_rdata_T_110 = { _GEN_599[31], 2'h0, _GEN_599[28:23], 2'h0, _GEN_599[20:15], 2'h0, _GEN_599[12:7], 2'h0, _GEN_599[4:0] };
  assign _io_rw_rdata_T_113 = _GEN_600[29:0];
  assign _io_rw_rdata_T_114 = _GEN_601[29:0];
  assign _io_rw_rdata_T_115 = _GEN_602[29:0];
  assign _io_rw_rdata_T_116 = _GEN_603[29:0];
  assign _io_rw_rdata_T_117 = _GEN_604[29:0];
  assign _io_rw_rdata_T_118 = _GEN_605[29:0];
  assign _io_rw_rdata_T_119 = _GEN_606[29:0];
  assign _io_rw_rdata_T_120 = _GEN_607[29:0];
  assign _io_rw_rdata_T_129 = { 28'h0000000, _GEN_608[3], 3'h0 };
  assign _io_rw_rdata_T_13 = _GEN_593[0];
  assign _io_rw_rdata_T_130 = { 31'h00000000, _GEN_609[0] };
  assign _io_rw_rdata_T_132 = { 2'h0, _GEN_610[29], 8'h00, _GEN_610[29], _GEN_610[29], 6'h00, _GEN_610[29], 9'h000, _GEN_610[29], 2'h0 };
  assign { _io_rw_rdata_T_14[31], _io_rw_rdata_T_14[29:16], _io_rw_rdata_T_14[14:9], _io_rw_rdata_T_14[5:3] } = 24'h000000;
  assign { _io_rw_rdata_T_148[31:3], _io_rw_rdata_T_148[1] } = { _GEN_595[31:3], _GEN_595[1] };
  assign _io_rw_rdata_T_149 = _GEN_595[31:0];
  assign _io_rw_rdata_T_15[0] = 1'h0;
  assign _io_rw_rdata_T_17 = { _GEN_594[2], 1'h0, _GEN_594[0] };
  assign _io_rw_rdata_T_240[30] = io_rw_rdata[30];
  assign { _io_rw_rdata_T_241[30:29], _io_rw_rdata_T_241[22:21], _io_rw_rdata_T_241[14:13], _io_rw_rdata_T_241[6:5] } = { io_rw_rdata[30], _io_rw_rdata_T_240[29], _io_rw_rdata_T_240[22:21], _io_rw_rdata_T_240[14:13], _io_rw_rdata_T_240[6:5] };
  assign { _io_rw_rdata_T_242[31:29], _io_rw_rdata_T_242[22:21], _io_rw_rdata_T_242[14:13], _io_rw_rdata_T_242[6:5] } = { io_rw_rdata[31:30], _io_rw_rdata_T_240[29], _io_rw_rdata_T_240[22:21], _io_rw_rdata_T_240[14:13], _io_rw_rdata_T_240[6:5] };
  assign _io_rw_rdata_T_245[31:30] = io_rw_rdata[31:30];
  assign _io_rw_rdata_T_246[31:30] = io_rw_rdata[31:30];
  assign _io_rw_rdata_T_247[31:30] = io_rw_rdata[31:30];
  assign _io_rw_rdata_T_248[31:30] = io_rw_rdata[31:30];
  assign _io_rw_rdata_T_249[31:30] = io_rw_rdata[31:30];
  assign _io_rw_rdata_T_250[31:30] = io_rw_rdata[31:30];
  assign _io_rw_rdata_T_251[31:30] = io_rw_rdata[31:30];
  assign { _io_rw_rdata_T_252[31:30], _io_rw_rdata_T_252[28:21], _io_rw_rdata_T_252[18:13], _io_rw_rdata_T_252[11:4], _io_rw_rdata_T_252[1] } = { io_rw_rdata[31:30], io_rw_rdata[28:21], io_rw_rdata[18:13], io_rw_rdata[11:4], io_rw_rdata[1] };
  assign _io_rw_rdata_T_261[31:0] = { io_rw_rdata[31:30], _io_rw_rdata_T_252[29], io_rw_rdata[28:21], _io_rw_rdata_T_252[20:19], io_rw_rdata[18:13], _io_rw_rdata_T_252[12], io_rw_rdata[11:3], _io_rw_rdata_T_252[2], io_rw_rdata[1], _io_rw_rdata_T_252[0] };
  assign _io_rw_rdata_T_262[31:0] = { io_rw_rdata[31:30], _io_rw_rdata_T_252[29], io_rw_rdata[28:21], _io_rw_rdata_T_252[20:19], io_rw_rdata[18:13], _io_rw_rdata_T_252[12], io_rw_rdata[11:3], _io_rw_rdata_T_252[2], io_rw_rdata[1:0] };
  assign _io_rw_rdata_T_264[31:0] = io_rw_rdata;
  assign { _io_rw_rdata_T_4[31], _io_rw_rdata_T_4[29:24], _io_rw_rdata_T_4[22:13], _io_rw_rdata_T_4[11:9], _io_rw_rdata_T_4[7:3], _io_rw_rdata_T_4[1] } = 26'h0000000;
  assign { _io_rw_rdata_T_5[31:13], _io_rw_rdata_T_5[10:8], _io_rw_rdata_T_5[6:4], _io_rw_rdata_T_5[2:0] } = 28'h0000000;
  assign _io_rw_rdata_T_6[1] = 1'h0;
  assign _io_rw_rdata_T_7 = { 4'h0, _GEN_592[11], 3'h0, _GEN_592[7], 3'h0, _GEN_592[3], 3'h0 };
  assign { _io_rw_rdata_T_8[31:12], _io_rw_rdata_T_8[10:8], _io_rw_rdata_T_8[6:4], _io_rw_rdata_T_8[2:0] } = 29'h00000000;
  assign { _m_interrupts_T_3[31:12], _m_interrupts_T_3[10:8], _m_interrupts_T_3[6:4], _m_interrupts_T_3[2:0] } = 29'h1fffffff;
  assign { _m_interrupts_T_5[31:12], _m_interrupts_T_5[10:8], _m_interrupts_T_5[6:4], _m_interrupts_T_5[2:0] } = 29'h00000000;
  assign { _newBPC_T_2[31:28], _newBPC_T_2[26:13], _newBPC_T_2[11:9], _newBPC_T_2[6:3] } = { 2'h0, io_rw_cmd[1], 4'h0, io_rw_cmd[1], 13'h0000, io_rw_cmd[1], 3'h0 };
  assign { _newBPC_T_3[31:30], _newBPC_T_3[28], _newBPC_T_3[26:24], _newBPC_T_3[22:13], _newBPC_T_3[11:9], _newBPC_T_3[5:3] } = { io_rw_wdata[31:30], io_rw_wdata[28], io_rw_wdata[26:24], io_rw_wdata[22:13], io_rw_wdata[11:9], io_rw_wdata[5:3] };
  assign _new_mstatus_WIRE = { 73'h0000000000000000000, _T_2000[31:0] };
  assign { _notDebugTVec_T_1[31:7], _notDebugTVec_T_1[1:0] } = { reg_mtvec[31:7], 2'h0 };
  assign _pmp_mask_T_12[0] = reg_pmp_2_cfg_a[0];
  assign _pmp_mask_T_13[29:0] = { io_pmp_2_mask[31:3], reg_pmp_2_cfg_a[0] };
  assign _pmp_mask_T_14 = { _pmp_mask_T_13[30], io_pmp_2_mask[31:3], reg_pmp_2_cfg_a[0], 2'h3 };
  assign _pmp_mask_T_17[0] = reg_pmp_3_cfg_a[0];
  assign _pmp_mask_T_18[29:0] = { io_pmp_3_mask[31:3], reg_pmp_3_cfg_a[0] };
  assign _pmp_mask_T_19 = { _pmp_mask_T_18[30], io_pmp_3_mask[31:3], reg_pmp_3_cfg_a[0], 2'h3 };
  assign _pmp_mask_T_2[0] = reg_pmp_0_cfg_a[0];
  assign _pmp_mask_T_22[0] = reg_pmp_4_cfg_a[0];
  assign _pmp_mask_T_23[29:0] = { io_pmp_4_mask[31:3], reg_pmp_4_cfg_a[0] };
  assign _pmp_mask_T_24 = { _pmp_mask_T_23[30], io_pmp_4_mask[31:3], reg_pmp_4_cfg_a[0], 2'h3 };
  assign _pmp_mask_T_27[0] = reg_pmp_5_cfg_a[0];
  assign _pmp_mask_T_28[29:0] = { io_pmp_5_mask[31:3], reg_pmp_5_cfg_a[0] };
  assign _pmp_mask_T_29 = { _pmp_mask_T_28[30], io_pmp_5_mask[31:3], reg_pmp_5_cfg_a[0], 2'h3 };
  assign _pmp_mask_T_3[29:0] = { io_pmp_0_mask[31:3], reg_pmp_0_cfg_a[0] };
  assign _pmp_mask_T_32[0] = reg_pmp_6_cfg_a[0];
  assign _pmp_mask_T_33[29:0] = { io_pmp_6_mask[31:3], reg_pmp_6_cfg_a[0] };
  assign _pmp_mask_T_34 = { _pmp_mask_T_33[30], io_pmp_6_mask[31:3], reg_pmp_6_cfg_a[0], 2'h3 };
  assign _pmp_mask_T_37[0] = reg_pmp_7_cfg_a[0];
  assign _pmp_mask_T_38[29:0] = { io_pmp_7_mask[31:3], reg_pmp_7_cfg_a[0] };
  assign _pmp_mask_T_39 = { _pmp_mask_T_38[30], io_pmp_7_mask[31:3], reg_pmp_7_cfg_a[0], 2'h3 };
  assign _pmp_mask_T_4 = { _pmp_mask_T_3[30], io_pmp_0_mask[31:3], reg_pmp_0_cfg_a[0], 2'h3 };
  assign _pmp_mask_T_7[0] = reg_pmp_1_cfg_a[0];
  assign _pmp_mask_T_8[29:0] = { io_pmp_1_mask[31:3], reg_pmp_1_cfg_a[0] };
  assign _pmp_mask_T_9 = { _pmp_mask_T_8[30], io_pmp_1_mask[31:3], reg_pmp_1_cfg_a[0], 2'h3 };
  assign _read_mip_T = { 4'h0, io_interrupts_meip, 3'h0, io_interrupts_mtip, 3'h0, io_interrupts_msip, 3'h0 };
  assign _read_mstatus_T = { reg_debug, io_status_cease_r, reg_wfi, 19'h20400, reg_misa[12], 9'h020, reg_misa[2], 1'h0, reg_misa[0], 31'h6c000000, reg_mstatus_gva, 30'h00000018, reg_mstatus_mpie, 3'h0, reg_mstatus_mie, 3'h0 };
  assign _read_mtvec_T_1 = { reg_mtvec[0], reg_mtvec[0], reg_mtvec[0], reg_mtvec[0], reg_mtvec[0], 2'h2 };
  assign _read_mtvec_T_3 = { 25'h0000000, reg_mtvec[0], reg_mtvec[0], reg_mtvec[0], reg_mtvec[0], reg_mtvec[0], 2'h2 };
  assign { _read_mtvec_T_4[31:7], _read_mtvec_T_4[5:0] } = { 25'h1ffffff, _read_mtvec_T_4[6], _read_mtvec_T_4[6], _read_mtvec_T_4[6], _read_mtvec_T_4[6], 2'h1 };
  assign _reg_custom_0_T = { 28'h0000000, _T_2000[3], 3'h0 };
  assign _reg_custom_0_T_2 = 32'd0;
  assign _reg_custom_0_T_3 = { 28'h0000000, _T_2000[3], 3'h0 };
  assign _reg_dcsr_cause_T_2[2] = reg_singleStepped;
  assign _reg_mcause_T = { _T_2000[31], 27'h0000000, _T_2000[3:0] };
  assign _reg_mcountinhibit_T_1 = { _T_2000[31:2], 1'h0, _T_2000[0] };
  assign { _reg_mepc_T_1[5], _reg_mepc_T_1[0] } = { _GEN_611[3], 1'h1 };
  assign _reg_mepc_T_2 = { _T_2000[31:1], 1'h0 };
  assign _reg_mie_T = { 20'h00000, _T_2000[11], 3'h0, _T_2000[7], 3'h0, _T_2000[3], 3'h0 };
  assign _reg_misa_T[31:1] = { _reg_mepc_T_1[31:6], _GEN_611[3], _reg_mepc_T_1[4:1] };
  assign _reg_misa_T_1 = _GEN_611[3];
  assign _reg_misa_T_2 = { _GEN_611[3], 3'h0 };
  assign { _reg_misa_T_3[31:4], _reg_misa_T_3[2:0] } = { _reg_mepc_T_1[31:6], _GEN_611[3], _reg_mepc_T_1[4], _reg_mepc_T_1[2:1], _reg_misa_T[0] };
  assign { _reg_misa_T_4[31:4], _reg_misa_T_4[2:0] } = { _T_2000[31:4], _T_2000[2:0] };
  assign _reg_misa_T_5 = { 19'h00000, _T_2000[12], 9'h000, _T_2000[2], 1'h0, _T_2000[0] };
  assign _reg_misa_T_7 = 32'd1082130688;
  assign _reg_misa_T_8 = { 19'h20400, _T_2000[12], 9'h020, _T_2000[2], 1'h0, _T_2000[0] };
  assign _which_T_100 = 4'h4;
  assign _which_T_101 = 4'h4;
  assign _which_T_102 = 4'h4;
  assign { _which_T_103[3:2], _which_T_103[0] } = { 2'h1, _which_T_103[1] };
  assign { _which_T_104[3], _which_T_104[0] } = { 1'h0, _which_T_104[1] };
  assign _which_T_105[0] = _which_T_105[1];
  assign _which_T_106 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_107 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_108 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_109 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_111 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_112 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_113 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_114 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_115 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_116 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_117 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_118 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_119 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_120 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_121 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_122 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_123 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_124 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_95 = 4'h4;
  assign _which_T_96 = 4'h4;
  assign _which_T_97 = 4'h4;
  assign _which_T_98 = 4'h4;
  assign _which_T_99 = 4'h4;
  assign addr = { 1'h0, io_rw_addr };
  assign addr_1 = io_decode_0_inst[31:20];
  assign d_interrupts = { io_interrupts_debug, 14'h0000 };
  assign { debugTVec[11:4], debugTVec[2:0] } = 11'h400;
  assign decoded_130 = _GEN_609[0];
  assign decoded_132 = _GEN_610[29];
  assign decoded_andMatrixInput_0_1 = io_rw_addr[0];
  assign decoded_andMatrixInput_0_10 = io_decode_0_inst[22];
  assign decoded_andMatrixInput_0_11 = io_decode_0_inst[30];
  assign decoded_andMatrixInput_0_2 = io_rw_addr[8];
  assign decoded_andMatrixInput_0_4 = io_rw_addr[2];
  assign decoded_andMatrixInput_0_5 = io_rw_addr[10];
  assign decoded_andMatrixInput_0_7 = io_decode_0_inst[20];
  assign decoded_andMatrixInput_0_8 = io_decode_0_inst[28];
  assign decoded_andMatrixInput_7_2 = io_rw_addr[9];
  assign decoded_andMatrixInput_7_6 = io_decode_0_inst[29];
  assign decoded_decoded_andMatrixInput_0_1 = io_rw_addr[0];
  assign decoded_decoded_andMatrixInput_0_5 = io_rw_addr[1];
  assign decoded_decoded_andMatrixInput_10_58 = io_rw_addr[10];
  assign decoded_decoded_andMatrixInput_10_65 = io_rw_addr[11];
  assign decoded_decoded_andMatrixInput_2_2 = io_rw_addr[2];
  assign decoded_decoded_andMatrixInput_3_10 = io_rw_addr[3];
  assign decoded_decoded_andMatrixInput_4_18 = io_rw_addr[4];
  assign decoded_decoded_andMatrixInput_4_4 = io_rw_addr[5];
  assign decoded_decoded_andMatrixInput_6_34 = io_rw_addr[6];
  assign decoded_decoded_andMatrixInput_7_39 = io_rw_addr[7];
  assign decoded_decoded_andMatrixInput_8 = io_rw_addr[8];
  assign decoded_decoded_andMatrixInput_9 = io_rw_addr[9];
  assign { decoded_decoded_invMatrixOutputs[2], decoded_decoded_invMatrixOutputs[0] } = { _GEN_609[0], _GEN_610[29] };
  assign { decoded_decoded_invMatrixOutputs_lo_lo[2], decoded_decoded_invMatrixOutputs_lo_lo[0] } = { _GEN_609[0], _GEN_610[29] };
  assign { decoded_decoded_invMatrixOutputs_lo_lo_lo_lo[2], decoded_decoded_invMatrixOutputs_lo_lo_lo_lo[0] } = { _GEN_609[0], _GEN_610[29] };
  assign decoded_decoded_lo[3:2] = { io_rw_addr[8], io_rw_addr[9] };
  assign decoded_decoded_lo_129[3:0] = { io_rw_addr[8], io_rw_addr[9], io_rw_addr[10], io_rw_addr[11] };
  assign decoded_decoded_lo_130[3:0] = { io_rw_addr[8], io_rw_addr[9], io_rw_addr[10], io_rw_addr[11] };
  assign { decoded_decoded_lo_34[5], decoded_decoded_lo_34[3:2] } = { io_rw_addr[6], io_rw_addr[8], io_rw_addr[9] };
  assign decoded_decoded_lo_39[4:2] = { io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign decoded_decoded_lo_4[3:2] = { io_rw_addr[8], io_rw_addr[9] };
  assign decoded_decoded_lo_59[4:1] = { io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[10] };
  assign decoded_decoded_lo_65[4:1] = { io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[10] };
  assign { decoded_decoded_lo_67[3:2], decoded_decoded_lo_67[0] } = { io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { decoded_decoded_lo_68[3:2], decoded_decoded_lo_68[0] } = { io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { decoded_decoded_lo_98[4:2], decoded_decoded_lo_98[0] } = { io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { decoded_decoded_lo_99[4:2], decoded_decoded_lo_99[0] } = { io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { decoded_decoded_orMatrixOutputs[2], decoded_decoded_orMatrixOutputs[0] } = { _GEN_609[0], _GEN_610[29] };
  assign { decoded_decoded_orMatrixOutputs_lo_lo[2], decoded_decoded_orMatrixOutputs_lo_lo[0] } = { _GEN_609[0], _GEN_610[29] };
  assign { decoded_decoded_orMatrixOutputs_lo_lo_lo_lo[2], decoded_decoded_orMatrixOutputs_lo_lo_lo_lo[0] } = { _GEN_609[0], _GEN_610[29] };
  assign decoded_decoded_plaInput = io_rw_addr;
  assign decoded_invInputs[19:0] = 20'hfff8c;
  assign decoded_invMatrixOutputs[3:0] = 4'h0;
  assign decoded_invMatrixOutputs_1[3:0] = 4'h0;
  assign decoded_orMatrixOutputs[3:0] = 4'h0;
  assign decoded_orMatrixOutputs_1[3:0] = 4'h0;
  assign decoded_plaInput = { io_rw_addr, 20'h00073 };
  assign epc = { io_pc[31:1], 1'h0 };
  assign exception = io_trace_0_exception;
  assign f = _T_2000[5];
  assign io_bp_0_address = reg_bp_0_address;
  assign io_bp_0_control_action = reg_bp_0_control_action;
  assign io_bp_0_control_r = reg_bp_0_control_r;
  assign io_bp_0_control_tmatch = reg_bp_0_control_tmatch;
  assign io_bp_0_control_w = reg_bp_0_control_w;
  assign io_bp_0_control_x = reg_bp_0_control_x;
  assign io_customCSRs_0_value = { 28'h0000000, reg_custom_0[3], 3'h0 };
  assign io_decode_0_fp_csr = 1'h0;
  assign io_decode_0_fp_illegal = 1'h1;
  assign io_decode_0_read_illegal_andMatrixInput_0 = io_decode_0_inst[24];
  assign io_decode_0_read_illegal_andMatrixInput_1 = io_decode_0_inst[25];
  assign io_decode_0_read_illegal_andMatrixInput_3 = io_decode_0_inst[27];
  assign io_decode_0_read_illegal_andMatrixInput_4 = io_decode_0_inst[28];
  assign io_decode_0_read_illegal_andMatrixInput_5 = io_decode_0_inst[29];
  assign io_decode_0_read_illegal_andMatrixInput_6 = io_decode_0_inst[30];
  assign io_decode_0_rocc_illegal = 1'h1;
  assign io_decode_0_write_flush_addr_m = { io_decode_0_inst[31:30], 2'h3, io_decode_0_inst[27:20] };
  assign io_evec[0] = 1'h0;
  assign io_inhibit_cycle = reg_mcountinhibit[0];
  assign io_interrupt_cause[31:4] = 28'h8000000;
  assign io_pmp_0_addr = reg_pmp_0_addr;
  assign io_pmp_0_cfg_a = reg_pmp_0_cfg_a;
  assign io_pmp_0_cfg_l = reg_pmp_0_cfg_l;
  assign io_pmp_0_cfg_r = reg_pmp_0_cfg_r;
  assign io_pmp_0_cfg_w = reg_pmp_0_cfg_w;
  assign io_pmp_0_cfg_x = reg_pmp_0_cfg_x;
  assign io_pmp_0_mask[2:0] = { reg_pmp_0_cfg_a[0], 2'h3 };
  assign io_pmp_1_addr = reg_pmp_1_addr;
  assign io_pmp_1_cfg_a = reg_pmp_1_cfg_a;
  assign io_pmp_1_cfg_l = reg_pmp_1_cfg_l;
  assign io_pmp_1_cfg_r = reg_pmp_1_cfg_r;
  assign io_pmp_1_cfg_w = reg_pmp_1_cfg_w;
  assign io_pmp_1_cfg_x = reg_pmp_1_cfg_x;
  assign io_pmp_1_mask[2:0] = { reg_pmp_1_cfg_a[0], 2'h3 };
  assign io_pmp_2_addr = reg_pmp_2_addr;
  assign io_pmp_2_cfg_a = reg_pmp_2_cfg_a;
  assign io_pmp_2_cfg_l = reg_pmp_2_cfg_l;
  assign io_pmp_2_cfg_r = reg_pmp_2_cfg_r;
  assign io_pmp_2_cfg_w = reg_pmp_2_cfg_w;
  assign io_pmp_2_cfg_x = reg_pmp_2_cfg_x;
  assign io_pmp_2_mask[2:0] = { reg_pmp_2_cfg_a[0], 2'h3 };
  assign io_pmp_3_addr = reg_pmp_3_addr;
  assign io_pmp_3_cfg_a = reg_pmp_3_cfg_a;
  assign io_pmp_3_cfg_l = reg_pmp_3_cfg_l;
  assign io_pmp_3_cfg_r = reg_pmp_3_cfg_r;
  assign io_pmp_3_cfg_w = reg_pmp_3_cfg_w;
  assign io_pmp_3_cfg_x = reg_pmp_3_cfg_x;
  assign io_pmp_3_mask[2:0] = { reg_pmp_3_cfg_a[0], 2'h3 };
  assign io_pmp_4_addr = reg_pmp_4_addr;
  assign io_pmp_4_cfg_a = reg_pmp_4_cfg_a;
  assign io_pmp_4_cfg_l = reg_pmp_4_cfg_l;
  assign io_pmp_4_cfg_r = reg_pmp_4_cfg_r;
  assign io_pmp_4_cfg_w = reg_pmp_4_cfg_w;
  assign io_pmp_4_cfg_x = reg_pmp_4_cfg_x;
  assign io_pmp_4_mask[2:0] = { reg_pmp_4_cfg_a[0], 2'h3 };
  assign io_pmp_5_addr = reg_pmp_5_addr;
  assign io_pmp_5_cfg_a = reg_pmp_5_cfg_a;
  assign io_pmp_5_cfg_l = reg_pmp_5_cfg_l;
  assign io_pmp_5_cfg_r = reg_pmp_5_cfg_r;
  assign io_pmp_5_cfg_w = reg_pmp_5_cfg_w;
  assign io_pmp_5_cfg_x = reg_pmp_5_cfg_x;
  assign io_pmp_5_mask[2:0] = { reg_pmp_5_cfg_a[0], 2'h3 };
  assign io_pmp_6_addr = reg_pmp_6_addr;
  assign io_pmp_6_cfg_a = reg_pmp_6_cfg_a;
  assign io_pmp_6_cfg_l = reg_pmp_6_cfg_l;
  assign io_pmp_6_cfg_r = reg_pmp_6_cfg_r;
  assign io_pmp_6_cfg_w = reg_pmp_6_cfg_w;
  assign io_pmp_6_cfg_x = reg_pmp_6_cfg_x;
  assign io_pmp_6_mask[2:0] = { reg_pmp_6_cfg_a[0], 2'h3 };
  assign io_pmp_7_addr = reg_pmp_7_addr;
  assign io_pmp_7_cfg_a = reg_pmp_7_cfg_a;
  assign io_pmp_7_cfg_l = reg_pmp_7_cfg_l;
  assign io_pmp_7_cfg_r = reg_pmp_7_cfg_r;
  assign io_pmp_7_cfg_w = reg_pmp_7_cfg_w;
  assign io_pmp_7_cfg_x = reg_pmp_7_cfg_x;
  assign io_pmp_7_mask[2:0] = { reg_pmp_7_cfg_a[0], 2'h3 };
  assign io_status_cease = io_status_cease_r;
  assign io_status_debug = reg_debug;
  assign io_status_dprv = 2'h3;
  assign io_status_dv = 1'h0;
  assign io_status_fs = 2'h0;
  assign io_status_gva = reg_mstatus_gva;
  assign io_status_hie = 1'h0;
  assign io_status_isa = { 19'h20400, reg_misa[12], 9'h020, reg_misa[2], 1'h0, reg_misa[0] };
  assign io_status_mbe = 1'h0;
  assign io_status_mie = reg_mstatus_mie;
  assign io_status_mpie = reg_mstatus_mpie;
  assign io_status_mpp = 2'h3;
  assign io_status_mprv = 1'h0;
  assign io_status_mpv = 1'h0;
  assign io_status_mxr = 1'h0;
  assign io_status_prv = 2'h3;
  assign io_status_sbe = 1'h0;
  assign io_status_sd = 1'h0;
  assign io_status_sd_rv32 = 1'h0;
  assign io_status_sie = 1'h0;
  assign io_status_spie = 1'h0;
  assign io_status_spp = 1'h0;
  assign io_status_sum = 1'h0;
  assign io_status_sxl = 2'h0;
  assign io_status_tsr = 1'h0;
  assign io_status_tvm = 1'h0;
  assign io_status_tw = 1'h0;
  assign io_status_ube = 1'h0;
  assign io_status_uie = 1'h0;
  assign io_status_upie = 1'h0;
  assign io_status_uxl = 2'h0;
  assign io_status_v = 1'h0;
  assign io_status_vs = 2'h0;
  assign io_status_wfi = reg_wfi;
  assign io_status_xs = 2'h0;
  assign io_status_zero1 = 8'h00;
  assign io_status_zero2 = 23'h000000;
  assign io_time = { large_1[25:0], small_1 };
  assign io_trace_0_iaddr = io_pc;
  assign io_trace_0_insn = io_inst_0;
  assign lo_11 = { reg_pmp_1_cfg_l, 2'h0, reg_pmp_1_cfg_a, reg_pmp_1_cfg_x, reg_pmp_1_cfg_w, reg_pmp_1_cfg_r, reg_pmp_0_cfg_l, 2'h0, reg_pmp_0_cfg_a, reg_pmp_0_cfg_x, reg_pmp_0_cfg_w, reg_pmp_0_cfg_r };
  assign lo_16 = { reg_pmp_5_cfg_l, 2'h0, reg_pmp_5_cfg_a, reg_pmp_5_cfg_x, reg_pmp_5_cfg_w, reg_pmp_5_cfg_r, reg_pmp_4_cfg_l, 2'h0, reg_pmp_4_cfg_a, reg_pmp_4_cfg_x, reg_pmp_4_cfg_w, reg_pmp_4_cfg_r };
  assign lo_4 = { 4'h8, reg_bp_0_control_x, reg_bp_0_control_w, reg_bp_0_control_r };
  assign { m_interrupts[31:4], m_interrupts[2:0] } = { 20'h00000, _which_T_105[3], 3'h0, _which_T_103[1], 6'h00 };
  assign newCfg_1_a = _T_2000[12:11];
  assign newCfg_1_l = _T_2000[15];
  assign newCfg_1_r = _T_2000[8];
  assign newCfg_1_w = _T_2000[9];
  assign newCfg_1_x = _T_2000[10];
  assign newCfg_2_a = _T_2000[20:19];
  assign newCfg_2_l = _T_2000[23];
  assign newCfg_2_r = _T_2000[16];
  assign newCfg_2_w = _T_2000[17];
  assign newCfg_2_x = _T_2000[18];
  assign newCfg_3_a = _T_2000[28:27];
  assign newCfg_3_l = _T_2000[31];
  assign newCfg_3_r = _T_2000[24];
  assign newCfg_3_w = _T_2000[25];
  assign newCfg_3_x = _T_2000[26];
  assign newCfg_a = _T_2000[4:3];
  assign newCfg_l = _T_2000[7];
  assign newCfg_r = _T_2000[0];
  assign newCfg_w = _T_2000[1];
  assign newCfg_x = _T_2000[2];
  assign new_dcsr_ebreakm = _T_2000[15];
  assign new_mstatus_mie = _T_2000[3];
  assign new_mstatus_mpie = _T_2000[7];
  assign { notDebugTVec[31:7], notDebugTVec[1:0] } = { reg_mtvec[31:7], 2'h0 };
  assign notDebugTVec_interruptOffset[1:0] = 2'h0;
  assign { notDebugTVec_interruptVec[31:7], notDebugTVec_interruptVec[1:0] } = { reg_mtvec[31:7], 2'h0 };
  assign pending_interrupts = { 20'h00000, _m_interrupts_T_5[11], 3'h0, _m_interrupts_T_5[7], 3'h0, _m_interrupts_T_5[3], 3'h0 };
  assign pmp_mask_base = { reg_pmp_0_addr, reg_pmp_0_cfg_a[0] };
  assign pmp_mask_base_1 = { reg_pmp_1_addr, reg_pmp_1_cfg_a[0] };
  assign pmp_mask_base_2 = { reg_pmp_2_addr, reg_pmp_2_cfg_a[0] };
  assign pmp_mask_base_3 = { reg_pmp_3_addr, reg_pmp_3_cfg_a[0] };
  assign pmp_mask_base_4 = { reg_pmp_4_addr, reg_pmp_4_cfg_a[0] };
  assign pmp_mask_base_5 = { reg_pmp_5_addr, reg_pmp_5_cfg_a[0] };
  assign pmp_mask_base_6 = { reg_pmp_6_addr, reg_pmp_6_cfg_a[0] };
  assign pmp_mask_base_7 = { reg_pmp_7_addr, reg_pmp_7_cfg_a[0] };
  assign read_mip = { 4'h0, io_interrupts_meip, 3'h0, io_interrupts_mtip, 3'h0, io_interrupts_msip, 3'h0 };
  assign read_mstatus = { 24'h000018, reg_mstatus_mpie, 3'h0, reg_mstatus_mie, 3'h0 };
  assign read_mstatus_hi = { reg_debug, io_status_cease_r, reg_wfi, 19'h20400, reg_misa[12], 9'h020, reg_misa[2], 1'h0, reg_misa[0], 31'h6c000000, reg_mstatus_gva, 16'h0000 };
  assign read_mstatus_hi_hi = { reg_debug, io_status_cease_r, reg_wfi, 19'h20400, reg_misa[12], 9'h020, reg_misa[2], 1'h0, reg_misa[0], 30'h36000000 };
  assign read_mstatus_lo = { 14'h0018, reg_mstatus_mpie, 3'h0, reg_mstatus_mie, 3'h0 };
  assign read_mstatus_lo_lo = { 1'h0, reg_mstatus_mpie, 3'h0, reg_mstatus_mie, 3'h0 };
  assign read_mtvec = { reg_mtvec[31:7], _notDebugTVec_T_1[6:2], 1'h0, reg_mtvec[0] };
  assign { reg_custom_0[31:4], reg_custom_0[2:0] } = 31'h00000000;
  assign reg_mcountinhibit[1] = 1'h0;
  assign { reg_mie[31:12], reg_mie[10:8], reg_mie[6:4], reg_mie[2:0] } = 29'h00000000;
  assign { reg_misa[31:13], reg_misa[11:3], reg_misa[1] } = 29'h08100040;
  assign reg_mstatus_spp = 1'h0;
  assign tvec[1:0] = 2'h0;
  assign value = { large_, small_ };
  assign value_1 = { large_1, small_1 };
  assign wdata = _T_2000[31:0];
  assign whichInterrupt = io_interrupt_cause[3:0];
  assign x79 = reg_mcountinhibit[2];
  assign x86 = _GEN_35[0];
endmodule
module IBuf(clock, reset, io_imem_ready, io_imem_valid, io_imem_bits_pc, io_imem_bits_data, io_imem_bits_xcpt_ae_inst, io_imem_bits_replay, io_kill, io_pc, io_inst_0_ready, io_inst_0_valid, io_inst_0_bits_xcpt0_ae_inst, io_inst_0_bits_xcpt1_pf_inst, io_inst_0_bits_xcpt1_gf_inst, io_inst_0_bits_xcpt1_ae_inst, io_inst_0_bits_replay, io_inst_0_bits_rvc, io_inst_0_bits_inst_bits, io_inst_0_bits_inst_rd, io_inst_0_bits_inst_rs1
, io_inst_0_bits_inst_rs2, io_inst_0_bits_raw);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  wire _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire _272_;
  wire _273_;
  wire _274_;
  wire _275_;
  wire _276_;
  wire _277_;
  wire _278_;
  wire _279_;
  wire _280_;
  wire _281_;
  wire _282_;
  wire _283_;
  wire _284_;
  wire _285_;
  wire _286_;
  wire _287_;
  wire _288_;
  wire _289_;
  wire _290_;
  wire _291_;
  wire _292_;
  wire _293_;
  wire _294_;
  wire _295_;
  wire _296_;
  wire _297_;
  wire _298_;
  wire _299_;
  wire _300_;
  wire _301_;
  wire _302_;
  wire _303_;
  wire _304_;
  wire _305_;
  wire _306_;
  wire _307_;
  wire _308_;
  wire _309_;
  wire _310_;
  wire _311_;
  wire _312_;
  wire _313_;
  wire _314_;
  wire _315_;
  wire _316_;
  wire _317_;
  wire _318_;
  wire _319_;
  wire _320_;
  wire _321_;
  wire _322_;
  wire _323_;
  wire _324_;
  wire _325_;
  wire _326_;
  wire _327_;
  wire _328_;
  wire _329_;
  wire _330_;
  wire _331_;
  wire _332_;
  wire _333_;
  wire _334_;
  wire _335_;
  wire _336_;
  wire _337_;
  wire _338_;
  wire _339_;
  wire _340_;
  wire _341_;
  wire _342_;
  wire _343_;
  wire _344_;
  wire _345_;
  wire _346_;
  wire _347_;
  wire _348_;
  wire _349_;
  wire _350_;
  wire _351_;
  wire _352_;
  wire _353_;
  wire _354_;
  wire _355_;
  wire _356_;
  wire _357_;
  wire _358_;
  wire _359_;
  wire _360_;
  wire _361_;
  wire _362_;
  wire _363_;
  wire _364_;
  wire _365_;
  wire _366_;
  wire _367_;
  wire _368_;
  wire _369_;
  wire _370_;
  wire _371_;
  wire _372_;
  wire [190:0] _GEN_1;
  wire [1:0] _GEN_58;
  wire [1:0] _GEN_59;
  wire [31:0] _GEN_67;
  wire [1:0] _bufMask_T;
  wire [5:0] _buf_data_T;
  wire [31:0] _buf_pc_T_1;
  wire [2:0] _buf_pc_T_2;
  wire [31:0] _buf_pc_T_4;
  wire [31:0] _buf_pc_T_5;
  wire [31:0] _buf_pc_T_6;
  wire [1:0] _full_insn_T_2;
  wire [63:0] _icData_T_2;
  wire [5:0] _icData_T_3;
  wire [190:0] _icData_T_4;
  wire [4:0] _icMask_T_1;
  wire [62:0] _icMask_T_2;
  wire [1:0] _icShiftAmt_T_1;
  wire [1:0] _ic_replay_T;
  wire [1:0] _ic_replay_T_1;
  wire [31:0] _inst_T;
  wire [31:0] _inst_T_1;
  wire [31:0] _inst_T_2;
  wire [2:0] _io_inst_0_bits_xcpt1_T_4;
  wire [2:0] _io_inst_0_bits_xcpt1_T_5;
  wire [1:0] _nReady_T_4;
  wire [1:0] _replay_T_5;
  wire [3:0] _valid_T_2;
  wire [1:0] bufMask;
  wire [31:0] buf__data;
  wire [31:0] buf__pc;
  wire buf__replay;
  wire buf__xcpt_ae_inst;
  wire [63:0] buf_data_data;
  wire [1:0] buf_replay;
  input clock;
  wire clock;
  wire [31:0] exp_io_in;
  wire [31:0] exp_io_out_bits;
  wire [4:0] exp_io_out_rd;
  wire [4:0] exp_io_out_rs1;
  wire [4:0] exp_io_out_rs2;
  wire exp_io_rvc;
  wire [31:0] icData;
  wire [127:0] icData_data;
  wire [31:0] icMask;
  wire [1:0] icShiftAmt;
  input [31:0] io_imem_bits_data;
  wire [31:0] io_imem_bits_data;
  input [31:0] io_imem_bits_pc;
  wire [31:0] io_imem_bits_pc;
  input io_imem_bits_replay;
  wire io_imem_bits_replay;
  input io_imem_bits_xcpt_ae_inst;
  wire io_imem_bits_xcpt_ae_inst;
  output io_imem_ready;
  wire io_imem_ready;
  input io_imem_valid;
  wire io_imem_valid;
  output [31:0] io_inst_0_bits_inst_bits;
  wire [31:0] io_inst_0_bits_inst_bits;
  output [4:0] io_inst_0_bits_inst_rd;
  wire [4:0] io_inst_0_bits_inst_rd;
  output [4:0] io_inst_0_bits_inst_rs1;
  wire [4:0] io_inst_0_bits_inst_rs1;
  output [4:0] io_inst_0_bits_inst_rs2;
  wire [4:0] io_inst_0_bits_inst_rs2;
  output [31:0] io_inst_0_bits_raw;
  wire [31:0] io_inst_0_bits_raw;
  output io_inst_0_bits_replay;
  wire io_inst_0_bits_replay;
  output io_inst_0_bits_rvc;
  wire io_inst_0_bits_rvc;
  output io_inst_0_bits_xcpt0_ae_inst;
  wire io_inst_0_bits_xcpt0_ae_inst;
  output io_inst_0_bits_xcpt1_ae_inst;
  wire io_inst_0_bits_xcpt1_ae_inst;
  output io_inst_0_bits_xcpt1_gf_inst;
  wire io_inst_0_bits_xcpt1_gf_inst;
  output io_inst_0_bits_xcpt1_pf_inst;
  wire io_inst_0_bits_xcpt1_pf_inst;
  input io_inst_0_ready;
  wire io_inst_0_ready;
  output io_inst_0_valid;
  wire io_inst_0_valid;
  input io_kill;
  wire io_kill;
  output [31:0] io_pc;
  wire [31:0] io_pc;
  wire nBufValid;
  wire [1:0] nIC;
  wire [1:0] nICReady;
  wire pcWordBits;
  input reset;
  wire reset;
  wire [1:0] shamt;
  wire [1:0] valid;
  wire xcpt_1_ae_inst;
  INV_X1 _373_ (
    .A(nBufValid),
    .ZN(_051_)
  );
  INV_X1 _374_ (
    .A(buf__pc[1]),
    .ZN(_052_)
  );
  INV_X1 _375_ (
    .A(reset),
    .ZN(_053_)
  );
  INV_X1 _376_ (
    .A(io_kill),
    .ZN(_054_)
  );
  INV_X1 _377_ (
    .A(io_imem_bits_pc[1]),
    .ZN(_055_)
  );
  INV_X1 _378_ (
    .A(io_imem_valid),
    .ZN(_056_)
  );
  INV_X1 _379_ (
    .A(exp_io_rvc),
    .ZN(_057_)
  );
  INV_X1 _380_ (
    .A(_bufMask_T[0]),
    .ZN(_058_)
  );
  INV_X1 _381_ (
    .A(io_imem_bits_data[0]),
    .ZN(_059_)
  );
  INV_X1 _382_ (
    .A(io_imem_bits_data[16]),
    .ZN(_060_)
  );
  INV_X1 _383_ (
    .A(io_imem_bits_data[1]),
    .ZN(_061_)
  );
  INV_X1 _384_ (
    .A(io_imem_bits_data[17]),
    .ZN(_062_)
  );
  INV_X1 _385_ (
    .A(io_imem_bits_data[2]),
    .ZN(_063_)
  );
  INV_X1 _386_ (
    .A(io_imem_bits_data[18]),
    .ZN(_064_)
  );
  INV_X1 _387_ (
    .A(io_imem_bits_data[3]),
    .ZN(_065_)
  );
  INV_X1 _388_ (
    .A(io_imem_bits_data[19]),
    .ZN(_066_)
  );
  INV_X1 _389_ (
    .A(io_imem_bits_data[4]),
    .ZN(_067_)
  );
  INV_X1 _390_ (
    .A(io_imem_bits_data[20]),
    .ZN(_068_)
  );
  INV_X1 _391_ (
    .A(io_imem_bits_data[5]),
    .ZN(_069_)
  );
  INV_X1 _392_ (
    .A(io_imem_bits_data[21]),
    .ZN(_070_)
  );
  INV_X1 _393_ (
    .A(io_imem_bits_data[6]),
    .ZN(_071_)
  );
  INV_X1 _394_ (
    .A(io_imem_bits_data[22]),
    .ZN(_072_)
  );
  INV_X1 _395_ (
    .A(io_imem_bits_data[7]),
    .ZN(_073_)
  );
  INV_X1 _396_ (
    .A(io_imem_bits_data[23]),
    .ZN(_074_)
  );
  INV_X1 _397_ (
    .A(io_imem_bits_data[8]),
    .ZN(_075_)
  );
  INV_X1 _398_ (
    .A(io_imem_bits_data[24]),
    .ZN(_076_)
  );
  INV_X1 _399_ (
    .A(io_imem_bits_data[9]),
    .ZN(_077_)
  );
  INV_X1 _400_ (
    .A(io_imem_bits_data[25]),
    .ZN(_078_)
  );
  INV_X1 _401_ (
    .A(io_imem_bits_data[10]),
    .ZN(_079_)
  );
  INV_X1 _402_ (
    .A(io_imem_bits_data[26]),
    .ZN(_080_)
  );
  INV_X1 _403_ (
    .A(io_imem_bits_data[11]),
    .ZN(_081_)
  );
  INV_X1 _404_ (
    .A(io_imem_bits_data[27]),
    .ZN(_082_)
  );
  INV_X1 _405_ (
    .A(io_imem_bits_data[12]),
    .ZN(_083_)
  );
  INV_X1 _406_ (
    .A(io_imem_bits_data[28]),
    .ZN(_084_)
  );
  INV_X1 _407_ (
    .A(io_imem_bits_data[13]),
    .ZN(_085_)
  );
  INV_X1 _408_ (
    .A(io_imem_bits_data[29]),
    .ZN(_086_)
  );
  INV_X1 _409_ (
    .A(io_imem_bits_data[14]),
    .ZN(_087_)
  );
  INV_X1 _410_ (
    .A(io_imem_bits_data[30]),
    .ZN(_088_)
  );
  INV_X1 _411_ (
    .A(io_imem_bits_data[15]),
    .ZN(_089_)
  );
  INV_X1 _412_ (
    .A(io_imem_bits_data[31]),
    .ZN(_090_)
  );
  AND2_X1 _413_ (
    .A1(_051_),
    .A2(io_imem_bits_pc[1]),
    .ZN(_091_)
  );
  INV_X1 _414_ (
    .A(_091_),
    .ZN(_092_)
  );
  AND2_X1 _415_ (
    .A1(io_imem_valid),
    .A2(_092_),
    .ZN(_093_)
  );
  INV_X1 _416_ (
    .A(_093_),
    .ZN(_094_)
  );
  AND2_X1 _417_ (
    .A1(nBufValid),
    .A2(buf__replay),
    .ZN(_095_)
  );
  INV_X1 _418_ (
    .A(_095_),
    .ZN(_096_)
  );
  AND2_X1 _419_ (
    .A1(_057_),
    .A2(_096_),
    .ZN(_097_)
  );
  AND2_X1 _420_ (
    .A1(_094_),
    .A2(_097_),
    .ZN(_098_)
  );
  INV_X1 _421_ (
    .A(_098_),
    .ZN(_099_)
  );
  AND2_X1 _422_ (
    .A1(_058_),
    .A2(_098_),
    .ZN(_100_)
  );
  INV_X1 _423_ (
    .A(_100_),
    .ZN(_101_)
  );
  AND2_X1 _424_ (
    .A1(_057_),
    .A2(_bufMask_T[0]),
    .ZN(_102_)
  );
  INV_X1 _425_ (
    .A(_102_),
    .ZN(_103_)
  );
  MUX2_X1 _426_ (
    .A(_103_),
    .B(_bufMask_T[0]),
    .S(_098_),
    .Z(_104_)
  );
  AND2_X1 _427_ (
    .A1(exp_io_rvc),
    .A2(_058_),
    .ZN(_105_)
  );
  INV_X1 _428_ (
    .A(_105_),
    .ZN(_106_)
  );
  AND2_X1 _429_ (
    .A1(_103_),
    .A2(_106_),
    .ZN(_107_)
  );
  INV_X1 _430_ (
    .A(_107_),
    .ZN(_108_)
  );
  AND2_X1 _431_ (
    .A1(_055_),
    .A2(_108_),
    .ZN(_109_)
  );
  INV_X1 _432_ (
    .A(_109_),
    .ZN(_110_)
  );
  AND2_X1 _433_ (
    .A1(_104_),
    .A2(_109_),
    .ZN(_111_)
  );
  INV_X1 _434_ (
    .A(_111_),
    .ZN(_112_)
  );
  AND2_X1 _435_ (
    .A1(io_inst_0_ready),
    .A2(_101_),
    .ZN(_113_)
  );
  INV_X1 _436_ (
    .A(_113_),
    .ZN(_114_)
  );
  AND2_X1 _437_ (
    .A1(_112_),
    .A2(_113_),
    .ZN(io_imem_ready)
  );
  AND2_X1 _438_ (
    .A1(io_imem_bits_pc[1]),
    .A2(_107_),
    .ZN(_115_)
  );
  INV_X1 _439_ (
    .A(_115_),
    .ZN(_116_)
  );
  AND2_X1 _440_ (
    .A1(io_imem_valid),
    .A2(_116_),
    .ZN(_117_)
  );
  AND2_X1 _441_ (
    .A1(_104_),
    .A2(_117_),
    .ZN(_118_)
  );
  AND2_X1 _442_ (
    .A1(io_imem_ready),
    .A2(_118_),
    .ZN(_119_)
  );
  INV_X1 _443_ (
    .A(_119_),
    .ZN(_120_)
  );
  MUX2_X1 _444_ (
    .A(buf__replay),
    .B(io_imem_bits_replay),
    .S(_119_),
    .Z(_000_)
  );
  MUX2_X1 _445_ (
    .A(_116_),
    .B(_110_),
    .S(_104_),
    .Z(_121_)
  );
  AND2_X1 _446_ (
    .A1(io_imem_bits_data[16]),
    .A2(_121_),
    .ZN(_122_)
  );
  MUX2_X1 _447_ (
    .A(buf__data[0]),
    .B(_122_),
    .S(_119_),
    .Z(_001_)
  );
  AND2_X1 _448_ (
    .A1(io_imem_bits_data[17]),
    .A2(_121_),
    .ZN(_123_)
  );
  MUX2_X1 _449_ (
    .A(buf__data[1]),
    .B(_123_),
    .S(_119_),
    .Z(_002_)
  );
  AND2_X1 _450_ (
    .A1(io_imem_bits_data[18]),
    .A2(_121_),
    .ZN(_124_)
  );
  MUX2_X1 _451_ (
    .A(buf__data[2]),
    .B(_124_),
    .S(_119_),
    .Z(_003_)
  );
  AND2_X1 _452_ (
    .A1(io_imem_bits_data[19]),
    .A2(_121_),
    .ZN(_125_)
  );
  MUX2_X1 _453_ (
    .A(buf__data[3]),
    .B(_125_),
    .S(_119_),
    .Z(_004_)
  );
  AND2_X1 _454_ (
    .A1(io_imem_bits_data[20]),
    .A2(_121_),
    .ZN(_126_)
  );
  MUX2_X1 _455_ (
    .A(buf__data[4]),
    .B(_126_),
    .S(_119_),
    .Z(_005_)
  );
  AND2_X1 _456_ (
    .A1(io_imem_bits_data[21]),
    .A2(_121_),
    .ZN(_127_)
  );
  MUX2_X1 _457_ (
    .A(buf__data[5]),
    .B(_127_),
    .S(_119_),
    .Z(_006_)
  );
  AND2_X1 _458_ (
    .A1(io_imem_bits_data[22]),
    .A2(_121_),
    .ZN(_128_)
  );
  MUX2_X1 _459_ (
    .A(buf__data[6]),
    .B(_128_),
    .S(_119_),
    .Z(_007_)
  );
  AND2_X1 _460_ (
    .A1(io_imem_bits_data[23]),
    .A2(_121_),
    .ZN(_129_)
  );
  MUX2_X1 _461_ (
    .A(buf__data[7]),
    .B(_129_),
    .S(_119_),
    .Z(_008_)
  );
  AND2_X1 _462_ (
    .A1(io_imem_bits_data[24]),
    .A2(_121_),
    .ZN(_130_)
  );
  MUX2_X1 _463_ (
    .A(buf__data[8]),
    .B(_130_),
    .S(_119_),
    .Z(_009_)
  );
  AND2_X1 _464_ (
    .A1(io_imem_bits_data[25]),
    .A2(_121_),
    .ZN(_131_)
  );
  MUX2_X1 _465_ (
    .A(buf__data[9]),
    .B(_131_),
    .S(_119_),
    .Z(_010_)
  );
  AND2_X1 _466_ (
    .A1(io_imem_bits_data[26]),
    .A2(_121_),
    .ZN(_132_)
  );
  MUX2_X1 _467_ (
    .A(buf__data[10]),
    .B(_132_),
    .S(_119_),
    .Z(_011_)
  );
  AND2_X1 _468_ (
    .A1(io_imem_bits_data[27]),
    .A2(_121_),
    .ZN(_133_)
  );
  MUX2_X1 _469_ (
    .A(buf__data[11]),
    .B(_133_),
    .S(_119_),
    .Z(_012_)
  );
  AND2_X1 _470_ (
    .A1(io_imem_bits_data[28]),
    .A2(_121_),
    .ZN(_134_)
  );
  MUX2_X1 _471_ (
    .A(buf__data[12]),
    .B(_134_),
    .S(_119_),
    .Z(_013_)
  );
  AND2_X1 _472_ (
    .A1(io_imem_bits_data[29]),
    .A2(_121_),
    .ZN(_135_)
  );
  MUX2_X1 _473_ (
    .A(buf__data[13]),
    .B(_135_),
    .S(_119_),
    .Z(_014_)
  );
  AND2_X1 _474_ (
    .A1(io_imem_bits_data[30]),
    .A2(_121_),
    .ZN(_136_)
  );
  MUX2_X1 _475_ (
    .A(buf__data[14]),
    .B(_136_),
    .S(_119_),
    .Z(_015_)
  );
  AND2_X1 _476_ (
    .A1(io_imem_bits_data[31]),
    .A2(_121_),
    .ZN(_137_)
  );
  MUX2_X1 _477_ (
    .A(buf__data[15]),
    .B(_137_),
    .S(_119_),
    .Z(_016_)
  );
  MUX2_X1 _478_ (
    .A(buf__pc[0]),
    .B(io_imem_bits_pc[0]),
    .S(_119_),
    .Z(_017_)
  );
  AND2_X1 _479_ (
    .A1(_052_),
    .A2(_120_),
    .ZN(_138_)
  );
  INV_X1 _480_ (
    .A(_138_),
    .ZN(_018_)
  );
  MUX2_X1 _481_ (
    .A(buf__pc[2]),
    .B(io_imem_bits_pc[2]),
    .S(_119_),
    .Z(_019_)
  );
  MUX2_X1 _482_ (
    .A(buf__pc[3]),
    .B(io_imem_bits_pc[3]),
    .S(_119_),
    .Z(_020_)
  );
  MUX2_X1 _483_ (
    .A(buf__pc[4]),
    .B(io_imem_bits_pc[4]),
    .S(_119_),
    .Z(_021_)
  );
  MUX2_X1 _484_ (
    .A(buf__pc[5]),
    .B(io_imem_bits_pc[5]),
    .S(_119_),
    .Z(_022_)
  );
  MUX2_X1 _485_ (
    .A(buf__pc[6]),
    .B(io_imem_bits_pc[6]),
    .S(_119_),
    .Z(_023_)
  );
  MUX2_X1 _486_ (
    .A(buf__pc[7]),
    .B(io_imem_bits_pc[7]),
    .S(_119_),
    .Z(_024_)
  );
  MUX2_X1 _487_ (
    .A(buf__pc[8]),
    .B(io_imem_bits_pc[8]),
    .S(_119_),
    .Z(_025_)
  );
  MUX2_X1 _488_ (
    .A(buf__pc[9]),
    .B(io_imem_bits_pc[9]),
    .S(_119_),
    .Z(_026_)
  );
  MUX2_X1 _489_ (
    .A(buf__pc[10]),
    .B(io_imem_bits_pc[10]),
    .S(_119_),
    .Z(_027_)
  );
  MUX2_X1 _490_ (
    .A(buf__pc[11]),
    .B(io_imem_bits_pc[11]),
    .S(_119_),
    .Z(_028_)
  );
  MUX2_X1 _491_ (
    .A(buf__pc[12]),
    .B(io_imem_bits_pc[12]),
    .S(_119_),
    .Z(_029_)
  );
  MUX2_X1 _492_ (
    .A(buf__pc[13]),
    .B(io_imem_bits_pc[13]),
    .S(_119_),
    .Z(_030_)
  );
  MUX2_X1 _493_ (
    .A(buf__pc[14]),
    .B(io_imem_bits_pc[14]),
    .S(_119_),
    .Z(_031_)
  );
  MUX2_X1 _494_ (
    .A(buf__pc[15]),
    .B(io_imem_bits_pc[15]),
    .S(_119_),
    .Z(_032_)
  );
  MUX2_X1 _495_ (
    .A(buf__pc[16]),
    .B(io_imem_bits_pc[16]),
    .S(_119_),
    .Z(_033_)
  );
  MUX2_X1 _496_ (
    .A(buf__pc[17]),
    .B(io_imem_bits_pc[17]),
    .S(_119_),
    .Z(_034_)
  );
  MUX2_X1 _497_ (
    .A(buf__pc[18]),
    .B(io_imem_bits_pc[18]),
    .S(_119_),
    .Z(_035_)
  );
  MUX2_X1 _498_ (
    .A(buf__pc[19]),
    .B(io_imem_bits_pc[19]),
    .S(_119_),
    .Z(_036_)
  );
  MUX2_X1 _499_ (
    .A(buf__pc[20]),
    .B(io_imem_bits_pc[20]),
    .S(_119_),
    .Z(_037_)
  );
  MUX2_X1 _500_ (
    .A(buf__pc[21]),
    .B(io_imem_bits_pc[21]),
    .S(_119_),
    .Z(_038_)
  );
  MUX2_X1 _501_ (
    .A(buf__pc[22]),
    .B(io_imem_bits_pc[22]),
    .S(_119_),
    .Z(_039_)
  );
  MUX2_X1 _502_ (
    .A(buf__pc[23]),
    .B(io_imem_bits_pc[23]),
    .S(_119_),
    .Z(_040_)
  );
  MUX2_X1 _503_ (
    .A(buf__pc[24]),
    .B(io_imem_bits_pc[24]),
    .S(_119_),
    .Z(_041_)
  );
  MUX2_X1 _504_ (
    .A(buf__pc[25]),
    .B(io_imem_bits_pc[25]),
    .S(_119_),
    .Z(_042_)
  );
  MUX2_X1 _505_ (
    .A(buf__pc[26]),
    .B(io_imem_bits_pc[26]),
    .S(_119_),
    .Z(_043_)
  );
  MUX2_X1 _506_ (
    .A(buf__pc[27]),
    .B(io_imem_bits_pc[27]),
    .S(_119_),
    .Z(_044_)
  );
  MUX2_X1 _507_ (
    .A(buf__pc[28]),
    .B(io_imem_bits_pc[28]),
    .S(_119_),
    .Z(_045_)
  );
  MUX2_X1 _508_ (
    .A(buf__pc[29]),
    .B(io_imem_bits_pc[29]),
    .S(_119_),
    .Z(_046_)
  );
  MUX2_X1 _509_ (
    .A(buf__pc[30]),
    .B(io_imem_bits_pc[30]),
    .S(_119_),
    .Z(_047_)
  );
  MUX2_X1 _510_ (
    .A(buf__pc[31]),
    .B(io_imem_bits_pc[31]),
    .S(_119_),
    .Z(_048_)
  );
  AND2_X1 _511_ (
    .A1(io_inst_0_ready),
    .A2(exp_io_rvc),
    .ZN(_139_)
  );
  INV_X1 _512_ (
    .A(_139_),
    .ZN(_140_)
  );
  AND2_X1 _513_ (
    .A1(_051_),
    .A2(_140_),
    .ZN(_141_)
  );
  INV_X1 _514_ (
    .A(_141_),
    .ZN(_142_)
  );
  AND2_X1 _515_ (
    .A1(nBufValid),
    .A2(_139_),
    .ZN(_143_)
  );
  INV_X1 _516_ (
    .A(_143_),
    .ZN(_144_)
  );
  AND2_X1 _517_ (
    .A1(_142_),
    .A2(_144_),
    .ZN(_145_)
  );
  AND2_X1 _518_ (
    .A1(_114_),
    .A2(_145_),
    .ZN(_146_)
  );
  INV_X1 _519_ (
    .A(_146_),
    .ZN(_147_)
  );
  AND2_X1 _520_ (
    .A1(_120_),
    .A2(_147_),
    .ZN(_148_)
  );
  INV_X1 _521_ (
    .A(_148_),
    .ZN(_149_)
  );
  AND2_X1 _522_ (
    .A1(_053_),
    .A2(_054_),
    .ZN(_150_)
  );
  AND2_X1 _523_ (
    .A1(_149_),
    .A2(_150_),
    .ZN(_049_)
  );
  MUX2_X1 _524_ (
    .A(buf__xcpt_ae_inst),
    .B(io_imem_bits_xcpt_ae_inst),
    .S(_119_),
    .Z(_050_)
  );
  AND2_X1 _525_ (
    .A1(io_imem_bits_xcpt_ae_inst),
    .A2(_057_),
    .ZN(io_inst_0_bits_xcpt1_ae_inst)
  );
  MUX2_X1 _526_ (
    .A(io_imem_bits_pc[0]),
    .B(buf__pc[0]),
    .S(nBufValid),
    .Z(io_pc[0])
  );
  MUX2_X1 _527_ (
    .A(io_imem_bits_pc[1]),
    .B(buf__pc[1]),
    .S(nBufValid),
    .Z(io_pc[1])
  );
  MUX2_X1 _528_ (
    .A(io_imem_bits_pc[2]),
    .B(buf__pc[2]),
    .S(nBufValid),
    .Z(io_pc[2])
  );
  MUX2_X1 _529_ (
    .A(io_imem_bits_pc[3]),
    .B(buf__pc[3]),
    .S(nBufValid),
    .Z(io_pc[3])
  );
  MUX2_X1 _530_ (
    .A(io_imem_bits_pc[4]),
    .B(buf__pc[4]),
    .S(nBufValid),
    .Z(io_pc[4])
  );
  MUX2_X1 _531_ (
    .A(io_imem_bits_pc[5]),
    .B(buf__pc[5]),
    .S(nBufValid),
    .Z(io_pc[5])
  );
  MUX2_X1 _532_ (
    .A(io_imem_bits_pc[6]),
    .B(buf__pc[6]),
    .S(nBufValid),
    .Z(io_pc[6])
  );
  MUX2_X1 _533_ (
    .A(io_imem_bits_pc[7]),
    .B(buf__pc[7]),
    .S(nBufValid),
    .Z(io_pc[7])
  );
  MUX2_X1 _534_ (
    .A(io_imem_bits_pc[8]),
    .B(buf__pc[8]),
    .S(nBufValid),
    .Z(io_pc[8])
  );
  MUX2_X1 _535_ (
    .A(io_imem_bits_pc[9]),
    .B(buf__pc[9]),
    .S(nBufValid),
    .Z(io_pc[9])
  );
  MUX2_X1 _536_ (
    .A(io_imem_bits_pc[10]),
    .B(buf__pc[10]),
    .S(nBufValid),
    .Z(io_pc[10])
  );
  MUX2_X1 _537_ (
    .A(io_imem_bits_pc[11]),
    .B(buf__pc[11]),
    .S(nBufValid),
    .Z(io_pc[11])
  );
  MUX2_X1 _538_ (
    .A(io_imem_bits_pc[12]),
    .B(buf__pc[12]),
    .S(nBufValid),
    .Z(io_pc[12])
  );
  MUX2_X1 _539_ (
    .A(io_imem_bits_pc[13]),
    .B(buf__pc[13]),
    .S(nBufValid),
    .Z(io_pc[13])
  );
  MUX2_X1 _540_ (
    .A(io_imem_bits_pc[14]),
    .B(buf__pc[14]),
    .S(nBufValid),
    .Z(io_pc[14])
  );
  MUX2_X1 _541_ (
    .A(io_imem_bits_pc[15]),
    .B(buf__pc[15]),
    .S(nBufValid),
    .Z(io_pc[15])
  );
  MUX2_X1 _542_ (
    .A(io_imem_bits_pc[16]),
    .B(buf__pc[16]),
    .S(nBufValid),
    .Z(io_pc[16])
  );
  MUX2_X1 _543_ (
    .A(io_imem_bits_pc[17]),
    .B(buf__pc[17]),
    .S(nBufValid),
    .Z(io_pc[17])
  );
  MUX2_X1 _544_ (
    .A(io_imem_bits_pc[18]),
    .B(buf__pc[18]),
    .S(nBufValid),
    .Z(io_pc[18])
  );
  MUX2_X1 _545_ (
    .A(io_imem_bits_pc[19]),
    .B(buf__pc[19]),
    .S(nBufValid),
    .Z(io_pc[19])
  );
  MUX2_X1 _546_ (
    .A(io_imem_bits_pc[20]),
    .B(buf__pc[20]),
    .S(nBufValid),
    .Z(io_pc[20])
  );
  MUX2_X1 _547_ (
    .A(io_imem_bits_pc[21]),
    .B(buf__pc[21]),
    .S(nBufValid),
    .Z(io_pc[21])
  );
  MUX2_X1 _548_ (
    .A(io_imem_bits_pc[22]),
    .B(buf__pc[22]),
    .S(nBufValid),
    .Z(io_pc[22])
  );
  MUX2_X1 _549_ (
    .A(io_imem_bits_pc[23]),
    .B(buf__pc[23]),
    .S(nBufValid),
    .Z(io_pc[23])
  );
  MUX2_X1 _550_ (
    .A(io_imem_bits_pc[24]),
    .B(buf__pc[24]),
    .S(nBufValid),
    .Z(io_pc[24])
  );
  MUX2_X1 _551_ (
    .A(io_imem_bits_pc[25]),
    .B(buf__pc[25]),
    .S(nBufValid),
    .Z(io_pc[25])
  );
  MUX2_X1 _552_ (
    .A(io_imem_bits_pc[26]),
    .B(buf__pc[26]),
    .S(nBufValid),
    .Z(io_pc[26])
  );
  MUX2_X1 _553_ (
    .A(io_imem_bits_pc[27]),
    .B(buf__pc[27]),
    .S(nBufValid),
    .Z(io_pc[27])
  );
  MUX2_X1 _554_ (
    .A(io_imem_bits_pc[28]),
    .B(buf__pc[28]),
    .S(nBufValid),
    .Z(io_pc[28])
  );
  MUX2_X1 _555_ (
    .A(io_imem_bits_pc[29]),
    .B(buf__pc[29]),
    .S(nBufValid),
    .Z(io_pc[29])
  );
  MUX2_X1 _556_ (
    .A(io_imem_bits_pc[30]),
    .B(buf__pc[30]),
    .S(nBufValid),
    .Z(io_pc[30])
  );
  MUX2_X1 _557_ (
    .A(io_imem_bits_pc[31]),
    .B(buf__pc[31]),
    .S(nBufValid),
    .Z(io_pc[31])
  );
  MUX2_X1 _558_ (
    .A(io_imem_bits_xcpt_ae_inst),
    .B(buf__xcpt_ae_inst),
    .S(nBufValid),
    .Z(io_inst_0_bits_xcpt0_ae_inst)
  );
  AND2_X1 _559_ (
    .A1(_051_),
    .A2(_056_),
    .ZN(_151_)
  );
  INV_X1 _560_ (
    .A(_151_),
    .ZN(_152_)
  );
  AND2_X1 _561_ (
    .A1(_099_),
    .A2(_152_),
    .ZN(io_inst_0_valid)
  );
  AND2_X1 _562_ (
    .A1(_bufMask_T[0]),
    .A2(_152_),
    .ZN(_153_)
  );
  INV_X1 _563_ (
    .A(_153_),
    .ZN(_154_)
  );
  AND2_X1 _564_ (
    .A1(_057_),
    .A2(_093_),
    .ZN(_155_)
  );
  INV_X1 _565_ (
    .A(_155_),
    .ZN(_156_)
  );
  AND2_X1 _566_ (
    .A1(_154_),
    .A2(_156_),
    .ZN(_157_)
  );
  INV_X1 _567_ (
    .A(_157_),
    .ZN(_158_)
  );
  AND2_X1 _568_ (
    .A1(io_imem_bits_replay),
    .A2(_158_),
    .ZN(_159_)
  );
  INV_X1 _569_ (
    .A(_159_),
    .ZN(_160_)
  );
  AND2_X1 _570_ (
    .A1(_096_),
    .A2(_160_),
    .ZN(_161_)
  );
  INV_X1 _571_ (
    .A(_161_),
    .ZN(io_inst_0_bits_replay)
  );
  AND2_X1 _572_ (
    .A1(nBufValid),
    .A2(buf__data[0]),
    .ZN(_162_)
  );
  INV_X1 _573_ (
    .A(_162_),
    .ZN(_163_)
  );
  AND2_X1 _574_ (
    .A1(_059_),
    .A2(_092_),
    .ZN(_164_)
  );
  INV_X1 _575_ (
    .A(_164_),
    .ZN(_165_)
  );
  AND2_X1 _576_ (
    .A1(_060_),
    .A2(_091_),
    .ZN(_166_)
  );
  INV_X1 _577_ (
    .A(_166_),
    .ZN(_167_)
  );
  AND2_X1 _578_ (
    .A1(_bufMask_T[0]),
    .A2(_167_),
    .ZN(_168_)
  );
  AND2_X1 _579_ (
    .A1(_165_),
    .A2(_168_),
    .ZN(_169_)
  );
  INV_X1 _580_ (
    .A(_169_),
    .ZN(_170_)
  );
  AND2_X1 _581_ (
    .A1(_163_),
    .A2(_170_),
    .ZN(_171_)
  );
  INV_X1 _582_ (
    .A(_171_),
    .ZN(exp_io_in[0])
  );
  AND2_X1 _583_ (
    .A1(nBufValid),
    .A2(buf__data[1]),
    .ZN(_172_)
  );
  INV_X1 _584_ (
    .A(_172_),
    .ZN(_173_)
  );
  AND2_X1 _585_ (
    .A1(_061_),
    .A2(_092_),
    .ZN(_174_)
  );
  INV_X1 _586_ (
    .A(_174_),
    .ZN(_175_)
  );
  AND2_X1 _587_ (
    .A1(_062_),
    .A2(_091_),
    .ZN(_176_)
  );
  INV_X1 _588_ (
    .A(_176_),
    .ZN(_177_)
  );
  AND2_X1 _589_ (
    .A1(_bufMask_T[0]),
    .A2(_177_),
    .ZN(_178_)
  );
  AND2_X1 _590_ (
    .A1(_175_),
    .A2(_178_),
    .ZN(_179_)
  );
  INV_X1 _591_ (
    .A(_179_),
    .ZN(_180_)
  );
  AND2_X1 _592_ (
    .A1(_173_),
    .A2(_180_),
    .ZN(_181_)
  );
  INV_X1 _593_ (
    .A(_181_),
    .ZN(exp_io_in[1])
  );
  AND2_X1 _594_ (
    .A1(nBufValid),
    .A2(buf__data[2]),
    .ZN(_182_)
  );
  INV_X1 _595_ (
    .A(_182_),
    .ZN(_183_)
  );
  AND2_X1 _596_ (
    .A1(_063_),
    .A2(_092_),
    .ZN(_184_)
  );
  INV_X1 _597_ (
    .A(_184_),
    .ZN(_185_)
  );
  AND2_X1 _598_ (
    .A1(_064_),
    .A2(_091_),
    .ZN(_186_)
  );
  INV_X1 _599_ (
    .A(_186_),
    .ZN(_187_)
  );
  AND2_X1 _600_ (
    .A1(_bufMask_T[0]),
    .A2(_187_),
    .ZN(_188_)
  );
  AND2_X1 _601_ (
    .A1(_185_),
    .A2(_188_),
    .ZN(_189_)
  );
  INV_X1 _602_ (
    .A(_189_),
    .ZN(_190_)
  );
  AND2_X1 _603_ (
    .A1(_183_),
    .A2(_190_),
    .ZN(_191_)
  );
  INV_X1 _604_ (
    .A(_191_),
    .ZN(exp_io_in[2])
  );
  AND2_X1 _605_ (
    .A1(nBufValid),
    .A2(buf__data[3]),
    .ZN(_192_)
  );
  INV_X1 _606_ (
    .A(_192_),
    .ZN(_193_)
  );
  AND2_X1 _607_ (
    .A1(_066_),
    .A2(_091_),
    .ZN(_194_)
  );
  INV_X1 _608_ (
    .A(_194_),
    .ZN(_195_)
  );
  AND2_X1 _609_ (
    .A1(_065_),
    .A2(_092_),
    .ZN(_196_)
  );
  INV_X1 _610_ (
    .A(_196_),
    .ZN(_197_)
  );
  AND2_X1 _611_ (
    .A1(_bufMask_T[0]),
    .A2(_195_),
    .ZN(_198_)
  );
  AND2_X1 _612_ (
    .A1(_197_),
    .A2(_198_),
    .ZN(_199_)
  );
  INV_X1 _613_ (
    .A(_199_),
    .ZN(_200_)
  );
  AND2_X1 _614_ (
    .A1(_193_),
    .A2(_200_),
    .ZN(_201_)
  );
  INV_X1 _615_ (
    .A(_201_),
    .ZN(exp_io_in[3])
  );
  AND2_X1 _616_ (
    .A1(nBufValid),
    .A2(buf__data[4]),
    .ZN(_202_)
  );
  INV_X1 _617_ (
    .A(_202_),
    .ZN(_203_)
  );
  AND2_X1 _618_ (
    .A1(_067_),
    .A2(_092_),
    .ZN(_204_)
  );
  INV_X1 _619_ (
    .A(_204_),
    .ZN(_205_)
  );
  AND2_X1 _620_ (
    .A1(_068_),
    .A2(_091_),
    .ZN(_206_)
  );
  INV_X1 _621_ (
    .A(_206_),
    .ZN(_207_)
  );
  AND2_X1 _622_ (
    .A1(_bufMask_T[0]),
    .A2(_207_),
    .ZN(_208_)
  );
  AND2_X1 _623_ (
    .A1(_205_),
    .A2(_208_),
    .ZN(_209_)
  );
  INV_X1 _624_ (
    .A(_209_),
    .ZN(_210_)
  );
  AND2_X1 _625_ (
    .A1(_203_),
    .A2(_210_),
    .ZN(_211_)
  );
  INV_X1 _626_ (
    .A(_211_),
    .ZN(exp_io_in[4])
  );
  AND2_X1 _627_ (
    .A1(nBufValid),
    .A2(buf__data[5]),
    .ZN(_212_)
  );
  INV_X1 _628_ (
    .A(_212_),
    .ZN(_213_)
  );
  AND2_X1 _629_ (
    .A1(_070_),
    .A2(_091_),
    .ZN(_214_)
  );
  INV_X1 _630_ (
    .A(_214_),
    .ZN(_215_)
  );
  AND2_X1 _631_ (
    .A1(_069_),
    .A2(_092_),
    .ZN(_216_)
  );
  INV_X1 _632_ (
    .A(_216_),
    .ZN(_217_)
  );
  AND2_X1 _633_ (
    .A1(_bufMask_T[0]),
    .A2(_215_),
    .ZN(_218_)
  );
  AND2_X1 _634_ (
    .A1(_217_),
    .A2(_218_),
    .ZN(_219_)
  );
  INV_X1 _635_ (
    .A(_219_),
    .ZN(_220_)
  );
  AND2_X1 _636_ (
    .A1(_213_),
    .A2(_220_),
    .ZN(_221_)
  );
  INV_X1 _637_ (
    .A(_221_),
    .ZN(exp_io_in[5])
  );
  AND2_X1 _638_ (
    .A1(nBufValid),
    .A2(buf__data[6]),
    .ZN(_222_)
  );
  INV_X1 _639_ (
    .A(_222_),
    .ZN(_223_)
  );
  AND2_X1 _640_ (
    .A1(_071_),
    .A2(_092_),
    .ZN(_224_)
  );
  INV_X1 _641_ (
    .A(_224_),
    .ZN(_225_)
  );
  AND2_X1 _642_ (
    .A1(_072_),
    .A2(_091_),
    .ZN(_226_)
  );
  INV_X1 _643_ (
    .A(_226_),
    .ZN(_227_)
  );
  AND2_X1 _644_ (
    .A1(_bufMask_T[0]),
    .A2(_227_),
    .ZN(_228_)
  );
  AND2_X1 _645_ (
    .A1(_225_),
    .A2(_228_),
    .ZN(_229_)
  );
  INV_X1 _646_ (
    .A(_229_),
    .ZN(_230_)
  );
  AND2_X1 _647_ (
    .A1(_223_),
    .A2(_230_),
    .ZN(_231_)
  );
  INV_X1 _648_ (
    .A(_231_),
    .ZN(exp_io_in[6])
  );
  AND2_X1 _649_ (
    .A1(nBufValid),
    .A2(buf__data[7]),
    .ZN(_232_)
  );
  INV_X1 _650_ (
    .A(_232_),
    .ZN(_233_)
  );
  AND2_X1 _651_ (
    .A1(_073_),
    .A2(_092_),
    .ZN(_234_)
  );
  INV_X1 _652_ (
    .A(_234_),
    .ZN(_235_)
  );
  AND2_X1 _653_ (
    .A1(_074_),
    .A2(_091_),
    .ZN(_236_)
  );
  INV_X1 _654_ (
    .A(_236_),
    .ZN(_237_)
  );
  AND2_X1 _655_ (
    .A1(_bufMask_T[0]),
    .A2(_237_),
    .ZN(_238_)
  );
  AND2_X1 _656_ (
    .A1(_235_),
    .A2(_238_),
    .ZN(_239_)
  );
  INV_X1 _657_ (
    .A(_239_),
    .ZN(_240_)
  );
  AND2_X1 _658_ (
    .A1(_233_),
    .A2(_240_),
    .ZN(_241_)
  );
  INV_X1 _659_ (
    .A(_241_),
    .ZN(exp_io_in[7])
  );
  AND2_X1 _660_ (
    .A1(nBufValid),
    .A2(buf__data[8]),
    .ZN(_242_)
  );
  INV_X1 _661_ (
    .A(_242_),
    .ZN(_243_)
  );
  AND2_X1 _662_ (
    .A1(_075_),
    .A2(_092_),
    .ZN(_244_)
  );
  INV_X1 _663_ (
    .A(_244_),
    .ZN(_245_)
  );
  AND2_X1 _664_ (
    .A1(_076_),
    .A2(_091_),
    .ZN(_246_)
  );
  INV_X1 _665_ (
    .A(_246_),
    .ZN(_247_)
  );
  AND2_X1 _666_ (
    .A1(_bufMask_T[0]),
    .A2(_247_),
    .ZN(_248_)
  );
  AND2_X1 _667_ (
    .A1(_245_),
    .A2(_248_),
    .ZN(_249_)
  );
  INV_X1 _668_ (
    .A(_249_),
    .ZN(_250_)
  );
  AND2_X1 _669_ (
    .A1(_243_),
    .A2(_250_),
    .ZN(_251_)
  );
  INV_X1 _670_ (
    .A(_251_),
    .ZN(exp_io_in[8])
  );
  AND2_X1 _671_ (
    .A1(nBufValid),
    .A2(buf__data[9]),
    .ZN(_252_)
  );
  INV_X1 _672_ (
    .A(_252_),
    .ZN(_253_)
  );
  AND2_X1 _673_ (
    .A1(_077_),
    .A2(_092_),
    .ZN(_254_)
  );
  INV_X1 _674_ (
    .A(_254_),
    .ZN(_255_)
  );
  AND2_X1 _675_ (
    .A1(_078_),
    .A2(_091_),
    .ZN(_256_)
  );
  INV_X1 _676_ (
    .A(_256_),
    .ZN(_257_)
  );
  AND2_X1 _677_ (
    .A1(_bufMask_T[0]),
    .A2(_257_),
    .ZN(_258_)
  );
  AND2_X1 _678_ (
    .A1(_255_),
    .A2(_258_),
    .ZN(_259_)
  );
  INV_X1 _679_ (
    .A(_259_),
    .ZN(_260_)
  );
  AND2_X1 _680_ (
    .A1(_253_),
    .A2(_260_),
    .ZN(_261_)
  );
  INV_X1 _681_ (
    .A(_261_),
    .ZN(exp_io_in[9])
  );
  AND2_X1 _682_ (
    .A1(nBufValid),
    .A2(buf__data[10]),
    .ZN(_262_)
  );
  INV_X1 _683_ (
    .A(_262_),
    .ZN(_263_)
  );
  AND2_X1 _684_ (
    .A1(_079_),
    .A2(_092_),
    .ZN(_264_)
  );
  INV_X1 _685_ (
    .A(_264_),
    .ZN(_265_)
  );
  AND2_X1 _686_ (
    .A1(_080_),
    .A2(_091_),
    .ZN(_266_)
  );
  INV_X1 _687_ (
    .A(_266_),
    .ZN(_267_)
  );
  AND2_X1 _688_ (
    .A1(_bufMask_T[0]),
    .A2(_267_),
    .ZN(_268_)
  );
  AND2_X1 _689_ (
    .A1(_265_),
    .A2(_268_),
    .ZN(_269_)
  );
  INV_X1 _690_ (
    .A(_269_),
    .ZN(_270_)
  );
  AND2_X1 _691_ (
    .A1(_263_),
    .A2(_270_),
    .ZN(_271_)
  );
  INV_X1 _692_ (
    .A(_271_),
    .ZN(exp_io_in[10])
  );
  AND2_X1 _693_ (
    .A1(nBufValid),
    .A2(buf__data[11]),
    .ZN(_272_)
  );
  INV_X1 _694_ (
    .A(_272_),
    .ZN(_273_)
  );
  AND2_X1 _695_ (
    .A1(_081_),
    .A2(_092_),
    .ZN(_274_)
  );
  INV_X1 _696_ (
    .A(_274_),
    .ZN(_275_)
  );
  AND2_X1 _697_ (
    .A1(_082_),
    .A2(_091_),
    .ZN(_276_)
  );
  INV_X1 _698_ (
    .A(_276_),
    .ZN(_277_)
  );
  AND2_X1 _699_ (
    .A1(_bufMask_T[0]),
    .A2(_277_),
    .ZN(_278_)
  );
  AND2_X1 _700_ (
    .A1(_275_),
    .A2(_278_),
    .ZN(_279_)
  );
  INV_X1 _701_ (
    .A(_279_),
    .ZN(_280_)
  );
  AND2_X1 _702_ (
    .A1(_273_),
    .A2(_280_),
    .ZN(_281_)
  );
  INV_X1 _703_ (
    .A(_281_),
    .ZN(exp_io_in[11])
  );
  AND2_X1 _704_ (
    .A1(nBufValid),
    .A2(buf__data[12]),
    .ZN(_282_)
  );
  INV_X1 _705_ (
    .A(_282_),
    .ZN(_283_)
  );
  AND2_X1 _706_ (
    .A1(_083_),
    .A2(_092_),
    .ZN(_284_)
  );
  INV_X1 _707_ (
    .A(_284_),
    .ZN(_285_)
  );
  AND2_X1 _708_ (
    .A1(_084_),
    .A2(_091_),
    .ZN(_286_)
  );
  INV_X1 _709_ (
    .A(_286_),
    .ZN(_287_)
  );
  AND2_X1 _710_ (
    .A1(_bufMask_T[0]),
    .A2(_287_),
    .ZN(_288_)
  );
  AND2_X1 _711_ (
    .A1(_285_),
    .A2(_288_),
    .ZN(_289_)
  );
  INV_X1 _712_ (
    .A(_289_),
    .ZN(_290_)
  );
  AND2_X1 _713_ (
    .A1(_283_),
    .A2(_290_),
    .ZN(_291_)
  );
  INV_X1 _714_ (
    .A(_291_),
    .ZN(exp_io_in[12])
  );
  AND2_X1 _715_ (
    .A1(nBufValid),
    .A2(buf__data[13]),
    .ZN(_292_)
  );
  INV_X1 _716_ (
    .A(_292_),
    .ZN(_293_)
  );
  AND2_X1 _717_ (
    .A1(_086_),
    .A2(_091_),
    .ZN(_294_)
  );
  INV_X1 _718_ (
    .A(_294_),
    .ZN(_295_)
  );
  AND2_X1 _719_ (
    .A1(_085_),
    .A2(_092_),
    .ZN(_296_)
  );
  INV_X1 _720_ (
    .A(_296_),
    .ZN(_297_)
  );
  AND2_X1 _721_ (
    .A1(_bufMask_T[0]),
    .A2(_295_),
    .ZN(_298_)
  );
  AND2_X1 _722_ (
    .A1(_297_),
    .A2(_298_),
    .ZN(_299_)
  );
  INV_X1 _723_ (
    .A(_299_),
    .ZN(_300_)
  );
  AND2_X1 _724_ (
    .A1(_293_),
    .A2(_300_),
    .ZN(_301_)
  );
  INV_X1 _725_ (
    .A(_301_),
    .ZN(exp_io_in[13])
  );
  AND2_X1 _726_ (
    .A1(nBufValid),
    .A2(buf__data[14]),
    .ZN(_302_)
  );
  INV_X1 _727_ (
    .A(_302_),
    .ZN(_303_)
  );
  AND2_X1 _728_ (
    .A1(_087_),
    .A2(_092_),
    .ZN(_304_)
  );
  INV_X1 _729_ (
    .A(_304_),
    .ZN(_305_)
  );
  AND2_X1 _730_ (
    .A1(_088_),
    .A2(_091_),
    .ZN(_306_)
  );
  INV_X1 _731_ (
    .A(_306_),
    .ZN(_307_)
  );
  AND2_X1 _732_ (
    .A1(_bufMask_T[0]),
    .A2(_307_),
    .ZN(_308_)
  );
  AND2_X1 _733_ (
    .A1(_305_),
    .A2(_308_),
    .ZN(_309_)
  );
  INV_X1 _734_ (
    .A(_309_),
    .ZN(_310_)
  );
  AND2_X1 _735_ (
    .A1(_303_),
    .A2(_310_),
    .ZN(_311_)
  );
  INV_X1 _736_ (
    .A(_311_),
    .ZN(exp_io_in[14])
  );
  AND2_X1 _737_ (
    .A1(nBufValid),
    .A2(buf__data[15]),
    .ZN(_312_)
  );
  INV_X1 _738_ (
    .A(_312_),
    .ZN(_313_)
  );
  AND2_X1 _739_ (
    .A1(_089_),
    .A2(_092_),
    .ZN(_314_)
  );
  INV_X1 _740_ (
    .A(_314_),
    .ZN(_315_)
  );
  AND2_X1 _741_ (
    .A1(_090_),
    .A2(_091_),
    .ZN(_316_)
  );
  INV_X1 _742_ (
    .A(_316_),
    .ZN(_317_)
  );
  AND2_X1 _743_ (
    .A1(_bufMask_T[0]),
    .A2(_317_),
    .ZN(_318_)
  );
  AND2_X1 _744_ (
    .A1(_315_),
    .A2(_318_),
    .ZN(_319_)
  );
  INV_X1 _745_ (
    .A(_319_),
    .ZN(_320_)
  );
  AND2_X1 _746_ (
    .A1(_313_),
    .A2(_320_),
    .ZN(_321_)
  );
  INV_X1 _747_ (
    .A(_321_),
    .ZN(exp_io_in[15])
  );
  AND2_X1 _748_ (
    .A1(nBufValid),
    .A2(_055_),
    .ZN(_322_)
  );
  MUX2_X1 _749_ (
    .A(io_imem_bits_data[16]),
    .B(io_imem_bits_data[0]),
    .S(_322_),
    .Z(_icData_T_4[80])
  );
  MUX2_X1 _750_ (
    .A(io_imem_bits_data[17]),
    .B(io_imem_bits_data[1]),
    .S(_322_),
    .Z(_icData_T_4[81])
  );
  MUX2_X1 _751_ (
    .A(io_imem_bits_data[18]),
    .B(io_imem_bits_data[2]),
    .S(_322_),
    .Z(_icData_T_4[82])
  );
  MUX2_X1 _752_ (
    .A(io_imem_bits_data[19]),
    .B(io_imem_bits_data[3]),
    .S(_322_),
    .Z(_icData_T_4[83])
  );
  MUX2_X1 _753_ (
    .A(io_imem_bits_data[20]),
    .B(io_imem_bits_data[4]),
    .S(_322_),
    .Z(_icData_T_4[84])
  );
  MUX2_X1 _754_ (
    .A(io_imem_bits_data[21]),
    .B(io_imem_bits_data[5]),
    .S(_322_),
    .Z(_icData_T_4[85])
  );
  MUX2_X1 _755_ (
    .A(io_imem_bits_data[22]),
    .B(io_imem_bits_data[6]),
    .S(_322_),
    .Z(_icData_T_4[86])
  );
  MUX2_X1 _756_ (
    .A(io_imem_bits_data[23]),
    .B(io_imem_bits_data[7]),
    .S(_322_),
    .Z(_icData_T_4[87])
  );
  MUX2_X1 _757_ (
    .A(io_imem_bits_data[24]),
    .B(io_imem_bits_data[8]),
    .S(_322_),
    .Z(_icData_T_4[88])
  );
  MUX2_X1 _758_ (
    .A(io_imem_bits_data[25]),
    .B(io_imem_bits_data[9]),
    .S(_322_),
    .Z(_icData_T_4[89])
  );
  MUX2_X1 _759_ (
    .A(io_imem_bits_data[26]),
    .B(io_imem_bits_data[10]),
    .S(_322_),
    .Z(_icData_T_4[90])
  );
  MUX2_X1 _760_ (
    .A(io_imem_bits_data[27]),
    .B(io_imem_bits_data[11]),
    .S(_322_),
    .Z(_icData_T_4[91])
  );
  MUX2_X1 _761_ (
    .A(io_imem_bits_data[28]),
    .B(io_imem_bits_data[12]),
    .S(_322_),
    .Z(_icData_T_4[92])
  );
  MUX2_X1 _762_ (
    .A(io_imem_bits_data[29]),
    .B(io_imem_bits_data[13]),
    .S(_322_),
    .Z(_icData_T_4[93])
  );
  MUX2_X1 _763_ (
    .A(io_imem_bits_data[30]),
    .B(io_imem_bits_data[14]),
    .S(_322_),
    .Z(_icData_T_4[94])
  );
  MUX2_X1 _764_ (
    .A(io_imem_bits_data[31]),
    .B(io_imem_bits_data[15]),
    .S(_322_),
    .Z(_icData_T_4[95])
  );
  DFF_X1 \buf__data[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_001_),
    .Q(buf__data[0]),
    .QN(_371_)
  );
  DFF_X1 \buf__data[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_011_),
    .Q(buf__data[10]),
    .QN(_361_)
  );
  DFF_X1 \buf__data[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_012_),
    .Q(buf__data[11]),
    .QN(_360_)
  );
  DFF_X1 \buf__data[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_013_),
    .Q(buf__data[12]),
    .QN(_359_)
  );
  DFF_X1 \buf__data[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_014_),
    .Q(buf__data[13]),
    .QN(_358_)
  );
  DFF_X1 \buf__data[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_015_),
    .Q(buf__data[14]),
    .QN(_357_)
  );
  DFF_X1 \buf__data[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_016_),
    .Q(buf__data[15]),
    .QN(_356_)
  );
  DFF_X1 \buf__data[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_002_),
    .Q(buf__data[1]),
    .QN(_370_)
  );
  DFF_X1 \buf__data[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_003_),
    .Q(buf__data[2]),
    .QN(_369_)
  );
  DFF_X1 \buf__data[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_004_),
    .Q(buf__data[3]),
    .QN(_368_)
  );
  DFF_X1 \buf__data[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_005_),
    .Q(buf__data[4]),
    .QN(_367_)
  );
  DFF_X1 \buf__data[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_006_),
    .Q(buf__data[5]),
    .QN(_366_)
  );
  DFF_X1 \buf__data[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_007_),
    .Q(buf__data[6]),
    .QN(_365_)
  );
  DFF_X1 \buf__data[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_008_),
    .Q(buf__data[7]),
    .QN(_364_)
  );
  DFF_X1 \buf__data[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_009_),
    .Q(buf__data[8]),
    .QN(_363_)
  );
  DFF_X1 \buf__data[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_010_),
    .Q(buf__data[9]),
    .QN(_362_)
  );
  DFF_X1 \buf__pc[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_017_),
    .Q(buf__pc[0]),
    .QN(_355_)
  );
  DFF_X1 \buf__pc[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_027_),
    .Q(buf__pc[10]),
    .QN(_345_)
  );
  DFF_X1 \buf__pc[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_028_),
    .Q(buf__pc[11]),
    .QN(_344_)
  );
  DFF_X1 \buf__pc[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_029_),
    .Q(buf__pc[12]),
    .QN(_343_)
  );
  DFF_X1 \buf__pc[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_030_),
    .Q(buf__pc[13]),
    .QN(_342_)
  );
  DFF_X1 \buf__pc[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_031_),
    .Q(buf__pc[14]),
    .QN(_341_)
  );
  DFF_X1 \buf__pc[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_032_),
    .Q(buf__pc[15]),
    .QN(_340_)
  );
  DFF_X1 \buf__pc[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_033_),
    .Q(buf__pc[16]),
    .QN(_339_)
  );
  DFF_X1 \buf__pc[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_034_),
    .Q(buf__pc[17]),
    .QN(_338_)
  );
  DFF_X1 \buf__pc[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_035_),
    .Q(buf__pc[18]),
    .QN(_337_)
  );
  DFF_X1 \buf__pc[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_036_),
    .Q(buf__pc[19]),
    .QN(_336_)
  );
  DFF_X1 \buf__pc[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_018_),
    .Q(buf__pc[1]),
    .QN(_354_)
  );
  DFF_X1 \buf__pc[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_037_),
    .Q(buf__pc[20]),
    .QN(_335_)
  );
  DFF_X1 \buf__pc[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_038_),
    .Q(buf__pc[21]),
    .QN(_334_)
  );
  DFF_X1 \buf__pc[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_039_),
    .Q(buf__pc[22]),
    .QN(_333_)
  );
  DFF_X1 \buf__pc[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_040_),
    .Q(buf__pc[23]),
    .QN(_332_)
  );
  DFF_X1 \buf__pc[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_041_),
    .Q(buf__pc[24]),
    .QN(_331_)
  );
  DFF_X1 \buf__pc[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_042_),
    .Q(buf__pc[25]),
    .QN(_330_)
  );
  DFF_X1 \buf__pc[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_043_),
    .Q(buf__pc[26]),
    .QN(_329_)
  );
  DFF_X1 \buf__pc[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_044_),
    .Q(buf__pc[27]),
    .QN(_328_)
  );
  DFF_X1 \buf__pc[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_045_),
    .Q(buf__pc[28]),
    .QN(_327_)
  );
  DFF_X1 \buf__pc[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_046_),
    .Q(buf__pc[29]),
    .QN(_326_)
  );
  DFF_X1 \buf__pc[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_019_),
    .Q(buf__pc[2]),
    .QN(_353_)
  );
  DFF_X1 \buf__pc[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_047_),
    .Q(buf__pc[30]),
    .QN(_325_)
  );
  DFF_X1 \buf__pc[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_048_),
    .Q(buf__pc[31]),
    .QN(_324_)
  );
  DFF_X1 \buf__pc[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_020_),
    .Q(buf__pc[3]),
    .QN(_352_)
  );
  DFF_X1 \buf__pc[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_021_),
    .Q(buf__pc[4]),
    .QN(_351_)
  );
  DFF_X1 \buf__pc[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_022_),
    .Q(buf__pc[5]),
    .QN(_350_)
  );
  DFF_X1 \buf__pc[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_023_),
    .Q(buf__pc[6]),
    .QN(_349_)
  );
  DFF_X1 \buf__pc[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_024_),
    .Q(buf__pc[7]),
    .QN(_348_)
  );
  DFF_X1 \buf__pc[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_025_),
    .Q(buf__pc[8]),
    .QN(_347_)
  );
  DFF_X1 \buf__pc[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_026_),
    .Q(buf__pc[9]),
    .QN(_346_)
  );
  DFF_X1 \buf__replay$_DFFE_PP_  (
    .CK(clock),
    .D(_000_),
    .Q(buf__replay),
    .QN(_372_)
  );
  DFF_X1 \buf__xcpt_ae_inst$_DFFE_PP_  (
    .CK(clock),
    .D(_050_),
    .Q(buf__xcpt_ae_inst),
    .QN(_323_)
  );
  RVCExpander exp (
    .io_in({ _icData_T_4[95:80], exp_io_in[15:0] }),
    .io_out_bits(exp_io_out_bits),
    .io_out_rd(exp_io_out_rd),
    .io_out_rs1(exp_io_out_rs1),
    .io_out_rs2(exp_io_out_rs2),
    .io_rvc(exp_io_rvc)
  );
  DFF_X1 \nBufValid$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_049_),
    .Q(nBufValid),
    .QN(_bufMask_T[0])
  );
  assign _GEN_1 = { 63'h0000000000000000, io_imem_bits_data[31:16], io_imem_bits_data[31:16], io_imem_bits_data[31:16], io_imem_bits_data[31:16], io_imem_bits_data, io_imem_bits_data[15:0], io_imem_bits_data[15:0] };
  assign _GEN_58 = { 1'h0, io_imem_bits_pc[1] };
  assign _GEN_59 = { 1'h0, nBufValid };
  assign { _GEN_67[31:3], _GEN_67[0] } = 30'h00000000;
  assign _bufMask_T[1] = nBufValid;
  assign _buf_data_T[3:0] = 4'h0;
  assign _buf_pc_T_1 = { io_imem_bits_pc[31:2], 2'h0 };
  assign _buf_pc_T_2 = { _GEN_67[2:1], 1'h0 };
  assign _buf_pc_T_4[1:0] = { _buf_data_T[4], io_imem_bits_pc[0] };
  assign _buf_pc_T_5 = { 30'h00000000, _buf_data_T[4], io_imem_bits_pc[0] };
  assign _buf_pc_T_6 = { io_imem_bits_pc[31:2], _buf_data_T[4], io_imem_bits_pc[0] };
  assign _full_insn_T_2[1] = 1'h0;
  assign _icData_T_2 = { io_imem_bits_data, io_imem_bits_data[15:0], io_imem_bits_data[15:0] };
  assign _icData_T_3[3:0] = 4'h0;
  assign { _icData_T_4[190:176], _icData_T_4[127:96] } = { 15'h0000, io_imem_bits_data[31:16], io_imem_bits_data[31:16] };
  assign _icMask_T_1 = { nBufValid, 4'h0 };
  assign _icMask_T_2 = { 15'h0000, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, 16'hffff, _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0] };
  assign _icShiftAmt_T_1 = { 1'h1, nBufValid };
  assign _ic_replay_T = { 1'h1, _bufMask_T[0] };
  assign _ic_replay_T_1[1] = _full_insn_T_2[0];
  assign _inst_T[31:16] = _icData_T_4[95:80];
  assign _inst_T_1 = { 16'h0000, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid };
  assign _inst_T_2[31:16] = 16'h0000;
  assign _io_inst_0_bits_xcpt1_T_4 = { 2'h0, io_imem_bits_xcpt_ae_inst };
  assign _io_inst_0_bits_xcpt1_T_5 = { 2'h0, io_inst_0_bits_xcpt1_ae_inst };
  assign _nReady_T_4[0] = exp_io_rvc;
  assign _replay_T_5[1] = 1'h0;
  assign _valid_T_2[1] = _full_insn_T_2[0];
  assign bufMask = { 1'h0, nBufValid };
  assign buf__data[31:16] = 16'h0000;
  assign buf_data_data = { io_imem_bits_data[31:16], io_imem_bits_data[31:16], io_imem_bits_data };
  assign buf_replay[1] = 1'h0;
  assign exp_io_in[31:16] = _icData_T_4[95:80];
  assign icData = _icData_T_4[95:64];
  assign icData_data = { io_imem_bits_data[31:16], io_imem_bits_data[31:16], io_imem_bits_data[31:16], io_imem_bits_data[31:16], io_imem_bits_data, io_imem_bits_data[15:0], io_imem_bits_data[15:0] };
  assign icMask = { 16'hffff, _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0] };
  assign icShiftAmt = _icData_T_3[5:4];
  assign io_inst_0_bits_inst_bits = exp_io_out_bits;
  assign io_inst_0_bits_inst_rd = exp_io_out_rd;
  assign io_inst_0_bits_inst_rs1 = exp_io_out_rs1;
  assign io_inst_0_bits_inst_rs2 = exp_io_out_rs2;
  assign io_inst_0_bits_raw = { _icData_T_4[95:80], exp_io_in[15:0] };
  assign io_inst_0_bits_rvc = exp_io_rvc;
  assign io_inst_0_bits_xcpt1_gf_inst = 1'h0;
  assign io_inst_0_bits_xcpt1_pf_inst = 1'h0;
  assign nIC[0] = io_imem_bits_pc[1];
  assign nICReady = _GEN_67[2:1];
  assign pcWordBits = io_imem_bits_pc[1];
  assign shamt = _buf_data_T[5:4];
  assign valid = { _full_insn_T_2[0], _valid_T_2[0] };
  assign xcpt_1_ae_inst = io_imem_bits_xcpt_ae_inst;
endmodule
module MulDiv(clock, reset, io_req_ready, io_req_valid, io_req_bits_fn, io_req_bits_in1, io_req_bits_in2, io_req_bits_tag, io_kill, io_resp_ready, io_resp_valid, io_resp_bits_data, io_resp_bits_tag);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire [32:0] _11217_;
  wire [65:0] _GEN_0;
  wire [65:0] _GEN_2;
  wire [41:0] _GEN_35;
  wire [5:0] _count_T_1;
  wire [1:0] _decoded_T_4;
  wire _decoded_T_6;
  wire [1:0] _decoded_T_7;
  wire [1:0] _decoded_orMatrixOutputs_T_4;
  wire [32:0] _divisor_T;
  wire _eOut_T_4;
  wire [8:0] _prod_T_2;
  wire [65:0] _remainder_T_2;
  wire [2:0] _state_T;
  wire [32:0] accum;
  input clock;
  wire clock;
  wire [5:0] count;
  wire decoded_andMatrixInput_0_3;
  wire decoded_andMatrixInput_0_4;
  wire decoded_andMatrixInput_1_2;
  wire [2:0] decoded_plaInput;
  wire [32:0] divisor;
  wire [15:0] hi;
  wire [15:0] hi_1;
  input io_kill;
  wire io_kill;
  input [3:0] io_req_bits_fn;
  wire [3:0] io_req_bits_fn;
  input [31:0] io_req_bits_in1;
  wire [31:0] io_req_bits_in1;
  input [31:0] io_req_bits_in2;
  wire [31:0] io_req_bits_in2;
  input [4:0] io_req_bits_tag;
  wire [4:0] io_req_bits_tag;
  output io_req_ready;
  wire io_req_ready;
  input io_req_valid;
  wire io_req_valid;
  output [31:0] io_resp_bits_data;
  wire [31:0] io_resp_bits_data;
  output [4:0] io_resp_bits_tag;
  wire [4:0] io_resp_bits_tag;
  input io_resp_ready;
  wire io_resp_ready;
  output io_resp_valid;
  wire io_resp_valid;
  wire isHi;
  wire [31:0] lhs_in;
  wire [15:0] loOut;
  wire [31:0] mplier;
  wire mplierSign;
  wire [64:0] mulReg;
  wire neg_out;
  wire [31:0] negated_remainder;
  wire nextMplierSign;
  wire [65:0] nextMulReg;
  wire [64:0] nextMulReg1;
  wire [41:0] nextMulReg_hi;
  wire [65:0] remainder;
  wire [4:0] req_tag;
  wire resHi;
  input reset;
  wire reset;
  wire [31:0] result;
  wire rhs_sign;
  wire [2:0] state;
  wire [64:0] unrolls_0;
  INV_X1 _11218_ (
    .A(remainder[65]),
    .ZN(_04404_)
  );
  INV_X1 _11219_ (
    .A(remainder[64]),
    .ZN(_04415_)
  );
  INV_X1 _11220_ (
    .A(remainder[63]),
    .ZN(_04426_)
  );
  INV_X1 _11221_ (
    .A(remainder[62]),
    .ZN(_04437_)
  );
  INV_X1 _11222_ (
    .A(remainder[61]),
    .ZN(_04448_)
  );
  INV_X1 _11223_ (
    .A(remainder[60]),
    .ZN(_04459_)
  );
  INV_X1 _11224_ (
    .A(remainder[59]),
    .ZN(_04470_)
  );
  INV_X1 _11225_ (
    .A(remainder[58]),
    .ZN(_04481_)
  );
  INV_X1 _11226_ (
    .A(remainder[57]),
    .ZN(_04492_)
  );
  INV_X1 _11227_ (
    .A(remainder[56]),
    .ZN(_04503_)
  );
  INV_X1 _11228_ (
    .A(remainder[55]),
    .ZN(_04514_)
  );
  INV_X1 _11229_ (
    .A(remainder[54]),
    .ZN(_04525_)
  );
  INV_X1 _11230_ (
    .A(remainder[53]),
    .ZN(_04536_)
  );
  INV_X1 _11231_ (
    .A(remainder[52]),
    .ZN(_04546_)
  );
  INV_X1 _11232_ (
    .A(remainder[51]),
    .ZN(_04557_)
  );
  INV_X1 _11233_ (
    .A(remainder[50]),
    .ZN(_04568_)
  );
  INV_X1 _11234_ (
    .A(remainder[49]),
    .ZN(_04579_)
  );
  INV_X1 _11235_ (
    .A(remainder[48]),
    .ZN(_04590_)
  );
  INV_X1 _11236_ (
    .A(remainder[47]),
    .ZN(_04601_)
  );
  INV_X1 _11237_ (
    .A(remainder[46]),
    .ZN(_04612_)
  );
  INV_X1 _11238_ (
    .A(remainder[45]),
    .ZN(_04623_)
  );
  INV_X1 _11239_ (
    .A(remainder[44]),
    .ZN(_04634_)
  );
  INV_X1 _11240_ (
    .A(remainder[43]),
    .ZN(_04645_)
  );
  INV_X1 _11241_ (
    .A(remainder[42]),
    .ZN(_04656_)
  );
  INV_X1 _11242_ (
    .A(remainder[41]),
    .ZN(_04667_)
  );
  INV_X1 _11243_ (
    .A(remainder[40]),
    .ZN(_04678_)
  );
  INV_X1 _11244_ (
    .A(remainder[39]),
    .ZN(_04689_)
  );
  INV_X1 _11245_ (
    .A(remainder[38]),
    .ZN(_04700_)
  );
  INV_X1 _11246_ (
    .A(remainder[37]),
    .ZN(_04711_)
  );
  INV_X1 _11247_ (
    .A(remainder[36]),
    .ZN(_04722_)
  );
  INV_X1 _11248_ (
    .A(remainder[35]),
    .ZN(_04733_)
  );
  INV_X1 _11249_ (
    .A(remainder[34]),
    .ZN(_04744_)
  );
  INV_X1 _11250_ (
    .A(remainder[33]),
    .ZN(_04755_)
  );
  INV_X1 _11251_ (
    .A(remainder[32]),
    .ZN(_04766_)
  );
  INV_X1 _11252_ (
    .A(count[5]),
    .ZN(_04777_)
  );
  INV_X1 _11253_ (
    .A(count[4]),
    .ZN(_04788_)
  );
  INV_X1 _11254_ (
    .A(count[3]),
    .ZN(_04799_)
  );
  INV_X1 _11255_ (
    .A(count[2]),
    .ZN(_04810_)
  );
  INV_X1 _11256_ (
    .A(count[1]),
    .ZN(_04820_)
  );
  INV_X1 _11257_ (
    .A(count[0]),
    .ZN(_04831_)
  );
  INV_X1 _11258_ (
    .A(reset),
    .ZN(_04842_)
  );
  INV_X1 _11259_ (
    .A(divisor[0]),
    .ZN(_04853_)
  );
  INV_X1 _11260_ (
    .A(divisor[2]),
    .ZN(_04864_)
  );
  INV_X1 _11261_ (
    .A(divisor[4]),
    .ZN(_04875_)
  );
  INV_X1 _11262_ (
    .A(divisor[5]),
    .ZN(_04886_)
  );
  INV_X1 _11263_ (
    .A(divisor[7]),
    .ZN(_04897_)
  );
  INV_X1 _11264_ (
    .A(divisor[8]),
    .ZN(_04908_)
  );
  INV_X1 _11265_ (
    .A(divisor[10]),
    .ZN(_04919_)
  );
  INV_X1 _11266_ (
    .A(divisor[11]),
    .ZN(_04930_)
  );
  INV_X1 _11267_ (
    .A(divisor[13]),
    .ZN(_04941_)
  );
  INV_X1 _11268_ (
    .A(divisor[14]),
    .ZN(_04952_)
  );
  INV_X1 _11269_ (
    .A(divisor[16]),
    .ZN(_04963_)
  );
  INV_X1 _11270_ (
    .A(divisor[17]),
    .ZN(_04974_)
  );
  INV_X1 _11271_ (
    .A(divisor[19]),
    .ZN(_04985_)
  );
  INV_X1 _11272_ (
    .A(divisor[20]),
    .ZN(_04996_)
  );
  INV_X1 _11273_ (
    .A(divisor[22]),
    .ZN(_05007_)
  );
  INV_X1 _11274_ (
    .A(divisor[23]),
    .ZN(_05018_)
  );
  INV_X1 _11275_ (
    .A(divisor[25]),
    .ZN(_05029_)
  );
  INV_X1 _11276_ (
    .A(divisor[26]),
    .ZN(_05040_)
  );
  INV_X1 _11277_ (
    .A(divisor[28]),
    .ZN(_05051_)
  );
  INV_X1 _11278_ (
    .A(divisor[29]),
    .ZN(_05062_)
  );
  INV_X1 _11279_ (
    .A(remainder[0]),
    .ZN(_05073_)
  );
  INV_X1 _11280_ (
    .A(remainder[1]),
    .ZN(_05084_)
  );
  INV_X1 _11281_ (
    .A(remainder[2]),
    .ZN(_05095_)
  );
  INV_X1 _11282_ (
    .A(remainder[3]),
    .ZN(_05105_)
  );
  INV_X1 _11283_ (
    .A(remainder[4]),
    .ZN(_05116_)
  );
  INV_X1 _11284_ (
    .A(remainder[5]),
    .ZN(_05127_)
  );
  INV_X1 _11285_ (
    .A(remainder[6]),
    .ZN(_05138_)
  );
  INV_X1 _11286_ (
    .A(remainder[7]),
    .ZN(_05149_)
  );
  INV_X1 _11287_ (
    .A(remainder[8]),
    .ZN(_05160_)
  );
  INV_X1 _11288_ (
    .A(remainder[9]),
    .ZN(_05171_)
  );
  INV_X1 _11289_ (
    .A(remainder[10]),
    .ZN(_05182_)
  );
  INV_X1 _11290_ (
    .A(remainder[11]),
    .ZN(_05193_)
  );
  INV_X1 _11291_ (
    .A(remainder[12]),
    .ZN(_05204_)
  );
  INV_X1 _11292_ (
    .A(remainder[13]),
    .ZN(_05215_)
  );
  INV_X1 _11293_ (
    .A(remainder[14]),
    .ZN(_05226_)
  );
  INV_X1 _11294_ (
    .A(remainder[15]),
    .ZN(_05237_)
  );
  INV_X1 _11295_ (
    .A(remainder[16]),
    .ZN(_05248_)
  );
  INV_X1 _11296_ (
    .A(remainder[17]),
    .ZN(_05259_)
  );
  INV_X1 _11297_ (
    .A(remainder[18]),
    .ZN(_05270_)
  );
  INV_X1 _11298_ (
    .A(remainder[19]),
    .ZN(_05281_)
  );
  INV_X1 _11299_ (
    .A(remainder[20]),
    .ZN(_05292_)
  );
  INV_X1 _11300_ (
    .A(remainder[21]),
    .ZN(_05303_)
  );
  INV_X1 _11301_ (
    .A(remainder[22]),
    .ZN(_05314_)
  );
  INV_X1 _11302_ (
    .A(remainder[23]),
    .ZN(_05325_)
  );
  INV_X1 _11303_ (
    .A(remainder[24]),
    .ZN(_05336_)
  );
  INV_X1 _11304_ (
    .A(remainder[25]),
    .ZN(_05347_)
  );
  INV_X1 _11305_ (
    .A(remainder[26]),
    .ZN(_05358_)
  );
  INV_X1 _11306_ (
    .A(remainder[27]),
    .ZN(_05369_)
  );
  INV_X1 _11307_ (
    .A(remainder[28]),
    .ZN(_05380_)
  );
  INV_X1 _11308_ (
    .A(remainder[29]),
    .ZN(_05391_)
  );
  INV_X1 _11309_ (
    .A(remainder[30]),
    .ZN(_05402_)
  );
  INV_X1 _11310_ (
    .A(state[1]),
    .ZN(_05412_)
  );
  INV_X1 _11311_ (
    .A(state[0]),
    .ZN(_05423_)
  );
  INV_X1 _11312_ (
    .A(state[2]),
    .ZN(_05434_)
  );
  INV_X1 _11313_ (
    .A(io_req_bits_fn[2]),
    .ZN(_05445_)
  );
  INV_X1 _11314_ (
    .A(io_req_bits_fn[1]),
    .ZN(_05456_)
  );
  INV_X1 _11315_ (
    .A(_00002_),
    .ZN(_05467_)
  );
  INV_X1 _11316_ (
    .A(_count_T_1[0]),
    .ZN(_05478_)
  );
  INV_X1 _11317_ (
    .A(_00000_),
    .ZN(_05489_)
  );
  INV_X1 _11318_ (
    .A(_00001_),
    .ZN(_05500_)
  );
  INV_X1 _11319_ (
    .A(_00004_),
    .ZN(_05511_)
  );
  INV_X1 _11320_ (
    .A(_00003_),
    .ZN(_05522_)
  );
  INV_X1 _11321_ (
    .A(io_req_bits_in1[1]),
    .ZN(_05533_)
  );
  INV_X1 _11322_ (
    .A(_state_T[1]),
    .ZN(_05544_)
  );
  INV_X1 _11323_ (
    .A(io_kill),
    .ZN(_05555_)
  );
  INV_X1 _11324_ (
    .A(_11217_[0]),
    .ZN(_05566_)
  );
  INV_X1 _11325_ (
    .A(_11217_[1]),
    .ZN(_05577_)
  );
  INV_X1 _11326_ (
    .A(_11217_[2]),
    .ZN(_05588_)
  );
  INV_X1 _11327_ (
    .A(_11217_[3]),
    .ZN(_05599_)
  );
  INV_X1 _11328_ (
    .A(_11217_[4]),
    .ZN(_05610_)
  );
  INV_X1 _11329_ (
    .A(_11217_[5]),
    .ZN(_05621_)
  );
  INV_X1 _11330_ (
    .A(_11217_[6]),
    .ZN(_05632_)
  );
  INV_X1 _11331_ (
    .A(_11217_[7]),
    .ZN(_05643_)
  );
  INV_X1 _11332_ (
    .A(_11217_[8]),
    .ZN(_05654_)
  );
  INV_X1 _11333_ (
    .A(_11217_[9]),
    .ZN(_05665_)
  );
  INV_X1 _11334_ (
    .A(_11217_[10]),
    .ZN(_05676_)
  );
  INV_X1 _11335_ (
    .A(_11217_[11]),
    .ZN(_05687_)
  );
  INV_X1 _11336_ (
    .A(_11217_[12]),
    .ZN(_05698_)
  );
  INV_X1 _11337_ (
    .A(_11217_[13]),
    .ZN(_05709_)
  );
  INV_X1 _11338_ (
    .A(_11217_[14]),
    .ZN(_05720_)
  );
  INV_X1 _11339_ (
    .A(_11217_[15]),
    .ZN(_05730_)
  );
  INV_X1 _11340_ (
    .A(_11217_[16]),
    .ZN(_05741_)
  );
  INV_X1 _11341_ (
    .A(_11217_[17]),
    .ZN(_05752_)
  );
  INV_X1 _11342_ (
    .A(_11217_[18]),
    .ZN(_05763_)
  );
  INV_X1 _11343_ (
    .A(_11217_[19]),
    .ZN(_05774_)
  );
  INV_X1 _11344_ (
    .A(_11217_[20]),
    .ZN(_05785_)
  );
  INV_X1 _11345_ (
    .A(_11217_[21]),
    .ZN(_05796_)
  );
  INV_X1 _11346_ (
    .A(_11217_[22]),
    .ZN(_05807_)
  );
  INV_X1 _11347_ (
    .A(_11217_[23]),
    .ZN(_05818_)
  );
  INV_X1 _11348_ (
    .A(_11217_[24]),
    .ZN(_05829_)
  );
  INV_X1 _11349_ (
    .A(_11217_[25]),
    .ZN(_05840_)
  );
  INV_X1 _11350_ (
    .A(_11217_[26]),
    .ZN(_05851_)
  );
  INV_X1 _11351_ (
    .A(_11217_[27]),
    .ZN(_05862_)
  );
  INV_X1 _11352_ (
    .A(_11217_[28]),
    .ZN(_05873_)
  );
  INV_X1 _11353_ (
    .A(_11217_[29]),
    .ZN(_05884_)
  );
  INV_X1 _11354_ (
    .A(_11217_[30]),
    .ZN(_05895_)
  );
  INV_X1 _11355_ (
    .A(_11217_[31]),
    .ZN(_05906_)
  );
  INV_X1 _11356_ (
    .A(_11217_[32]),
    .ZN(_05917_)
  );
  AND2_X1 _11357_ (
    .A1(_04799_),
    .A2(_04810_),
    .ZN(_05928_)
  );
  AND2_X1 _11358_ (
    .A1(_04820_),
    .A2(_04831_),
    .ZN(_05939_)
  );
  AND2_X1 _11359_ (
    .A1(_05928_),
    .A2(_05939_),
    .ZN(_05950_)
  );
  AND2_X1 _11360_ (
    .A1(_05511_),
    .A2(_05522_),
    .ZN(_05961_)
  );
  INV_X1 _11361_ (
    .A(_05961_),
    .ZN(_05972_)
  );
  AND2_X1 _11362_ (
    .A1(_05434_),
    .A2(_05961_),
    .ZN(_05983_)
  );
  INV_X1 _11363_ (
    .A(_05983_),
    .ZN(_05994_)
  );
  AND2_X1 _11364_ (
    .A1(_04788_),
    .A2(_05500_),
    .ZN(_06005_)
  );
  AND2_X1 _11365_ (
    .A1(_05983_),
    .A2(_06005_),
    .ZN(_06016_)
  );
  AND2_X1 _11366_ (
    .A1(_05950_),
    .A2(_06016_),
    .ZN(_06027_)
  );
  INV_X1 _11367_ (
    .A(_06027_),
    .ZN(_06038_)
  );
  AND2_X1 _11368_ (
    .A1(_04777_),
    .A2(_04788_),
    .ZN(_06048_)
  );
  AND2_X1 _11369_ (
    .A1(_05928_),
    .A2(_06048_),
    .ZN(_06059_)
  );
  AND2_X1 _11370_ (
    .A1(_05467_),
    .A2(_06059_),
    .ZN(_06070_)
  );
  AND2_X1 _11371_ (
    .A1(_05423_),
    .A2(_05522_),
    .ZN(_06081_)
  );
  INV_X1 _11372_ (
    .A(_06081_),
    .ZN(_06092_)
  );
  AND2_X1 _11373_ (
    .A1(_05434_),
    .A2(_06081_),
    .ZN(_06103_)
  );
  INV_X1 _11374_ (
    .A(_06103_),
    .ZN(_06114_)
  );
  AND2_X1 _11375_ (
    .A1(_05478_),
    .A2(_06103_),
    .ZN(_06125_)
  );
  AND2_X1 _11376_ (
    .A1(_06070_),
    .A2(_06125_),
    .ZN(_06136_)
  );
  INV_X1 _11377_ (
    .A(_06136_),
    .ZN(_06147_)
  );
  AND2_X1 _11378_ (
    .A1(_06038_),
    .A2(_06147_),
    .ZN(_06158_)
  );
  AND2_X1 _11379_ (
    .A1(_05412_),
    .A2(_05434_),
    .ZN(_06169_)
  );
  AND2_X1 _11380_ (
    .A1(_05423_),
    .A2(_06169_),
    .ZN(io_req_ready)
  );
  AND2_X1 _11381_ (
    .A1(io_req_valid),
    .A2(io_req_ready),
    .ZN(_06190_)
  );
  INV_X1 _11382_ (
    .A(_06190_),
    .ZN(_06201_)
  );
  AND2_X1 _11383_ (
    .A1(isHi),
    .A2(_06201_),
    .ZN(_06212_)
  );
  AND2_X1 _11384_ (
    .A1(resHi),
    .A2(_06201_),
    .ZN(_06223_)
  );
  AND2_X1 _11385_ (
    .A1(_05412_),
    .A2(_05511_),
    .ZN(_06234_)
  );
  AND2_X1 _11386_ (
    .A1(_05489_),
    .A2(_06234_),
    .ZN(_06245_)
  );
  INV_X1 _11387_ (
    .A(_06245_),
    .ZN(_06256_)
  );
  AND2_X1 _11388_ (
    .A1(_06158_),
    .A2(_06256_),
    .ZN(_06267_)
  );
  AND2_X1 _11389_ (
    .A1(_06223_),
    .A2(_06256_),
    .ZN(_06278_)
  );
  MUX2_X1 _11390_ (
    .A(_06212_),
    .B(_06278_),
    .S(_06158_),
    .Z(_00005_)
  );
  AND2_X1 _11391_ (
    .A1(_05434_),
    .A2(_06234_),
    .ZN(_06299_)
  );
  INV_X1 _11392_ (
    .A(_06299_),
    .ZN(_06310_)
  );
  AND2_X1 _11393_ (
    .A1(_06256_),
    .A2(_06310_),
    .ZN(_06321_)
  );
  AND2_X1 _11394_ (
    .A1(_05423_),
    .A2(_06321_),
    .ZN(_06332_)
  );
  INV_X1 _11395_ (
    .A(_06332_),
    .ZN(_06343_)
  );
  AND2_X1 _11396_ (
    .A1(_06147_),
    .A2(_06343_),
    .ZN(_06354_)
  );
  INV_X1 _11397_ (
    .A(_06354_),
    .ZN(_06365_)
  );
  AND2_X1 _11398_ (
    .A1(_06038_),
    .A2(_06365_),
    .ZN(_06375_)
  );
  INV_X1 _11399_ (
    .A(_06375_),
    .ZN(_06386_)
  );
  AND2_X1 _11400_ (
    .A1(_05972_),
    .A2(_06092_),
    .ZN(_06397_)
  );
  INV_X1 _11401_ (
    .A(_06397_),
    .ZN(_06408_)
  );
  AND2_X1 _11402_ (
    .A1(_05489_),
    .A2(_06408_),
    .ZN(io_resp_valid)
  );
  AND2_X1 _11403_ (
    .A1(io_resp_ready),
    .A2(io_resp_valid),
    .ZN(_06429_)
  );
  INV_X1 _11404_ (
    .A(_06429_),
    .ZN(_06440_)
  );
  AND2_X1 _11405_ (
    .A1(_05555_),
    .A2(_06440_),
    .ZN(_06451_)
  );
  AND2_X1 _11406_ (
    .A1(_06201_),
    .A2(_06451_),
    .ZN(_06462_)
  );
  AND2_X1 _11407_ (
    .A1(_06386_),
    .A2(_06462_),
    .ZN(_06473_)
  );
  INV_X1 _11408_ (
    .A(_06473_),
    .ZN(_06484_)
  );
  AND2_X1 _11409_ (
    .A1(io_req_bits_fn[2]),
    .A2(_06190_),
    .ZN(_06495_)
  );
  INV_X1 _11410_ (
    .A(_06495_),
    .ZN(_06506_)
  );
  AND2_X1 _11411_ (
    .A1(_06484_),
    .A2(_06506_),
    .ZN(_06517_)
  );
  INV_X1 _11412_ (
    .A(_06517_),
    .ZN(_06528_)
  );
  AND2_X1 _11413_ (
    .A1(_04842_),
    .A2(_06528_),
    .ZN(_00006_)
  );
  AND2_X1 _11414_ (
    .A1(_05412_),
    .A2(_06321_),
    .ZN(_06549_)
  );
  AND2_X1 _11415_ (
    .A1(_06158_),
    .A2(_06549_),
    .ZN(_06560_)
  );
  INV_X1 _11416_ (
    .A(_06560_),
    .ZN(_06571_)
  );
  AND2_X1 _11417_ (
    .A1(_05544_),
    .A2(_06027_),
    .ZN(_06582_)
  );
  INV_X1 _11418_ (
    .A(_06582_),
    .ZN(_06593_)
  );
  AND2_X1 _11419_ (
    .A1(_06451_),
    .A2(_06593_),
    .ZN(_06604_)
  );
  AND2_X1 _11420_ (
    .A1(_06571_),
    .A2(_06604_),
    .ZN(_06615_)
  );
  INV_X1 _11421_ (
    .A(_06615_),
    .ZN(_06626_)
  );
  AND2_X1 _11422_ (
    .A1(_06201_),
    .A2(_06626_),
    .ZN(_06637_)
  );
  INV_X1 _11423_ (
    .A(_06637_),
    .ZN(_06648_)
  );
  AND2_X1 _11424_ (
    .A1(_05445_),
    .A2(_05456_),
    .ZN(_06659_)
  );
  INV_X1 _11425_ (
    .A(_06659_),
    .ZN(_06670_)
  );
  AND2_X1 _11426_ (
    .A1(io_req_bits_fn[0]),
    .A2(_06670_),
    .ZN(_06681_)
  );
  INV_X1 _11427_ (
    .A(_06681_),
    .ZN(_06691_)
  );
  AND2_X1 _11428_ (
    .A1(io_req_bits_in1[31]),
    .A2(_06691_),
    .ZN(_06702_)
  );
  INV_X1 _11429_ (
    .A(_06702_),
    .ZN(_06713_)
  );
  MUX2_X1 _11430_ (
    .A(io_req_bits_fn[1]),
    .B(io_req_bits_fn[0]),
    .S(io_req_bits_fn[2]),
    .Z(_06724_)
  );
  INV_X1 _11431_ (
    .A(_06724_),
    .ZN(_06735_)
  );
  AND2_X1 _11432_ (
    .A1(io_req_bits_in2[31]),
    .A2(_06735_),
    .ZN(_06746_)
  );
  INV_X1 _11433_ (
    .A(_06746_),
    .ZN(_06757_)
  );
  AND2_X1 _11434_ (
    .A1(_06713_),
    .A2(_06757_),
    .ZN(_06768_)
  );
  INV_X1 _11435_ (
    .A(_06768_),
    .ZN(_06779_)
  );
  AND2_X1 _11436_ (
    .A1(_06495_),
    .A2(_06779_),
    .ZN(_06790_)
  );
  INV_X1 _11437_ (
    .A(_06790_),
    .ZN(_06801_)
  );
  AND2_X1 _11438_ (
    .A1(_04842_),
    .A2(_06801_),
    .ZN(_06812_)
  );
  AND2_X1 _11439_ (
    .A1(_06648_),
    .A2(_06812_),
    .ZN(_00007_)
  );
  AND2_X1 _11440_ (
    .A1(_04426_),
    .A2(_05906_),
    .ZN(_06833_)
  );
  INV_X1 _11441_ (
    .A(_06833_),
    .ZN(_06844_)
  );
  AND2_X1 _11442_ (
    .A1(remainder[63]),
    .A2(_11217_[31]),
    .ZN(_06855_)
  );
  INV_X1 _11443_ (
    .A(_06855_),
    .ZN(_06866_)
  );
  AND2_X1 _11444_ (
    .A1(remainder[62]),
    .A2(_11217_[30]),
    .ZN(_06877_)
  );
  INV_X1 _11445_ (
    .A(_06877_),
    .ZN(_06888_)
  );
  AND2_X1 _11446_ (
    .A1(_04437_),
    .A2(_05895_),
    .ZN(_06899_)
  );
  INV_X1 _11447_ (
    .A(_06899_),
    .ZN(_06910_)
  );
  AND2_X1 _11448_ (
    .A1(_06888_),
    .A2(_06910_),
    .ZN(_06921_)
  );
  INV_X1 _11449_ (
    .A(_06921_),
    .ZN(_06932_)
  );
  AND2_X1 _11450_ (
    .A1(_04448_),
    .A2(_05884_),
    .ZN(_06943_)
  );
  INV_X1 _11451_ (
    .A(_06943_),
    .ZN(_06954_)
  );
  AND2_X1 _11452_ (
    .A1(remainder[61]),
    .A2(_11217_[29]),
    .ZN(_06965_)
  );
  INV_X1 _11453_ (
    .A(_06965_),
    .ZN(_06976_)
  );
  AND2_X1 _11454_ (
    .A1(remainder[60]),
    .A2(_11217_[28]),
    .ZN(_06987_)
  );
  INV_X1 _11455_ (
    .A(_06987_),
    .ZN(_06997_)
  );
  AND2_X1 _11456_ (
    .A1(_04459_),
    .A2(_05873_),
    .ZN(_07008_)
  );
  INV_X1 _11457_ (
    .A(_07008_),
    .ZN(_07019_)
  );
  AND2_X1 _11458_ (
    .A1(_06997_),
    .A2(_07019_),
    .ZN(_07030_)
  );
  INV_X1 _11459_ (
    .A(_07030_),
    .ZN(_07041_)
  );
  AND2_X1 _11460_ (
    .A1(remainder[59]),
    .A2(_11217_[27]),
    .ZN(_07052_)
  );
  INV_X1 _11461_ (
    .A(_07052_),
    .ZN(_07063_)
  );
  AND2_X1 _11462_ (
    .A1(_04470_),
    .A2(_05862_),
    .ZN(_07074_)
  );
  INV_X1 _11463_ (
    .A(_07074_),
    .ZN(_07085_)
  );
  AND2_X1 _11464_ (
    .A1(remainder[58]),
    .A2(_11217_[26]),
    .ZN(_07096_)
  );
  INV_X1 _11465_ (
    .A(_07096_),
    .ZN(_07107_)
  );
  AND2_X1 _11466_ (
    .A1(_04481_),
    .A2(_05851_),
    .ZN(_07118_)
  );
  INV_X1 _11467_ (
    .A(_07118_),
    .ZN(_07129_)
  );
  AND2_X1 _11468_ (
    .A1(_07107_),
    .A2(_07129_),
    .ZN(_07140_)
  );
  INV_X1 _11469_ (
    .A(_07140_),
    .ZN(_07151_)
  );
  AND2_X1 _11470_ (
    .A1(_04492_),
    .A2(_05840_),
    .ZN(_07162_)
  );
  INV_X1 _11471_ (
    .A(_07162_),
    .ZN(_07173_)
  );
  AND2_X1 _11472_ (
    .A1(remainder[57]),
    .A2(_11217_[25]),
    .ZN(_07184_)
  );
  INV_X1 _11473_ (
    .A(_07184_),
    .ZN(_07195_)
  );
  AND2_X1 _11474_ (
    .A1(remainder[56]),
    .A2(_11217_[24]),
    .ZN(_07206_)
  );
  INV_X1 _11475_ (
    .A(_07206_),
    .ZN(_07217_)
  );
  AND2_X1 _11476_ (
    .A1(_04503_),
    .A2(_05829_),
    .ZN(_07228_)
  );
  INV_X1 _11477_ (
    .A(_07228_),
    .ZN(_07239_)
  );
  AND2_X1 _11478_ (
    .A1(_07217_),
    .A2(_07239_),
    .ZN(_07250_)
  );
  INV_X1 _11479_ (
    .A(_07250_),
    .ZN(_07261_)
  );
  AND2_X1 _11480_ (
    .A1(remainder[55]),
    .A2(_11217_[23]),
    .ZN(_07272_)
  );
  INV_X1 _11481_ (
    .A(_07272_),
    .ZN(_07283_)
  );
  AND2_X1 _11482_ (
    .A1(_04514_),
    .A2(_05818_),
    .ZN(_07293_)
  );
  INV_X1 _11483_ (
    .A(_07293_),
    .ZN(_07304_)
  );
  AND2_X1 _11484_ (
    .A1(remainder[54]),
    .A2(_11217_[22]),
    .ZN(_07315_)
  );
  INV_X1 _11485_ (
    .A(_07315_),
    .ZN(_07326_)
  );
  AND2_X1 _11486_ (
    .A1(_04525_),
    .A2(_05807_),
    .ZN(_07337_)
  );
  INV_X1 _11487_ (
    .A(_07337_),
    .ZN(_07348_)
  );
  AND2_X1 _11488_ (
    .A1(_07326_),
    .A2(_07348_),
    .ZN(_07359_)
  );
  INV_X1 _11489_ (
    .A(_07359_),
    .ZN(_07370_)
  );
  AND2_X1 _11490_ (
    .A1(remainder[53]),
    .A2(_11217_[21]),
    .ZN(_07381_)
  );
  INV_X1 _11491_ (
    .A(_07381_),
    .ZN(_07392_)
  );
  AND2_X1 _11492_ (
    .A1(_04536_),
    .A2(_05796_),
    .ZN(_07403_)
  );
  INV_X1 _11493_ (
    .A(_07403_),
    .ZN(_07414_)
  );
  AND2_X1 _11494_ (
    .A1(remainder[52]),
    .A2(_11217_[20]),
    .ZN(_07425_)
  );
  INV_X1 _11495_ (
    .A(_07425_),
    .ZN(_07436_)
  );
  AND2_X1 _11496_ (
    .A1(_04546_),
    .A2(_05785_),
    .ZN(_07447_)
  );
  INV_X1 _11497_ (
    .A(_07447_),
    .ZN(_07458_)
  );
  AND2_X1 _11498_ (
    .A1(_07436_),
    .A2(_07458_),
    .ZN(_07469_)
  );
  INV_X1 _11499_ (
    .A(_07469_),
    .ZN(_07480_)
  );
  AND2_X1 _11500_ (
    .A1(remainder[51]),
    .A2(_11217_[19]),
    .ZN(_07491_)
  );
  INV_X1 _11501_ (
    .A(_07491_),
    .ZN(_07502_)
  );
  AND2_X1 _11502_ (
    .A1(_04557_),
    .A2(_05774_),
    .ZN(_07513_)
  );
  INV_X1 _11503_ (
    .A(_07513_),
    .ZN(_07524_)
  );
  AND2_X1 _11504_ (
    .A1(remainder[50]),
    .A2(_11217_[18]),
    .ZN(_07535_)
  );
  INV_X1 _11505_ (
    .A(_07535_),
    .ZN(_07546_)
  );
  AND2_X1 _11506_ (
    .A1(_04568_),
    .A2(_05763_),
    .ZN(_07557_)
  );
  INV_X1 _11507_ (
    .A(_07557_),
    .ZN(_07568_)
  );
  AND2_X1 _11508_ (
    .A1(_07546_),
    .A2(_07568_),
    .ZN(_07579_)
  );
  INV_X1 _11509_ (
    .A(_07579_),
    .ZN(_07590_)
  );
  AND2_X1 _11510_ (
    .A1(remainder[49]),
    .A2(_11217_[17]),
    .ZN(_07600_)
  );
  INV_X1 _11511_ (
    .A(_07600_),
    .ZN(_07611_)
  );
  AND2_X1 _11512_ (
    .A1(_04579_),
    .A2(_05752_),
    .ZN(_07622_)
  );
  INV_X1 _11513_ (
    .A(_07622_),
    .ZN(_07633_)
  );
  AND2_X1 _11514_ (
    .A1(remainder[48]),
    .A2(_11217_[16]),
    .ZN(_07644_)
  );
  INV_X1 _11515_ (
    .A(_07644_),
    .ZN(_07655_)
  );
  AND2_X1 _11516_ (
    .A1(_04590_),
    .A2(_05741_),
    .ZN(_07666_)
  );
  INV_X1 _11517_ (
    .A(_07666_),
    .ZN(_07677_)
  );
  AND2_X1 _11518_ (
    .A1(_07655_),
    .A2(_07677_),
    .ZN(_07688_)
  );
  INV_X1 _11519_ (
    .A(_07688_),
    .ZN(_07699_)
  );
  AND2_X1 _11520_ (
    .A1(remainder[47]),
    .A2(_11217_[15]),
    .ZN(_07710_)
  );
  INV_X1 _11521_ (
    .A(_07710_),
    .ZN(_07721_)
  );
  AND2_X1 _11522_ (
    .A1(_04601_),
    .A2(_05730_),
    .ZN(_07732_)
  );
  INV_X1 _11523_ (
    .A(_07732_),
    .ZN(_07743_)
  );
  AND2_X1 _11524_ (
    .A1(remainder[46]),
    .A2(_11217_[14]),
    .ZN(_07754_)
  );
  INV_X1 _11525_ (
    .A(_07754_),
    .ZN(_07765_)
  );
  AND2_X1 _11526_ (
    .A1(_04612_),
    .A2(_05720_),
    .ZN(_07776_)
  );
  INV_X1 _11527_ (
    .A(_07776_),
    .ZN(_07787_)
  );
  AND2_X1 _11528_ (
    .A1(_07765_),
    .A2(_07787_),
    .ZN(_07798_)
  );
  INV_X1 _11529_ (
    .A(_07798_),
    .ZN(_07809_)
  );
  AND2_X1 _11530_ (
    .A1(remainder[45]),
    .A2(_11217_[13]),
    .ZN(_07820_)
  );
  INV_X1 _11531_ (
    .A(_07820_),
    .ZN(_07831_)
  );
  AND2_X1 _11532_ (
    .A1(_04623_),
    .A2(_05709_),
    .ZN(_07842_)
  );
  INV_X1 _11533_ (
    .A(_07842_),
    .ZN(_07853_)
  );
  AND2_X1 _11534_ (
    .A1(remainder[44]),
    .A2(_11217_[12]),
    .ZN(_07864_)
  );
  INV_X1 _11535_ (
    .A(_07864_),
    .ZN(_07875_)
  );
  AND2_X1 _11536_ (
    .A1(_04634_),
    .A2(_05698_),
    .ZN(_07886_)
  );
  INV_X1 _11537_ (
    .A(_07886_),
    .ZN(_07896_)
  );
  AND2_X1 _11538_ (
    .A1(_07875_),
    .A2(_07896_),
    .ZN(_07907_)
  );
  INV_X1 _11539_ (
    .A(_07907_),
    .ZN(_07918_)
  );
  AND2_X1 _11540_ (
    .A1(remainder[43]),
    .A2(_11217_[11]),
    .ZN(_07929_)
  );
  INV_X1 _11541_ (
    .A(_07929_),
    .ZN(_07940_)
  );
  AND2_X1 _11542_ (
    .A1(_04645_),
    .A2(_05687_),
    .ZN(_07951_)
  );
  INV_X1 _11543_ (
    .A(_07951_),
    .ZN(_07962_)
  );
  AND2_X1 _11544_ (
    .A1(remainder[42]),
    .A2(_11217_[10]),
    .ZN(_07973_)
  );
  INV_X1 _11545_ (
    .A(_07973_),
    .ZN(_07984_)
  );
  AND2_X1 _11546_ (
    .A1(_04656_),
    .A2(_05676_),
    .ZN(_07995_)
  );
  INV_X1 _11547_ (
    .A(_07995_),
    .ZN(_08006_)
  );
  AND2_X1 _11548_ (
    .A1(_07984_),
    .A2(_08006_),
    .ZN(_08017_)
  );
  INV_X1 _11549_ (
    .A(_08017_),
    .ZN(_08028_)
  );
  AND2_X1 _11550_ (
    .A1(remainder[41]),
    .A2(_11217_[9]),
    .ZN(_08039_)
  );
  INV_X1 _11551_ (
    .A(_08039_),
    .ZN(_08050_)
  );
  AND2_X1 _11552_ (
    .A1(_04667_),
    .A2(_05665_),
    .ZN(_08061_)
  );
  INV_X1 _11553_ (
    .A(_08061_),
    .ZN(_08072_)
  );
  AND2_X1 _11554_ (
    .A1(remainder[40]),
    .A2(_11217_[8]),
    .ZN(_08083_)
  );
  INV_X1 _11555_ (
    .A(_08083_),
    .ZN(_08094_)
  );
  AND2_X1 _11556_ (
    .A1(_04678_),
    .A2(_05654_),
    .ZN(_08105_)
  );
  INV_X1 _11557_ (
    .A(_08105_),
    .ZN(_08116_)
  );
  AND2_X1 _11558_ (
    .A1(_08094_),
    .A2(_08116_),
    .ZN(_08127_)
  );
  INV_X1 _11559_ (
    .A(_08127_),
    .ZN(_08138_)
  );
  AND2_X1 _11560_ (
    .A1(remainder[39]),
    .A2(_11217_[7]),
    .ZN(_08149_)
  );
  INV_X1 _11561_ (
    .A(_08149_),
    .ZN(_08160_)
  );
  AND2_X1 _11562_ (
    .A1(_04689_),
    .A2(_05643_),
    .ZN(_08171_)
  );
  INV_X1 _11563_ (
    .A(_08171_),
    .ZN(_08182_)
  );
  AND2_X1 _11564_ (
    .A1(remainder[38]),
    .A2(_11217_[6]),
    .ZN(_08193_)
  );
  INV_X1 _11565_ (
    .A(_08193_),
    .ZN(_08203_)
  );
  AND2_X1 _11566_ (
    .A1(_04700_),
    .A2(_05632_),
    .ZN(_08214_)
  );
  INV_X1 _11567_ (
    .A(_08214_),
    .ZN(_08225_)
  );
  AND2_X1 _11568_ (
    .A1(_08203_),
    .A2(_08225_),
    .ZN(_08236_)
  );
  INV_X1 _11569_ (
    .A(_08236_),
    .ZN(_08247_)
  );
  AND2_X1 _11570_ (
    .A1(remainder[37]),
    .A2(_11217_[5]),
    .ZN(_08258_)
  );
  INV_X1 _11571_ (
    .A(_08258_),
    .ZN(_08269_)
  );
  AND2_X1 _11572_ (
    .A1(remainder[36]),
    .A2(_11217_[4]),
    .ZN(_08280_)
  );
  INV_X1 _11573_ (
    .A(_08280_),
    .ZN(_08291_)
  );
  AND2_X1 _11574_ (
    .A1(_04722_),
    .A2(_05610_),
    .ZN(_08302_)
  );
  INV_X1 _11575_ (
    .A(_08302_),
    .ZN(_08313_)
  );
  AND2_X1 _11576_ (
    .A1(_08291_),
    .A2(_08313_),
    .ZN(_08324_)
  );
  INV_X1 _11577_ (
    .A(_08324_),
    .ZN(_08335_)
  );
  AND2_X1 _11578_ (
    .A1(remainder[35]),
    .A2(_11217_[3]),
    .ZN(_08346_)
  );
  INV_X1 _11579_ (
    .A(_08346_),
    .ZN(_08357_)
  );
  AND2_X1 _11580_ (
    .A1(_04733_),
    .A2(_05599_),
    .ZN(_08368_)
  );
  INV_X1 _11581_ (
    .A(_08368_),
    .ZN(_08379_)
  );
  AND2_X1 _11582_ (
    .A1(remainder[34]),
    .A2(_11217_[2]),
    .ZN(_08390_)
  );
  INV_X1 _11583_ (
    .A(_08390_),
    .ZN(_08401_)
  );
  AND2_X1 _11584_ (
    .A1(remainder[33]),
    .A2(_11217_[1]),
    .ZN(_08412_)
  );
  INV_X1 _11585_ (
    .A(_08412_),
    .ZN(_08423_)
  );
  AND2_X1 _11586_ (
    .A1(_04766_),
    .A2(_05566_),
    .ZN(_08434_)
  );
  INV_X1 _11587_ (
    .A(_08434_),
    .ZN(_08445_)
  );
  AND2_X1 _11588_ (
    .A1(_04755_),
    .A2(_05577_),
    .ZN(_08456_)
  );
  INV_X1 _11589_ (
    .A(_08456_),
    .ZN(_08467_)
  );
  AND2_X1 _11590_ (
    .A1(_08423_),
    .A2(_08467_),
    .ZN(_08478_)
  );
  INV_X1 _11591_ (
    .A(_08478_),
    .ZN(_08489_)
  );
  AND2_X1 _11592_ (
    .A1(_08445_),
    .A2(_08478_),
    .ZN(_08500_)
  );
  INV_X1 _11593_ (
    .A(_08500_),
    .ZN(_08510_)
  );
  AND2_X1 _11594_ (
    .A1(_08423_),
    .A2(_08510_),
    .ZN(_08521_)
  );
  INV_X1 _11595_ (
    .A(_08521_),
    .ZN(_08532_)
  );
  AND2_X1 _11596_ (
    .A1(_04744_),
    .A2(_05588_),
    .ZN(_08543_)
  );
  INV_X1 _11597_ (
    .A(_08543_),
    .ZN(_08554_)
  );
  AND2_X1 _11598_ (
    .A1(_08401_),
    .A2(_08554_),
    .ZN(_08565_)
  );
  INV_X1 _11599_ (
    .A(_08565_),
    .ZN(_08576_)
  );
  AND2_X1 _11600_ (
    .A1(_08532_),
    .A2(_08565_),
    .ZN(_08587_)
  );
  INV_X1 _11601_ (
    .A(_08587_),
    .ZN(_08598_)
  );
  AND2_X1 _11602_ (
    .A1(_08401_),
    .A2(_08598_),
    .ZN(_08609_)
  );
  INV_X1 _11603_ (
    .A(_08609_),
    .ZN(_08620_)
  );
  AND2_X1 _11604_ (
    .A1(_08379_),
    .A2(_08620_),
    .ZN(_08631_)
  );
  INV_X1 _11605_ (
    .A(_08631_),
    .ZN(_08642_)
  );
  AND2_X1 _11606_ (
    .A1(_08357_),
    .A2(_08609_),
    .ZN(_08653_)
  );
  INV_X1 _11607_ (
    .A(_08653_),
    .ZN(_08664_)
  );
  AND2_X1 _11608_ (
    .A1(_08357_),
    .A2(_08642_),
    .ZN(_08675_)
  );
  AND2_X1 _11609_ (
    .A1(_08379_),
    .A2(_08664_),
    .ZN(_08686_)
  );
  AND2_X1 _11610_ (
    .A1(_08324_),
    .A2(_08686_),
    .ZN(_08697_)
  );
  INV_X1 _11611_ (
    .A(_08697_),
    .ZN(_08708_)
  );
  AND2_X1 _11612_ (
    .A1(_08291_),
    .A2(_08708_),
    .ZN(_08719_)
  );
  INV_X1 _11613_ (
    .A(_08719_),
    .ZN(_08730_)
  );
  AND2_X1 _11614_ (
    .A1(_04711_),
    .A2(_05621_),
    .ZN(_08741_)
  );
  INV_X1 _11615_ (
    .A(_08741_),
    .ZN(_08752_)
  );
  AND2_X1 _11616_ (
    .A1(_08269_),
    .A2(_08752_),
    .ZN(_08763_)
  );
  INV_X1 _11617_ (
    .A(_08763_),
    .ZN(_08774_)
  );
  AND2_X1 _11618_ (
    .A1(_08730_),
    .A2(_08763_),
    .ZN(_08785_)
  );
  INV_X1 _11619_ (
    .A(_08785_),
    .ZN(_08796_)
  );
  AND2_X1 _11620_ (
    .A1(_08269_),
    .A2(_08796_),
    .ZN(_08807_)
  );
  INV_X1 _11621_ (
    .A(_08807_),
    .ZN(_08818_)
  );
  AND2_X1 _11622_ (
    .A1(_08236_),
    .A2(_08818_),
    .ZN(_08828_)
  );
  INV_X1 _11623_ (
    .A(_08828_),
    .ZN(_08839_)
  );
  AND2_X1 _11624_ (
    .A1(_08203_),
    .A2(_08839_),
    .ZN(_08850_)
  );
  INV_X1 _11625_ (
    .A(_08850_),
    .ZN(_08861_)
  );
  AND2_X1 _11626_ (
    .A1(_08182_),
    .A2(_08861_),
    .ZN(_08872_)
  );
  INV_X1 _11627_ (
    .A(_08872_),
    .ZN(_08883_)
  );
  AND2_X1 _11628_ (
    .A1(_08160_),
    .A2(_08850_),
    .ZN(_08894_)
  );
  INV_X1 _11629_ (
    .A(_08894_),
    .ZN(_08905_)
  );
  AND2_X1 _11630_ (
    .A1(_08160_),
    .A2(_08883_),
    .ZN(_08916_)
  );
  AND2_X1 _11631_ (
    .A1(_08182_),
    .A2(_08905_),
    .ZN(_08927_)
  );
  AND2_X1 _11632_ (
    .A1(_08127_),
    .A2(_08927_),
    .ZN(_08938_)
  );
  INV_X1 _11633_ (
    .A(_08938_),
    .ZN(_08949_)
  );
  AND2_X1 _11634_ (
    .A1(_08094_),
    .A2(_08949_),
    .ZN(_08960_)
  );
  INV_X1 _11635_ (
    .A(_08960_),
    .ZN(_08971_)
  );
  AND2_X1 _11636_ (
    .A1(_08072_),
    .A2(_08971_),
    .ZN(_08982_)
  );
  INV_X1 _11637_ (
    .A(_08982_),
    .ZN(_08993_)
  );
  AND2_X1 _11638_ (
    .A1(_08050_),
    .A2(_08960_),
    .ZN(_09004_)
  );
  INV_X1 _11639_ (
    .A(_09004_),
    .ZN(_09015_)
  );
  AND2_X1 _11640_ (
    .A1(_08050_),
    .A2(_08993_),
    .ZN(_09026_)
  );
  AND2_X1 _11641_ (
    .A1(_08072_),
    .A2(_09015_),
    .ZN(_09037_)
  );
  AND2_X1 _11642_ (
    .A1(_08017_),
    .A2(_09037_),
    .ZN(_09048_)
  );
  INV_X1 _11643_ (
    .A(_09048_),
    .ZN(_09059_)
  );
  AND2_X1 _11644_ (
    .A1(_07984_),
    .A2(_09059_),
    .ZN(_09070_)
  );
  INV_X1 _11645_ (
    .A(_09070_),
    .ZN(_09081_)
  );
  AND2_X1 _11646_ (
    .A1(_07962_),
    .A2(_09081_),
    .ZN(_09092_)
  );
  INV_X1 _11647_ (
    .A(_09092_),
    .ZN(_09103_)
  );
  AND2_X1 _11648_ (
    .A1(_07940_),
    .A2(_09070_),
    .ZN(_09114_)
  );
  INV_X1 _11649_ (
    .A(_09114_),
    .ZN(_09125_)
  );
  AND2_X1 _11650_ (
    .A1(_07940_),
    .A2(_09103_),
    .ZN(_09135_)
  );
  AND2_X1 _11651_ (
    .A1(_07962_),
    .A2(_09125_),
    .ZN(_09146_)
  );
  AND2_X1 _11652_ (
    .A1(_07907_),
    .A2(_09146_),
    .ZN(_09157_)
  );
  INV_X1 _11653_ (
    .A(_09157_),
    .ZN(_09168_)
  );
  AND2_X1 _11654_ (
    .A1(_07875_),
    .A2(_09168_),
    .ZN(_09179_)
  );
  INV_X1 _11655_ (
    .A(_09179_),
    .ZN(_09190_)
  );
  AND2_X1 _11656_ (
    .A1(_07853_),
    .A2(_09190_),
    .ZN(_09201_)
  );
  INV_X1 _11657_ (
    .A(_09201_),
    .ZN(_09212_)
  );
  AND2_X1 _11658_ (
    .A1(_07831_),
    .A2(_09179_),
    .ZN(_09223_)
  );
  INV_X1 _11659_ (
    .A(_09223_),
    .ZN(_09234_)
  );
  AND2_X1 _11660_ (
    .A1(_07831_),
    .A2(_09212_),
    .ZN(_09245_)
  );
  AND2_X1 _11661_ (
    .A1(_07853_),
    .A2(_09234_),
    .ZN(_09256_)
  );
  AND2_X1 _11662_ (
    .A1(_07798_),
    .A2(_09256_),
    .ZN(_09267_)
  );
  INV_X1 _11663_ (
    .A(_09267_),
    .ZN(_09278_)
  );
  AND2_X1 _11664_ (
    .A1(_07765_),
    .A2(_09278_),
    .ZN(_09289_)
  );
  INV_X1 _11665_ (
    .A(_09289_),
    .ZN(_09300_)
  );
  AND2_X1 _11666_ (
    .A1(_07743_),
    .A2(_09300_),
    .ZN(_09311_)
  );
  INV_X1 _11667_ (
    .A(_09311_),
    .ZN(_09322_)
  );
  AND2_X1 _11668_ (
    .A1(_07721_),
    .A2(_09289_),
    .ZN(_09333_)
  );
  INV_X1 _11669_ (
    .A(_09333_),
    .ZN(_09344_)
  );
  AND2_X1 _11670_ (
    .A1(_07721_),
    .A2(_09322_),
    .ZN(_09355_)
  );
  AND2_X1 _11671_ (
    .A1(_07743_),
    .A2(_09344_),
    .ZN(_09366_)
  );
  AND2_X1 _11672_ (
    .A1(_07688_),
    .A2(_09366_),
    .ZN(_09377_)
  );
  INV_X1 _11673_ (
    .A(_09377_),
    .ZN(_09388_)
  );
  AND2_X1 _11674_ (
    .A1(_07655_),
    .A2(_09388_),
    .ZN(_09399_)
  );
  INV_X1 _11675_ (
    .A(_09399_),
    .ZN(_09410_)
  );
  AND2_X1 _11676_ (
    .A1(_07633_),
    .A2(_09410_),
    .ZN(_09421_)
  );
  INV_X1 _11677_ (
    .A(_09421_),
    .ZN(_09432_)
  );
  AND2_X1 _11678_ (
    .A1(_07611_),
    .A2(_09399_),
    .ZN(_09443_)
  );
  INV_X1 _11679_ (
    .A(_09443_),
    .ZN(_09453_)
  );
  AND2_X1 _11680_ (
    .A1(_07611_),
    .A2(_09432_),
    .ZN(_09464_)
  );
  AND2_X1 _11681_ (
    .A1(_07633_),
    .A2(_09453_),
    .ZN(_09475_)
  );
  AND2_X1 _11682_ (
    .A1(_07579_),
    .A2(_09475_),
    .ZN(_09486_)
  );
  INV_X1 _11683_ (
    .A(_09486_),
    .ZN(_09497_)
  );
  AND2_X1 _11684_ (
    .A1(_07546_),
    .A2(_09497_),
    .ZN(_09508_)
  );
  INV_X1 _11685_ (
    .A(_09508_),
    .ZN(_09519_)
  );
  AND2_X1 _11686_ (
    .A1(_07524_),
    .A2(_09519_),
    .ZN(_09530_)
  );
  INV_X1 _11687_ (
    .A(_09530_),
    .ZN(_09541_)
  );
  AND2_X1 _11688_ (
    .A1(_07502_),
    .A2(_09508_),
    .ZN(_09552_)
  );
  INV_X1 _11689_ (
    .A(_09552_),
    .ZN(_09563_)
  );
  AND2_X1 _11690_ (
    .A1(_07502_),
    .A2(_09541_),
    .ZN(_09574_)
  );
  AND2_X1 _11691_ (
    .A1(_07524_),
    .A2(_09563_),
    .ZN(_09585_)
  );
  AND2_X1 _11692_ (
    .A1(_07469_),
    .A2(_09585_),
    .ZN(_09596_)
  );
  INV_X1 _11693_ (
    .A(_09596_),
    .ZN(_09607_)
  );
  AND2_X1 _11694_ (
    .A1(_07436_),
    .A2(_09607_),
    .ZN(_09618_)
  );
  INV_X1 _11695_ (
    .A(_09618_),
    .ZN(_09629_)
  );
  AND2_X1 _11696_ (
    .A1(_07414_),
    .A2(_09629_),
    .ZN(_09640_)
  );
  INV_X1 _11697_ (
    .A(_09640_),
    .ZN(_09651_)
  );
  AND2_X1 _11698_ (
    .A1(_07392_),
    .A2(_09618_),
    .ZN(_09662_)
  );
  INV_X1 _11699_ (
    .A(_09662_),
    .ZN(_09673_)
  );
  AND2_X1 _11700_ (
    .A1(_07392_),
    .A2(_09651_),
    .ZN(_09684_)
  );
  AND2_X1 _11701_ (
    .A1(_07414_),
    .A2(_09673_),
    .ZN(_09695_)
  );
  AND2_X1 _11702_ (
    .A1(_07359_),
    .A2(_09695_),
    .ZN(_09706_)
  );
  INV_X1 _11703_ (
    .A(_09706_),
    .ZN(_09717_)
  );
  AND2_X1 _11704_ (
    .A1(_07326_),
    .A2(_09717_),
    .ZN(_09728_)
  );
  INV_X1 _11705_ (
    .A(_09728_),
    .ZN(_09739_)
  );
  AND2_X1 _11706_ (
    .A1(_07304_),
    .A2(_09739_),
    .ZN(_09750_)
  );
  INV_X1 _11707_ (
    .A(_09750_),
    .ZN(_09760_)
  );
  AND2_X1 _11708_ (
    .A1(_07283_),
    .A2(_09728_),
    .ZN(_09771_)
  );
  INV_X1 _11709_ (
    .A(_09771_),
    .ZN(_09782_)
  );
  AND2_X1 _11710_ (
    .A1(_07283_),
    .A2(_09760_),
    .ZN(_09793_)
  );
  AND2_X1 _11711_ (
    .A1(_07304_),
    .A2(_09782_),
    .ZN(_09804_)
  );
  AND2_X1 _11712_ (
    .A1(_07250_),
    .A2(_09804_),
    .ZN(_09815_)
  );
  INV_X1 _11713_ (
    .A(_09815_),
    .ZN(_09826_)
  );
  AND2_X1 _11714_ (
    .A1(_07217_),
    .A2(_09826_),
    .ZN(_09837_)
  );
  INV_X1 _11715_ (
    .A(_09837_),
    .ZN(_09848_)
  );
  AND2_X1 _11716_ (
    .A1(_07195_),
    .A2(_09837_),
    .ZN(_09859_)
  );
  INV_X1 _11717_ (
    .A(_09859_),
    .ZN(_09870_)
  );
  AND2_X1 _11718_ (
    .A1(_07173_),
    .A2(_09848_),
    .ZN(_09881_)
  );
  INV_X1 _11719_ (
    .A(_09881_),
    .ZN(_09892_)
  );
  AND2_X1 _11720_ (
    .A1(_07173_),
    .A2(_09870_),
    .ZN(_09903_)
  );
  AND2_X1 _11721_ (
    .A1(_07195_),
    .A2(_09892_),
    .ZN(_09914_)
  );
  AND2_X1 _11722_ (
    .A1(_07140_),
    .A2(_09903_),
    .ZN(_09925_)
  );
  INV_X1 _11723_ (
    .A(_09925_),
    .ZN(_09936_)
  );
  AND2_X1 _11724_ (
    .A1(_07107_),
    .A2(_09936_),
    .ZN(_09947_)
  );
  INV_X1 _11725_ (
    .A(_09947_),
    .ZN(_09958_)
  );
  AND2_X1 _11726_ (
    .A1(_07085_),
    .A2(_09958_),
    .ZN(_09969_)
  );
  INV_X1 _11727_ (
    .A(_09969_),
    .ZN(_09980_)
  );
  AND2_X1 _11728_ (
    .A1(_07063_),
    .A2(_09947_),
    .ZN(_09991_)
  );
  INV_X1 _11729_ (
    .A(_09991_),
    .ZN(_10002_)
  );
  AND2_X1 _11730_ (
    .A1(_07063_),
    .A2(_09980_),
    .ZN(_10013_)
  );
  AND2_X1 _11731_ (
    .A1(_07085_),
    .A2(_10002_),
    .ZN(_10024_)
  );
  AND2_X1 _11732_ (
    .A1(_07030_),
    .A2(_10024_),
    .ZN(_10035_)
  );
  INV_X1 _11733_ (
    .A(_10035_),
    .ZN(_10046_)
  );
  AND2_X1 _11734_ (
    .A1(_06997_),
    .A2(_10046_),
    .ZN(_10057_)
  );
  INV_X1 _11735_ (
    .A(_10057_),
    .ZN(_10068_)
  );
  AND2_X1 _11736_ (
    .A1(_06976_),
    .A2(_10057_),
    .ZN(_10079_)
  );
  INV_X1 _11737_ (
    .A(_10079_),
    .ZN(_10090_)
  );
  AND2_X1 _11738_ (
    .A1(_06954_),
    .A2(_10068_),
    .ZN(_10100_)
  );
  INV_X1 _11739_ (
    .A(_10100_),
    .ZN(_10111_)
  );
  AND2_X1 _11740_ (
    .A1(_06954_),
    .A2(_10090_),
    .ZN(_10122_)
  );
  AND2_X1 _11741_ (
    .A1(_06976_),
    .A2(_10111_),
    .ZN(_10133_)
  );
  AND2_X1 _11742_ (
    .A1(_06921_),
    .A2(_10122_),
    .ZN(_10144_)
  );
  INV_X1 _11743_ (
    .A(_10144_),
    .ZN(_10155_)
  );
  AND2_X1 _11744_ (
    .A1(_06888_),
    .A2(_10155_),
    .ZN(_10166_)
  );
  INV_X1 _11745_ (
    .A(_10166_),
    .ZN(_10177_)
  );
  AND2_X1 _11746_ (
    .A1(_06866_),
    .A2(_10166_),
    .ZN(_10188_)
  );
  INV_X1 _11747_ (
    .A(_10188_),
    .ZN(_10199_)
  );
  AND2_X1 _11748_ (
    .A1(_06844_),
    .A2(_10177_),
    .ZN(_10210_)
  );
  INV_X1 _11749_ (
    .A(_10210_),
    .ZN(_10221_)
  );
  AND2_X1 _11750_ (
    .A1(_06844_),
    .A2(_10199_),
    .ZN(_10232_)
  );
  AND2_X1 _11751_ (
    .A1(_06866_),
    .A2(_10221_),
    .ZN(_10243_)
  );
  AND2_X1 _11752_ (
    .A1(_04415_),
    .A2(_05917_),
    .ZN(_10254_)
  );
  INV_X1 _11753_ (
    .A(_10254_),
    .ZN(_10265_)
  );
  AND2_X1 _11754_ (
    .A1(remainder[64]),
    .A2(_11217_[32]),
    .ZN(_10276_)
  );
  INV_X1 _11755_ (
    .A(_10276_),
    .ZN(_10287_)
  );
  AND2_X1 _11756_ (
    .A1(_04415_),
    .A2(_11217_[32]),
    .ZN(_10298_)
  );
  INV_X1 _11757_ (
    .A(_10298_),
    .ZN(_10309_)
  );
  AND2_X1 _11758_ (
    .A1(remainder[64]),
    .A2(_05917_),
    .ZN(_10320_)
  );
  INV_X1 _11759_ (
    .A(_10320_),
    .ZN(_10331_)
  );
  AND2_X1 _11760_ (
    .A1(_10265_),
    .A2(_10287_),
    .ZN(_10342_)
  );
  AND2_X1 _11761_ (
    .A1(_10309_),
    .A2(_10331_),
    .ZN(_10353_)
  );
  AND2_X1 _11762_ (
    .A1(_10232_),
    .A2(_10342_),
    .ZN(_10364_)
  );
  INV_X1 _11763_ (
    .A(_10364_),
    .ZN(_10375_)
  );
  AND2_X1 _11764_ (
    .A1(_10243_),
    .A2(_10353_),
    .ZN(_10385_)
  );
  INV_X1 _11765_ (
    .A(_10385_),
    .ZN(_10396_)
  );
  AND2_X1 _11766_ (
    .A1(_10243_),
    .A2(_10342_),
    .ZN(_10407_)
  );
  INV_X1 _11767_ (
    .A(_10407_),
    .ZN(_10418_)
  );
  AND2_X1 _11768_ (
    .A1(_10232_),
    .A2(_10353_),
    .ZN(_10429_)
  );
  INV_X1 _11769_ (
    .A(_10429_),
    .ZN(_10440_)
  );
  AND2_X1 _11770_ (
    .A1(_10375_),
    .A2(_10396_),
    .ZN(_10451_)
  );
  AND2_X1 _11771_ (
    .A1(_10418_),
    .A2(_10440_),
    .ZN(_10462_)
  );
  AND2_X1 _11772_ (
    .A1(_05983_),
    .A2(_10462_),
    .ZN(_10473_)
  );
  AND2_X1 _11773_ (
    .A1(_eOut_T_4),
    .A2(_06048_),
    .ZN(_10484_)
  );
  AND2_X1 _11774_ (
    .A1(_05950_),
    .A2(_10484_),
    .ZN(_10495_)
  );
  AND2_X1 _11775_ (
    .A1(_10473_),
    .A2(_10495_),
    .ZN(_10506_)
  );
  INV_X1 _11776_ (
    .A(_10506_),
    .ZN(_10517_)
  );
  AND2_X1 _11777_ (
    .A1(neg_out),
    .A2(_06201_),
    .ZN(_10528_)
  );
  AND2_X1 _11778_ (
    .A1(_10517_),
    .A2(_10528_),
    .ZN(_10539_)
  );
  INV_X1 _11779_ (
    .A(_10539_),
    .ZN(_10550_)
  );
  AND2_X1 _11780_ (
    .A1(io_req_bits_fn[0]),
    .A2(_05445_),
    .ZN(_10561_)
  );
  INV_X1 _11781_ (
    .A(_10561_),
    .ZN(_10572_)
  );
  AND2_X1 _11782_ (
    .A1(_05456_),
    .A2(_10572_),
    .ZN(_10583_)
  );
  INV_X1 _11783_ (
    .A(_10583_),
    .ZN(_10594_)
  );
  AND2_X1 _11784_ (
    .A1(_06746_),
    .A2(_10583_),
    .ZN(_10605_)
  );
  INV_X1 _11785_ (
    .A(_10605_),
    .ZN(_10616_)
  );
  AND2_X1 _11786_ (
    .A1(_06702_),
    .A2(_10605_),
    .ZN(_10627_)
  );
  INV_X1 _11787_ (
    .A(_10627_),
    .ZN(_10638_)
  );
  AND2_X1 _11788_ (
    .A1(_06713_),
    .A2(_10616_),
    .ZN(_10649_)
  );
  INV_X1 _11789_ (
    .A(_10649_),
    .ZN(_10660_)
  );
  AND2_X1 _11790_ (
    .A1(_10638_),
    .A2(_10660_),
    .ZN(_10670_)
  );
  AND2_X1 _11791_ (
    .A1(_06190_),
    .A2(_10670_),
    .ZN(_10681_)
  );
  INV_X1 _11792_ (
    .A(_10681_),
    .ZN(_10692_)
  );
  AND2_X1 _11793_ (
    .A1(_10550_),
    .A2(_10692_),
    .ZN(_10703_)
  );
  INV_X1 _11794_ (
    .A(_10703_),
    .ZN(_00008_)
  );
  MUX2_X1 _11795_ (
    .A(req_tag[0]),
    .B(io_req_bits_tag[0]),
    .S(_06190_),
    .Z(_00009_)
  );
  MUX2_X1 _11796_ (
    .A(req_tag[1]),
    .B(io_req_bits_tag[1]),
    .S(_06190_),
    .Z(_00010_)
  );
  MUX2_X1 _11797_ (
    .A(req_tag[2]),
    .B(io_req_bits_tag[2]),
    .S(_06190_),
    .Z(_00011_)
  );
  MUX2_X1 _11798_ (
    .A(req_tag[3]),
    .B(io_req_bits_tag[3]),
    .S(_06190_),
    .Z(_00012_)
  );
  MUX2_X1 _11799_ (
    .A(req_tag[4]),
    .B(io_req_bits_tag[4]),
    .S(_06190_),
    .Z(_00013_)
  );
  AND2_X1 _11800_ (
    .A1(_05994_),
    .A2(_06114_),
    .ZN(_10774_)
  );
  INV_X1 _11801_ (
    .A(_10774_),
    .ZN(_10785_)
  );
  MUX2_X1 _11802_ (
    .A(_count_T_1[0]),
    .B(count[0]),
    .S(_10774_),
    .Z(_10796_)
  );
  AND2_X1 _11803_ (
    .A1(_06201_),
    .A2(_10796_),
    .ZN(_00014_)
  );
  AND2_X1 _11804_ (
    .A1(count[0]),
    .A2(_10785_),
    .ZN(_10817_)
  );
  INV_X1 _11805_ (
    .A(_10817_),
    .ZN(_10828_)
  );
  AND2_X1 _11806_ (
    .A1(count[1]),
    .A2(_10817_),
    .ZN(_10839_)
  );
  INV_X1 _11807_ (
    .A(_10839_),
    .ZN(_10850_)
  );
  AND2_X1 _11808_ (
    .A1(_04820_),
    .A2(_10828_),
    .ZN(_10861_)
  );
  INV_X1 _11809_ (
    .A(_10861_),
    .ZN(_10872_)
  );
  AND2_X1 _11810_ (
    .A1(_06201_),
    .A2(_10872_),
    .ZN(_10883_)
  );
  AND2_X1 _11811_ (
    .A1(_10850_),
    .A2(_10883_),
    .ZN(_00015_)
  );
  AND2_X1 _11812_ (
    .A1(count[2]),
    .A2(_10839_),
    .ZN(_10904_)
  );
  INV_X1 _11813_ (
    .A(_10904_),
    .ZN(_10915_)
  );
  AND2_X1 _11814_ (
    .A1(_04810_),
    .A2(_10850_),
    .ZN(_10926_)
  );
  INV_X1 _11815_ (
    .A(_10926_),
    .ZN(_10937_)
  );
  AND2_X1 _11816_ (
    .A1(_06201_),
    .A2(_10937_),
    .ZN(_10948_)
  );
  AND2_X1 _11817_ (
    .A1(_10915_),
    .A2(_10948_),
    .ZN(_00016_)
  );
  AND2_X1 _11818_ (
    .A1(count[3]),
    .A2(_10904_),
    .ZN(_10968_)
  );
  INV_X1 _11819_ (
    .A(_10968_),
    .ZN(_10979_)
  );
  AND2_X1 _11820_ (
    .A1(_04799_),
    .A2(_10915_),
    .ZN(_10990_)
  );
  INV_X1 _11821_ (
    .A(_10990_),
    .ZN(_11001_)
  );
  AND2_X1 _11822_ (
    .A1(_06201_),
    .A2(_11001_),
    .ZN(_11012_)
  );
  AND2_X1 _11823_ (
    .A1(_10979_),
    .A2(_11012_),
    .ZN(_00017_)
  );
  AND2_X1 _11824_ (
    .A1(count[4]),
    .A2(_10968_),
    .ZN(_11033_)
  );
  INV_X1 _11825_ (
    .A(_11033_),
    .ZN(_11044_)
  );
  AND2_X1 _11826_ (
    .A1(_04788_),
    .A2(_10979_),
    .ZN(_11055_)
  );
  INV_X1 _11827_ (
    .A(_11055_),
    .ZN(_11066_)
  );
  AND2_X1 _11828_ (
    .A1(_06201_),
    .A2(_11066_),
    .ZN(_11077_)
  );
  AND2_X1 _11829_ (
    .A1(_11044_),
    .A2(_11077_),
    .ZN(_00018_)
  );
  AND2_X1 _11830_ (
    .A1(count[5]),
    .A2(_11033_),
    .ZN(_11098_)
  );
  INV_X1 _11831_ (
    .A(_11098_),
    .ZN(_11109_)
  );
  AND2_X1 _11832_ (
    .A1(_04777_),
    .A2(_11044_),
    .ZN(_11120_)
  );
  INV_X1 _11833_ (
    .A(_11120_),
    .ZN(_11131_)
  );
  AND2_X1 _11834_ (
    .A1(_11109_),
    .A2(_11131_),
    .ZN(_00121_)
  );
  AND2_X1 _11835_ (
    .A1(_06201_),
    .A2(_00121_),
    .ZN(_00019_)
  );
  AND2_X1 _11836_ (
    .A1(divisor[31]),
    .A2(_06299_),
    .ZN(_00142_)
  );
  INV_X1 _11837_ (
    .A(_00142_),
    .ZN(_00153_)
  );
  AND2_X1 _11838_ (
    .A1(_06201_),
    .A2(_00153_),
    .ZN(_00164_)
  );
  AND2_X1 _11839_ (
    .A1(divisor[0]),
    .A2(_00164_),
    .ZN(_00175_)
  );
  INV_X1 _11840_ (
    .A(_00175_),
    .ZN(_00186_)
  );
  AND2_X1 _11841_ (
    .A1(io_req_bits_in2[0]),
    .A2(_06190_),
    .ZN(_00197_)
  );
  INV_X1 _11842_ (
    .A(_00197_),
    .ZN(_00208_)
  );
  AND2_X1 _11843_ (
    .A1(remainder[32]),
    .A2(_11217_[0]),
    .ZN(_00219_)
  );
  INV_X1 _11844_ (
    .A(_00219_),
    .ZN(_00229_)
  );
  AND2_X1 _11845_ (
    .A1(_08445_),
    .A2(_00229_),
    .ZN(_00240_)
  );
  INV_X1 _11846_ (
    .A(_00240_),
    .ZN(_00251_)
  );
  AND2_X1 _11847_ (
    .A1(_06201_),
    .A2(_00142_),
    .ZN(_00262_)
  );
  AND2_X1 _11848_ (
    .A1(_00251_),
    .A2(_00262_),
    .ZN(_00273_)
  );
  INV_X1 _11849_ (
    .A(_00273_),
    .ZN(_00284_)
  );
  AND2_X1 _11850_ (
    .A1(_00186_),
    .A2(_00284_),
    .ZN(_00295_)
  );
  AND2_X1 _11851_ (
    .A1(_00208_),
    .A2(_00295_),
    .ZN(_00306_)
  );
  INV_X1 _11852_ (
    .A(_00306_),
    .ZN(_00020_)
  );
  AND2_X1 _11853_ (
    .A1(divisor[1]),
    .A2(_00164_),
    .ZN(_00327_)
  );
  INV_X1 _11854_ (
    .A(_00327_),
    .ZN(_00338_)
  );
  AND2_X1 _11855_ (
    .A1(io_req_bits_in2[1]),
    .A2(_06190_),
    .ZN(_00349_)
  );
  INV_X1 _11856_ (
    .A(_00349_),
    .ZN(_00360_)
  );
  AND2_X1 _11857_ (
    .A1(_08434_),
    .A2(_08489_),
    .ZN(_00371_)
  );
  INV_X1 _11858_ (
    .A(_00371_),
    .ZN(_00382_)
  );
  AND2_X1 _11859_ (
    .A1(_08510_),
    .A2(_00382_),
    .ZN(_00393_)
  );
  INV_X1 _11860_ (
    .A(_00393_),
    .ZN(_00404_)
  );
  AND2_X1 _11861_ (
    .A1(_00262_),
    .A2(_00393_),
    .ZN(_00415_)
  );
  INV_X1 _11862_ (
    .A(_00415_),
    .ZN(_00426_)
  );
  AND2_X1 _11863_ (
    .A1(_00338_),
    .A2(_00426_),
    .ZN(_00437_)
  );
  AND2_X1 _11864_ (
    .A1(_00360_),
    .A2(_00437_),
    .ZN(_00448_)
  );
  INV_X1 _11865_ (
    .A(_00448_),
    .ZN(_00021_)
  );
  AND2_X1 _11866_ (
    .A1(_08521_),
    .A2(_08576_),
    .ZN(_00469_)
  );
  INV_X1 _11867_ (
    .A(_00469_),
    .ZN(_00480_)
  );
  AND2_X1 _11868_ (
    .A1(_08598_),
    .A2(_00480_),
    .ZN(_00491_)
  );
  INV_X1 _11869_ (
    .A(_00491_),
    .ZN(_00502_)
  );
  AND2_X1 _11870_ (
    .A1(_00262_),
    .A2(_00491_),
    .ZN(_00513_)
  );
  INV_X1 _11871_ (
    .A(_00513_),
    .ZN(_00523_)
  );
  AND2_X1 _11872_ (
    .A1(io_req_bits_in2[2]),
    .A2(_06190_),
    .ZN(_00534_)
  );
  INV_X1 _11873_ (
    .A(_00534_),
    .ZN(_00545_)
  );
  AND2_X1 _11874_ (
    .A1(divisor[2]),
    .A2(_00164_),
    .ZN(_00556_)
  );
  INV_X1 _11875_ (
    .A(_00556_),
    .ZN(_00567_)
  );
  AND2_X1 _11876_ (
    .A1(_00545_),
    .A2(_00567_),
    .ZN(_00578_)
  );
  AND2_X1 _11877_ (
    .A1(_00523_),
    .A2(_00578_),
    .ZN(_00589_)
  );
  INV_X1 _11878_ (
    .A(_00589_),
    .ZN(_00022_)
  );
  AND2_X1 _11879_ (
    .A1(_08357_),
    .A2(_08379_),
    .ZN(_00610_)
  );
  INV_X1 _11880_ (
    .A(_00610_),
    .ZN(_00621_)
  );
  AND2_X1 _11881_ (
    .A1(_08609_),
    .A2(_00621_),
    .ZN(_00632_)
  );
  INV_X1 _11882_ (
    .A(_00632_),
    .ZN(_00643_)
  );
  AND2_X1 _11883_ (
    .A1(_08620_),
    .A2(_00610_),
    .ZN(_00654_)
  );
  INV_X1 _11884_ (
    .A(_00654_),
    .ZN(_00665_)
  );
  AND2_X1 _11885_ (
    .A1(_08609_),
    .A2(_00610_),
    .ZN(_00676_)
  );
  INV_X1 _11886_ (
    .A(_00676_),
    .ZN(_00687_)
  );
  AND2_X1 _11887_ (
    .A1(_08620_),
    .A2(_00621_),
    .ZN(_00698_)
  );
  INV_X1 _11888_ (
    .A(_00698_),
    .ZN(_00709_)
  );
  AND2_X1 _11889_ (
    .A1(_00643_),
    .A2(_00665_),
    .ZN(_00720_)
  );
  AND2_X1 _11890_ (
    .A1(_00687_),
    .A2(_00709_),
    .ZN(_00731_)
  );
  AND2_X1 _11891_ (
    .A1(_00262_),
    .A2(_00720_),
    .ZN(_00742_)
  );
  INV_X1 _11892_ (
    .A(_00742_),
    .ZN(_00753_)
  );
  AND2_X1 _11893_ (
    .A1(io_req_bits_in2[3]),
    .A2(_06190_),
    .ZN(_00764_)
  );
  INV_X1 _11894_ (
    .A(_00764_),
    .ZN(_00775_)
  );
  AND2_X1 _11895_ (
    .A1(divisor[3]),
    .A2(_00164_),
    .ZN(_00786_)
  );
  INV_X1 _11896_ (
    .A(_00786_),
    .ZN(_00797_)
  );
  AND2_X1 _11897_ (
    .A1(_00775_),
    .A2(_00797_),
    .ZN(_00808_)
  );
  AND2_X1 _11898_ (
    .A1(_00753_),
    .A2(_00808_),
    .ZN(_00819_)
  );
  INV_X1 _11899_ (
    .A(_00819_),
    .ZN(_00023_)
  );
  AND2_X1 _11900_ (
    .A1(_08335_),
    .A2(_08675_),
    .ZN(_00840_)
  );
  INV_X1 _11901_ (
    .A(_00840_),
    .ZN(_00851_)
  );
  AND2_X1 _11902_ (
    .A1(_08708_),
    .A2(_00851_),
    .ZN(_00862_)
  );
  INV_X1 _11903_ (
    .A(_00862_),
    .ZN(_00873_)
  );
  AND2_X1 _11904_ (
    .A1(_00262_),
    .A2(_00862_),
    .ZN(_00884_)
  );
  INV_X1 _11905_ (
    .A(_00884_),
    .ZN(_00895_)
  );
  AND2_X1 _11906_ (
    .A1(divisor[4]),
    .A2(_00164_),
    .ZN(_00905_)
  );
  INV_X1 _11907_ (
    .A(_00905_),
    .ZN(_00915_)
  );
  AND2_X1 _11908_ (
    .A1(io_req_bits_in2[4]),
    .A2(_06190_),
    .ZN(_00925_)
  );
  INV_X1 _11909_ (
    .A(_00925_),
    .ZN(_00935_)
  );
  AND2_X1 _11910_ (
    .A1(_00915_),
    .A2(_00935_),
    .ZN(_00945_)
  );
  AND2_X1 _11911_ (
    .A1(_00895_),
    .A2(_00945_),
    .ZN(_00955_)
  );
  INV_X1 _11912_ (
    .A(_00955_),
    .ZN(_00024_)
  );
  AND2_X1 _11913_ (
    .A1(_08719_),
    .A2(_08774_),
    .ZN(_00974_)
  );
  INV_X1 _11914_ (
    .A(_00974_),
    .ZN(_00985_)
  );
  AND2_X1 _11915_ (
    .A1(_08796_),
    .A2(_00985_),
    .ZN(_00994_)
  );
  INV_X1 _11916_ (
    .A(_00994_),
    .ZN(_01005_)
  );
  AND2_X1 _11917_ (
    .A1(_00262_),
    .A2(_00994_),
    .ZN(_01015_)
  );
  INV_X1 _11918_ (
    .A(_01015_),
    .ZN(_01025_)
  );
  AND2_X1 _11919_ (
    .A1(io_req_bits_in2[5]),
    .A2(_06190_),
    .ZN(_01035_)
  );
  INV_X1 _11920_ (
    .A(_01035_),
    .ZN(_01045_)
  );
  AND2_X1 _11921_ (
    .A1(divisor[5]),
    .A2(_00164_),
    .ZN(_01056_)
  );
  INV_X1 _11922_ (
    .A(_01056_),
    .ZN(_01065_)
  );
  AND2_X1 _11923_ (
    .A1(_01045_),
    .A2(_01065_),
    .ZN(_01076_)
  );
  AND2_X1 _11924_ (
    .A1(_01025_),
    .A2(_01076_),
    .ZN(_01086_)
  );
  INV_X1 _11925_ (
    .A(_01086_),
    .ZN(_00025_)
  );
  AND2_X1 _11926_ (
    .A1(_08247_),
    .A2(_08807_),
    .ZN(_01106_)
  );
  INV_X1 _11927_ (
    .A(_01106_),
    .ZN(_01115_)
  );
  AND2_X1 _11928_ (
    .A1(_08839_),
    .A2(_01115_),
    .ZN(_01126_)
  );
  INV_X1 _11929_ (
    .A(_01126_),
    .ZN(_01136_)
  );
  AND2_X1 _11930_ (
    .A1(_00262_),
    .A2(_01126_),
    .ZN(_01146_)
  );
  INV_X1 _11931_ (
    .A(_01146_),
    .ZN(_01157_)
  );
  AND2_X1 _11932_ (
    .A1(io_req_bits_in2[6]),
    .A2(_06190_),
    .ZN(_01166_)
  );
  INV_X1 _11933_ (
    .A(_01166_),
    .ZN(_01177_)
  );
  AND2_X1 _11934_ (
    .A1(divisor[6]),
    .A2(_00164_),
    .ZN(_01188_)
  );
  INV_X1 _11935_ (
    .A(_01188_),
    .ZN(_01197_)
  );
  AND2_X1 _11936_ (
    .A1(_01177_),
    .A2(_01197_),
    .ZN(_01208_)
  );
  AND2_X1 _11937_ (
    .A1(_01157_),
    .A2(_01208_),
    .ZN(_01218_)
  );
  INV_X1 _11938_ (
    .A(_01218_),
    .ZN(_00026_)
  );
  AND2_X1 _11939_ (
    .A1(_08160_),
    .A2(_08182_),
    .ZN(_01238_)
  );
  INV_X1 _11940_ (
    .A(_01238_),
    .ZN(_01247_)
  );
  AND2_X1 _11941_ (
    .A1(_08861_),
    .A2(_01247_),
    .ZN(_01258_)
  );
  INV_X1 _11942_ (
    .A(_01258_),
    .ZN(_01268_)
  );
  AND2_X1 _11943_ (
    .A1(_08850_),
    .A2(_01238_),
    .ZN(_01278_)
  );
  INV_X1 _11944_ (
    .A(_01278_),
    .ZN(_01289_)
  );
  AND2_X1 _11945_ (
    .A1(_01268_),
    .A2(_01289_),
    .ZN(_01298_)
  );
  INV_X1 _11946_ (
    .A(_01298_),
    .ZN(_01309_)
  );
  AND2_X1 _11947_ (
    .A1(_00262_),
    .A2(_01309_),
    .ZN(_01320_)
  );
  INV_X1 _11948_ (
    .A(_01320_),
    .ZN(_01329_)
  );
  AND2_X1 _11949_ (
    .A1(io_req_bits_in2[7]),
    .A2(_06190_),
    .ZN(_01340_)
  );
  INV_X1 _11950_ (
    .A(_01340_),
    .ZN(_01350_)
  );
  AND2_X1 _11951_ (
    .A1(divisor[7]),
    .A2(_00164_),
    .ZN(_01360_)
  );
  INV_X1 _11952_ (
    .A(_01360_),
    .ZN(_01371_)
  );
  AND2_X1 _11953_ (
    .A1(_01350_),
    .A2(_01371_),
    .ZN(_01380_)
  );
  AND2_X1 _11954_ (
    .A1(_01329_),
    .A2(_01380_),
    .ZN(_01391_)
  );
  INV_X1 _11955_ (
    .A(_01391_),
    .ZN(_00027_)
  );
  AND2_X1 _11956_ (
    .A1(_08138_),
    .A2(_08916_),
    .ZN(_01410_)
  );
  INV_X1 _11957_ (
    .A(_01410_),
    .ZN(_01421_)
  );
  AND2_X1 _11958_ (
    .A1(_08949_),
    .A2(_01421_),
    .ZN(_01430_)
  );
  INV_X1 _11959_ (
    .A(_01430_),
    .ZN(_01441_)
  );
  AND2_X1 _11960_ (
    .A1(_00262_),
    .A2(_01430_),
    .ZN(_01452_)
  );
  INV_X1 _11961_ (
    .A(_01452_),
    .ZN(_01461_)
  );
  AND2_X1 _11962_ (
    .A1(divisor[8]),
    .A2(_00164_),
    .ZN(_01472_)
  );
  INV_X1 _11963_ (
    .A(_01472_),
    .ZN(_01482_)
  );
  AND2_X1 _11964_ (
    .A1(io_req_bits_in2[8]),
    .A2(_06190_),
    .ZN(_01492_)
  );
  INV_X1 _11965_ (
    .A(_01492_),
    .ZN(_01503_)
  );
  AND2_X1 _11966_ (
    .A1(_01482_),
    .A2(_01503_),
    .ZN(_01512_)
  );
  AND2_X1 _11967_ (
    .A1(_01461_),
    .A2(_01512_),
    .ZN(_01523_)
  );
  INV_X1 _11968_ (
    .A(_01523_),
    .ZN(_00028_)
  );
  AND2_X1 _11969_ (
    .A1(_08050_),
    .A2(_08072_),
    .ZN(_01542_)
  );
  INV_X1 _11970_ (
    .A(_01542_),
    .ZN(_01553_)
  );
  AND2_X1 _11971_ (
    .A1(_08971_),
    .A2(_01553_),
    .ZN(_01564_)
  );
  INV_X1 _11972_ (
    .A(_01564_),
    .ZN(_01573_)
  );
  AND2_X1 _11973_ (
    .A1(_08960_),
    .A2(_01542_),
    .ZN(_01584_)
  );
  INV_X1 _11974_ (
    .A(_01584_),
    .ZN(_01595_)
  );
  AND2_X1 _11975_ (
    .A1(_01573_),
    .A2(_01595_),
    .ZN(_01604_)
  );
  INV_X1 _11976_ (
    .A(_01604_),
    .ZN(_01615_)
  );
  AND2_X1 _11977_ (
    .A1(_00262_),
    .A2(_01615_),
    .ZN(_01626_)
  );
  INV_X1 _11978_ (
    .A(_01626_),
    .ZN(_01635_)
  );
  AND2_X1 _11979_ (
    .A1(io_req_bits_in2[9]),
    .A2(_06190_),
    .ZN(_01646_)
  );
  INV_X1 _11980_ (
    .A(_01646_),
    .ZN(_01657_)
  );
  AND2_X1 _11981_ (
    .A1(divisor[9]),
    .A2(_00164_),
    .ZN(_01666_)
  );
  INV_X1 _11982_ (
    .A(_01666_),
    .ZN(_01677_)
  );
  AND2_X1 _11983_ (
    .A1(_01657_),
    .A2(_01677_),
    .ZN(_01688_)
  );
  AND2_X1 _11984_ (
    .A1(_01635_),
    .A2(_01688_),
    .ZN(_01697_)
  );
  INV_X1 _11985_ (
    .A(_01697_),
    .ZN(_00029_)
  );
  AND2_X1 _11986_ (
    .A1(_08028_),
    .A2(_09026_),
    .ZN(_01718_)
  );
  INV_X1 _11987_ (
    .A(_01718_),
    .ZN(_01727_)
  );
  AND2_X1 _11988_ (
    .A1(_09059_),
    .A2(_01727_),
    .ZN(_01738_)
  );
  INV_X1 _11989_ (
    .A(_01738_),
    .ZN(_01748_)
  );
  AND2_X1 _11990_ (
    .A1(_00262_),
    .A2(_01738_),
    .ZN(_01752_)
  );
  INV_X1 _11991_ (
    .A(_01752_),
    .ZN(_01753_)
  );
  AND2_X1 _11992_ (
    .A1(io_req_bits_in2[10]),
    .A2(_06190_),
    .ZN(_01754_)
  );
  INV_X1 _11993_ (
    .A(_01754_),
    .ZN(_01755_)
  );
  AND2_X1 _11994_ (
    .A1(divisor[10]),
    .A2(_00164_),
    .ZN(_01756_)
  );
  INV_X1 _11995_ (
    .A(_01756_),
    .ZN(_01757_)
  );
  AND2_X1 _11996_ (
    .A1(_01755_),
    .A2(_01757_),
    .ZN(_01758_)
  );
  AND2_X1 _11997_ (
    .A1(_01753_),
    .A2(_01758_),
    .ZN(_01759_)
  );
  INV_X1 _11998_ (
    .A(_01759_),
    .ZN(_00030_)
  );
  AND2_X1 _11999_ (
    .A1(_07940_),
    .A2(_07962_),
    .ZN(_01760_)
  );
  INV_X1 _12000_ (
    .A(_01760_),
    .ZN(_01761_)
  );
  AND2_X1 _12001_ (
    .A1(_09081_),
    .A2(_01761_),
    .ZN(_01762_)
  );
  INV_X1 _12002_ (
    .A(_01762_),
    .ZN(_01763_)
  );
  AND2_X1 _12003_ (
    .A1(_09070_),
    .A2(_01760_),
    .ZN(_01764_)
  );
  INV_X1 _12004_ (
    .A(_01764_),
    .ZN(_01765_)
  );
  AND2_X1 _12005_ (
    .A1(_09070_),
    .A2(_01761_),
    .ZN(_01766_)
  );
  INV_X1 _12006_ (
    .A(_01766_),
    .ZN(_01767_)
  );
  AND2_X1 _12007_ (
    .A1(_09081_),
    .A2(_01760_),
    .ZN(_01768_)
  );
  INV_X1 _12008_ (
    .A(_01768_),
    .ZN(_01769_)
  );
  AND2_X1 _12009_ (
    .A1(_01763_),
    .A2(_01765_),
    .ZN(_01770_)
  );
  AND2_X1 _12010_ (
    .A1(_01767_),
    .A2(_01769_),
    .ZN(_01771_)
  );
  AND2_X1 _12011_ (
    .A1(_00262_),
    .A2(_01771_),
    .ZN(_01772_)
  );
  INV_X1 _12012_ (
    .A(_01772_),
    .ZN(_01773_)
  );
  AND2_X1 _12013_ (
    .A1(io_req_bits_in2[11]),
    .A2(_06190_),
    .ZN(_01774_)
  );
  INV_X1 _12014_ (
    .A(_01774_),
    .ZN(_01775_)
  );
  AND2_X1 _12015_ (
    .A1(divisor[11]),
    .A2(_00164_),
    .ZN(_01776_)
  );
  INV_X1 _12016_ (
    .A(_01776_),
    .ZN(_01777_)
  );
  AND2_X1 _12017_ (
    .A1(_01775_),
    .A2(_01777_),
    .ZN(_01778_)
  );
  AND2_X1 _12018_ (
    .A1(_01773_),
    .A2(_01778_),
    .ZN(_01779_)
  );
  INV_X1 _12019_ (
    .A(_01779_),
    .ZN(_00031_)
  );
  AND2_X1 _12020_ (
    .A1(_07918_),
    .A2(_09135_),
    .ZN(_01780_)
  );
  INV_X1 _12021_ (
    .A(_01780_),
    .ZN(_01781_)
  );
  AND2_X1 _12022_ (
    .A1(_09168_),
    .A2(_01781_),
    .ZN(_01782_)
  );
  INV_X1 _12023_ (
    .A(_01782_),
    .ZN(_01783_)
  );
  AND2_X1 _12024_ (
    .A1(_00262_),
    .A2(_01782_),
    .ZN(_01784_)
  );
  INV_X1 _12025_ (
    .A(_01784_),
    .ZN(_01785_)
  );
  AND2_X1 _12026_ (
    .A1(divisor[12]),
    .A2(_00164_),
    .ZN(_01786_)
  );
  INV_X1 _12027_ (
    .A(_01786_),
    .ZN(_01787_)
  );
  AND2_X1 _12028_ (
    .A1(io_req_bits_in2[12]),
    .A2(_06190_),
    .ZN(_01788_)
  );
  INV_X1 _12029_ (
    .A(_01788_),
    .ZN(_01789_)
  );
  AND2_X1 _12030_ (
    .A1(_01787_),
    .A2(_01789_),
    .ZN(_01790_)
  );
  AND2_X1 _12031_ (
    .A1(_01785_),
    .A2(_01790_),
    .ZN(_01791_)
  );
  INV_X1 _12032_ (
    .A(_01791_),
    .ZN(_00032_)
  );
  AND2_X1 _12033_ (
    .A1(_07831_),
    .A2(_07853_),
    .ZN(_01792_)
  );
  INV_X1 _12034_ (
    .A(_01792_),
    .ZN(_01793_)
  );
  AND2_X1 _12035_ (
    .A1(_09190_),
    .A2(_01793_),
    .ZN(_01794_)
  );
  INV_X1 _12036_ (
    .A(_01794_),
    .ZN(_01795_)
  );
  AND2_X1 _12037_ (
    .A1(_09179_),
    .A2(_01792_),
    .ZN(_01796_)
  );
  INV_X1 _12038_ (
    .A(_01796_),
    .ZN(_01797_)
  );
  AND2_X1 _12039_ (
    .A1(_09179_),
    .A2(_01793_),
    .ZN(_01798_)
  );
  INV_X1 _12040_ (
    .A(_01798_),
    .ZN(_01799_)
  );
  AND2_X1 _12041_ (
    .A1(_09190_),
    .A2(_01792_),
    .ZN(_01800_)
  );
  INV_X1 _12042_ (
    .A(_01800_),
    .ZN(_01801_)
  );
  AND2_X1 _12043_ (
    .A1(_01795_),
    .A2(_01797_),
    .ZN(_01802_)
  );
  AND2_X1 _12044_ (
    .A1(_01799_),
    .A2(_01801_),
    .ZN(_01803_)
  );
  AND2_X1 _12045_ (
    .A1(_00262_),
    .A2(_01803_),
    .ZN(_01804_)
  );
  INV_X1 _12046_ (
    .A(_01804_),
    .ZN(_01805_)
  );
  AND2_X1 _12047_ (
    .A1(divisor[13]),
    .A2(_00164_),
    .ZN(_01806_)
  );
  INV_X1 _12048_ (
    .A(_01806_),
    .ZN(_01807_)
  );
  AND2_X1 _12049_ (
    .A1(io_req_bits_in2[13]),
    .A2(_06190_),
    .ZN(_01808_)
  );
  INV_X1 _12050_ (
    .A(_01808_),
    .ZN(_01809_)
  );
  AND2_X1 _12051_ (
    .A1(_01807_),
    .A2(_01809_),
    .ZN(_01810_)
  );
  AND2_X1 _12052_ (
    .A1(_01805_),
    .A2(_01810_),
    .ZN(_01811_)
  );
  INV_X1 _12053_ (
    .A(_01811_),
    .ZN(_00033_)
  );
  AND2_X1 _12054_ (
    .A1(_07809_),
    .A2(_09245_),
    .ZN(_01812_)
  );
  INV_X1 _12055_ (
    .A(_01812_),
    .ZN(_01813_)
  );
  AND2_X1 _12056_ (
    .A1(_09278_),
    .A2(_01813_),
    .ZN(_01814_)
  );
  INV_X1 _12057_ (
    .A(_01814_),
    .ZN(_01815_)
  );
  AND2_X1 _12058_ (
    .A1(_00262_),
    .A2(_01814_),
    .ZN(_01816_)
  );
  INV_X1 _12059_ (
    .A(_01816_),
    .ZN(_01817_)
  );
  AND2_X1 _12060_ (
    .A1(io_req_bits_in2[14]),
    .A2(_06190_),
    .ZN(_01818_)
  );
  INV_X1 _12061_ (
    .A(_01818_),
    .ZN(_01819_)
  );
  AND2_X1 _12062_ (
    .A1(divisor[14]),
    .A2(_00164_),
    .ZN(_01820_)
  );
  INV_X1 _12063_ (
    .A(_01820_),
    .ZN(_01821_)
  );
  AND2_X1 _12064_ (
    .A1(_01819_),
    .A2(_01821_),
    .ZN(_01822_)
  );
  AND2_X1 _12065_ (
    .A1(_01817_),
    .A2(_01822_),
    .ZN(_01823_)
  );
  INV_X1 _12066_ (
    .A(_01823_),
    .ZN(_00034_)
  );
  AND2_X1 _12067_ (
    .A1(_07721_),
    .A2(_07743_),
    .ZN(_01824_)
  );
  INV_X1 _12068_ (
    .A(_01824_),
    .ZN(_01825_)
  );
  AND2_X1 _12069_ (
    .A1(_09300_),
    .A2(_01825_),
    .ZN(_01826_)
  );
  INV_X1 _12070_ (
    .A(_01826_),
    .ZN(_01827_)
  );
  AND2_X1 _12071_ (
    .A1(_09289_),
    .A2(_01824_),
    .ZN(_01828_)
  );
  INV_X1 _12072_ (
    .A(_01828_),
    .ZN(_01829_)
  );
  AND2_X1 _12073_ (
    .A1(_09289_),
    .A2(_01825_),
    .ZN(_01830_)
  );
  INV_X1 _12074_ (
    .A(_01830_),
    .ZN(_01831_)
  );
  AND2_X1 _12075_ (
    .A1(_09300_),
    .A2(_01824_),
    .ZN(_01832_)
  );
  INV_X1 _12076_ (
    .A(_01832_),
    .ZN(_01833_)
  );
  AND2_X1 _12077_ (
    .A1(_01827_),
    .A2(_01829_),
    .ZN(_01834_)
  );
  AND2_X1 _12078_ (
    .A1(_01831_),
    .A2(_01833_),
    .ZN(_01835_)
  );
  AND2_X1 _12079_ (
    .A1(_00262_),
    .A2(_01835_),
    .ZN(_01836_)
  );
  INV_X1 _12080_ (
    .A(_01836_),
    .ZN(_01837_)
  );
  AND2_X1 _12081_ (
    .A1(divisor[15]),
    .A2(_00164_),
    .ZN(_01838_)
  );
  INV_X1 _12082_ (
    .A(_01838_),
    .ZN(_01839_)
  );
  AND2_X1 _12083_ (
    .A1(io_req_bits_in2[15]),
    .A2(_06190_),
    .ZN(_01840_)
  );
  INV_X1 _12084_ (
    .A(_01840_),
    .ZN(_01841_)
  );
  AND2_X1 _12085_ (
    .A1(_01839_),
    .A2(_01841_),
    .ZN(_01842_)
  );
  AND2_X1 _12086_ (
    .A1(_01837_),
    .A2(_01842_),
    .ZN(_01843_)
  );
  INV_X1 _12087_ (
    .A(_01843_),
    .ZN(_00035_)
  );
  AND2_X1 _12088_ (
    .A1(_07699_),
    .A2(_09355_),
    .ZN(_01844_)
  );
  INV_X1 _12089_ (
    .A(_01844_),
    .ZN(_01845_)
  );
  AND2_X1 _12090_ (
    .A1(_09388_),
    .A2(_01845_),
    .ZN(_01846_)
  );
  INV_X1 _12091_ (
    .A(_01846_),
    .ZN(_01847_)
  );
  AND2_X1 _12092_ (
    .A1(_00262_),
    .A2(_01846_),
    .ZN(_01848_)
  );
  INV_X1 _12093_ (
    .A(_01848_),
    .ZN(_01849_)
  );
  AND2_X1 _12094_ (
    .A1(io_req_bits_in2[16]),
    .A2(_06190_),
    .ZN(_01850_)
  );
  INV_X1 _12095_ (
    .A(_01850_),
    .ZN(_01851_)
  );
  AND2_X1 _12096_ (
    .A1(divisor[16]),
    .A2(_00164_),
    .ZN(_01852_)
  );
  INV_X1 _12097_ (
    .A(_01852_),
    .ZN(_01853_)
  );
  AND2_X1 _12098_ (
    .A1(_01851_),
    .A2(_01853_),
    .ZN(_01854_)
  );
  AND2_X1 _12099_ (
    .A1(_01849_),
    .A2(_01854_),
    .ZN(_01855_)
  );
  INV_X1 _12100_ (
    .A(_01855_),
    .ZN(_00036_)
  );
  AND2_X1 _12101_ (
    .A1(_07611_),
    .A2(_07633_),
    .ZN(_01856_)
  );
  INV_X1 _12102_ (
    .A(_01856_),
    .ZN(_01857_)
  );
  AND2_X1 _12103_ (
    .A1(_09399_),
    .A2(_01857_),
    .ZN(_01858_)
  );
  INV_X1 _12104_ (
    .A(_01858_),
    .ZN(_01859_)
  );
  AND2_X1 _12105_ (
    .A1(_09410_),
    .A2(_01856_),
    .ZN(_01860_)
  );
  INV_X1 _12106_ (
    .A(_01860_),
    .ZN(_01861_)
  );
  AND2_X1 _12107_ (
    .A1(_01859_),
    .A2(_01861_),
    .ZN(_01862_)
  );
  AND2_X1 _12108_ (
    .A1(_00262_),
    .A2(_01862_),
    .ZN(_01863_)
  );
  INV_X1 _12109_ (
    .A(_01863_),
    .ZN(_01864_)
  );
  AND2_X1 _12110_ (
    .A1(io_req_bits_in2[17]),
    .A2(_06190_),
    .ZN(_01865_)
  );
  INV_X1 _12111_ (
    .A(_01865_),
    .ZN(_01866_)
  );
  AND2_X1 _12112_ (
    .A1(divisor[17]),
    .A2(_00164_),
    .ZN(_01867_)
  );
  INV_X1 _12113_ (
    .A(_01867_),
    .ZN(_01868_)
  );
  AND2_X1 _12114_ (
    .A1(_01866_),
    .A2(_01868_),
    .ZN(_01869_)
  );
  AND2_X1 _12115_ (
    .A1(_01864_),
    .A2(_01869_),
    .ZN(_01870_)
  );
  INV_X1 _12116_ (
    .A(_01870_),
    .ZN(_00037_)
  );
  AND2_X1 _12117_ (
    .A1(_07590_),
    .A2(_09464_),
    .ZN(_01871_)
  );
  INV_X1 _12118_ (
    .A(_01871_),
    .ZN(_01872_)
  );
  AND2_X1 _12119_ (
    .A1(_09497_),
    .A2(_01872_),
    .ZN(_01873_)
  );
  AND2_X1 _12120_ (
    .A1(_00262_),
    .A2(_01873_),
    .ZN(_01874_)
  );
  INV_X1 _12121_ (
    .A(_01874_),
    .ZN(_01875_)
  );
  AND2_X1 _12122_ (
    .A1(io_req_bits_in2[18]),
    .A2(_06190_),
    .ZN(_01876_)
  );
  INV_X1 _12123_ (
    .A(_01876_),
    .ZN(_01877_)
  );
  AND2_X1 _12124_ (
    .A1(divisor[18]),
    .A2(_00164_),
    .ZN(_01878_)
  );
  INV_X1 _12125_ (
    .A(_01878_),
    .ZN(_01879_)
  );
  AND2_X1 _12126_ (
    .A1(_01877_),
    .A2(_01879_),
    .ZN(_01880_)
  );
  AND2_X1 _12127_ (
    .A1(_01875_),
    .A2(_01880_),
    .ZN(_01881_)
  );
  INV_X1 _12128_ (
    .A(_01881_),
    .ZN(_00038_)
  );
  AND2_X1 _12129_ (
    .A1(_07502_),
    .A2(_07524_),
    .ZN(_01882_)
  );
  INV_X1 _12130_ (
    .A(_01882_),
    .ZN(_01883_)
  );
  AND2_X1 _12131_ (
    .A1(_09519_),
    .A2(_01883_),
    .ZN(_01884_)
  );
  INV_X1 _12132_ (
    .A(_01884_),
    .ZN(_01885_)
  );
  AND2_X1 _12133_ (
    .A1(_09508_),
    .A2(_01882_),
    .ZN(_01886_)
  );
  INV_X1 _12134_ (
    .A(_01886_),
    .ZN(_01887_)
  );
  AND2_X1 _12135_ (
    .A1(_09508_),
    .A2(_01883_),
    .ZN(_01888_)
  );
  INV_X1 _12136_ (
    .A(_01888_),
    .ZN(_01889_)
  );
  AND2_X1 _12137_ (
    .A1(_09519_),
    .A2(_01882_),
    .ZN(_01890_)
  );
  INV_X1 _12138_ (
    .A(_01890_),
    .ZN(_01891_)
  );
  AND2_X1 _12139_ (
    .A1(_01885_),
    .A2(_01887_),
    .ZN(_01892_)
  );
  AND2_X1 _12140_ (
    .A1(_01889_),
    .A2(_01891_),
    .ZN(_01893_)
  );
  AND2_X1 _12141_ (
    .A1(_00262_),
    .A2(_01893_),
    .ZN(_01894_)
  );
  INV_X1 _12142_ (
    .A(_01894_),
    .ZN(_01895_)
  );
  AND2_X1 _12143_ (
    .A1(io_req_bits_in2[19]),
    .A2(_06190_),
    .ZN(_01896_)
  );
  INV_X1 _12144_ (
    .A(_01896_),
    .ZN(_01897_)
  );
  AND2_X1 _12145_ (
    .A1(divisor[19]),
    .A2(_00164_),
    .ZN(_01898_)
  );
  INV_X1 _12146_ (
    .A(_01898_),
    .ZN(_01899_)
  );
  AND2_X1 _12147_ (
    .A1(_01897_),
    .A2(_01899_),
    .ZN(_01900_)
  );
  AND2_X1 _12148_ (
    .A1(_01895_),
    .A2(_01900_),
    .ZN(_01901_)
  );
  INV_X1 _12149_ (
    .A(_01901_),
    .ZN(_00039_)
  );
  AND2_X1 _12150_ (
    .A1(_07480_),
    .A2(_09574_),
    .ZN(_01902_)
  );
  INV_X1 _12151_ (
    .A(_01902_),
    .ZN(_01903_)
  );
  AND2_X1 _12152_ (
    .A1(_09607_),
    .A2(_01903_),
    .ZN(_01904_)
  );
  INV_X1 _12153_ (
    .A(_01904_),
    .ZN(_01905_)
  );
  AND2_X1 _12154_ (
    .A1(_00262_),
    .A2(_01904_),
    .ZN(_01906_)
  );
  INV_X1 _12155_ (
    .A(_01906_),
    .ZN(_01907_)
  );
  AND2_X1 _12156_ (
    .A1(divisor[20]),
    .A2(_00164_),
    .ZN(_01908_)
  );
  INV_X1 _12157_ (
    .A(_01908_),
    .ZN(_01909_)
  );
  AND2_X1 _12158_ (
    .A1(io_req_bits_in2[20]),
    .A2(_06190_),
    .ZN(_01910_)
  );
  INV_X1 _12159_ (
    .A(_01910_),
    .ZN(_01911_)
  );
  AND2_X1 _12160_ (
    .A1(_01909_),
    .A2(_01911_),
    .ZN(_01912_)
  );
  AND2_X1 _12161_ (
    .A1(_01907_),
    .A2(_01912_),
    .ZN(_01913_)
  );
  INV_X1 _12162_ (
    .A(_01913_),
    .ZN(_00040_)
  );
  AND2_X1 _12163_ (
    .A1(_07392_),
    .A2(_07414_),
    .ZN(_01914_)
  );
  INV_X1 _12164_ (
    .A(_01914_),
    .ZN(_01915_)
  );
  AND2_X1 _12165_ (
    .A1(_09629_),
    .A2(_01915_),
    .ZN(_01916_)
  );
  INV_X1 _12166_ (
    .A(_01916_),
    .ZN(_01917_)
  );
  AND2_X1 _12167_ (
    .A1(_09618_),
    .A2(_01914_),
    .ZN(_01918_)
  );
  INV_X1 _12168_ (
    .A(_01918_),
    .ZN(_01919_)
  );
  AND2_X1 _12169_ (
    .A1(_09618_),
    .A2(_01915_),
    .ZN(_01920_)
  );
  INV_X1 _12170_ (
    .A(_01920_),
    .ZN(_01921_)
  );
  AND2_X1 _12171_ (
    .A1(_09629_),
    .A2(_01914_),
    .ZN(_01922_)
  );
  INV_X1 _12172_ (
    .A(_01922_),
    .ZN(_01923_)
  );
  AND2_X1 _12173_ (
    .A1(_01917_),
    .A2(_01919_),
    .ZN(_01924_)
  );
  AND2_X1 _12174_ (
    .A1(_01921_),
    .A2(_01923_),
    .ZN(_01925_)
  );
  AND2_X1 _12175_ (
    .A1(_00262_),
    .A2(_01925_),
    .ZN(_01926_)
  );
  INV_X1 _12176_ (
    .A(_01926_),
    .ZN(_01927_)
  );
  AND2_X1 _12177_ (
    .A1(io_req_bits_in2[21]),
    .A2(_06190_),
    .ZN(_01928_)
  );
  INV_X1 _12178_ (
    .A(_01928_),
    .ZN(_01929_)
  );
  AND2_X1 _12179_ (
    .A1(divisor[21]),
    .A2(_00164_),
    .ZN(_01930_)
  );
  INV_X1 _12180_ (
    .A(_01930_),
    .ZN(_01931_)
  );
  AND2_X1 _12181_ (
    .A1(_01929_),
    .A2(_01931_),
    .ZN(_01932_)
  );
  AND2_X1 _12182_ (
    .A1(_01927_),
    .A2(_01932_),
    .ZN(_01933_)
  );
  INV_X1 _12183_ (
    .A(_01933_),
    .ZN(_00041_)
  );
  AND2_X1 _12184_ (
    .A1(_07370_),
    .A2(_09684_),
    .ZN(_01934_)
  );
  INV_X1 _12185_ (
    .A(_01934_),
    .ZN(_01935_)
  );
  AND2_X1 _12186_ (
    .A1(_09717_),
    .A2(_01935_),
    .ZN(_01936_)
  );
  INV_X1 _12187_ (
    .A(_01936_),
    .ZN(_01937_)
  );
  AND2_X1 _12188_ (
    .A1(_00262_),
    .A2(_01936_),
    .ZN(_01938_)
  );
  INV_X1 _12189_ (
    .A(_01938_),
    .ZN(_01939_)
  );
  AND2_X1 _12190_ (
    .A1(divisor[22]),
    .A2(_00164_),
    .ZN(_01940_)
  );
  INV_X1 _12191_ (
    .A(_01940_),
    .ZN(_01941_)
  );
  AND2_X1 _12192_ (
    .A1(io_req_bits_in2[22]),
    .A2(_06190_),
    .ZN(_01942_)
  );
  INV_X1 _12193_ (
    .A(_01942_),
    .ZN(_01943_)
  );
  AND2_X1 _12194_ (
    .A1(_01941_),
    .A2(_01943_),
    .ZN(_01944_)
  );
  AND2_X1 _12195_ (
    .A1(_01939_),
    .A2(_01944_),
    .ZN(_01945_)
  );
  INV_X1 _12196_ (
    .A(_01945_),
    .ZN(_00042_)
  );
  AND2_X1 _12197_ (
    .A1(_07283_),
    .A2(_07304_),
    .ZN(_01946_)
  );
  INV_X1 _12198_ (
    .A(_01946_),
    .ZN(_01947_)
  );
  AND2_X1 _12199_ (
    .A1(_09728_),
    .A2(_01947_),
    .ZN(_01948_)
  );
  INV_X1 _12200_ (
    .A(_01948_),
    .ZN(_01949_)
  );
  AND2_X1 _12201_ (
    .A1(_09739_),
    .A2(_01946_),
    .ZN(_01950_)
  );
  INV_X1 _12202_ (
    .A(_01950_),
    .ZN(_01951_)
  );
  AND2_X1 _12203_ (
    .A1(_01949_),
    .A2(_01951_),
    .ZN(_01952_)
  );
  AND2_X1 _12204_ (
    .A1(_00262_),
    .A2(_01952_),
    .ZN(_01953_)
  );
  INV_X1 _12205_ (
    .A(_01953_),
    .ZN(_01954_)
  );
  AND2_X1 _12206_ (
    .A1(io_req_bits_in2[23]),
    .A2(_06190_),
    .ZN(_01955_)
  );
  INV_X1 _12207_ (
    .A(_01955_),
    .ZN(_01956_)
  );
  AND2_X1 _12208_ (
    .A1(divisor[23]),
    .A2(_00164_),
    .ZN(_01957_)
  );
  INV_X1 _12209_ (
    .A(_01957_),
    .ZN(_01958_)
  );
  AND2_X1 _12210_ (
    .A1(_01956_),
    .A2(_01958_),
    .ZN(_01959_)
  );
  AND2_X1 _12211_ (
    .A1(_01954_),
    .A2(_01959_),
    .ZN(_01960_)
  );
  INV_X1 _12212_ (
    .A(_01960_),
    .ZN(_00043_)
  );
  AND2_X1 _12213_ (
    .A1(_07261_),
    .A2(_09793_),
    .ZN(_01961_)
  );
  INV_X1 _12214_ (
    .A(_01961_),
    .ZN(_01962_)
  );
  AND2_X1 _12215_ (
    .A1(_09826_),
    .A2(_01962_),
    .ZN(_01963_)
  );
  INV_X1 _12216_ (
    .A(_01963_),
    .ZN(_01964_)
  );
  AND2_X1 _12217_ (
    .A1(_00262_),
    .A2(_01963_),
    .ZN(_01965_)
  );
  INV_X1 _12218_ (
    .A(_01965_),
    .ZN(_01966_)
  );
  AND2_X1 _12219_ (
    .A1(io_req_bits_in2[24]),
    .A2(_06190_),
    .ZN(_01967_)
  );
  INV_X1 _12220_ (
    .A(_01967_),
    .ZN(_01968_)
  );
  AND2_X1 _12221_ (
    .A1(divisor[24]),
    .A2(_00164_),
    .ZN(_01969_)
  );
  INV_X1 _12222_ (
    .A(_01969_),
    .ZN(_01970_)
  );
  AND2_X1 _12223_ (
    .A1(_01968_),
    .A2(_01970_),
    .ZN(_01971_)
  );
  AND2_X1 _12224_ (
    .A1(_01966_),
    .A2(_01971_),
    .ZN(_01972_)
  );
  INV_X1 _12225_ (
    .A(_01972_),
    .ZN(_00044_)
  );
  AND2_X1 _12226_ (
    .A1(_07173_),
    .A2(_07195_),
    .ZN(_01973_)
  );
  INV_X1 _12227_ (
    .A(_01973_),
    .ZN(_01974_)
  );
  AND2_X1 _12228_ (
    .A1(_09837_),
    .A2(_01974_),
    .ZN(_01975_)
  );
  INV_X1 _12229_ (
    .A(_01975_),
    .ZN(_01976_)
  );
  AND2_X1 _12230_ (
    .A1(_09848_),
    .A2(_01973_),
    .ZN(_01977_)
  );
  INV_X1 _12231_ (
    .A(_01977_),
    .ZN(_01978_)
  );
  AND2_X1 _12232_ (
    .A1(_01976_),
    .A2(_01978_),
    .ZN(_01979_)
  );
  AND2_X1 _12233_ (
    .A1(_00262_),
    .A2(_01979_),
    .ZN(_01980_)
  );
  INV_X1 _12234_ (
    .A(_01980_),
    .ZN(_01981_)
  );
  AND2_X1 _12235_ (
    .A1(divisor[25]),
    .A2(_00164_),
    .ZN(_01982_)
  );
  INV_X1 _12236_ (
    .A(_01982_),
    .ZN(_01983_)
  );
  AND2_X1 _12237_ (
    .A1(io_req_bits_in2[25]),
    .A2(_06190_),
    .ZN(_01984_)
  );
  INV_X1 _12238_ (
    .A(_01984_),
    .ZN(_01985_)
  );
  AND2_X1 _12239_ (
    .A1(_01983_),
    .A2(_01985_),
    .ZN(_01986_)
  );
  AND2_X1 _12240_ (
    .A1(_01981_),
    .A2(_01986_),
    .ZN(_01987_)
  );
  INV_X1 _12241_ (
    .A(_01987_),
    .ZN(_00045_)
  );
  AND2_X1 _12242_ (
    .A1(_07151_),
    .A2(_09914_),
    .ZN(_01988_)
  );
  INV_X1 _12243_ (
    .A(_01988_),
    .ZN(_01989_)
  );
  AND2_X1 _12244_ (
    .A1(_09936_),
    .A2(_01989_),
    .ZN(_01990_)
  );
  INV_X1 _12245_ (
    .A(_01990_),
    .ZN(_01991_)
  );
  AND2_X1 _12246_ (
    .A1(_00262_),
    .A2(_01990_),
    .ZN(_01992_)
  );
  INV_X1 _12247_ (
    .A(_01992_),
    .ZN(_01993_)
  );
  AND2_X1 _12248_ (
    .A1(divisor[26]),
    .A2(_00164_),
    .ZN(_01994_)
  );
  INV_X1 _12249_ (
    .A(_01994_),
    .ZN(_01995_)
  );
  AND2_X1 _12250_ (
    .A1(io_req_bits_in2[26]),
    .A2(_06190_),
    .ZN(_01996_)
  );
  INV_X1 _12251_ (
    .A(_01996_),
    .ZN(_01997_)
  );
  AND2_X1 _12252_ (
    .A1(_01995_),
    .A2(_01997_),
    .ZN(_01998_)
  );
  AND2_X1 _12253_ (
    .A1(_01993_),
    .A2(_01998_),
    .ZN(_01999_)
  );
  INV_X1 _12254_ (
    .A(_01999_),
    .ZN(_00046_)
  );
  AND2_X1 _12255_ (
    .A1(_07063_),
    .A2(_07085_),
    .ZN(_02000_)
  );
  INV_X1 _12256_ (
    .A(_02000_),
    .ZN(_02001_)
  );
  AND2_X1 _12257_ (
    .A1(_09947_),
    .A2(_02001_),
    .ZN(_02002_)
  );
  INV_X1 _12258_ (
    .A(_02002_),
    .ZN(_02003_)
  );
  AND2_X1 _12259_ (
    .A1(_09958_),
    .A2(_02000_),
    .ZN(_02004_)
  );
  INV_X1 _12260_ (
    .A(_02004_),
    .ZN(_02005_)
  );
  AND2_X1 _12261_ (
    .A1(_02003_),
    .A2(_02005_),
    .ZN(_02006_)
  );
  AND2_X1 _12262_ (
    .A1(_00262_),
    .A2(_02006_),
    .ZN(_02007_)
  );
  INV_X1 _12263_ (
    .A(_02007_),
    .ZN(_02008_)
  );
  AND2_X1 _12264_ (
    .A1(io_req_bits_in2[27]),
    .A2(_06190_),
    .ZN(_02009_)
  );
  INV_X1 _12265_ (
    .A(_02009_),
    .ZN(_02010_)
  );
  AND2_X1 _12266_ (
    .A1(divisor[27]),
    .A2(_00164_),
    .ZN(_02011_)
  );
  INV_X1 _12267_ (
    .A(_02011_),
    .ZN(_02012_)
  );
  AND2_X1 _12268_ (
    .A1(_02010_),
    .A2(_02012_),
    .ZN(_02013_)
  );
  AND2_X1 _12269_ (
    .A1(_02008_),
    .A2(_02013_),
    .ZN(_02014_)
  );
  INV_X1 _12270_ (
    .A(_02014_),
    .ZN(_00047_)
  );
  AND2_X1 _12271_ (
    .A1(_07041_),
    .A2(_10013_),
    .ZN(_02015_)
  );
  INV_X1 _12272_ (
    .A(_02015_),
    .ZN(_02016_)
  );
  AND2_X1 _12273_ (
    .A1(_10046_),
    .A2(_02016_),
    .ZN(_02017_)
  );
  INV_X1 _12274_ (
    .A(_02017_),
    .ZN(_02018_)
  );
  AND2_X1 _12275_ (
    .A1(_00262_),
    .A2(_02017_),
    .ZN(_02019_)
  );
  INV_X1 _12276_ (
    .A(_02019_),
    .ZN(_02020_)
  );
  AND2_X1 _12277_ (
    .A1(io_req_bits_in2[28]),
    .A2(_06190_),
    .ZN(_02021_)
  );
  INV_X1 _12278_ (
    .A(_02021_),
    .ZN(_02022_)
  );
  AND2_X1 _12279_ (
    .A1(divisor[28]),
    .A2(_00164_),
    .ZN(_02023_)
  );
  INV_X1 _12280_ (
    .A(_02023_),
    .ZN(_02024_)
  );
  AND2_X1 _12281_ (
    .A1(_02022_),
    .A2(_02024_),
    .ZN(_02025_)
  );
  AND2_X1 _12282_ (
    .A1(_02020_),
    .A2(_02025_),
    .ZN(_02026_)
  );
  INV_X1 _12283_ (
    .A(_02026_),
    .ZN(_00048_)
  );
  AND2_X1 _12284_ (
    .A1(_06954_),
    .A2(_06976_),
    .ZN(_02027_)
  );
  INV_X1 _12285_ (
    .A(_02027_),
    .ZN(_02028_)
  );
  AND2_X1 _12286_ (
    .A1(_10057_),
    .A2(_02028_),
    .ZN(_02029_)
  );
  INV_X1 _12287_ (
    .A(_02029_),
    .ZN(_02030_)
  );
  AND2_X1 _12288_ (
    .A1(_10068_),
    .A2(_02027_),
    .ZN(_02031_)
  );
  INV_X1 _12289_ (
    .A(_02031_),
    .ZN(_02032_)
  );
  AND2_X1 _12290_ (
    .A1(_02030_),
    .A2(_02032_),
    .ZN(_02033_)
  );
  INV_X1 _12291_ (
    .A(_02033_),
    .ZN(_02034_)
  );
  AND2_X1 _12292_ (
    .A1(_00262_),
    .A2(_02033_),
    .ZN(_02035_)
  );
  INV_X1 _12293_ (
    .A(_02035_),
    .ZN(_02036_)
  );
  AND2_X1 _12294_ (
    .A1(divisor[29]),
    .A2(_00164_),
    .ZN(_02037_)
  );
  INV_X1 _12295_ (
    .A(_02037_),
    .ZN(_02038_)
  );
  AND2_X1 _12296_ (
    .A1(io_req_bits_in2[29]),
    .A2(_06190_),
    .ZN(_02039_)
  );
  INV_X1 _12297_ (
    .A(_02039_),
    .ZN(_02040_)
  );
  AND2_X1 _12298_ (
    .A1(_02038_),
    .A2(_02040_),
    .ZN(_02041_)
  );
  AND2_X1 _12299_ (
    .A1(_02036_),
    .A2(_02041_),
    .ZN(_02042_)
  );
  INV_X1 _12300_ (
    .A(_02042_),
    .ZN(_00049_)
  );
  AND2_X1 _12301_ (
    .A1(_06932_),
    .A2(_10133_),
    .ZN(_02043_)
  );
  INV_X1 _12302_ (
    .A(_02043_),
    .ZN(_02044_)
  );
  AND2_X1 _12303_ (
    .A1(_10155_),
    .A2(_02044_),
    .ZN(_02045_)
  );
  INV_X1 _12304_ (
    .A(_02045_),
    .ZN(_02046_)
  );
  AND2_X1 _12305_ (
    .A1(_00262_),
    .A2(_02045_),
    .ZN(_02047_)
  );
  INV_X1 _12306_ (
    .A(_02047_),
    .ZN(_02048_)
  );
  AND2_X1 _12307_ (
    .A1(divisor[30]),
    .A2(_00164_),
    .ZN(_02049_)
  );
  INV_X1 _12308_ (
    .A(_02049_),
    .ZN(_02050_)
  );
  AND2_X1 _12309_ (
    .A1(io_req_bits_in2[30]),
    .A2(_06190_),
    .ZN(_02051_)
  );
  INV_X1 _12310_ (
    .A(_02051_),
    .ZN(_02052_)
  );
  AND2_X1 _12311_ (
    .A1(_02050_),
    .A2(_02052_),
    .ZN(_02053_)
  );
  AND2_X1 _12312_ (
    .A1(_02048_),
    .A2(_02053_),
    .ZN(_02054_)
  );
  INV_X1 _12313_ (
    .A(_02054_),
    .ZN(_00050_)
  );
  AND2_X1 _12314_ (
    .A1(_06844_),
    .A2(_06866_),
    .ZN(_02055_)
  );
  INV_X1 _12315_ (
    .A(_02055_),
    .ZN(_02056_)
  );
  AND2_X1 _12316_ (
    .A1(_10177_),
    .A2(_02056_),
    .ZN(_02057_)
  );
  INV_X1 _12317_ (
    .A(_02057_),
    .ZN(_02058_)
  );
  AND2_X1 _12318_ (
    .A1(_10166_),
    .A2(_02055_),
    .ZN(_02059_)
  );
  INV_X1 _12319_ (
    .A(_02059_),
    .ZN(_02060_)
  );
  AND2_X1 _12320_ (
    .A1(_02058_),
    .A2(_02060_),
    .ZN(_02061_)
  );
  AND2_X1 _12321_ (
    .A1(_06299_),
    .A2(_02061_),
    .ZN(_02062_)
  );
  INV_X1 _12322_ (
    .A(_02062_),
    .ZN(_02063_)
  );
  AND2_X1 _12323_ (
    .A1(divisor[31]),
    .A2(_02063_),
    .ZN(_02064_)
  );
  MUX2_X1 _12324_ (
    .A(io_req_bits_in2[31]),
    .B(_02064_),
    .S(_06201_),
    .Z(_00051_)
  );
  AND2_X1 _12325_ (
    .A1(_10451_),
    .A2(_00262_),
    .ZN(_02065_)
  );
  INV_X1 _12326_ (
    .A(_02065_),
    .ZN(_02066_)
  );
  AND2_X1 _12327_ (
    .A1(_06190_),
    .A2(_06746_),
    .ZN(_02067_)
  );
  INV_X1 _12328_ (
    .A(_02067_),
    .ZN(_02068_)
  );
  AND2_X1 _12329_ (
    .A1(divisor[32]),
    .A2(_00164_),
    .ZN(_02069_)
  );
  INV_X1 _12330_ (
    .A(_02069_),
    .ZN(_02070_)
  );
  AND2_X1 _12331_ (
    .A1(_02068_),
    .A2(_02070_),
    .ZN(_02071_)
  );
  AND2_X1 _12332_ (
    .A1(_02066_),
    .A2(_02071_),
    .ZN(_02072_)
  );
  INV_X1 _12333_ (
    .A(_02072_),
    .ZN(_00052_)
  );
  AND2_X1 _12334_ (
    .A1(remainder[31]),
    .A2(_06299_),
    .ZN(_02073_)
  );
  INV_X1 _12335_ (
    .A(_02073_),
    .ZN(_02074_)
  );
  AND2_X1 _12336_ (
    .A1(_06256_),
    .A2(_02074_),
    .ZN(_02075_)
  );
  INV_X1 _12337_ (
    .A(_02075_),
    .ZN(_02076_)
  );
  AND2_X1 _12338_ (
    .A1(_10774_),
    .A2(_02075_),
    .ZN(_02077_)
  );
  AND2_X1 _12339_ (
    .A1(remainder[32]),
    .A2(_02077_),
    .ZN(_02078_)
  );
  INV_X1 _12340_ (
    .A(_02078_),
    .ZN(_02079_)
  );
  AND2_X1 _12341_ (
    .A1(remainder[31]),
    .A2(_05983_),
    .ZN(_02080_)
  );
  INV_X1 _12342_ (
    .A(_02080_),
    .ZN(_02081_)
  );
  AND2_X1 _12343_ (
    .A1(_00004_),
    .A2(_06103_),
    .ZN(_02082_)
  );
  AND2_X1 _12344_ (
    .A1(_04831_),
    .A2(neg_out),
    .ZN(_02083_)
  );
  AND2_X1 _12345_ (
    .A1(_06070_),
    .A2(_02083_),
    .ZN(_02084_)
  );
  AND2_X1 _12346_ (
    .A1(_02082_),
    .A2(_02084_),
    .ZN(_02085_)
  );
  INV_X1 _12347_ (
    .A(_02085_),
    .ZN(_02086_)
  );
  AND2_X1 _12348_ (
    .A1(_02081_),
    .A2(_02086_),
    .ZN(_02087_)
  );
  AND2_X1 _12349_ (
    .A1(_02079_),
    .A2(_02087_),
    .ZN(_02088_)
  );
  INV_X1 _12350_ (
    .A(_02088_),
    .ZN(_02089_)
  );
  AND2_X1 _12351_ (
    .A1(_06201_),
    .A2(_02089_),
    .ZN(_00053_)
  );
  MUX2_X1 _12352_ (
    .A(remainder[32]),
    .B(_00251_),
    .S(_10462_),
    .Z(_02090_)
  );
  AND2_X1 _12353_ (
    .A1(_05983_),
    .A2(_02090_),
    .ZN(_02091_)
  );
  INV_X1 _12354_ (
    .A(_02091_),
    .ZN(_02092_)
  );
  AND2_X1 _12355_ (
    .A1(remainder[33]),
    .A2(_02077_),
    .ZN(_02093_)
  );
  INV_X1 _12356_ (
    .A(_02093_),
    .ZN(_02094_)
  );
  AND2_X1 _12357_ (
    .A1(divisor[3]),
    .A2(remainder[3]),
    .ZN(_02095_)
  );
  INV_X1 _12358_ (
    .A(_02095_),
    .ZN(_02096_)
  );
  AND2_X1 _12359_ (
    .A1(divisor[0]),
    .A2(remainder[4]),
    .ZN(_02097_)
  );
  INV_X1 _12360_ (
    .A(_02097_),
    .ZN(_02098_)
  );
  AND2_X1 _12361_ (
    .A1(divisor[1]),
    .A2(remainder[3]),
    .ZN(_02099_)
  );
  INV_X1 _12362_ (
    .A(_02099_),
    .ZN(_02100_)
  );
  AND2_X1 _12363_ (
    .A1(divisor[1]),
    .A2(remainder[4]),
    .ZN(_02101_)
  );
  INV_X1 _12364_ (
    .A(_02101_),
    .ZN(_02102_)
  );
  AND2_X1 _12365_ (
    .A1(divisor[0]),
    .A2(remainder[3]),
    .ZN(_02103_)
  );
  INV_X1 _12366_ (
    .A(_02103_),
    .ZN(_02104_)
  );
  AND2_X1 _12367_ (
    .A1(_02097_),
    .A2(_02099_),
    .ZN(_02105_)
  );
  INV_X1 _12368_ (
    .A(_02105_),
    .ZN(_02106_)
  );
  AND2_X1 _12369_ (
    .A1(divisor[2]),
    .A2(remainder[2]),
    .ZN(_02107_)
  );
  INV_X1 _12370_ (
    .A(_02107_),
    .ZN(_02108_)
  );
  AND2_X1 _12371_ (
    .A1(_02098_),
    .A2(_02100_),
    .ZN(_02109_)
  );
  INV_X1 _12372_ (
    .A(_02109_),
    .ZN(_02110_)
  );
  AND2_X1 _12373_ (
    .A1(_02106_),
    .A2(_02110_),
    .ZN(_02111_)
  );
  INV_X1 _12374_ (
    .A(_02111_),
    .ZN(_02112_)
  );
  AND2_X1 _12375_ (
    .A1(_02107_),
    .A2(_02111_),
    .ZN(_02113_)
  );
  INV_X1 _12376_ (
    .A(_02113_),
    .ZN(_02114_)
  );
  AND2_X1 _12377_ (
    .A1(_02106_),
    .A2(_02114_),
    .ZN(_02115_)
  );
  INV_X1 _12378_ (
    .A(_02115_),
    .ZN(_02116_)
  );
  AND2_X1 _12379_ (
    .A1(divisor[4]),
    .A2(remainder[0]),
    .ZN(_02117_)
  );
  INV_X1 _12380_ (
    .A(_02117_),
    .ZN(_02118_)
  );
  AND2_X1 _12381_ (
    .A1(_02108_),
    .A2(_02112_),
    .ZN(_02119_)
  );
  INV_X1 _12382_ (
    .A(_02119_),
    .ZN(_02120_)
  );
  AND2_X1 _12383_ (
    .A1(_02114_),
    .A2(_02120_),
    .ZN(_02121_)
  );
  INV_X1 _12384_ (
    .A(_02121_),
    .ZN(_02122_)
  );
  AND2_X1 _12385_ (
    .A1(_02117_),
    .A2(_02121_),
    .ZN(_02123_)
  );
  INV_X1 _12386_ (
    .A(_02123_),
    .ZN(_02124_)
  );
  AND2_X1 _12387_ (
    .A1(divisor[2]),
    .A2(remainder[3]),
    .ZN(_02125_)
  );
  INV_X1 _12388_ (
    .A(_02125_),
    .ZN(_02126_)
  );
  AND2_X1 _12389_ (
    .A1(divisor[0]),
    .A2(remainder[5]),
    .ZN(_02127_)
  );
  INV_X1 _12390_ (
    .A(_02127_),
    .ZN(_02128_)
  );
  AND2_X1 _12391_ (
    .A1(divisor[1]),
    .A2(remainder[5]),
    .ZN(_02129_)
  );
  INV_X1 _12392_ (
    .A(_02129_),
    .ZN(_02130_)
  );
  AND2_X1 _12393_ (
    .A1(_02101_),
    .A2(_02127_),
    .ZN(_02131_)
  );
  INV_X1 _12394_ (
    .A(_02131_),
    .ZN(_02132_)
  );
  AND2_X1 _12395_ (
    .A1(_02102_),
    .A2(_02128_),
    .ZN(_02133_)
  );
  INV_X1 _12396_ (
    .A(_02133_),
    .ZN(_02134_)
  );
  AND2_X1 _12397_ (
    .A1(_02132_),
    .A2(_02134_),
    .ZN(_02135_)
  );
  INV_X1 _12398_ (
    .A(_02135_),
    .ZN(_02136_)
  );
  AND2_X1 _12399_ (
    .A1(_02125_),
    .A2(_02135_),
    .ZN(_02137_)
  );
  INV_X1 _12400_ (
    .A(_02137_),
    .ZN(_02138_)
  );
  AND2_X1 _12401_ (
    .A1(_02126_),
    .A2(_02136_),
    .ZN(_02139_)
  );
  INV_X1 _12402_ (
    .A(_02139_),
    .ZN(_02140_)
  );
  AND2_X1 _12403_ (
    .A1(_02138_),
    .A2(_02140_),
    .ZN(_02141_)
  );
  INV_X1 _12404_ (
    .A(_02141_),
    .ZN(_02142_)
  );
  AND2_X1 _12405_ (
    .A1(divisor[4]),
    .A2(remainder[1]),
    .ZN(_02143_)
  );
  INV_X1 _12406_ (
    .A(_02143_),
    .ZN(_02144_)
  );
  AND2_X1 _12407_ (
    .A1(divisor[5]),
    .A2(remainder[0]),
    .ZN(_02145_)
  );
  INV_X1 _12408_ (
    .A(_02145_),
    .ZN(_02146_)
  );
  AND2_X1 _12409_ (
    .A1(divisor[5]),
    .A2(remainder[1]),
    .ZN(_02147_)
  );
  INV_X1 _12410_ (
    .A(_02147_),
    .ZN(_02148_)
  );
  AND2_X1 _12411_ (
    .A1(_02117_),
    .A2(_02147_),
    .ZN(_02149_)
  );
  INV_X1 _12412_ (
    .A(_02149_),
    .ZN(_02150_)
  );
  AND2_X1 _12413_ (
    .A1(_02144_),
    .A2(_02146_),
    .ZN(_02151_)
  );
  INV_X1 _12414_ (
    .A(_02151_),
    .ZN(_02152_)
  );
  AND2_X1 _12415_ (
    .A1(_02150_),
    .A2(_02152_),
    .ZN(_02153_)
  );
  INV_X1 _12416_ (
    .A(_02153_),
    .ZN(_02154_)
  );
  AND2_X1 _12417_ (
    .A1(_02141_),
    .A2(_02153_),
    .ZN(_02155_)
  );
  INV_X1 _12418_ (
    .A(_02155_),
    .ZN(_02156_)
  );
  AND2_X1 _12419_ (
    .A1(_02142_),
    .A2(_02154_),
    .ZN(_02157_)
  );
  INV_X1 _12420_ (
    .A(_02157_),
    .ZN(_02158_)
  );
  AND2_X1 _12421_ (
    .A1(_02156_),
    .A2(_02158_),
    .ZN(_02159_)
  );
  INV_X1 _12422_ (
    .A(_02159_),
    .ZN(_02160_)
  );
  AND2_X1 _12423_ (
    .A1(_02123_),
    .A2(_02159_),
    .ZN(_02161_)
  );
  INV_X1 _12424_ (
    .A(_02161_),
    .ZN(_02162_)
  );
  AND2_X1 _12425_ (
    .A1(_02124_),
    .A2(_02160_),
    .ZN(_02163_)
  );
  INV_X1 _12426_ (
    .A(_02163_),
    .ZN(_02164_)
  );
  AND2_X1 _12427_ (
    .A1(_02162_),
    .A2(_02164_),
    .ZN(_02165_)
  );
  INV_X1 _12428_ (
    .A(_02165_),
    .ZN(_02166_)
  );
  AND2_X1 _12429_ (
    .A1(_02116_),
    .A2(_02165_),
    .ZN(_02167_)
  );
  INV_X1 _12430_ (
    .A(_02167_),
    .ZN(_02168_)
  );
  AND2_X1 _12431_ (
    .A1(_02132_),
    .A2(_02138_),
    .ZN(_02169_)
  );
  INV_X1 _12432_ (
    .A(_02169_),
    .ZN(_02170_)
  );
  AND2_X1 _12433_ (
    .A1(divisor[2]),
    .A2(remainder[4]),
    .ZN(_02171_)
  );
  INV_X1 _12434_ (
    .A(_02171_),
    .ZN(_02172_)
  );
  AND2_X1 _12435_ (
    .A1(divisor[0]),
    .A2(remainder[6]),
    .ZN(_02173_)
  );
  INV_X1 _12436_ (
    .A(_02173_),
    .ZN(_02174_)
  );
  AND2_X1 _12437_ (
    .A1(divisor[1]),
    .A2(remainder[6]),
    .ZN(_02175_)
  );
  INV_X1 _12438_ (
    .A(_02175_),
    .ZN(_02176_)
  );
  AND2_X1 _12439_ (
    .A1(_02129_),
    .A2(_02173_),
    .ZN(_02177_)
  );
  INV_X1 _12440_ (
    .A(_02177_),
    .ZN(_02178_)
  );
  AND2_X1 _12441_ (
    .A1(_02130_),
    .A2(_02174_),
    .ZN(_02179_)
  );
  INV_X1 _12442_ (
    .A(_02179_),
    .ZN(_02180_)
  );
  AND2_X1 _12443_ (
    .A1(_02178_),
    .A2(_02180_),
    .ZN(_02181_)
  );
  INV_X1 _12444_ (
    .A(_02181_),
    .ZN(_02182_)
  );
  AND2_X1 _12445_ (
    .A1(_02171_),
    .A2(_02181_),
    .ZN(_02183_)
  );
  INV_X1 _12446_ (
    .A(_02183_),
    .ZN(_02184_)
  );
  AND2_X1 _12447_ (
    .A1(_02172_),
    .A2(_02182_),
    .ZN(_02185_)
  );
  INV_X1 _12448_ (
    .A(_02185_),
    .ZN(_02186_)
  );
  AND2_X1 _12449_ (
    .A1(_02184_),
    .A2(_02186_),
    .ZN(_02187_)
  );
  INV_X1 _12450_ (
    .A(_02187_),
    .ZN(_02188_)
  );
  AND2_X1 _12451_ (
    .A1(divisor[4]),
    .A2(remainder[2]),
    .ZN(_02189_)
  );
  INV_X1 _12452_ (
    .A(_02189_),
    .ZN(_02190_)
  );
  AND2_X1 _12453_ (
    .A1(divisor[6]),
    .A2(remainder[0]),
    .ZN(_02191_)
  );
  INV_X1 _12454_ (
    .A(_02191_),
    .ZN(_02192_)
  );
  AND2_X1 _12455_ (
    .A1(divisor[6]),
    .A2(remainder[1]),
    .ZN(_02193_)
  );
  INV_X1 _12456_ (
    .A(_02193_),
    .ZN(_02194_)
  );
  AND2_X1 _12457_ (
    .A1(_02145_),
    .A2(_02193_),
    .ZN(_02195_)
  );
  INV_X1 _12458_ (
    .A(_02195_),
    .ZN(_02196_)
  );
  AND2_X1 _12459_ (
    .A1(_02148_),
    .A2(_02192_),
    .ZN(_02197_)
  );
  INV_X1 _12460_ (
    .A(_02197_),
    .ZN(_02198_)
  );
  AND2_X1 _12461_ (
    .A1(_02196_),
    .A2(_02198_),
    .ZN(_02199_)
  );
  INV_X1 _12462_ (
    .A(_02199_),
    .ZN(_02200_)
  );
  AND2_X1 _12463_ (
    .A1(_02189_),
    .A2(_02199_),
    .ZN(_02201_)
  );
  INV_X1 _12464_ (
    .A(_02201_),
    .ZN(_02202_)
  );
  AND2_X1 _12465_ (
    .A1(_02190_),
    .A2(_02200_),
    .ZN(_02203_)
  );
  INV_X1 _12466_ (
    .A(_02203_),
    .ZN(_02204_)
  );
  AND2_X1 _12467_ (
    .A1(_02202_),
    .A2(_02204_),
    .ZN(_02205_)
  );
  INV_X1 _12468_ (
    .A(_02205_),
    .ZN(_02206_)
  );
  AND2_X1 _12469_ (
    .A1(_02149_),
    .A2(_02205_),
    .ZN(_02207_)
  );
  INV_X1 _12470_ (
    .A(_02207_),
    .ZN(_02208_)
  );
  AND2_X1 _12471_ (
    .A1(_02150_),
    .A2(_02206_),
    .ZN(_02209_)
  );
  INV_X1 _12472_ (
    .A(_02209_),
    .ZN(_02210_)
  );
  AND2_X1 _12473_ (
    .A1(_02208_),
    .A2(_02210_),
    .ZN(_02211_)
  );
  INV_X1 _12474_ (
    .A(_02211_),
    .ZN(_02212_)
  );
  AND2_X1 _12475_ (
    .A1(_02187_),
    .A2(_02211_),
    .ZN(_02213_)
  );
  INV_X1 _12476_ (
    .A(_02213_),
    .ZN(_02214_)
  );
  AND2_X1 _12477_ (
    .A1(_02188_),
    .A2(_02212_),
    .ZN(_02215_)
  );
  INV_X1 _12478_ (
    .A(_02215_),
    .ZN(_02216_)
  );
  AND2_X1 _12479_ (
    .A1(_02214_),
    .A2(_02216_),
    .ZN(_02217_)
  );
  INV_X1 _12480_ (
    .A(_02217_),
    .ZN(_02218_)
  );
  AND2_X1 _12481_ (
    .A1(_02155_),
    .A2(_02217_),
    .ZN(_02219_)
  );
  INV_X1 _12482_ (
    .A(_02219_),
    .ZN(_02220_)
  );
  AND2_X1 _12483_ (
    .A1(_02156_),
    .A2(_02218_),
    .ZN(_02221_)
  );
  INV_X1 _12484_ (
    .A(_02221_),
    .ZN(_02222_)
  );
  AND2_X1 _12485_ (
    .A1(_02220_),
    .A2(_02222_),
    .ZN(_02223_)
  );
  INV_X1 _12486_ (
    .A(_02223_),
    .ZN(_02224_)
  );
  AND2_X1 _12487_ (
    .A1(_02161_),
    .A2(_02223_),
    .ZN(_02225_)
  );
  INV_X1 _12488_ (
    .A(_02225_),
    .ZN(_02226_)
  );
  AND2_X1 _12489_ (
    .A1(_02162_),
    .A2(_02224_),
    .ZN(_02227_)
  );
  INV_X1 _12490_ (
    .A(_02227_),
    .ZN(_02228_)
  );
  AND2_X1 _12491_ (
    .A1(_02226_),
    .A2(_02228_),
    .ZN(_02229_)
  );
  INV_X1 _12492_ (
    .A(_02229_),
    .ZN(_02230_)
  );
  AND2_X1 _12493_ (
    .A1(_02170_),
    .A2(_02229_),
    .ZN(_02231_)
  );
  INV_X1 _12494_ (
    .A(_02231_),
    .ZN(_02232_)
  );
  AND2_X1 _12495_ (
    .A1(_02169_),
    .A2(_02230_),
    .ZN(_02233_)
  );
  INV_X1 _12496_ (
    .A(_02233_),
    .ZN(_02234_)
  );
  AND2_X1 _12497_ (
    .A1(_02232_),
    .A2(_02234_),
    .ZN(_02235_)
  );
  INV_X1 _12498_ (
    .A(_02235_),
    .ZN(_02236_)
  );
  AND2_X1 _12499_ (
    .A1(_02167_),
    .A2(_02235_),
    .ZN(_02237_)
  );
  INV_X1 _12500_ (
    .A(_02237_),
    .ZN(_02238_)
  );
  AND2_X1 _12501_ (
    .A1(_02168_),
    .A2(_02236_),
    .ZN(_02239_)
  );
  INV_X1 _12502_ (
    .A(_02239_),
    .ZN(_02240_)
  );
  AND2_X1 _12503_ (
    .A1(_02238_),
    .A2(_02240_),
    .ZN(_02241_)
  );
  INV_X1 _12504_ (
    .A(_02241_),
    .ZN(_02242_)
  );
  AND2_X1 _12505_ (
    .A1(_02095_),
    .A2(_02241_),
    .ZN(_02243_)
  );
  INV_X1 _12506_ (
    .A(_02243_),
    .ZN(_02244_)
  );
  AND2_X1 _12507_ (
    .A1(_02096_),
    .A2(_02242_),
    .ZN(_02245_)
  );
  INV_X1 _12508_ (
    .A(_02245_),
    .ZN(_02246_)
  );
  AND2_X1 _12509_ (
    .A1(_02244_),
    .A2(_02246_),
    .ZN(_02247_)
  );
  INV_X1 _12510_ (
    .A(_02247_),
    .ZN(_02248_)
  );
  AND2_X1 _12511_ (
    .A1(divisor[1]),
    .A2(remainder[2]),
    .ZN(_02249_)
  );
  INV_X1 _12512_ (
    .A(_02249_),
    .ZN(_02250_)
  );
  AND2_X1 _12513_ (
    .A1(divisor[0]),
    .A2(remainder[2]),
    .ZN(_02251_)
  );
  INV_X1 _12514_ (
    .A(_02251_),
    .ZN(_02252_)
  );
  AND2_X1 _12515_ (
    .A1(_02103_),
    .A2(_02249_),
    .ZN(_02253_)
  );
  INV_X1 _12516_ (
    .A(_02253_),
    .ZN(_02254_)
  );
  AND2_X1 _12517_ (
    .A1(divisor[2]),
    .A2(remainder[1]),
    .ZN(_02255_)
  );
  INV_X1 _12518_ (
    .A(_02255_),
    .ZN(_02256_)
  );
  AND2_X1 _12519_ (
    .A1(_02104_),
    .A2(_02250_),
    .ZN(_02257_)
  );
  INV_X1 _12520_ (
    .A(_02257_),
    .ZN(_02258_)
  );
  AND2_X1 _12521_ (
    .A1(_02254_),
    .A2(_02258_),
    .ZN(_02259_)
  );
  INV_X1 _12522_ (
    .A(_02259_),
    .ZN(_02260_)
  );
  AND2_X1 _12523_ (
    .A1(_02255_),
    .A2(_02259_),
    .ZN(_02261_)
  );
  INV_X1 _12524_ (
    .A(_02261_),
    .ZN(_02262_)
  );
  AND2_X1 _12525_ (
    .A1(_02254_),
    .A2(_02262_),
    .ZN(_02263_)
  );
  INV_X1 _12526_ (
    .A(_02263_),
    .ZN(_02264_)
  );
  AND2_X1 _12527_ (
    .A1(_02118_),
    .A2(_02122_),
    .ZN(_02265_)
  );
  INV_X1 _12528_ (
    .A(_02265_),
    .ZN(_02266_)
  );
  AND2_X1 _12529_ (
    .A1(_02124_),
    .A2(_02266_),
    .ZN(_02267_)
  );
  INV_X1 _12530_ (
    .A(_02267_),
    .ZN(_02268_)
  );
  AND2_X1 _12531_ (
    .A1(_02264_),
    .A2(_02267_),
    .ZN(_02269_)
  );
  INV_X1 _12532_ (
    .A(_02269_),
    .ZN(_02270_)
  );
  AND2_X1 _12533_ (
    .A1(_02115_),
    .A2(_02166_),
    .ZN(_02271_)
  );
  INV_X1 _12534_ (
    .A(_02271_),
    .ZN(_02272_)
  );
  AND2_X1 _12535_ (
    .A1(_02168_),
    .A2(_02272_),
    .ZN(_02273_)
  );
  INV_X1 _12536_ (
    .A(_02273_),
    .ZN(_02274_)
  );
  AND2_X1 _12537_ (
    .A1(_02269_),
    .A2(_02273_),
    .ZN(_02275_)
  );
  INV_X1 _12538_ (
    .A(_02275_),
    .ZN(_02276_)
  );
  AND2_X1 _12539_ (
    .A1(divisor[3]),
    .A2(remainder[2]),
    .ZN(_02277_)
  );
  INV_X1 _12540_ (
    .A(_02277_),
    .ZN(_02278_)
  );
  AND2_X1 _12541_ (
    .A1(_02270_),
    .A2(_02274_),
    .ZN(_02279_)
  );
  INV_X1 _12542_ (
    .A(_02279_),
    .ZN(_02280_)
  );
  AND2_X1 _12543_ (
    .A1(_02276_),
    .A2(_02280_),
    .ZN(_02281_)
  );
  INV_X1 _12544_ (
    .A(_02281_),
    .ZN(_02282_)
  );
  AND2_X1 _12545_ (
    .A1(_02277_),
    .A2(_02281_),
    .ZN(_02283_)
  );
  INV_X1 _12546_ (
    .A(_02283_),
    .ZN(_02284_)
  );
  AND2_X1 _12547_ (
    .A1(_02276_),
    .A2(_02284_),
    .ZN(_02285_)
  );
  INV_X1 _12548_ (
    .A(_02285_),
    .ZN(_02286_)
  );
  AND2_X1 _12549_ (
    .A1(_02247_),
    .A2(_02286_),
    .ZN(_02287_)
  );
  INV_X1 _12550_ (
    .A(_02287_),
    .ZN(_02288_)
  );
  AND2_X1 _12551_ (
    .A1(_02178_),
    .A2(_02184_),
    .ZN(_02289_)
  );
  INV_X1 _12552_ (
    .A(_02289_),
    .ZN(_02290_)
  );
  AND2_X1 _12553_ (
    .A1(_02208_),
    .A2(_02214_),
    .ZN(_02291_)
  );
  INV_X1 _12554_ (
    .A(_02291_),
    .ZN(_02292_)
  );
  AND2_X1 _12555_ (
    .A1(divisor[2]),
    .A2(remainder[5]),
    .ZN(_02293_)
  );
  INV_X1 _12556_ (
    .A(_02293_),
    .ZN(_02294_)
  );
  AND2_X1 _12557_ (
    .A1(divisor[0]),
    .A2(remainder[7]),
    .ZN(_02295_)
  );
  INV_X1 _12558_ (
    .A(_02295_),
    .ZN(_02296_)
  );
  AND2_X1 _12559_ (
    .A1(divisor[1]),
    .A2(remainder[7]),
    .ZN(_02297_)
  );
  INV_X1 _12560_ (
    .A(_02297_),
    .ZN(_02298_)
  );
  AND2_X1 _12561_ (
    .A1(_02173_),
    .A2(_02297_),
    .ZN(_02299_)
  );
  INV_X1 _12562_ (
    .A(_02299_),
    .ZN(_02300_)
  );
  AND2_X1 _12563_ (
    .A1(_02176_),
    .A2(_02296_),
    .ZN(_02301_)
  );
  INV_X1 _12564_ (
    .A(_02301_),
    .ZN(_02302_)
  );
  AND2_X1 _12565_ (
    .A1(_02300_),
    .A2(_02302_),
    .ZN(_02303_)
  );
  INV_X1 _12566_ (
    .A(_02303_),
    .ZN(_02304_)
  );
  AND2_X1 _12567_ (
    .A1(_02293_),
    .A2(_02303_),
    .ZN(_02305_)
  );
  INV_X1 _12568_ (
    .A(_02305_),
    .ZN(_02306_)
  );
  AND2_X1 _12569_ (
    .A1(_02294_),
    .A2(_02304_),
    .ZN(_02307_)
  );
  INV_X1 _12570_ (
    .A(_02307_),
    .ZN(_02308_)
  );
  AND2_X1 _12571_ (
    .A1(_02306_),
    .A2(_02308_),
    .ZN(_02309_)
  );
  INV_X1 _12572_ (
    .A(_02309_),
    .ZN(_02310_)
  );
  AND2_X1 _12573_ (
    .A1(_02196_),
    .A2(_02202_),
    .ZN(_02311_)
  );
  INV_X1 _12574_ (
    .A(_02311_),
    .ZN(_02312_)
  );
  AND2_X1 _12575_ (
    .A1(divisor[4]),
    .A2(remainder[3]),
    .ZN(_02313_)
  );
  INV_X1 _12576_ (
    .A(_02313_),
    .ZN(_02314_)
  );
  AND2_X1 _12577_ (
    .A1(divisor[5]),
    .A2(remainder[2]),
    .ZN(_02315_)
  );
  INV_X1 _12578_ (
    .A(_02315_),
    .ZN(_02316_)
  );
  AND2_X1 _12579_ (
    .A1(divisor[6]),
    .A2(remainder[2]),
    .ZN(_02317_)
  );
  INV_X1 _12580_ (
    .A(_02317_),
    .ZN(_02318_)
  );
  AND2_X1 _12581_ (
    .A1(_02147_),
    .A2(_02317_),
    .ZN(_02319_)
  );
  INV_X1 _12582_ (
    .A(_02319_),
    .ZN(_02320_)
  );
  AND2_X1 _12583_ (
    .A1(_02194_),
    .A2(_02316_),
    .ZN(_02321_)
  );
  INV_X1 _12584_ (
    .A(_02321_),
    .ZN(_02322_)
  );
  AND2_X1 _12585_ (
    .A1(_02320_),
    .A2(_02322_),
    .ZN(_02323_)
  );
  INV_X1 _12586_ (
    .A(_02323_),
    .ZN(_02324_)
  );
  AND2_X1 _12587_ (
    .A1(_02313_),
    .A2(_02323_),
    .ZN(_02325_)
  );
  INV_X1 _12588_ (
    .A(_02325_),
    .ZN(_02326_)
  );
  AND2_X1 _12589_ (
    .A1(_02314_),
    .A2(_02324_),
    .ZN(_02327_)
  );
  INV_X1 _12590_ (
    .A(_02327_),
    .ZN(_02328_)
  );
  AND2_X1 _12591_ (
    .A1(_02326_),
    .A2(_02328_),
    .ZN(_02329_)
  );
  INV_X1 _12592_ (
    .A(_02329_),
    .ZN(_02330_)
  );
  AND2_X1 _12593_ (
    .A1(_02312_),
    .A2(_02329_),
    .ZN(_02331_)
  );
  INV_X1 _12594_ (
    .A(_02331_),
    .ZN(_02332_)
  );
  AND2_X1 _12595_ (
    .A1(_02311_),
    .A2(_02330_),
    .ZN(_02333_)
  );
  INV_X1 _12596_ (
    .A(_02333_),
    .ZN(_02334_)
  );
  AND2_X1 _12597_ (
    .A1(_02332_),
    .A2(_02334_),
    .ZN(_02335_)
  );
  INV_X1 _12598_ (
    .A(_02335_),
    .ZN(_02336_)
  );
  AND2_X1 _12599_ (
    .A1(_02309_),
    .A2(_02335_),
    .ZN(_02337_)
  );
  INV_X1 _12600_ (
    .A(_02337_),
    .ZN(_02338_)
  );
  AND2_X1 _12601_ (
    .A1(_02310_),
    .A2(_02336_),
    .ZN(_02339_)
  );
  INV_X1 _12602_ (
    .A(_02339_),
    .ZN(_02340_)
  );
  AND2_X1 _12603_ (
    .A1(_02338_),
    .A2(_02340_),
    .ZN(_02341_)
  );
  INV_X1 _12604_ (
    .A(_02341_),
    .ZN(_02342_)
  );
  AND2_X1 _12605_ (
    .A1(_02292_),
    .A2(_02341_),
    .ZN(_02343_)
  );
  INV_X1 _12606_ (
    .A(_02343_),
    .ZN(_02344_)
  );
  AND2_X1 _12607_ (
    .A1(_02291_),
    .A2(_02342_),
    .ZN(_02345_)
  );
  INV_X1 _12608_ (
    .A(_02345_),
    .ZN(_02346_)
  );
  AND2_X1 _12609_ (
    .A1(_02344_),
    .A2(_02346_),
    .ZN(_02347_)
  );
  INV_X1 _12610_ (
    .A(_02347_),
    .ZN(_02348_)
  );
  AND2_X1 _12611_ (
    .A1(_02220_),
    .A2(_02226_),
    .ZN(_02349_)
  );
  INV_X1 _12612_ (
    .A(_02349_),
    .ZN(_02350_)
  );
  AND2_X1 _12613_ (
    .A1(_02348_),
    .A2(_02349_),
    .ZN(_02351_)
  );
  INV_X1 _12614_ (
    .A(_02351_),
    .ZN(_02352_)
  );
  AND2_X1 _12615_ (
    .A1(_02347_),
    .A2(_02350_),
    .ZN(_02353_)
  );
  INV_X1 _12616_ (
    .A(_02353_),
    .ZN(_02354_)
  );
  AND2_X1 _12617_ (
    .A1(_02347_),
    .A2(_02349_),
    .ZN(_02355_)
  );
  INV_X1 _12618_ (
    .A(_02355_),
    .ZN(_02356_)
  );
  AND2_X1 _12619_ (
    .A1(_02348_),
    .A2(_02350_),
    .ZN(_02357_)
  );
  INV_X1 _12620_ (
    .A(_02357_),
    .ZN(_02358_)
  );
  AND2_X1 _12621_ (
    .A1(_02352_),
    .A2(_02354_),
    .ZN(_02359_)
  );
  AND2_X1 _12622_ (
    .A1(_02356_),
    .A2(_02358_),
    .ZN(_02360_)
  );
  AND2_X1 _12623_ (
    .A1(_02290_),
    .A2(_02359_),
    .ZN(_02361_)
  );
  INV_X1 _12624_ (
    .A(_02361_),
    .ZN(_02362_)
  );
  AND2_X1 _12625_ (
    .A1(_02289_),
    .A2(_02360_),
    .ZN(_02363_)
  );
  INV_X1 _12626_ (
    .A(_02363_),
    .ZN(_02364_)
  );
  AND2_X1 _12627_ (
    .A1(_02362_),
    .A2(_02364_),
    .ZN(_02365_)
  );
  INV_X1 _12628_ (
    .A(_02365_),
    .ZN(_02366_)
  );
  AND2_X1 _12629_ (
    .A1(_02231_),
    .A2(_02365_),
    .ZN(_02367_)
  );
  INV_X1 _12630_ (
    .A(_02367_),
    .ZN(_02368_)
  );
  AND2_X1 _12631_ (
    .A1(_02232_),
    .A2(_02366_),
    .ZN(_02369_)
  );
  INV_X1 _12632_ (
    .A(_02369_),
    .ZN(_02370_)
  );
  AND2_X1 _12633_ (
    .A1(_02368_),
    .A2(_02370_),
    .ZN(_02371_)
  );
  INV_X1 _12634_ (
    .A(_02371_),
    .ZN(_02372_)
  );
  AND2_X1 _12635_ (
    .A1(divisor[7]),
    .A2(remainder[0]),
    .ZN(_02373_)
  );
  INV_X1 _12636_ (
    .A(_02373_),
    .ZN(_02374_)
  );
  AND2_X1 _12637_ (
    .A1(divisor[3]),
    .A2(remainder[4]),
    .ZN(_02375_)
  );
  INV_X1 _12638_ (
    .A(_02375_),
    .ZN(_02376_)
  );
  AND2_X1 _12639_ (
    .A1(divisor[3]),
    .A2(remainder[0]),
    .ZN(_02377_)
  );
  INV_X1 _12640_ (
    .A(_02377_),
    .ZN(_02378_)
  );
  AND2_X1 _12641_ (
    .A1(divisor[7]),
    .A2(remainder[4]),
    .ZN(_02379_)
  );
  INV_X1 _12642_ (
    .A(_02379_),
    .ZN(_02380_)
  );
  AND2_X1 _12643_ (
    .A1(_02377_),
    .A2(_02379_),
    .ZN(_02381_)
  );
  INV_X1 _12644_ (
    .A(_02381_),
    .ZN(_02382_)
  );
  AND2_X1 _12645_ (
    .A1(_02374_),
    .A2(_02376_),
    .ZN(_02383_)
  );
  INV_X1 _12646_ (
    .A(_02383_),
    .ZN(_02384_)
  );
  AND2_X1 _12647_ (
    .A1(_02382_),
    .A2(_02384_),
    .ZN(_02385_)
  );
  INV_X1 _12648_ (
    .A(_02385_),
    .ZN(_02386_)
  );
  AND2_X1 _12649_ (
    .A1(_02371_),
    .A2(_02385_),
    .ZN(_02387_)
  );
  INV_X1 _12650_ (
    .A(_02387_),
    .ZN(_02388_)
  );
  AND2_X1 _12651_ (
    .A1(_02372_),
    .A2(_02386_),
    .ZN(_02389_)
  );
  INV_X1 _12652_ (
    .A(_02389_),
    .ZN(_02390_)
  );
  AND2_X1 _12653_ (
    .A1(_02388_),
    .A2(_02390_),
    .ZN(_02391_)
  );
  INV_X1 _12654_ (
    .A(_02391_),
    .ZN(_02392_)
  );
  AND2_X1 _12655_ (
    .A1(_02238_),
    .A2(_02244_),
    .ZN(_02393_)
  );
  INV_X1 _12656_ (
    .A(_02393_),
    .ZN(_02394_)
  );
  AND2_X1 _12657_ (
    .A1(_02391_),
    .A2(_02394_),
    .ZN(_02395_)
  );
  INV_X1 _12658_ (
    .A(_02395_),
    .ZN(_02396_)
  );
  AND2_X1 _12659_ (
    .A1(_02392_),
    .A2(_02393_),
    .ZN(_02397_)
  );
  INV_X1 _12660_ (
    .A(_02397_),
    .ZN(_02398_)
  );
  AND2_X1 _12661_ (
    .A1(_02396_),
    .A2(_02398_),
    .ZN(_02399_)
  );
  INV_X1 _12662_ (
    .A(_02399_),
    .ZN(_02400_)
  );
  AND2_X1 _12663_ (
    .A1(_02287_),
    .A2(_02399_),
    .ZN(_02401_)
  );
  INV_X1 _12664_ (
    .A(_02401_),
    .ZN(_02402_)
  );
  AND2_X1 _12665_ (
    .A1(_02288_),
    .A2(_02400_),
    .ZN(_02403_)
  );
  INV_X1 _12666_ (
    .A(_02403_),
    .ZN(_02404_)
  );
  AND2_X1 _12667_ (
    .A1(_02402_),
    .A2(_02404_),
    .ZN(_02405_)
  );
  INV_X1 _12668_ (
    .A(_02405_),
    .ZN(_02406_)
  );
  AND2_X1 _12669_ (
    .A1(_02248_),
    .A2(_02285_),
    .ZN(_02407_)
  );
  INV_X1 _12670_ (
    .A(_02407_),
    .ZN(_02408_)
  );
  AND2_X1 _12671_ (
    .A1(_02288_),
    .A2(_02408_),
    .ZN(_02409_)
  );
  INV_X1 _12672_ (
    .A(_02409_),
    .ZN(_02410_)
  );
  AND2_X1 _12673_ (
    .A1(_02278_),
    .A2(_02282_),
    .ZN(_02411_)
  );
  INV_X1 _12674_ (
    .A(_02411_),
    .ZN(_02412_)
  );
  AND2_X1 _12675_ (
    .A1(_02284_),
    .A2(_02412_),
    .ZN(_02413_)
  );
  INV_X1 _12676_ (
    .A(_02413_),
    .ZN(_02414_)
  );
  AND2_X1 _12677_ (
    .A1(divisor[1]),
    .A2(remainder[1]),
    .ZN(_02415_)
  );
  INV_X1 _12678_ (
    .A(_02415_),
    .ZN(_02416_)
  );
  AND2_X1 _12679_ (
    .A1(divisor[0]),
    .A2(remainder[1]),
    .ZN(_02417_)
  );
  INV_X1 _12680_ (
    .A(_02417_),
    .ZN(_02418_)
  );
  AND2_X1 _12681_ (
    .A1(_02251_),
    .A2(_02415_),
    .ZN(_02419_)
  );
  INV_X1 _12682_ (
    .A(_02419_),
    .ZN(_02420_)
  );
  AND2_X1 _12683_ (
    .A1(divisor[2]),
    .A2(remainder[0]),
    .ZN(_02421_)
  );
  INV_X1 _12684_ (
    .A(_02421_),
    .ZN(_02422_)
  );
  AND2_X1 _12685_ (
    .A1(_02252_),
    .A2(_02416_),
    .ZN(_02423_)
  );
  INV_X1 _12686_ (
    .A(_02423_),
    .ZN(_02424_)
  );
  AND2_X1 _12687_ (
    .A1(_02420_),
    .A2(_02424_),
    .ZN(_02425_)
  );
  INV_X1 _12688_ (
    .A(_02425_),
    .ZN(_02426_)
  );
  AND2_X1 _12689_ (
    .A1(_02421_),
    .A2(_02425_),
    .ZN(_02427_)
  );
  INV_X1 _12690_ (
    .A(_02427_),
    .ZN(_02428_)
  );
  AND2_X1 _12691_ (
    .A1(_02420_),
    .A2(_02428_),
    .ZN(_02429_)
  );
  INV_X1 _12692_ (
    .A(_02429_),
    .ZN(_02430_)
  );
  AND2_X1 _12693_ (
    .A1(_02256_),
    .A2(_02260_),
    .ZN(_02431_)
  );
  INV_X1 _12694_ (
    .A(_02431_),
    .ZN(_02432_)
  );
  AND2_X1 _12695_ (
    .A1(_02262_),
    .A2(_02432_),
    .ZN(_02433_)
  );
  INV_X1 _12696_ (
    .A(_02433_),
    .ZN(_02434_)
  );
  AND2_X1 _12697_ (
    .A1(_02430_),
    .A2(_02433_),
    .ZN(_02435_)
  );
  INV_X1 _12698_ (
    .A(_02435_),
    .ZN(_02436_)
  );
  AND2_X1 _12699_ (
    .A1(_02263_),
    .A2(_02268_),
    .ZN(_02437_)
  );
  INV_X1 _12700_ (
    .A(_02437_),
    .ZN(_02438_)
  );
  AND2_X1 _12701_ (
    .A1(_02270_),
    .A2(_02438_),
    .ZN(_02439_)
  );
  INV_X1 _12702_ (
    .A(_02439_),
    .ZN(_02440_)
  );
  AND2_X1 _12703_ (
    .A1(_02435_),
    .A2(_02439_),
    .ZN(_02441_)
  );
  INV_X1 _12704_ (
    .A(_02441_),
    .ZN(_02442_)
  );
  AND2_X1 _12705_ (
    .A1(divisor[3]),
    .A2(remainder[1]),
    .ZN(_02443_)
  );
  INV_X1 _12706_ (
    .A(_02443_),
    .ZN(_02444_)
  );
  AND2_X1 _12707_ (
    .A1(_02436_),
    .A2(_02440_),
    .ZN(_02445_)
  );
  INV_X1 _12708_ (
    .A(_02445_),
    .ZN(_02446_)
  );
  AND2_X1 _12709_ (
    .A1(_02442_),
    .A2(_02446_),
    .ZN(_02447_)
  );
  INV_X1 _12710_ (
    .A(_02447_),
    .ZN(_02448_)
  );
  AND2_X1 _12711_ (
    .A1(_02443_),
    .A2(_02447_),
    .ZN(_02449_)
  );
  INV_X1 _12712_ (
    .A(_02449_),
    .ZN(_02450_)
  );
  AND2_X1 _12713_ (
    .A1(_02442_),
    .A2(_02450_),
    .ZN(_02451_)
  );
  INV_X1 _12714_ (
    .A(_02451_),
    .ZN(_02452_)
  );
  AND2_X1 _12715_ (
    .A1(_02413_),
    .A2(_02452_),
    .ZN(_02453_)
  );
  INV_X1 _12716_ (
    .A(_02453_),
    .ZN(_02454_)
  );
  AND2_X1 _12717_ (
    .A1(_02409_),
    .A2(_02453_),
    .ZN(_02455_)
  );
  INV_X1 _12718_ (
    .A(_02455_),
    .ZN(_02456_)
  );
  AND2_X1 _12719_ (
    .A1(_02414_),
    .A2(_02451_),
    .ZN(_02457_)
  );
  INV_X1 _12720_ (
    .A(_02457_),
    .ZN(_02458_)
  );
  AND2_X1 _12721_ (
    .A1(_02454_),
    .A2(_02458_),
    .ZN(_02459_)
  );
  INV_X1 _12722_ (
    .A(_02459_),
    .ZN(_02460_)
  );
  AND2_X1 _12723_ (
    .A1(_02444_),
    .A2(_02448_),
    .ZN(_02461_)
  );
  INV_X1 _12724_ (
    .A(_02461_),
    .ZN(_02462_)
  );
  AND2_X1 _12725_ (
    .A1(_02450_),
    .A2(_02462_),
    .ZN(_02463_)
  );
  INV_X1 _12726_ (
    .A(_02463_),
    .ZN(_02464_)
  );
  AND2_X1 _12727_ (
    .A1(divisor[1]),
    .A2(remainder[0]),
    .ZN(_02465_)
  );
  INV_X1 _12728_ (
    .A(_02465_),
    .ZN(_02466_)
  );
  AND2_X1 _12729_ (
    .A1(divisor[0]),
    .A2(remainder[0]),
    .ZN(_02467_)
  );
  INV_X1 _12730_ (
    .A(_02467_),
    .ZN(_02468_)
  );
  AND2_X1 _12731_ (
    .A1(_02415_),
    .A2(_02467_),
    .ZN(_02469_)
  );
  INV_X1 _12732_ (
    .A(_02469_),
    .ZN(_02470_)
  );
  AND2_X1 _12733_ (
    .A1(_02422_),
    .A2(_02426_),
    .ZN(_02471_)
  );
  INV_X1 _12734_ (
    .A(_02471_),
    .ZN(_02472_)
  );
  AND2_X1 _12735_ (
    .A1(_02428_),
    .A2(_02472_),
    .ZN(_02473_)
  );
  INV_X1 _12736_ (
    .A(_02473_),
    .ZN(_02474_)
  );
  AND2_X1 _12737_ (
    .A1(_02469_),
    .A2(_02473_),
    .ZN(_02475_)
  );
  INV_X1 _12738_ (
    .A(_02475_),
    .ZN(_02476_)
  );
  AND2_X1 _12739_ (
    .A1(_02429_),
    .A2(_02434_),
    .ZN(_02477_)
  );
  INV_X1 _12740_ (
    .A(_02477_),
    .ZN(_02478_)
  );
  AND2_X1 _12741_ (
    .A1(_02436_),
    .A2(_02478_),
    .ZN(_02479_)
  );
  INV_X1 _12742_ (
    .A(_02479_),
    .ZN(_02480_)
  );
  AND2_X1 _12743_ (
    .A1(_02475_),
    .A2(_02479_),
    .ZN(_02481_)
  );
  INV_X1 _12744_ (
    .A(_02481_),
    .ZN(_02482_)
  );
  AND2_X1 _12745_ (
    .A1(_02476_),
    .A2(_02480_),
    .ZN(_02483_)
  );
  INV_X1 _12746_ (
    .A(_02483_),
    .ZN(_02484_)
  );
  AND2_X1 _12747_ (
    .A1(_02482_),
    .A2(_02484_),
    .ZN(_02485_)
  );
  INV_X1 _12748_ (
    .A(_02485_),
    .ZN(_02486_)
  );
  AND2_X1 _12749_ (
    .A1(_02377_),
    .A2(_02485_),
    .ZN(_02487_)
  );
  INV_X1 _12750_ (
    .A(_02487_),
    .ZN(_02488_)
  );
  AND2_X1 _12751_ (
    .A1(_02482_),
    .A2(_02488_),
    .ZN(_02489_)
  );
  INV_X1 _12752_ (
    .A(_02489_),
    .ZN(_02490_)
  );
  AND2_X1 _12753_ (
    .A1(_02463_),
    .A2(_02490_),
    .ZN(_02491_)
  );
  INV_X1 _12754_ (
    .A(_02491_),
    .ZN(_02492_)
  );
  AND2_X1 _12755_ (
    .A1(_02459_),
    .A2(_02491_),
    .ZN(_02493_)
  );
  INV_X1 _12756_ (
    .A(_02493_),
    .ZN(_02494_)
  );
  AND2_X1 _12757_ (
    .A1(_02410_),
    .A2(_02454_),
    .ZN(_02495_)
  );
  INV_X1 _12758_ (
    .A(_02495_),
    .ZN(_02496_)
  );
  AND2_X1 _12759_ (
    .A1(_02456_),
    .A2(_02496_),
    .ZN(_02497_)
  );
  INV_X1 _12760_ (
    .A(_02497_),
    .ZN(_02498_)
  );
  AND2_X1 _12761_ (
    .A1(_02493_),
    .A2(_02497_),
    .ZN(_02499_)
  );
  INV_X1 _12762_ (
    .A(_02499_),
    .ZN(_02500_)
  );
  AND2_X1 _12763_ (
    .A1(_02456_),
    .A2(_02500_),
    .ZN(_02501_)
  );
  INV_X1 _12764_ (
    .A(_02501_),
    .ZN(_02502_)
  );
  AND2_X1 _12765_ (
    .A1(_02405_),
    .A2(_02502_),
    .ZN(_02503_)
  );
  INV_X1 _12766_ (
    .A(_02503_),
    .ZN(_02504_)
  );
  AND2_X1 _12767_ (
    .A1(_02406_),
    .A2(_02501_),
    .ZN(_02505_)
  );
  INV_X1 _12768_ (
    .A(_02505_),
    .ZN(_02506_)
  );
  AND2_X1 _12769_ (
    .A1(_02504_),
    .A2(_02506_),
    .ZN(_02507_)
  );
  INV_X1 _12770_ (
    .A(_02507_),
    .ZN(_02508_)
  );
  AND2_X1 _12771_ (
    .A1(remainder[40]),
    .A2(_02507_),
    .ZN(_02509_)
  );
  INV_X1 _12772_ (
    .A(_02509_),
    .ZN(_02510_)
  );
  AND2_X1 _12773_ (
    .A1(_02494_),
    .A2(_02498_),
    .ZN(_02511_)
  );
  INV_X1 _12774_ (
    .A(_02511_),
    .ZN(_02512_)
  );
  AND2_X1 _12775_ (
    .A1(_02500_),
    .A2(_02512_),
    .ZN(_02513_)
  );
  INV_X1 _12776_ (
    .A(_02513_),
    .ZN(_02514_)
  );
  AND2_X1 _12777_ (
    .A1(remainder[39]),
    .A2(_02513_),
    .ZN(_02515_)
  );
  INV_X1 _12778_ (
    .A(_02515_),
    .ZN(_02516_)
  );
  AND2_X1 _12779_ (
    .A1(_02460_),
    .A2(_02492_),
    .ZN(_02517_)
  );
  INV_X1 _12780_ (
    .A(_02517_),
    .ZN(_02518_)
  );
  AND2_X1 _12781_ (
    .A1(_02494_),
    .A2(_02518_),
    .ZN(_02519_)
  );
  INV_X1 _12782_ (
    .A(_02519_),
    .ZN(_02520_)
  );
  AND2_X1 _12783_ (
    .A1(remainder[38]),
    .A2(_02519_),
    .ZN(_02521_)
  );
  INV_X1 _12784_ (
    .A(_02521_),
    .ZN(_02522_)
  );
  AND2_X1 _12785_ (
    .A1(_04700_),
    .A2(_02520_),
    .ZN(_02523_)
  );
  INV_X1 _12786_ (
    .A(_02523_),
    .ZN(_02524_)
  );
  AND2_X1 _12787_ (
    .A1(_02522_),
    .A2(_02524_),
    .ZN(_02525_)
  );
  INV_X1 _12788_ (
    .A(_02525_),
    .ZN(_02526_)
  );
  AND2_X1 _12789_ (
    .A1(_02464_),
    .A2(_02489_),
    .ZN(_02527_)
  );
  INV_X1 _12790_ (
    .A(_02527_),
    .ZN(_02528_)
  );
  AND2_X1 _12791_ (
    .A1(_02492_),
    .A2(_02528_),
    .ZN(_02529_)
  );
  INV_X1 _12792_ (
    .A(_02529_),
    .ZN(_02530_)
  );
  AND2_X1 _12793_ (
    .A1(remainder[37]),
    .A2(_02529_),
    .ZN(_02531_)
  );
  INV_X1 _12794_ (
    .A(_02531_),
    .ZN(_02532_)
  );
  AND2_X1 _12795_ (
    .A1(_04711_),
    .A2(_02530_),
    .ZN(_02533_)
  );
  INV_X1 _12796_ (
    .A(_02533_),
    .ZN(_02534_)
  );
  AND2_X1 _12797_ (
    .A1(_02532_),
    .A2(_02534_),
    .ZN(_02535_)
  );
  INV_X1 _12798_ (
    .A(_02535_),
    .ZN(_02536_)
  );
  AND2_X1 _12799_ (
    .A1(_02378_),
    .A2(_02486_),
    .ZN(_02537_)
  );
  INV_X1 _12800_ (
    .A(_02537_),
    .ZN(_02538_)
  );
  AND2_X1 _12801_ (
    .A1(_02488_),
    .A2(_02538_),
    .ZN(_02539_)
  );
  INV_X1 _12802_ (
    .A(_02539_),
    .ZN(_02540_)
  );
  AND2_X1 _12803_ (
    .A1(remainder[36]),
    .A2(_02539_),
    .ZN(_02541_)
  );
  INV_X1 _12804_ (
    .A(_02541_),
    .ZN(_02542_)
  );
  AND2_X1 _12805_ (
    .A1(_04722_),
    .A2(_02540_),
    .ZN(_02543_)
  );
  INV_X1 _12806_ (
    .A(_02543_),
    .ZN(_02544_)
  );
  AND2_X1 _12807_ (
    .A1(_02470_),
    .A2(_02474_),
    .ZN(_02545_)
  );
  INV_X1 _12808_ (
    .A(_02545_),
    .ZN(_02546_)
  );
  AND2_X1 _12809_ (
    .A1(_02476_),
    .A2(_02546_),
    .ZN(_02547_)
  );
  INV_X1 _12810_ (
    .A(_02547_),
    .ZN(_02548_)
  );
  AND2_X1 _12811_ (
    .A1(remainder[35]),
    .A2(_02547_),
    .ZN(_02549_)
  );
  INV_X1 _12812_ (
    .A(_02549_),
    .ZN(_02550_)
  );
  AND2_X1 _12813_ (
    .A1(_02418_),
    .A2(_02466_),
    .ZN(_02551_)
  );
  INV_X1 _12814_ (
    .A(_02551_),
    .ZN(_02552_)
  );
  AND2_X1 _12815_ (
    .A1(_02470_),
    .A2(_02552_),
    .ZN(_02553_)
  );
  INV_X1 _12816_ (
    .A(_02553_),
    .ZN(_02554_)
  );
  AND2_X1 _12817_ (
    .A1(remainder[34]),
    .A2(_02553_),
    .ZN(_02555_)
  );
  INV_X1 _12818_ (
    .A(_02555_),
    .ZN(_02556_)
  );
  AND2_X1 _12819_ (
    .A1(remainder[33]),
    .A2(_02467_),
    .ZN(_02557_)
  );
  INV_X1 _12820_ (
    .A(_02557_),
    .ZN(_02558_)
  );
  AND2_X1 _12821_ (
    .A1(_04744_),
    .A2(_02554_),
    .ZN(_02559_)
  );
  INV_X1 _12822_ (
    .A(_02559_),
    .ZN(_02560_)
  );
  AND2_X1 _12823_ (
    .A1(_02556_),
    .A2(_02560_),
    .ZN(_02561_)
  );
  INV_X1 _12824_ (
    .A(_02561_),
    .ZN(_02562_)
  );
  AND2_X1 _12825_ (
    .A1(_02557_),
    .A2(_02561_),
    .ZN(_02563_)
  );
  INV_X1 _12826_ (
    .A(_02563_),
    .ZN(_02564_)
  );
  AND2_X1 _12827_ (
    .A1(_02556_),
    .A2(_02564_),
    .ZN(_02565_)
  );
  INV_X1 _12828_ (
    .A(_02565_),
    .ZN(_02566_)
  );
  AND2_X1 _12829_ (
    .A1(_04733_),
    .A2(_02548_),
    .ZN(_02567_)
  );
  INV_X1 _12830_ (
    .A(_02567_),
    .ZN(_02568_)
  );
  AND2_X1 _12831_ (
    .A1(_02550_),
    .A2(_02568_),
    .ZN(_02569_)
  );
  INV_X1 _12832_ (
    .A(_02569_),
    .ZN(_02570_)
  );
  AND2_X1 _12833_ (
    .A1(_02566_),
    .A2(_02569_),
    .ZN(_02571_)
  );
  INV_X1 _12834_ (
    .A(_02571_),
    .ZN(_02572_)
  );
  AND2_X1 _12835_ (
    .A1(_02550_),
    .A2(_02572_),
    .ZN(_02573_)
  );
  INV_X1 _12836_ (
    .A(_02573_),
    .ZN(_02574_)
  );
  AND2_X1 _12837_ (
    .A1(_02544_),
    .A2(_02574_),
    .ZN(_02575_)
  );
  INV_X1 _12838_ (
    .A(_02575_),
    .ZN(_02576_)
  );
  AND2_X1 _12839_ (
    .A1(_02542_),
    .A2(_02573_),
    .ZN(_02577_)
  );
  INV_X1 _12840_ (
    .A(_02577_),
    .ZN(_02578_)
  );
  AND2_X1 _12841_ (
    .A1(_02542_),
    .A2(_02576_),
    .ZN(_02579_)
  );
  AND2_X1 _12842_ (
    .A1(_02544_),
    .A2(_02578_),
    .ZN(_02580_)
  );
  AND2_X1 _12843_ (
    .A1(_02535_),
    .A2(_02580_),
    .ZN(_02581_)
  );
  INV_X1 _12844_ (
    .A(_02581_),
    .ZN(_02582_)
  );
  AND2_X1 _12845_ (
    .A1(_02532_),
    .A2(_02582_),
    .ZN(_02583_)
  );
  INV_X1 _12846_ (
    .A(_02583_),
    .ZN(_02584_)
  );
  AND2_X1 _12847_ (
    .A1(_02525_),
    .A2(_02584_),
    .ZN(_02585_)
  );
  INV_X1 _12848_ (
    .A(_02585_),
    .ZN(_02586_)
  );
  AND2_X1 _12849_ (
    .A1(_02522_),
    .A2(_02586_),
    .ZN(_02587_)
  );
  INV_X1 _12850_ (
    .A(_02587_),
    .ZN(_02588_)
  );
  AND2_X1 _12851_ (
    .A1(_04689_),
    .A2(_02514_),
    .ZN(_02589_)
  );
  INV_X1 _12852_ (
    .A(_02589_),
    .ZN(_02590_)
  );
  AND2_X1 _12853_ (
    .A1(_02516_),
    .A2(_02590_),
    .ZN(_02591_)
  );
  INV_X1 _12854_ (
    .A(_02591_),
    .ZN(_02592_)
  );
  AND2_X1 _12855_ (
    .A1(_02588_),
    .A2(_02591_),
    .ZN(_02593_)
  );
  INV_X1 _12856_ (
    .A(_02593_),
    .ZN(_02594_)
  );
  AND2_X1 _12857_ (
    .A1(_02516_),
    .A2(_02594_),
    .ZN(_02595_)
  );
  INV_X1 _12858_ (
    .A(_02595_),
    .ZN(_02596_)
  );
  AND2_X1 _12859_ (
    .A1(_04678_),
    .A2(_02508_),
    .ZN(_02597_)
  );
  INV_X1 _12860_ (
    .A(_02597_),
    .ZN(_02598_)
  );
  AND2_X1 _12861_ (
    .A1(_02510_),
    .A2(_02598_),
    .ZN(_02599_)
  );
  INV_X1 _12862_ (
    .A(_02599_),
    .ZN(_02600_)
  );
  AND2_X1 _12863_ (
    .A1(_02596_),
    .A2(_02599_),
    .ZN(_02601_)
  );
  INV_X1 _12864_ (
    .A(_02601_),
    .ZN(_02602_)
  );
  AND2_X1 _12865_ (
    .A1(_02510_),
    .A2(_02602_),
    .ZN(_02603_)
  );
  INV_X1 _12866_ (
    .A(_02603_),
    .ZN(_02604_)
  );
  AND2_X1 _12867_ (
    .A1(divisor[3]),
    .A2(remainder[5]),
    .ZN(_02605_)
  );
  INV_X1 _12868_ (
    .A(_02605_),
    .ZN(_02606_)
  );
  AND2_X1 _12869_ (
    .A1(divisor[8]),
    .A2(remainder[0]),
    .ZN(_02607_)
  );
  INV_X1 _12870_ (
    .A(_02607_),
    .ZN(_02608_)
  );
  AND2_X1 _12871_ (
    .A1(divisor[7]),
    .A2(remainder[1]),
    .ZN(_02609_)
  );
  INV_X1 _12872_ (
    .A(_02609_),
    .ZN(_02610_)
  );
  AND2_X1 _12873_ (
    .A1(divisor[8]),
    .A2(remainder[1]),
    .ZN(_02611_)
  );
  INV_X1 _12874_ (
    .A(_02611_),
    .ZN(_02612_)
  );
  AND2_X1 _12875_ (
    .A1(_02373_),
    .A2(_02611_),
    .ZN(_02613_)
  );
  INV_X1 _12876_ (
    .A(_02613_),
    .ZN(_02614_)
  );
  AND2_X1 _12877_ (
    .A1(_02608_),
    .A2(_02610_),
    .ZN(_02615_)
  );
  INV_X1 _12878_ (
    .A(_02615_),
    .ZN(_02616_)
  );
  AND2_X1 _12879_ (
    .A1(_02614_),
    .A2(_02616_),
    .ZN(_02617_)
  );
  INV_X1 _12880_ (
    .A(_02617_),
    .ZN(_02618_)
  );
  AND2_X1 _12881_ (
    .A1(_02605_),
    .A2(_02617_),
    .ZN(_02619_)
  );
  INV_X1 _12882_ (
    .A(_02619_),
    .ZN(_02620_)
  );
  AND2_X1 _12883_ (
    .A1(_02606_),
    .A2(_02618_),
    .ZN(_02621_)
  );
  INV_X1 _12884_ (
    .A(_02621_),
    .ZN(_02622_)
  );
  AND2_X1 _12885_ (
    .A1(_02620_),
    .A2(_02622_),
    .ZN(_02623_)
  );
  INV_X1 _12886_ (
    .A(_02623_),
    .ZN(_02624_)
  );
  AND2_X1 _12887_ (
    .A1(_02381_),
    .A2(_02623_),
    .ZN(_02625_)
  );
  INV_X1 _12888_ (
    .A(_02625_),
    .ZN(_02626_)
  );
  AND2_X1 _12889_ (
    .A1(_02382_),
    .A2(_02624_),
    .ZN(_02627_)
  );
  INV_X1 _12890_ (
    .A(_02627_),
    .ZN(_02628_)
  );
  AND2_X1 _12891_ (
    .A1(_02626_),
    .A2(_02628_),
    .ZN(_02629_)
  );
  INV_X1 _12892_ (
    .A(_02629_),
    .ZN(_02630_)
  );
  AND2_X1 _12893_ (
    .A1(_02225_),
    .A2(_02347_),
    .ZN(_02631_)
  );
  INV_X1 _12894_ (
    .A(_02631_),
    .ZN(_02632_)
  );
  AND2_X1 _12895_ (
    .A1(_02362_),
    .A2(_02632_),
    .ZN(_02633_)
  );
  INV_X1 _12896_ (
    .A(_02633_),
    .ZN(_02634_)
  );
  AND2_X1 _12897_ (
    .A1(_02300_),
    .A2(_02306_),
    .ZN(_02635_)
  );
  INV_X1 _12898_ (
    .A(_02635_),
    .ZN(_02636_)
  );
  AND2_X1 _12899_ (
    .A1(_02219_),
    .A2(_02347_),
    .ZN(_02637_)
  );
  INV_X1 _12900_ (
    .A(_02637_),
    .ZN(_02638_)
  );
  AND2_X1 _12901_ (
    .A1(_02332_),
    .A2(_02338_),
    .ZN(_02639_)
  );
  INV_X1 _12902_ (
    .A(_02639_),
    .ZN(_02640_)
  );
  AND2_X1 _12903_ (
    .A1(_02320_),
    .A2(_02326_),
    .ZN(_02641_)
  );
  INV_X1 _12904_ (
    .A(_02641_),
    .ZN(_02642_)
  );
  AND2_X1 _12905_ (
    .A1(divisor[4]),
    .A2(remainder[4]),
    .ZN(_02643_)
  );
  INV_X1 _12906_ (
    .A(_02643_),
    .ZN(_02644_)
  );
  AND2_X1 _12907_ (
    .A1(divisor[5]),
    .A2(remainder[3]),
    .ZN(_02645_)
  );
  INV_X1 _12908_ (
    .A(_02645_),
    .ZN(_02646_)
  );
  AND2_X1 _12909_ (
    .A1(divisor[6]),
    .A2(remainder[3]),
    .ZN(_02647_)
  );
  INV_X1 _12910_ (
    .A(_02647_),
    .ZN(_02648_)
  );
  AND2_X1 _12911_ (
    .A1(_02317_),
    .A2(_02645_),
    .ZN(_02649_)
  );
  INV_X1 _12912_ (
    .A(_02649_),
    .ZN(_02650_)
  );
  AND2_X1 _12913_ (
    .A1(_02318_),
    .A2(_02646_),
    .ZN(_02651_)
  );
  INV_X1 _12914_ (
    .A(_02651_),
    .ZN(_02652_)
  );
  AND2_X1 _12915_ (
    .A1(_02650_),
    .A2(_02652_),
    .ZN(_02653_)
  );
  INV_X1 _12916_ (
    .A(_02653_),
    .ZN(_02654_)
  );
  AND2_X1 _12917_ (
    .A1(_02643_),
    .A2(_02653_),
    .ZN(_02655_)
  );
  INV_X1 _12918_ (
    .A(_02655_),
    .ZN(_02656_)
  );
  AND2_X1 _12919_ (
    .A1(_02644_),
    .A2(_02654_),
    .ZN(_02657_)
  );
  INV_X1 _12920_ (
    .A(_02657_),
    .ZN(_02658_)
  );
  AND2_X1 _12921_ (
    .A1(_02656_),
    .A2(_02658_),
    .ZN(_02659_)
  );
  INV_X1 _12922_ (
    .A(_02659_),
    .ZN(_02660_)
  );
  AND2_X1 _12923_ (
    .A1(_02642_),
    .A2(_02659_),
    .ZN(_02661_)
  );
  INV_X1 _12924_ (
    .A(_02661_),
    .ZN(_02662_)
  );
  AND2_X1 _12925_ (
    .A1(_02641_),
    .A2(_02660_),
    .ZN(_02663_)
  );
  INV_X1 _12926_ (
    .A(_02663_),
    .ZN(_02664_)
  );
  AND2_X1 _12927_ (
    .A1(_02662_),
    .A2(_02664_),
    .ZN(_02665_)
  );
  INV_X1 _12928_ (
    .A(_02665_),
    .ZN(_02666_)
  );
  AND2_X1 _12929_ (
    .A1(divisor[2]),
    .A2(remainder[6]),
    .ZN(_02667_)
  );
  INV_X1 _12930_ (
    .A(_02667_),
    .ZN(_02668_)
  );
  AND2_X1 _12931_ (
    .A1(remainder[32]),
    .A2(divisor[1]),
    .ZN(_02669_)
  );
  AND2_X1 _12932_ (
    .A1(remainder[32]),
    .A2(divisor[0]),
    .ZN(_02670_)
  );
  INV_X1 _12933_ (
    .A(_02670_),
    .ZN(_02671_)
  );
  AND2_X1 _12934_ (
    .A1(divisor[1]),
    .A2(_02670_),
    .ZN(_02672_)
  );
  INV_X1 _12935_ (
    .A(_02672_),
    .ZN(_02673_)
  );
  AND2_X1 _12936_ (
    .A1(_02297_),
    .A2(_02670_),
    .ZN(_02674_)
  );
  INV_X1 _12937_ (
    .A(_02674_),
    .ZN(_02675_)
  );
  AND2_X1 _12938_ (
    .A1(_02298_),
    .A2(_02671_),
    .ZN(_02676_)
  );
  INV_X1 _12939_ (
    .A(_02676_),
    .ZN(_02677_)
  );
  AND2_X1 _12940_ (
    .A1(_02675_),
    .A2(_02677_),
    .ZN(_02678_)
  );
  INV_X1 _12941_ (
    .A(_02678_),
    .ZN(_02679_)
  );
  AND2_X1 _12942_ (
    .A1(_02667_),
    .A2(_02678_),
    .ZN(_02680_)
  );
  INV_X1 _12943_ (
    .A(_02680_),
    .ZN(_02681_)
  );
  AND2_X1 _12944_ (
    .A1(_02668_),
    .A2(_02679_),
    .ZN(_02682_)
  );
  INV_X1 _12945_ (
    .A(_02682_),
    .ZN(_02683_)
  );
  AND2_X1 _12946_ (
    .A1(_02681_),
    .A2(_02683_),
    .ZN(_02684_)
  );
  INV_X1 _12947_ (
    .A(_02684_),
    .ZN(_02685_)
  );
  AND2_X1 _12948_ (
    .A1(_02665_),
    .A2(_02684_),
    .ZN(_02686_)
  );
  INV_X1 _12949_ (
    .A(_02686_),
    .ZN(_02687_)
  );
  AND2_X1 _12950_ (
    .A1(_02666_),
    .A2(_02685_),
    .ZN(_02688_)
  );
  INV_X1 _12951_ (
    .A(_02688_),
    .ZN(_02689_)
  );
  AND2_X1 _12952_ (
    .A1(_02687_),
    .A2(_02689_),
    .ZN(_02690_)
  );
  INV_X1 _12953_ (
    .A(_02690_),
    .ZN(_02691_)
  );
  AND2_X1 _12954_ (
    .A1(_02640_),
    .A2(_02690_),
    .ZN(_02692_)
  );
  INV_X1 _12955_ (
    .A(_02692_),
    .ZN(_02693_)
  );
  AND2_X1 _12956_ (
    .A1(_02639_),
    .A2(_02691_),
    .ZN(_02694_)
  );
  INV_X1 _12957_ (
    .A(_02694_),
    .ZN(_02695_)
  );
  AND2_X1 _12958_ (
    .A1(_02693_),
    .A2(_02695_),
    .ZN(_02696_)
  );
  INV_X1 _12959_ (
    .A(_02696_),
    .ZN(_02697_)
  );
  AND2_X1 _12960_ (
    .A1(_02343_),
    .A2(_02696_),
    .ZN(_02698_)
  );
  INV_X1 _12961_ (
    .A(_02698_),
    .ZN(_02699_)
  );
  AND2_X1 _12962_ (
    .A1(_02344_),
    .A2(_02697_),
    .ZN(_02700_)
  );
  INV_X1 _12963_ (
    .A(_02700_),
    .ZN(_02701_)
  );
  AND2_X1 _12964_ (
    .A1(_02699_),
    .A2(_02701_),
    .ZN(_02702_)
  );
  INV_X1 _12965_ (
    .A(_02702_),
    .ZN(_02703_)
  );
  AND2_X1 _12966_ (
    .A1(_02637_),
    .A2(_02702_),
    .ZN(_02704_)
  );
  INV_X1 _12967_ (
    .A(_02704_),
    .ZN(_02705_)
  );
  AND2_X1 _12968_ (
    .A1(_02638_),
    .A2(_02703_),
    .ZN(_02706_)
  );
  INV_X1 _12969_ (
    .A(_02706_),
    .ZN(_02707_)
  );
  AND2_X1 _12970_ (
    .A1(_02705_),
    .A2(_02707_),
    .ZN(_02708_)
  );
  INV_X1 _12971_ (
    .A(_02708_),
    .ZN(_02709_)
  );
  AND2_X1 _12972_ (
    .A1(_02636_),
    .A2(_02708_),
    .ZN(_02710_)
  );
  INV_X1 _12973_ (
    .A(_02710_),
    .ZN(_02711_)
  );
  AND2_X1 _12974_ (
    .A1(_02635_),
    .A2(_02709_),
    .ZN(_02712_)
  );
  INV_X1 _12975_ (
    .A(_02712_),
    .ZN(_02713_)
  );
  AND2_X1 _12976_ (
    .A1(_02711_),
    .A2(_02713_),
    .ZN(_02714_)
  );
  INV_X1 _12977_ (
    .A(_02714_),
    .ZN(_02715_)
  );
  AND2_X1 _12978_ (
    .A1(_02634_),
    .A2(_02714_),
    .ZN(_02716_)
  );
  INV_X1 _12979_ (
    .A(_02716_),
    .ZN(_02717_)
  );
  AND2_X1 _12980_ (
    .A1(_02633_),
    .A2(_02715_),
    .ZN(_02718_)
  );
  INV_X1 _12981_ (
    .A(_02718_),
    .ZN(_02719_)
  );
  AND2_X1 _12982_ (
    .A1(_02717_),
    .A2(_02719_),
    .ZN(_02720_)
  );
  INV_X1 _12983_ (
    .A(_02720_),
    .ZN(_02721_)
  );
  AND2_X1 _12984_ (
    .A1(_02629_),
    .A2(_02720_),
    .ZN(_02722_)
  );
  INV_X1 _12985_ (
    .A(_02722_),
    .ZN(_02723_)
  );
  AND2_X1 _12986_ (
    .A1(_02630_),
    .A2(_02721_),
    .ZN(_02724_)
  );
  INV_X1 _12987_ (
    .A(_02724_),
    .ZN(_02725_)
  );
  AND2_X1 _12988_ (
    .A1(_02723_),
    .A2(_02725_),
    .ZN(_02726_)
  );
  INV_X1 _12989_ (
    .A(_02726_),
    .ZN(_02727_)
  );
  AND2_X1 _12990_ (
    .A1(_02368_),
    .A2(_02388_),
    .ZN(_02728_)
  );
  INV_X1 _12991_ (
    .A(_02728_),
    .ZN(_02729_)
  );
  AND2_X1 _12992_ (
    .A1(_02726_),
    .A2(_02729_),
    .ZN(_02730_)
  );
  INV_X1 _12993_ (
    .A(_02730_),
    .ZN(_02731_)
  );
  AND2_X1 _12994_ (
    .A1(_02727_),
    .A2(_02728_),
    .ZN(_02732_)
  );
  INV_X1 _12995_ (
    .A(_02732_),
    .ZN(_02733_)
  );
  AND2_X1 _12996_ (
    .A1(_02731_),
    .A2(_02733_),
    .ZN(_02734_)
  );
  AND2_X1 _12997_ (
    .A1(_02401_),
    .A2(_02734_),
    .ZN(_02735_)
  );
  INV_X1 _12998_ (
    .A(_02735_),
    .ZN(_02736_)
  );
  AND2_X1 _12999_ (
    .A1(_02395_),
    .A2(_02734_),
    .ZN(_02737_)
  );
  INV_X1 _13000_ (
    .A(_02737_),
    .ZN(_02738_)
  );
  AND2_X1 _13001_ (
    .A1(_02396_),
    .A2(_02402_),
    .ZN(_02739_)
  );
  INV_X1 _13002_ (
    .A(_02739_),
    .ZN(_02740_)
  );
  MUX2_X1 _13003_ (
    .A(_02740_),
    .B(_02396_),
    .S(_02734_),
    .Z(_02741_)
  );
  AND2_X1 _13004_ (
    .A1(_02736_),
    .A2(_02741_),
    .ZN(_02742_)
  );
  INV_X1 _13005_ (
    .A(_02742_),
    .ZN(_02743_)
  );
  AND2_X1 _13006_ (
    .A1(_02503_),
    .A2(_02742_),
    .ZN(_02744_)
  );
  INV_X1 _13007_ (
    .A(_02744_),
    .ZN(_02745_)
  );
  AND2_X1 _13008_ (
    .A1(_02504_),
    .A2(_02743_),
    .ZN(_02746_)
  );
  INV_X1 _13009_ (
    .A(_02746_),
    .ZN(_02747_)
  );
  AND2_X1 _13010_ (
    .A1(_02745_),
    .A2(_02747_),
    .ZN(_02748_)
  );
  INV_X1 _13011_ (
    .A(_02748_),
    .ZN(_02749_)
  );
  AND2_X1 _13012_ (
    .A1(remainder[41]),
    .A2(_02748_),
    .ZN(_02750_)
  );
  INV_X1 _13013_ (
    .A(_02750_),
    .ZN(_02751_)
  );
  AND2_X1 _13014_ (
    .A1(_04667_),
    .A2(_02749_),
    .ZN(_02752_)
  );
  INV_X1 _13015_ (
    .A(_02752_),
    .ZN(_02753_)
  );
  AND2_X1 _13016_ (
    .A1(_02751_),
    .A2(_02753_),
    .ZN(_02754_)
  );
  INV_X1 _13017_ (
    .A(_02754_),
    .ZN(_02755_)
  );
  AND2_X1 _13018_ (
    .A1(_02603_),
    .A2(_02755_),
    .ZN(_02756_)
  );
  INV_X1 _13019_ (
    .A(_02756_),
    .ZN(_02757_)
  );
  AND2_X1 _13020_ (
    .A1(_02604_),
    .A2(_02754_),
    .ZN(_02758_)
  );
  INV_X1 _13021_ (
    .A(_02758_),
    .ZN(_02759_)
  );
  AND2_X1 _13022_ (
    .A1(_02082_),
    .A2(_02757_),
    .ZN(_02760_)
  );
  AND2_X1 _13023_ (
    .A1(_02759_),
    .A2(_02760_),
    .ZN(_02761_)
  );
  INV_X1 _13024_ (
    .A(_02761_),
    .ZN(_02762_)
  );
  AND2_X1 _13025_ (
    .A1(_02094_),
    .A2(_02762_),
    .ZN(_02763_)
  );
  AND2_X1 _13026_ (
    .A1(_02092_),
    .A2(_02763_),
    .ZN(_02764_)
  );
  INV_X1 _13027_ (
    .A(_02764_),
    .ZN(_02765_)
  );
  AND2_X1 _13028_ (
    .A1(_06201_),
    .A2(_02765_),
    .ZN(_00054_)
  );
  AND2_X1 _13029_ (
    .A1(_04755_),
    .A2(_10451_),
    .ZN(_02766_)
  );
  INV_X1 _13030_ (
    .A(_02766_),
    .ZN(_02767_)
  );
  AND2_X1 _13031_ (
    .A1(_10462_),
    .A2(_00404_),
    .ZN(_02768_)
  );
  INV_X1 _13032_ (
    .A(_02768_),
    .ZN(_02769_)
  );
  AND2_X1 _13033_ (
    .A1(_05983_),
    .A2(_02769_),
    .ZN(_02770_)
  );
  AND2_X1 _13034_ (
    .A1(_02767_),
    .A2(_02770_),
    .ZN(_02771_)
  );
  INV_X1 _13035_ (
    .A(_02771_),
    .ZN(_02772_)
  );
  AND2_X1 _13036_ (
    .A1(remainder[34]),
    .A2(_02077_),
    .ZN(_02773_)
  );
  INV_X1 _13037_ (
    .A(_02773_),
    .ZN(_02774_)
  );
  AND2_X1 _13038_ (
    .A1(_02751_),
    .A2(_02759_),
    .ZN(_02775_)
  );
  INV_X1 _13039_ (
    .A(_02775_),
    .ZN(_02776_)
  );
  AND2_X1 _13040_ (
    .A1(_02736_),
    .A2(_02745_),
    .ZN(_02777_)
  );
  INV_X1 _13041_ (
    .A(_02777_),
    .ZN(_02778_)
  );
  AND2_X1 _13042_ (
    .A1(_02626_),
    .A2(_02723_),
    .ZN(_02779_)
  );
  INV_X1 _13043_ (
    .A(_02779_),
    .ZN(_02780_)
  );
  AND2_X1 _13044_ (
    .A1(divisor[3]),
    .A2(remainder[6]),
    .ZN(_02781_)
  );
  INV_X1 _13045_ (
    .A(_02781_),
    .ZN(_02782_)
  );
  AND2_X1 _13046_ (
    .A1(divisor[7]),
    .A2(remainder[2]),
    .ZN(_02783_)
  );
  INV_X1 _13047_ (
    .A(_02783_),
    .ZN(_02784_)
  );
  AND2_X1 _13048_ (
    .A1(divisor[9]),
    .A2(remainder[0]),
    .ZN(_02785_)
  );
  INV_X1 _13049_ (
    .A(_02785_),
    .ZN(_02786_)
  );
  AND2_X1 _13050_ (
    .A1(divisor[9]),
    .A2(remainder[1]),
    .ZN(_02787_)
  );
  INV_X1 _13051_ (
    .A(_02787_),
    .ZN(_02788_)
  );
  AND2_X1 _13052_ (
    .A1(_02607_),
    .A2(_02787_),
    .ZN(_02789_)
  );
  INV_X1 _13053_ (
    .A(_02789_),
    .ZN(_02790_)
  );
  AND2_X1 _13054_ (
    .A1(_02612_),
    .A2(_02786_),
    .ZN(_02791_)
  );
  INV_X1 _13055_ (
    .A(_02791_),
    .ZN(_02792_)
  );
  AND2_X1 _13056_ (
    .A1(_02790_),
    .A2(_02792_),
    .ZN(_02793_)
  );
  INV_X1 _13057_ (
    .A(_02793_),
    .ZN(_02794_)
  );
  AND2_X1 _13058_ (
    .A1(_02783_),
    .A2(_02793_),
    .ZN(_02795_)
  );
  INV_X1 _13059_ (
    .A(_02795_),
    .ZN(_02796_)
  );
  AND2_X1 _13060_ (
    .A1(_02784_),
    .A2(_02794_),
    .ZN(_02797_)
  );
  INV_X1 _13061_ (
    .A(_02797_),
    .ZN(_02798_)
  );
  AND2_X1 _13062_ (
    .A1(_02796_),
    .A2(_02798_),
    .ZN(_02799_)
  );
  INV_X1 _13063_ (
    .A(_02799_),
    .ZN(_02800_)
  );
  AND2_X1 _13064_ (
    .A1(_02613_),
    .A2(_02799_),
    .ZN(_02801_)
  );
  INV_X1 _13065_ (
    .A(_02801_),
    .ZN(_02802_)
  );
  AND2_X1 _13066_ (
    .A1(_02614_),
    .A2(_02800_),
    .ZN(_02803_)
  );
  INV_X1 _13067_ (
    .A(_02803_),
    .ZN(_02804_)
  );
  AND2_X1 _13068_ (
    .A1(_02802_),
    .A2(_02804_),
    .ZN(_02805_)
  );
  INV_X1 _13069_ (
    .A(_02805_),
    .ZN(_02806_)
  );
  AND2_X1 _13070_ (
    .A1(_02781_),
    .A2(_02805_),
    .ZN(_02807_)
  );
  INV_X1 _13071_ (
    .A(_02807_),
    .ZN(_02808_)
  );
  AND2_X1 _13072_ (
    .A1(_02782_),
    .A2(_02806_),
    .ZN(_02809_)
  );
  INV_X1 _13073_ (
    .A(_02809_),
    .ZN(_02810_)
  );
  AND2_X1 _13074_ (
    .A1(_02808_),
    .A2(_02810_),
    .ZN(_02811_)
  );
  INV_X1 _13075_ (
    .A(_02811_),
    .ZN(_02812_)
  );
  AND2_X1 _13076_ (
    .A1(_02619_),
    .A2(_02811_),
    .ZN(_02813_)
  );
  INV_X1 _13077_ (
    .A(_02813_),
    .ZN(_02814_)
  );
  AND2_X1 _13078_ (
    .A1(_02620_),
    .A2(_02812_),
    .ZN(_02815_)
  );
  INV_X1 _13079_ (
    .A(_02815_),
    .ZN(_02816_)
  );
  AND2_X1 _13080_ (
    .A1(_02814_),
    .A2(_02816_),
    .ZN(_02817_)
  );
  INV_X1 _13081_ (
    .A(_02817_),
    .ZN(_02818_)
  );
  AND2_X1 _13082_ (
    .A1(_02705_),
    .A2(_02711_),
    .ZN(_02819_)
  );
  INV_X1 _13083_ (
    .A(_02819_),
    .ZN(_02820_)
  );
  AND2_X1 _13084_ (
    .A1(_02675_),
    .A2(_02681_),
    .ZN(_02821_)
  );
  INV_X1 _13085_ (
    .A(_02821_),
    .ZN(_02822_)
  );
  AND2_X1 _13086_ (
    .A1(_02662_),
    .A2(_02687_),
    .ZN(_02823_)
  );
  INV_X1 _13087_ (
    .A(_02823_),
    .ZN(_02824_)
  );
  AND2_X1 _13088_ (
    .A1(_02650_),
    .A2(_02656_),
    .ZN(_02825_)
  );
  INV_X1 _13089_ (
    .A(_02825_),
    .ZN(_02826_)
  );
  AND2_X1 _13090_ (
    .A1(divisor[4]),
    .A2(remainder[5]),
    .ZN(_02827_)
  );
  INV_X1 _13091_ (
    .A(_02827_),
    .ZN(_02828_)
  );
  AND2_X1 _13092_ (
    .A1(divisor[5]),
    .A2(remainder[4]),
    .ZN(_02829_)
  );
  INV_X1 _13093_ (
    .A(_02829_),
    .ZN(_02830_)
  );
  AND2_X1 _13094_ (
    .A1(divisor[6]),
    .A2(remainder[4]),
    .ZN(_02831_)
  );
  INV_X1 _13095_ (
    .A(_02831_),
    .ZN(_02832_)
  );
  AND2_X1 _13096_ (
    .A1(_02647_),
    .A2(_02829_),
    .ZN(_02833_)
  );
  INV_X1 _13097_ (
    .A(_02833_),
    .ZN(_02834_)
  );
  AND2_X1 _13098_ (
    .A1(_02648_),
    .A2(_02830_),
    .ZN(_02835_)
  );
  INV_X1 _13099_ (
    .A(_02835_),
    .ZN(_02836_)
  );
  AND2_X1 _13100_ (
    .A1(_02834_),
    .A2(_02836_),
    .ZN(_02837_)
  );
  INV_X1 _13101_ (
    .A(_02837_),
    .ZN(_02838_)
  );
  AND2_X1 _13102_ (
    .A1(_02827_),
    .A2(_02837_),
    .ZN(_02839_)
  );
  INV_X1 _13103_ (
    .A(_02839_),
    .ZN(_02840_)
  );
  AND2_X1 _13104_ (
    .A1(_02828_),
    .A2(_02838_),
    .ZN(_02841_)
  );
  INV_X1 _13105_ (
    .A(_02841_),
    .ZN(_02842_)
  );
  AND2_X1 _13106_ (
    .A1(_02840_),
    .A2(_02842_),
    .ZN(_02843_)
  );
  INV_X1 _13107_ (
    .A(_02843_),
    .ZN(_02844_)
  );
  AND2_X1 _13108_ (
    .A1(_02826_),
    .A2(_02843_),
    .ZN(_02845_)
  );
  INV_X1 _13109_ (
    .A(_02845_),
    .ZN(_02846_)
  );
  AND2_X1 _13110_ (
    .A1(_02825_),
    .A2(_02844_),
    .ZN(_02847_)
  );
  INV_X1 _13111_ (
    .A(_02847_),
    .ZN(_02848_)
  );
  AND2_X1 _13112_ (
    .A1(_02846_),
    .A2(_02848_),
    .ZN(_02849_)
  );
  INV_X1 _13113_ (
    .A(_02849_),
    .ZN(_02850_)
  );
  MUX2_X1 _13114_ (
    .A(_02670_),
    .B(_04853_),
    .S(_02669_),
    .Z(_02851_)
  );
  INV_X1 _13115_ (
    .A(_02851_),
    .ZN(_02852_)
  );
  AND2_X1 _13116_ (
    .A1(divisor[2]),
    .A2(remainder[7]),
    .ZN(_02853_)
  );
  INV_X1 _13117_ (
    .A(_02853_),
    .ZN(_02854_)
  );
  AND2_X1 _13118_ (
    .A1(divisor[2]),
    .A2(_02851_),
    .ZN(_02855_)
  );
  INV_X1 _13119_ (
    .A(_02855_),
    .ZN(_02856_)
  );
  AND2_X1 _13120_ (
    .A1(_02851_),
    .A2(_02853_),
    .ZN(_02857_)
  );
  INV_X1 _13121_ (
    .A(_02857_),
    .ZN(_02858_)
  );
  AND2_X1 _13122_ (
    .A1(_02852_),
    .A2(_02854_),
    .ZN(_02859_)
  );
  INV_X1 _13123_ (
    .A(_02859_),
    .ZN(_02860_)
  );
  AND2_X1 _13124_ (
    .A1(_02858_),
    .A2(_02860_),
    .ZN(_02861_)
  );
  INV_X1 _13125_ (
    .A(_02861_),
    .ZN(_02862_)
  );
  AND2_X1 _13126_ (
    .A1(_02849_),
    .A2(_02861_),
    .ZN(_02863_)
  );
  INV_X1 _13127_ (
    .A(_02863_),
    .ZN(_02864_)
  );
  AND2_X1 _13128_ (
    .A1(_02850_),
    .A2(_02862_),
    .ZN(_02865_)
  );
  INV_X1 _13129_ (
    .A(_02865_),
    .ZN(_02866_)
  );
  AND2_X1 _13130_ (
    .A1(_02864_),
    .A2(_02866_),
    .ZN(_02867_)
  );
  INV_X1 _13131_ (
    .A(_02867_),
    .ZN(_02868_)
  );
  AND2_X1 _13132_ (
    .A1(_02824_),
    .A2(_02867_),
    .ZN(_02869_)
  );
  INV_X1 _13133_ (
    .A(_02869_),
    .ZN(_02870_)
  );
  AND2_X1 _13134_ (
    .A1(_02823_),
    .A2(_02868_),
    .ZN(_02871_)
  );
  INV_X1 _13135_ (
    .A(_02871_),
    .ZN(_02872_)
  );
  AND2_X1 _13136_ (
    .A1(_02870_),
    .A2(_02872_),
    .ZN(_02873_)
  );
  INV_X1 _13137_ (
    .A(_02873_),
    .ZN(_02874_)
  );
  AND2_X1 _13138_ (
    .A1(_02692_),
    .A2(_02873_),
    .ZN(_02875_)
  );
  INV_X1 _13139_ (
    .A(_02875_),
    .ZN(_02876_)
  );
  AND2_X1 _13140_ (
    .A1(_02693_),
    .A2(_02874_),
    .ZN(_02877_)
  );
  INV_X1 _13141_ (
    .A(_02877_),
    .ZN(_02878_)
  );
  AND2_X1 _13142_ (
    .A1(_02876_),
    .A2(_02878_),
    .ZN(_02879_)
  );
  INV_X1 _13143_ (
    .A(_02879_),
    .ZN(_02880_)
  );
  AND2_X1 _13144_ (
    .A1(_02698_),
    .A2(_02879_),
    .ZN(_02881_)
  );
  INV_X1 _13145_ (
    .A(_02881_),
    .ZN(_02882_)
  );
  AND2_X1 _13146_ (
    .A1(_02699_),
    .A2(_02880_),
    .ZN(_02883_)
  );
  INV_X1 _13147_ (
    .A(_02883_),
    .ZN(_02884_)
  );
  AND2_X1 _13148_ (
    .A1(_02882_),
    .A2(_02884_),
    .ZN(_02885_)
  );
  INV_X1 _13149_ (
    .A(_02885_),
    .ZN(_02886_)
  );
  AND2_X1 _13150_ (
    .A1(_02822_),
    .A2(_02885_),
    .ZN(_02887_)
  );
  INV_X1 _13151_ (
    .A(_02887_),
    .ZN(_02888_)
  );
  AND2_X1 _13152_ (
    .A1(_02821_),
    .A2(_02886_),
    .ZN(_02889_)
  );
  INV_X1 _13153_ (
    .A(_02889_),
    .ZN(_02890_)
  );
  AND2_X1 _13154_ (
    .A1(_02888_),
    .A2(_02890_),
    .ZN(_02891_)
  );
  INV_X1 _13155_ (
    .A(_02891_),
    .ZN(_02892_)
  );
  AND2_X1 _13156_ (
    .A1(_02820_),
    .A2(_02891_),
    .ZN(_02893_)
  );
  INV_X1 _13157_ (
    .A(_02893_),
    .ZN(_02894_)
  );
  AND2_X1 _13158_ (
    .A1(_02819_),
    .A2(_02892_),
    .ZN(_02895_)
  );
  INV_X1 _13159_ (
    .A(_02895_),
    .ZN(_02896_)
  );
  AND2_X1 _13160_ (
    .A1(_02894_),
    .A2(_02896_),
    .ZN(_02897_)
  );
  INV_X1 _13161_ (
    .A(_02897_),
    .ZN(_02898_)
  );
  AND2_X1 _13162_ (
    .A1(_02817_),
    .A2(_02897_),
    .ZN(_02899_)
  );
  INV_X1 _13163_ (
    .A(_02899_),
    .ZN(_02900_)
  );
  AND2_X1 _13164_ (
    .A1(_02818_),
    .A2(_02898_),
    .ZN(_02901_)
  );
  INV_X1 _13165_ (
    .A(_02901_),
    .ZN(_02902_)
  );
  AND2_X1 _13166_ (
    .A1(_02900_),
    .A2(_02902_),
    .ZN(_02903_)
  );
  INV_X1 _13167_ (
    .A(_02903_),
    .ZN(_02904_)
  );
  AND2_X1 _13168_ (
    .A1(_02780_),
    .A2(_02903_),
    .ZN(_02905_)
  );
  INV_X1 _13169_ (
    .A(_02905_),
    .ZN(_02906_)
  );
  AND2_X1 _13170_ (
    .A1(_02779_),
    .A2(_02904_),
    .ZN(_02907_)
  );
  INV_X1 _13171_ (
    .A(_02907_),
    .ZN(_02908_)
  );
  AND2_X1 _13172_ (
    .A1(_02906_),
    .A2(_02908_),
    .ZN(_02909_)
  );
  INV_X1 _13173_ (
    .A(_02909_),
    .ZN(_02910_)
  );
  AND2_X1 _13174_ (
    .A1(_02716_),
    .A2(_02909_),
    .ZN(_02911_)
  );
  INV_X1 _13175_ (
    .A(_02911_),
    .ZN(_02912_)
  );
  AND2_X1 _13176_ (
    .A1(_02717_),
    .A2(_02910_),
    .ZN(_02913_)
  );
  INV_X1 _13177_ (
    .A(_02913_),
    .ZN(_02914_)
  );
  AND2_X1 _13178_ (
    .A1(_02912_),
    .A2(_02914_),
    .ZN(_02915_)
  );
  INV_X1 _13179_ (
    .A(_02915_),
    .ZN(_02916_)
  );
  AND2_X1 _13180_ (
    .A1(_02730_),
    .A2(_02915_),
    .ZN(_02917_)
  );
  INV_X1 _13181_ (
    .A(_02917_),
    .ZN(_02918_)
  );
  AND2_X1 _13182_ (
    .A1(_02731_),
    .A2(_02916_),
    .ZN(_02919_)
  );
  INV_X1 _13183_ (
    .A(_02919_),
    .ZN(_02920_)
  );
  AND2_X1 _13184_ (
    .A1(_02918_),
    .A2(_02920_),
    .ZN(_02921_)
  );
  INV_X1 _13185_ (
    .A(_02921_),
    .ZN(_02922_)
  );
  AND2_X1 _13186_ (
    .A1(_02738_),
    .A2(_02922_),
    .ZN(_02923_)
  );
  INV_X1 _13187_ (
    .A(_02923_),
    .ZN(_02924_)
  );
  AND2_X1 _13188_ (
    .A1(_02737_),
    .A2(_02921_),
    .ZN(_02925_)
  );
  INV_X1 _13189_ (
    .A(_02925_),
    .ZN(_02926_)
  );
  AND2_X1 _13190_ (
    .A1(_02924_),
    .A2(_02926_),
    .ZN(_02927_)
  );
  INV_X1 _13191_ (
    .A(_02927_),
    .ZN(_02928_)
  );
  AND2_X1 _13192_ (
    .A1(_02778_),
    .A2(_02924_),
    .ZN(_02929_)
  );
  INV_X1 _13193_ (
    .A(_02929_),
    .ZN(_02930_)
  );
  AND2_X1 _13194_ (
    .A1(_02777_),
    .A2(_02928_),
    .ZN(_02931_)
  );
  INV_X1 _13195_ (
    .A(_02931_),
    .ZN(_02932_)
  );
  AND2_X1 _13196_ (
    .A1(_02930_),
    .A2(_02932_),
    .ZN(_02933_)
  );
  INV_X1 _13197_ (
    .A(_02933_),
    .ZN(_02934_)
  );
  AND2_X1 _13198_ (
    .A1(remainder[42]),
    .A2(_02933_),
    .ZN(_02935_)
  );
  INV_X1 _13199_ (
    .A(_02935_),
    .ZN(_02936_)
  );
  AND2_X1 _13200_ (
    .A1(_04656_),
    .A2(_02934_),
    .ZN(_02937_)
  );
  INV_X1 _13201_ (
    .A(_02937_),
    .ZN(_02938_)
  );
  AND2_X1 _13202_ (
    .A1(_02936_),
    .A2(_02938_),
    .ZN(_02939_)
  );
  INV_X1 _13203_ (
    .A(_02939_),
    .ZN(_02940_)
  );
  AND2_X1 _13204_ (
    .A1(_02776_),
    .A2(_02939_),
    .ZN(_02941_)
  );
  INV_X1 _13205_ (
    .A(_02941_),
    .ZN(_02942_)
  );
  AND2_X1 _13206_ (
    .A1(_02775_),
    .A2(_02940_),
    .ZN(_02943_)
  );
  INV_X1 _13207_ (
    .A(_02943_),
    .ZN(_02944_)
  );
  AND2_X1 _13208_ (
    .A1(_02942_),
    .A2(_02944_),
    .ZN(_02945_)
  );
  AND2_X1 _13209_ (
    .A1(_02082_),
    .A2(_02945_),
    .ZN(_02946_)
  );
  INV_X1 _13210_ (
    .A(_02946_),
    .ZN(_02947_)
  );
  AND2_X1 _13211_ (
    .A1(_02774_),
    .A2(_02947_),
    .ZN(_02948_)
  );
  AND2_X1 _13212_ (
    .A1(_02772_),
    .A2(_02948_),
    .ZN(_02949_)
  );
  INV_X1 _13213_ (
    .A(_02949_),
    .ZN(_02950_)
  );
  AND2_X1 _13214_ (
    .A1(_06201_),
    .A2(_02950_),
    .ZN(_00055_)
  );
  AND2_X1 _13215_ (
    .A1(_04744_),
    .A2(_10451_),
    .ZN(_02951_)
  );
  INV_X1 _13216_ (
    .A(_02951_),
    .ZN(_02952_)
  );
  AND2_X1 _13217_ (
    .A1(_10462_),
    .A2(_00502_),
    .ZN(_02953_)
  );
  INV_X1 _13218_ (
    .A(_02953_),
    .ZN(_02954_)
  );
  AND2_X1 _13219_ (
    .A1(_05983_),
    .A2(_02954_),
    .ZN(_02955_)
  );
  AND2_X1 _13220_ (
    .A1(_02952_),
    .A2(_02955_),
    .ZN(_02956_)
  );
  INV_X1 _13221_ (
    .A(_02956_),
    .ZN(_02957_)
  );
  AND2_X1 _13222_ (
    .A1(remainder[35]),
    .A2(_02077_),
    .ZN(_02958_)
  );
  INV_X1 _13223_ (
    .A(_02958_),
    .ZN(_02959_)
  );
  AND2_X1 _13224_ (
    .A1(_02906_),
    .A2(_02912_),
    .ZN(_02960_)
  );
  INV_X1 _13225_ (
    .A(_02960_),
    .ZN(_02961_)
  );
  AND2_X1 _13226_ (
    .A1(_02814_),
    .A2(_02900_),
    .ZN(_02962_)
  );
  INV_X1 _13227_ (
    .A(_02962_),
    .ZN(_02963_)
  );
  AND2_X1 _13228_ (
    .A1(divisor[3]),
    .A2(remainder[7]),
    .ZN(_02964_)
  );
  INV_X1 _13229_ (
    .A(_02964_),
    .ZN(_02965_)
  );
  AND2_X1 _13230_ (
    .A1(divisor[10]),
    .A2(remainder[0]),
    .ZN(_02966_)
  );
  INV_X1 _13231_ (
    .A(_02966_),
    .ZN(_02967_)
  );
  AND2_X1 _13232_ (
    .A1(_02790_),
    .A2(_02796_),
    .ZN(_02968_)
  );
  INV_X1 _13233_ (
    .A(_02968_),
    .ZN(_02969_)
  );
  AND2_X1 _13234_ (
    .A1(divisor[7]),
    .A2(remainder[3]),
    .ZN(_02970_)
  );
  INV_X1 _13235_ (
    .A(_02970_),
    .ZN(_02971_)
  );
  AND2_X1 _13236_ (
    .A1(divisor[8]),
    .A2(remainder[2]),
    .ZN(_02972_)
  );
  INV_X1 _13237_ (
    .A(_02972_),
    .ZN(_02973_)
  );
  AND2_X1 _13238_ (
    .A1(divisor[9]),
    .A2(remainder[2]),
    .ZN(_02974_)
  );
  INV_X1 _13239_ (
    .A(_02974_),
    .ZN(_02975_)
  );
  AND2_X1 _13240_ (
    .A1(_02611_),
    .A2(_02974_),
    .ZN(_02976_)
  );
  INV_X1 _13241_ (
    .A(_02976_),
    .ZN(_02977_)
  );
  AND2_X1 _13242_ (
    .A1(_02788_),
    .A2(_02973_),
    .ZN(_02978_)
  );
  INV_X1 _13243_ (
    .A(_02978_),
    .ZN(_02979_)
  );
  AND2_X1 _13244_ (
    .A1(_02977_),
    .A2(_02979_),
    .ZN(_02980_)
  );
  INV_X1 _13245_ (
    .A(_02980_),
    .ZN(_02981_)
  );
  AND2_X1 _13246_ (
    .A1(_02970_),
    .A2(_02980_),
    .ZN(_02982_)
  );
  INV_X1 _13247_ (
    .A(_02982_),
    .ZN(_02983_)
  );
  AND2_X1 _13248_ (
    .A1(_02971_),
    .A2(_02981_),
    .ZN(_02984_)
  );
  INV_X1 _13249_ (
    .A(_02984_),
    .ZN(_02985_)
  );
  AND2_X1 _13250_ (
    .A1(_02983_),
    .A2(_02985_),
    .ZN(_02986_)
  );
  INV_X1 _13251_ (
    .A(_02986_),
    .ZN(_02987_)
  );
  AND2_X1 _13252_ (
    .A1(_02969_),
    .A2(_02986_),
    .ZN(_02988_)
  );
  INV_X1 _13253_ (
    .A(_02988_),
    .ZN(_02989_)
  );
  AND2_X1 _13254_ (
    .A1(_02968_),
    .A2(_02987_),
    .ZN(_02990_)
  );
  INV_X1 _13255_ (
    .A(_02990_),
    .ZN(_02991_)
  );
  AND2_X1 _13256_ (
    .A1(_02989_),
    .A2(_02991_),
    .ZN(_02992_)
  );
  INV_X1 _13257_ (
    .A(_02992_),
    .ZN(_02993_)
  );
  AND2_X1 _13258_ (
    .A1(_02966_),
    .A2(_02992_),
    .ZN(_02994_)
  );
  INV_X1 _13259_ (
    .A(_02994_),
    .ZN(_02995_)
  );
  AND2_X1 _13260_ (
    .A1(_02967_),
    .A2(_02993_),
    .ZN(_02996_)
  );
  INV_X1 _13261_ (
    .A(_02996_),
    .ZN(_02997_)
  );
  AND2_X1 _13262_ (
    .A1(_02995_),
    .A2(_02997_),
    .ZN(_02998_)
  );
  INV_X1 _13263_ (
    .A(_02998_),
    .ZN(_02999_)
  );
  AND2_X1 _13264_ (
    .A1(_02964_),
    .A2(_02998_),
    .ZN(_03000_)
  );
  INV_X1 _13265_ (
    .A(_03000_),
    .ZN(_03001_)
  );
  AND2_X1 _13266_ (
    .A1(_02965_),
    .A2(_02999_),
    .ZN(_03002_)
  );
  INV_X1 _13267_ (
    .A(_03002_),
    .ZN(_03003_)
  );
  AND2_X1 _13268_ (
    .A1(_03001_),
    .A2(_03003_),
    .ZN(_03004_)
  );
  INV_X1 _13269_ (
    .A(_03004_),
    .ZN(_03005_)
  );
  AND2_X1 _13270_ (
    .A1(_02807_),
    .A2(_03004_),
    .ZN(_03006_)
  );
  INV_X1 _13271_ (
    .A(_03006_),
    .ZN(_03007_)
  );
  AND2_X1 _13272_ (
    .A1(_02808_),
    .A2(_03005_),
    .ZN(_03008_)
  );
  INV_X1 _13273_ (
    .A(_03008_),
    .ZN(_03009_)
  );
  AND2_X1 _13274_ (
    .A1(_03007_),
    .A2(_03009_),
    .ZN(_03010_)
  );
  INV_X1 _13275_ (
    .A(_03010_),
    .ZN(_03011_)
  );
  AND2_X1 _13276_ (
    .A1(_02882_),
    .A2(_02888_),
    .ZN(_03012_)
  );
  INV_X1 _13277_ (
    .A(_03012_),
    .ZN(_03013_)
  );
  AND2_X1 _13278_ (
    .A1(_02673_),
    .A2(_02858_),
    .ZN(_03014_)
  );
  INV_X1 _13279_ (
    .A(_03014_),
    .ZN(_03015_)
  );
  AND2_X1 _13280_ (
    .A1(_02846_),
    .A2(_02864_),
    .ZN(_03016_)
  );
  INV_X1 _13281_ (
    .A(_03016_),
    .ZN(_03017_)
  );
  AND2_X1 _13282_ (
    .A1(_02834_),
    .A2(_02840_),
    .ZN(_03018_)
  );
  INV_X1 _13283_ (
    .A(_03018_),
    .ZN(_03019_)
  );
  AND2_X1 _13284_ (
    .A1(divisor[4]),
    .A2(remainder[6]),
    .ZN(_03020_)
  );
  INV_X1 _13285_ (
    .A(_03020_),
    .ZN(_03021_)
  );
  AND2_X1 _13286_ (
    .A1(divisor[5]),
    .A2(remainder[5]),
    .ZN(_03022_)
  );
  INV_X1 _13287_ (
    .A(_03022_),
    .ZN(_03023_)
  );
  AND2_X1 _13288_ (
    .A1(divisor[6]),
    .A2(remainder[5]),
    .ZN(_03024_)
  );
  INV_X1 _13289_ (
    .A(_03024_),
    .ZN(_03025_)
  );
  AND2_X1 _13290_ (
    .A1(_02831_),
    .A2(_03022_),
    .ZN(_03026_)
  );
  INV_X1 _13291_ (
    .A(_03026_),
    .ZN(_03027_)
  );
  AND2_X1 _13292_ (
    .A1(_02832_),
    .A2(_03023_),
    .ZN(_03028_)
  );
  INV_X1 _13293_ (
    .A(_03028_),
    .ZN(_03029_)
  );
  AND2_X1 _13294_ (
    .A1(_03027_),
    .A2(_03029_),
    .ZN(_03030_)
  );
  INV_X1 _13295_ (
    .A(_03030_),
    .ZN(_03031_)
  );
  AND2_X1 _13296_ (
    .A1(_03020_),
    .A2(_03030_),
    .ZN(_03032_)
  );
  INV_X1 _13297_ (
    .A(_03032_),
    .ZN(_03033_)
  );
  AND2_X1 _13298_ (
    .A1(_03021_),
    .A2(_03031_),
    .ZN(_03034_)
  );
  INV_X1 _13299_ (
    .A(_03034_),
    .ZN(_03035_)
  );
  AND2_X1 _13300_ (
    .A1(_03033_),
    .A2(_03035_),
    .ZN(_03036_)
  );
  INV_X1 _13301_ (
    .A(_03036_),
    .ZN(_03037_)
  );
  AND2_X1 _13302_ (
    .A1(_03019_),
    .A2(_03036_),
    .ZN(_03038_)
  );
  INV_X1 _13303_ (
    .A(_03038_),
    .ZN(_03039_)
  );
  AND2_X1 _13304_ (
    .A1(_03018_),
    .A2(_03037_),
    .ZN(_03040_)
  );
  INV_X1 _13305_ (
    .A(_03040_),
    .ZN(_03041_)
  );
  AND2_X1 _13306_ (
    .A1(_03039_),
    .A2(_03041_),
    .ZN(_03042_)
  );
  INV_X1 _13307_ (
    .A(_03042_),
    .ZN(_03043_)
  );
  AND2_X1 _13308_ (
    .A1(remainder[32]),
    .A2(divisor[2]),
    .ZN(_03044_)
  );
  INV_X1 _13309_ (
    .A(_03044_),
    .ZN(_03045_)
  );
  MUX2_X1 _13310_ (
    .A(_03044_),
    .B(_04864_),
    .S(_02851_),
    .Z(_03046_)
  );
  MUX2_X1 _13311_ (
    .A(_03045_),
    .B(divisor[2]),
    .S(_02851_),
    .Z(_03047_)
  );
  AND2_X1 _13312_ (
    .A1(_03042_),
    .A2(_03046_),
    .ZN(_03048_)
  );
  INV_X1 _13313_ (
    .A(_03048_),
    .ZN(_03049_)
  );
  AND2_X1 _13314_ (
    .A1(_03043_),
    .A2(_03047_),
    .ZN(_03050_)
  );
  INV_X1 _13315_ (
    .A(_03050_),
    .ZN(_03051_)
  );
  AND2_X1 _13316_ (
    .A1(_03049_),
    .A2(_03051_),
    .ZN(_03052_)
  );
  INV_X1 _13317_ (
    .A(_03052_),
    .ZN(_03053_)
  );
  AND2_X1 _13318_ (
    .A1(_02801_),
    .A2(_03052_),
    .ZN(_03054_)
  );
  INV_X1 _13319_ (
    .A(_03054_),
    .ZN(_03055_)
  );
  AND2_X1 _13320_ (
    .A1(_02802_),
    .A2(_03053_),
    .ZN(_03056_)
  );
  INV_X1 _13321_ (
    .A(_03056_),
    .ZN(_03057_)
  );
  AND2_X1 _13322_ (
    .A1(_03055_),
    .A2(_03057_),
    .ZN(_03058_)
  );
  INV_X1 _13323_ (
    .A(_03058_),
    .ZN(_03059_)
  );
  AND2_X1 _13324_ (
    .A1(_03017_),
    .A2(_03058_),
    .ZN(_03060_)
  );
  INV_X1 _13325_ (
    .A(_03060_),
    .ZN(_03061_)
  );
  AND2_X1 _13326_ (
    .A1(_03016_),
    .A2(_03059_),
    .ZN(_03062_)
  );
  INV_X1 _13327_ (
    .A(_03062_),
    .ZN(_03063_)
  );
  AND2_X1 _13328_ (
    .A1(_03061_),
    .A2(_03063_),
    .ZN(_03064_)
  );
  INV_X1 _13329_ (
    .A(_03064_),
    .ZN(_03065_)
  );
  AND2_X1 _13330_ (
    .A1(_02869_),
    .A2(_03064_),
    .ZN(_03066_)
  );
  INV_X1 _13331_ (
    .A(_03066_),
    .ZN(_03067_)
  );
  AND2_X1 _13332_ (
    .A1(_02870_),
    .A2(_03065_),
    .ZN(_03068_)
  );
  INV_X1 _13333_ (
    .A(_03068_),
    .ZN(_03069_)
  );
  AND2_X1 _13334_ (
    .A1(_03067_),
    .A2(_03069_),
    .ZN(_03070_)
  );
  INV_X1 _13335_ (
    .A(_03070_),
    .ZN(_03071_)
  );
  AND2_X1 _13336_ (
    .A1(_02875_),
    .A2(_03070_),
    .ZN(_03072_)
  );
  INV_X1 _13337_ (
    .A(_03072_),
    .ZN(_03073_)
  );
  AND2_X1 _13338_ (
    .A1(_02876_),
    .A2(_03071_),
    .ZN(_03074_)
  );
  INV_X1 _13339_ (
    .A(_03074_),
    .ZN(_03075_)
  );
  AND2_X1 _13340_ (
    .A1(_03073_),
    .A2(_03075_),
    .ZN(_03076_)
  );
  INV_X1 _13341_ (
    .A(_03076_),
    .ZN(_03077_)
  );
  AND2_X1 _13342_ (
    .A1(_03015_),
    .A2(_03076_),
    .ZN(_03078_)
  );
  INV_X1 _13343_ (
    .A(_03078_),
    .ZN(_03079_)
  );
  AND2_X1 _13344_ (
    .A1(_03014_),
    .A2(_03077_),
    .ZN(_03080_)
  );
  INV_X1 _13345_ (
    .A(_03080_),
    .ZN(_03081_)
  );
  AND2_X1 _13346_ (
    .A1(_03079_),
    .A2(_03081_),
    .ZN(_03082_)
  );
  INV_X1 _13347_ (
    .A(_03082_),
    .ZN(_03083_)
  );
  AND2_X1 _13348_ (
    .A1(_03013_),
    .A2(_03082_),
    .ZN(_03084_)
  );
  INV_X1 _13349_ (
    .A(_03084_),
    .ZN(_03085_)
  );
  AND2_X1 _13350_ (
    .A1(_03012_),
    .A2(_03083_),
    .ZN(_03086_)
  );
  INV_X1 _13351_ (
    .A(_03086_),
    .ZN(_03087_)
  );
  AND2_X1 _13352_ (
    .A1(_03085_),
    .A2(_03087_),
    .ZN(_03088_)
  );
  INV_X1 _13353_ (
    .A(_03088_),
    .ZN(_03089_)
  );
  AND2_X1 _13354_ (
    .A1(_03010_),
    .A2(_03088_),
    .ZN(_03090_)
  );
  INV_X1 _13355_ (
    .A(_03090_),
    .ZN(_03091_)
  );
  AND2_X1 _13356_ (
    .A1(_03011_),
    .A2(_03089_),
    .ZN(_03092_)
  );
  INV_X1 _13357_ (
    .A(_03092_),
    .ZN(_03093_)
  );
  AND2_X1 _13358_ (
    .A1(_03091_),
    .A2(_03093_),
    .ZN(_03094_)
  );
  INV_X1 _13359_ (
    .A(_03094_),
    .ZN(_03095_)
  );
  AND2_X1 _13360_ (
    .A1(_02963_),
    .A2(_03094_),
    .ZN(_03096_)
  );
  INV_X1 _13361_ (
    .A(_03096_),
    .ZN(_03097_)
  );
  AND2_X1 _13362_ (
    .A1(_02962_),
    .A2(_03095_),
    .ZN(_03098_)
  );
  INV_X1 _13363_ (
    .A(_03098_),
    .ZN(_03099_)
  );
  AND2_X1 _13364_ (
    .A1(_03097_),
    .A2(_03099_),
    .ZN(_03100_)
  );
  INV_X1 _13365_ (
    .A(_03100_),
    .ZN(_03101_)
  );
  AND2_X1 _13366_ (
    .A1(_02893_),
    .A2(_03100_),
    .ZN(_03102_)
  );
  INV_X1 _13367_ (
    .A(_03102_),
    .ZN(_03103_)
  );
  AND2_X1 _13368_ (
    .A1(_02894_),
    .A2(_03101_),
    .ZN(_03104_)
  );
  INV_X1 _13369_ (
    .A(_03104_),
    .ZN(_03105_)
  );
  AND2_X1 _13370_ (
    .A1(_03103_),
    .A2(_03105_),
    .ZN(_03106_)
  );
  INV_X1 _13371_ (
    .A(_03106_),
    .ZN(_03107_)
  );
  AND2_X1 _13372_ (
    .A1(_02961_),
    .A2(_03106_),
    .ZN(_03108_)
  );
  INV_X1 _13373_ (
    .A(_03108_),
    .ZN(_03109_)
  );
  AND2_X1 _13374_ (
    .A1(_02960_),
    .A2(_03107_),
    .ZN(_03110_)
  );
  INV_X1 _13375_ (
    .A(_03110_),
    .ZN(_03111_)
  );
  AND2_X1 _13376_ (
    .A1(_03109_),
    .A2(_03111_),
    .ZN(_03112_)
  );
  INV_X1 _13377_ (
    .A(_03112_),
    .ZN(_03113_)
  );
  AND2_X1 _13378_ (
    .A1(_02917_),
    .A2(_03112_),
    .ZN(_03114_)
  );
  INV_X1 _13379_ (
    .A(_03114_),
    .ZN(_03115_)
  );
  AND2_X1 _13380_ (
    .A1(_02918_),
    .A2(_03113_),
    .ZN(_03116_)
  );
  INV_X1 _13381_ (
    .A(_03116_),
    .ZN(_03117_)
  );
  AND2_X1 _13382_ (
    .A1(_03115_),
    .A2(_03117_),
    .ZN(_03118_)
  );
  INV_X1 _13383_ (
    .A(_03118_),
    .ZN(_03119_)
  );
  AND2_X1 _13384_ (
    .A1(_02926_),
    .A2(_02930_),
    .ZN(_03120_)
  );
  INV_X1 _13385_ (
    .A(_03120_),
    .ZN(_03121_)
  );
  AND2_X1 _13386_ (
    .A1(_03118_),
    .A2(_03121_),
    .ZN(_03122_)
  );
  INV_X1 _13387_ (
    .A(_03122_),
    .ZN(_03123_)
  );
  AND2_X1 _13388_ (
    .A1(_03119_),
    .A2(_03120_),
    .ZN(_03124_)
  );
  INV_X1 _13389_ (
    .A(_03124_),
    .ZN(_03125_)
  );
  AND2_X1 _13390_ (
    .A1(_03123_),
    .A2(_03125_),
    .ZN(_03126_)
  );
  INV_X1 _13391_ (
    .A(_03126_),
    .ZN(_03127_)
  );
  AND2_X1 _13392_ (
    .A1(remainder[43]),
    .A2(_03126_),
    .ZN(_03128_)
  );
  INV_X1 _13393_ (
    .A(_03128_),
    .ZN(_03129_)
  );
  AND2_X1 _13394_ (
    .A1(_04645_),
    .A2(_03127_),
    .ZN(_03130_)
  );
  INV_X1 _13395_ (
    .A(_03130_),
    .ZN(_03131_)
  );
  AND2_X1 _13396_ (
    .A1(_03129_),
    .A2(_03131_),
    .ZN(_03132_)
  );
  INV_X1 _13397_ (
    .A(_03132_),
    .ZN(_03133_)
  );
  AND2_X1 _13398_ (
    .A1(_02775_),
    .A2(_02936_),
    .ZN(_03134_)
  );
  INV_X1 _13399_ (
    .A(_03134_),
    .ZN(_03135_)
  );
  AND2_X1 _13400_ (
    .A1(_02776_),
    .A2(_02938_),
    .ZN(_03136_)
  );
  INV_X1 _13401_ (
    .A(_03136_),
    .ZN(_03137_)
  );
  AND2_X1 _13402_ (
    .A1(_02938_),
    .A2(_03135_),
    .ZN(_03138_)
  );
  AND2_X1 _13403_ (
    .A1(_02936_),
    .A2(_03137_),
    .ZN(_03139_)
  );
  AND2_X1 _13404_ (
    .A1(_03132_),
    .A2(_03138_),
    .ZN(_03140_)
  );
  INV_X1 _13405_ (
    .A(_03140_),
    .ZN(_03141_)
  );
  AND2_X1 _13406_ (
    .A1(_03133_),
    .A2(_03139_),
    .ZN(_03142_)
  );
  INV_X1 _13407_ (
    .A(_03142_),
    .ZN(_03143_)
  );
  AND2_X1 _13408_ (
    .A1(_02082_),
    .A2(_03141_),
    .ZN(_03144_)
  );
  AND2_X1 _13409_ (
    .A1(_03143_),
    .A2(_03144_),
    .ZN(_03145_)
  );
  INV_X1 _13410_ (
    .A(_03145_),
    .ZN(_03146_)
  );
  AND2_X1 _13411_ (
    .A1(_02959_),
    .A2(_03146_),
    .ZN(_03147_)
  );
  AND2_X1 _13412_ (
    .A1(_02957_),
    .A2(_03147_),
    .ZN(_03148_)
  );
  INV_X1 _13413_ (
    .A(_03148_),
    .ZN(_03149_)
  );
  AND2_X1 _13414_ (
    .A1(_06201_),
    .A2(_03149_),
    .ZN(_00056_)
  );
  AND2_X1 _13415_ (
    .A1(_10462_),
    .A2(_00731_),
    .ZN(_03150_)
  );
  INV_X1 _13416_ (
    .A(_03150_),
    .ZN(_03151_)
  );
  AND2_X1 _13417_ (
    .A1(_04733_),
    .A2(_10451_),
    .ZN(_03152_)
  );
  INV_X1 _13418_ (
    .A(_03152_),
    .ZN(_03153_)
  );
  AND2_X1 _13419_ (
    .A1(_05983_),
    .A2(_03151_),
    .ZN(_03154_)
  );
  AND2_X1 _13420_ (
    .A1(_03153_),
    .A2(_03154_),
    .ZN(_03155_)
  );
  INV_X1 _13421_ (
    .A(_03155_),
    .ZN(_03156_)
  );
  AND2_X1 _13422_ (
    .A1(remainder[36]),
    .A2(_02077_),
    .ZN(_03157_)
  );
  INV_X1 _13423_ (
    .A(_03157_),
    .ZN(_03158_)
  );
  AND2_X1 _13424_ (
    .A1(_03129_),
    .A2(_03141_),
    .ZN(_03159_)
  );
  INV_X1 _13425_ (
    .A(_03159_),
    .ZN(_03160_)
  );
  AND2_X1 _13426_ (
    .A1(_03115_),
    .A2(_03123_),
    .ZN(_03161_)
  );
  INV_X1 _13427_ (
    .A(_03161_),
    .ZN(_03162_)
  );
  AND2_X1 _13428_ (
    .A1(_03097_),
    .A2(_03103_),
    .ZN(_03163_)
  );
  INV_X1 _13429_ (
    .A(_03163_),
    .ZN(_03164_)
  );
  AND2_X1 _13430_ (
    .A1(_03007_),
    .A2(_03091_),
    .ZN(_03165_)
  );
  INV_X1 _13431_ (
    .A(_03165_),
    .ZN(_03166_)
  );
  AND2_X1 _13432_ (
    .A1(_03073_),
    .A2(_03079_),
    .ZN(_03167_)
  );
  INV_X1 _13433_ (
    .A(_03167_),
    .ZN(_03168_)
  );
  AND2_X1 _13434_ (
    .A1(_02673_),
    .A2(_02856_),
    .ZN(_03169_)
  );
  INV_X1 _13435_ (
    .A(_03169_),
    .ZN(_03170_)
  );
  AND2_X1 _13436_ (
    .A1(_03055_),
    .A2(_03061_),
    .ZN(_03171_)
  );
  INV_X1 _13437_ (
    .A(_03171_),
    .ZN(_03172_)
  );
  AND2_X1 _13438_ (
    .A1(_03039_),
    .A2(_03049_),
    .ZN(_03173_)
  );
  INV_X1 _13439_ (
    .A(_03173_),
    .ZN(_03174_)
  );
  AND2_X1 _13440_ (
    .A1(_03027_),
    .A2(_03033_),
    .ZN(_03175_)
  );
  INV_X1 _13441_ (
    .A(_03175_),
    .ZN(_03176_)
  );
  AND2_X1 _13442_ (
    .A1(divisor[4]),
    .A2(remainder[7]),
    .ZN(_03177_)
  );
  INV_X1 _13443_ (
    .A(_03177_),
    .ZN(_03178_)
  );
  AND2_X1 _13444_ (
    .A1(divisor[5]),
    .A2(remainder[6]),
    .ZN(_03179_)
  );
  INV_X1 _13445_ (
    .A(_03179_),
    .ZN(_03180_)
  );
  AND2_X1 _13446_ (
    .A1(divisor[6]),
    .A2(remainder[6]),
    .ZN(_03181_)
  );
  INV_X1 _13447_ (
    .A(_03181_),
    .ZN(_03182_)
  );
  AND2_X1 _13448_ (
    .A1(_03024_),
    .A2(_03179_),
    .ZN(_03183_)
  );
  INV_X1 _13449_ (
    .A(_03183_),
    .ZN(_03184_)
  );
  AND2_X1 _13450_ (
    .A1(_03025_),
    .A2(_03180_),
    .ZN(_03185_)
  );
  INV_X1 _13451_ (
    .A(_03185_),
    .ZN(_03186_)
  );
  AND2_X1 _13452_ (
    .A1(_03184_),
    .A2(_03186_),
    .ZN(_03187_)
  );
  INV_X1 _13453_ (
    .A(_03187_),
    .ZN(_03188_)
  );
  AND2_X1 _13454_ (
    .A1(_03177_),
    .A2(_03187_),
    .ZN(_03189_)
  );
  INV_X1 _13455_ (
    .A(_03189_),
    .ZN(_03190_)
  );
  AND2_X1 _13456_ (
    .A1(_03178_),
    .A2(_03188_),
    .ZN(_03191_)
  );
  INV_X1 _13457_ (
    .A(_03191_),
    .ZN(_03192_)
  );
  AND2_X1 _13458_ (
    .A1(_03190_),
    .A2(_03192_),
    .ZN(_03193_)
  );
  INV_X1 _13459_ (
    .A(_03193_),
    .ZN(_03194_)
  );
  AND2_X1 _13460_ (
    .A1(_03176_),
    .A2(_03193_),
    .ZN(_03195_)
  );
  INV_X1 _13461_ (
    .A(_03195_),
    .ZN(_03196_)
  );
  AND2_X1 _13462_ (
    .A1(_03175_),
    .A2(_03194_),
    .ZN(_03197_)
  );
  INV_X1 _13463_ (
    .A(_03197_),
    .ZN(_03198_)
  );
  AND2_X1 _13464_ (
    .A1(_03196_),
    .A2(_03198_),
    .ZN(_03199_)
  );
  INV_X1 _13465_ (
    .A(_03199_),
    .ZN(_03200_)
  );
  AND2_X1 _13466_ (
    .A1(_03046_),
    .A2(_03199_),
    .ZN(_03201_)
  );
  INV_X1 _13467_ (
    .A(_03201_),
    .ZN(_03202_)
  );
  AND2_X1 _13468_ (
    .A1(_03047_),
    .A2(_03200_),
    .ZN(_03203_)
  );
  INV_X1 _13469_ (
    .A(_03203_),
    .ZN(_03204_)
  );
  AND2_X1 _13470_ (
    .A1(_03202_),
    .A2(_03204_),
    .ZN(_03205_)
  );
  INV_X1 _13471_ (
    .A(_03205_),
    .ZN(_03206_)
  );
  AND2_X1 _13472_ (
    .A1(_02988_),
    .A2(_03205_),
    .ZN(_03207_)
  );
  INV_X1 _13473_ (
    .A(_03207_),
    .ZN(_03208_)
  );
  AND2_X1 _13474_ (
    .A1(_02989_),
    .A2(_03206_),
    .ZN(_03209_)
  );
  INV_X1 _13475_ (
    .A(_03209_),
    .ZN(_03210_)
  );
  AND2_X1 _13476_ (
    .A1(_03208_),
    .A2(_03210_),
    .ZN(_03211_)
  );
  INV_X1 _13477_ (
    .A(_03211_),
    .ZN(_03212_)
  );
  AND2_X1 _13478_ (
    .A1(_03174_),
    .A2(_03211_),
    .ZN(_03213_)
  );
  INV_X1 _13479_ (
    .A(_03213_),
    .ZN(_03214_)
  );
  AND2_X1 _13480_ (
    .A1(_03173_),
    .A2(_03212_),
    .ZN(_03215_)
  );
  INV_X1 _13481_ (
    .A(_03215_),
    .ZN(_03216_)
  );
  AND2_X1 _13482_ (
    .A1(_03214_),
    .A2(_03216_),
    .ZN(_03217_)
  );
  INV_X1 _13483_ (
    .A(_03217_),
    .ZN(_03218_)
  );
  AND2_X1 _13484_ (
    .A1(_02994_),
    .A2(_03217_),
    .ZN(_03219_)
  );
  INV_X1 _13485_ (
    .A(_03219_),
    .ZN(_03220_)
  );
  AND2_X1 _13486_ (
    .A1(_02995_),
    .A2(_03218_),
    .ZN(_03221_)
  );
  INV_X1 _13487_ (
    .A(_03221_),
    .ZN(_03222_)
  );
  AND2_X1 _13488_ (
    .A1(_03220_),
    .A2(_03222_),
    .ZN(_03223_)
  );
  INV_X1 _13489_ (
    .A(_03223_),
    .ZN(_03224_)
  );
  AND2_X1 _13490_ (
    .A1(_03172_),
    .A2(_03223_),
    .ZN(_03225_)
  );
  INV_X1 _13491_ (
    .A(_03225_),
    .ZN(_03226_)
  );
  AND2_X1 _13492_ (
    .A1(_03171_),
    .A2(_03224_),
    .ZN(_03227_)
  );
  INV_X1 _13493_ (
    .A(_03227_),
    .ZN(_03228_)
  );
  AND2_X1 _13494_ (
    .A1(_03226_),
    .A2(_03228_),
    .ZN(_03229_)
  );
  INV_X1 _13495_ (
    .A(_03229_),
    .ZN(_03230_)
  );
  AND2_X1 _13496_ (
    .A1(_03066_),
    .A2(_03229_),
    .ZN(_03231_)
  );
  INV_X1 _13497_ (
    .A(_03231_),
    .ZN(_03232_)
  );
  AND2_X1 _13498_ (
    .A1(_03067_),
    .A2(_03230_),
    .ZN(_03233_)
  );
  INV_X1 _13499_ (
    .A(_03233_),
    .ZN(_03234_)
  );
  AND2_X1 _13500_ (
    .A1(_03232_),
    .A2(_03234_),
    .ZN(_03235_)
  );
  INV_X1 _13501_ (
    .A(_03235_),
    .ZN(_03236_)
  );
  AND2_X1 _13502_ (
    .A1(_03170_),
    .A2(_03235_),
    .ZN(_03237_)
  );
  INV_X1 _13503_ (
    .A(_03237_),
    .ZN(_03238_)
  );
  AND2_X1 _13504_ (
    .A1(_03169_),
    .A2(_03236_),
    .ZN(_03239_)
  );
  INV_X1 _13505_ (
    .A(_03239_),
    .ZN(_03240_)
  );
  AND2_X1 _13506_ (
    .A1(_03238_),
    .A2(_03240_),
    .ZN(_03241_)
  );
  INV_X1 _13507_ (
    .A(_03241_),
    .ZN(_03242_)
  );
  AND2_X1 _13508_ (
    .A1(_03168_),
    .A2(_03241_),
    .ZN(_03243_)
  );
  INV_X1 _13509_ (
    .A(_03243_),
    .ZN(_03244_)
  );
  AND2_X1 _13510_ (
    .A1(_03167_),
    .A2(_03242_),
    .ZN(_03245_)
  );
  INV_X1 _13511_ (
    .A(_03245_),
    .ZN(_03246_)
  );
  AND2_X1 _13512_ (
    .A1(_03244_),
    .A2(_03246_),
    .ZN(_03247_)
  );
  INV_X1 _13513_ (
    .A(_03247_),
    .ZN(_03248_)
  );
  AND2_X1 _13514_ (
    .A1(remainder[32]),
    .A2(divisor[3]),
    .ZN(_03249_)
  );
  INV_X1 _13515_ (
    .A(_03249_),
    .ZN(_03250_)
  );
  AND2_X1 _13516_ (
    .A1(divisor[11]),
    .A2(remainder[0]),
    .ZN(_03251_)
  );
  INV_X1 _13517_ (
    .A(_03251_),
    .ZN(_03252_)
  );
  AND2_X1 _13518_ (
    .A1(divisor[10]),
    .A2(remainder[1]),
    .ZN(_03253_)
  );
  INV_X1 _13519_ (
    .A(_03253_),
    .ZN(_03254_)
  );
  AND2_X1 _13520_ (
    .A1(divisor[11]),
    .A2(remainder[1]),
    .ZN(_03255_)
  );
  INV_X1 _13521_ (
    .A(_03255_),
    .ZN(_03256_)
  );
  AND2_X1 _13522_ (
    .A1(_02966_),
    .A2(_03255_),
    .ZN(_03257_)
  );
  INV_X1 _13523_ (
    .A(_03257_),
    .ZN(_03258_)
  );
  AND2_X1 _13524_ (
    .A1(_03252_),
    .A2(_03254_),
    .ZN(_03259_)
  );
  INV_X1 _13525_ (
    .A(_03259_),
    .ZN(_03260_)
  );
  AND2_X1 _13526_ (
    .A1(_03258_),
    .A2(_03260_),
    .ZN(_03261_)
  );
  INV_X1 _13527_ (
    .A(_03261_),
    .ZN(_03262_)
  );
  AND2_X1 _13528_ (
    .A1(_02977_),
    .A2(_02983_),
    .ZN(_03263_)
  );
  INV_X1 _13529_ (
    .A(_03263_),
    .ZN(_03264_)
  );
  AND2_X1 _13530_ (
    .A1(divisor[8]),
    .A2(remainder[3]),
    .ZN(_03265_)
  );
  INV_X1 _13531_ (
    .A(_03265_),
    .ZN(_03266_)
  );
  AND2_X1 _13532_ (
    .A1(divisor[9]),
    .A2(remainder[3]),
    .ZN(_03267_)
  );
  INV_X1 _13533_ (
    .A(_03267_),
    .ZN(_03268_)
  );
  AND2_X1 _13534_ (
    .A1(_02974_),
    .A2(_03265_),
    .ZN(_03269_)
  );
  INV_X1 _13535_ (
    .A(_03269_),
    .ZN(_03270_)
  );
  AND2_X1 _13536_ (
    .A1(_02975_),
    .A2(_03266_),
    .ZN(_03271_)
  );
  INV_X1 _13537_ (
    .A(_03271_),
    .ZN(_03272_)
  );
  AND2_X1 _13538_ (
    .A1(_03270_),
    .A2(_03272_),
    .ZN(_03273_)
  );
  INV_X1 _13539_ (
    .A(_03273_),
    .ZN(_03274_)
  );
  AND2_X1 _13540_ (
    .A1(_02379_),
    .A2(_03273_),
    .ZN(_03275_)
  );
  INV_X1 _13541_ (
    .A(_03275_),
    .ZN(_03276_)
  );
  AND2_X1 _13542_ (
    .A1(_02380_),
    .A2(_03274_),
    .ZN(_03277_)
  );
  INV_X1 _13543_ (
    .A(_03277_),
    .ZN(_03278_)
  );
  AND2_X1 _13544_ (
    .A1(_03276_),
    .A2(_03278_),
    .ZN(_03279_)
  );
  INV_X1 _13545_ (
    .A(_03279_),
    .ZN(_03280_)
  );
  AND2_X1 _13546_ (
    .A1(_03264_),
    .A2(_03279_),
    .ZN(_03281_)
  );
  INV_X1 _13547_ (
    .A(_03281_),
    .ZN(_03282_)
  );
  AND2_X1 _13548_ (
    .A1(_03263_),
    .A2(_03280_),
    .ZN(_03283_)
  );
  INV_X1 _13549_ (
    .A(_03283_),
    .ZN(_03284_)
  );
  AND2_X1 _13550_ (
    .A1(_03282_),
    .A2(_03284_),
    .ZN(_03285_)
  );
  INV_X1 _13551_ (
    .A(_03285_),
    .ZN(_03286_)
  );
  AND2_X1 _13552_ (
    .A1(_03261_),
    .A2(_03285_),
    .ZN(_03287_)
  );
  INV_X1 _13553_ (
    .A(_03287_),
    .ZN(_03288_)
  );
  AND2_X1 _13554_ (
    .A1(_03262_),
    .A2(_03286_),
    .ZN(_03289_)
  );
  INV_X1 _13555_ (
    .A(_03289_),
    .ZN(_03290_)
  );
  AND2_X1 _13556_ (
    .A1(_03288_),
    .A2(_03290_),
    .ZN(_03291_)
  );
  INV_X1 _13557_ (
    .A(_03291_),
    .ZN(_03292_)
  );
  AND2_X1 _13558_ (
    .A1(_03249_),
    .A2(_03292_),
    .ZN(_03293_)
  );
  INV_X1 _13559_ (
    .A(_03293_),
    .ZN(_03294_)
  );
  AND2_X1 _13560_ (
    .A1(_03250_),
    .A2(_03291_),
    .ZN(_03295_)
  );
  INV_X1 _13561_ (
    .A(_03295_),
    .ZN(_03296_)
  );
  AND2_X1 _13562_ (
    .A1(_03294_),
    .A2(_03296_),
    .ZN(_03297_)
  );
  INV_X1 _13563_ (
    .A(_03297_),
    .ZN(_03298_)
  );
  AND2_X1 _13564_ (
    .A1(_03000_),
    .A2(_03298_),
    .ZN(_03299_)
  );
  INV_X1 _13565_ (
    .A(_03299_),
    .ZN(_03300_)
  );
  AND2_X1 _13566_ (
    .A1(_03001_),
    .A2(_03297_),
    .ZN(_03301_)
  );
  INV_X1 _13567_ (
    .A(_03301_),
    .ZN(_03302_)
  );
  AND2_X1 _13568_ (
    .A1(_03300_),
    .A2(_03302_),
    .ZN(_03303_)
  );
  INV_X1 _13569_ (
    .A(_03303_),
    .ZN(_03304_)
  );
  AND2_X1 _13570_ (
    .A1(_03247_),
    .A2(_03303_),
    .ZN(_03305_)
  );
  INV_X1 _13571_ (
    .A(_03305_),
    .ZN(_03306_)
  );
  AND2_X1 _13572_ (
    .A1(_03248_),
    .A2(_03304_),
    .ZN(_03307_)
  );
  INV_X1 _13573_ (
    .A(_03307_),
    .ZN(_03308_)
  );
  AND2_X1 _13574_ (
    .A1(_03306_),
    .A2(_03308_),
    .ZN(_03309_)
  );
  INV_X1 _13575_ (
    .A(_03309_),
    .ZN(_03310_)
  );
  AND2_X1 _13576_ (
    .A1(_03166_),
    .A2(_03309_),
    .ZN(_03311_)
  );
  INV_X1 _13577_ (
    .A(_03311_),
    .ZN(_03312_)
  );
  AND2_X1 _13578_ (
    .A1(_03165_),
    .A2(_03310_),
    .ZN(_03313_)
  );
  INV_X1 _13579_ (
    .A(_03313_),
    .ZN(_03314_)
  );
  AND2_X1 _13580_ (
    .A1(_03312_),
    .A2(_03314_),
    .ZN(_03315_)
  );
  INV_X1 _13581_ (
    .A(_03315_),
    .ZN(_03316_)
  );
  AND2_X1 _13582_ (
    .A1(_03084_),
    .A2(_03315_),
    .ZN(_03317_)
  );
  INV_X1 _13583_ (
    .A(_03317_),
    .ZN(_03318_)
  );
  AND2_X1 _13584_ (
    .A1(_03085_),
    .A2(_03316_),
    .ZN(_03319_)
  );
  INV_X1 _13585_ (
    .A(_03319_),
    .ZN(_03320_)
  );
  AND2_X1 _13586_ (
    .A1(_03318_),
    .A2(_03320_),
    .ZN(_03321_)
  );
  INV_X1 _13587_ (
    .A(_03321_),
    .ZN(_03322_)
  );
  AND2_X1 _13588_ (
    .A1(_03164_),
    .A2(_03321_),
    .ZN(_03323_)
  );
  INV_X1 _13589_ (
    .A(_03323_),
    .ZN(_03324_)
  );
  AND2_X1 _13590_ (
    .A1(_03163_),
    .A2(_03322_),
    .ZN(_03325_)
  );
  INV_X1 _13591_ (
    .A(_03325_),
    .ZN(_03326_)
  );
  AND2_X1 _13592_ (
    .A1(_03324_),
    .A2(_03326_),
    .ZN(_03327_)
  );
  INV_X1 _13593_ (
    .A(_03327_),
    .ZN(_03328_)
  );
  AND2_X1 _13594_ (
    .A1(_03108_),
    .A2(_03327_),
    .ZN(_03329_)
  );
  INV_X1 _13595_ (
    .A(_03329_),
    .ZN(_03330_)
  );
  AND2_X1 _13596_ (
    .A1(_03109_),
    .A2(_03328_),
    .ZN(_03331_)
  );
  INV_X1 _13597_ (
    .A(_03331_),
    .ZN(_03332_)
  );
  AND2_X1 _13598_ (
    .A1(_03330_),
    .A2(_03332_),
    .ZN(_03333_)
  );
  INV_X1 _13599_ (
    .A(_03333_),
    .ZN(_03334_)
  );
  AND2_X1 _13600_ (
    .A1(_03162_),
    .A2(_03333_),
    .ZN(_03335_)
  );
  INV_X1 _13601_ (
    .A(_03335_),
    .ZN(_03336_)
  );
  AND2_X1 _13602_ (
    .A1(_03161_),
    .A2(_03334_),
    .ZN(_03337_)
  );
  INV_X1 _13603_ (
    .A(_03337_),
    .ZN(_03338_)
  );
  AND2_X1 _13604_ (
    .A1(_03336_),
    .A2(_03338_),
    .ZN(_03339_)
  );
  INV_X1 _13605_ (
    .A(_03339_),
    .ZN(_03340_)
  );
  AND2_X1 _13606_ (
    .A1(remainder[44]),
    .A2(_03339_),
    .ZN(_03341_)
  );
  INV_X1 _13607_ (
    .A(_03341_),
    .ZN(_03342_)
  );
  AND2_X1 _13608_ (
    .A1(_04634_),
    .A2(_03340_),
    .ZN(_03343_)
  );
  INV_X1 _13609_ (
    .A(_03343_),
    .ZN(_03344_)
  );
  AND2_X1 _13610_ (
    .A1(_03342_),
    .A2(_03344_),
    .ZN(_03345_)
  );
  INV_X1 _13611_ (
    .A(_03345_),
    .ZN(_03346_)
  );
  AND2_X1 _13612_ (
    .A1(_03160_),
    .A2(_03345_),
    .ZN(_03347_)
  );
  INV_X1 _13613_ (
    .A(_03347_),
    .ZN(_03348_)
  );
  AND2_X1 _13614_ (
    .A1(_03159_),
    .A2(_03346_),
    .ZN(_03349_)
  );
  INV_X1 _13615_ (
    .A(_03349_),
    .ZN(_03350_)
  );
  AND2_X1 _13616_ (
    .A1(_02082_),
    .A2(_03348_),
    .ZN(_03351_)
  );
  AND2_X1 _13617_ (
    .A1(_03350_),
    .A2(_03351_),
    .ZN(_03352_)
  );
  INV_X1 _13618_ (
    .A(_03352_),
    .ZN(_03353_)
  );
  AND2_X1 _13619_ (
    .A1(_03158_),
    .A2(_03353_),
    .ZN(_03354_)
  );
  AND2_X1 _13620_ (
    .A1(_03156_),
    .A2(_03354_),
    .ZN(_03355_)
  );
  INV_X1 _13621_ (
    .A(_03355_),
    .ZN(_03356_)
  );
  AND2_X1 _13622_ (
    .A1(_06201_),
    .A2(_03356_),
    .ZN(_00057_)
  );
  AND2_X1 _13623_ (
    .A1(_04722_),
    .A2(_10451_),
    .ZN(_03357_)
  );
  INV_X1 _13624_ (
    .A(_03357_),
    .ZN(_03358_)
  );
  AND2_X1 _13625_ (
    .A1(_10462_),
    .A2(_00873_),
    .ZN(_03359_)
  );
  INV_X1 _13626_ (
    .A(_03359_),
    .ZN(_03360_)
  );
  AND2_X1 _13627_ (
    .A1(_05983_),
    .A2(_03360_),
    .ZN(_03361_)
  );
  AND2_X1 _13628_ (
    .A1(_03358_),
    .A2(_03361_),
    .ZN(_03362_)
  );
  INV_X1 _13629_ (
    .A(_03362_),
    .ZN(_03363_)
  );
  AND2_X1 _13630_ (
    .A1(remainder[37]),
    .A2(_02077_),
    .ZN(_03364_)
  );
  INV_X1 _13631_ (
    .A(_03364_),
    .ZN(_03365_)
  );
  AND2_X1 _13632_ (
    .A1(_03342_),
    .A2(_03348_),
    .ZN(_03366_)
  );
  INV_X1 _13633_ (
    .A(_03366_),
    .ZN(_03367_)
  );
  AND2_X1 _13634_ (
    .A1(_03330_),
    .A2(_03336_),
    .ZN(_03368_)
  );
  INV_X1 _13635_ (
    .A(_03368_),
    .ZN(_03369_)
  );
  AND2_X1 _13636_ (
    .A1(_03312_),
    .A2(_03318_),
    .ZN(_03370_)
  );
  INV_X1 _13637_ (
    .A(_03370_),
    .ZN(_03371_)
  );
  AND2_X1 _13638_ (
    .A1(_03300_),
    .A2(_03306_),
    .ZN(_03372_)
  );
  INV_X1 _13639_ (
    .A(_03372_),
    .ZN(_03373_)
  );
  AND2_X1 _13640_ (
    .A1(_03232_),
    .A2(_03238_),
    .ZN(_03374_)
  );
  INV_X1 _13641_ (
    .A(_03374_),
    .ZN(_03375_)
  );
  AND2_X1 _13642_ (
    .A1(_03220_),
    .A2(_03226_),
    .ZN(_03376_)
  );
  INV_X1 _13643_ (
    .A(_03376_),
    .ZN(_03377_)
  );
  AND2_X1 _13644_ (
    .A1(_03208_),
    .A2(_03214_),
    .ZN(_03378_)
  );
  INV_X1 _13645_ (
    .A(_03378_),
    .ZN(_03379_)
  );
  AND2_X1 _13646_ (
    .A1(_03196_),
    .A2(_03202_),
    .ZN(_03380_)
  );
  INV_X1 _13647_ (
    .A(_03380_),
    .ZN(_03381_)
  );
  AND2_X1 _13648_ (
    .A1(_03184_),
    .A2(_03190_),
    .ZN(_03382_)
  );
  INV_X1 _13649_ (
    .A(_03382_),
    .ZN(_03383_)
  );
  AND2_X1 _13650_ (
    .A1(remainder[32]),
    .A2(divisor[4]),
    .ZN(_03384_)
  );
  INV_X1 _13651_ (
    .A(_03384_),
    .ZN(_03385_)
  );
  AND2_X1 _13652_ (
    .A1(divisor[5]),
    .A2(remainder[7]),
    .ZN(_03386_)
  );
  INV_X1 _13653_ (
    .A(_03386_),
    .ZN(_03387_)
  );
  AND2_X1 _13654_ (
    .A1(divisor[6]),
    .A2(remainder[7]),
    .ZN(_03388_)
  );
  INV_X1 _13655_ (
    .A(_03388_),
    .ZN(_03389_)
  );
  AND2_X1 _13656_ (
    .A1(_03179_),
    .A2(_03388_),
    .ZN(_03390_)
  );
  INV_X1 _13657_ (
    .A(_03390_),
    .ZN(_03391_)
  );
  AND2_X1 _13658_ (
    .A1(_03182_),
    .A2(_03387_),
    .ZN(_03392_)
  );
  INV_X1 _13659_ (
    .A(_03392_),
    .ZN(_03393_)
  );
  AND2_X1 _13660_ (
    .A1(_03391_),
    .A2(_03393_),
    .ZN(_03394_)
  );
  INV_X1 _13661_ (
    .A(_03394_),
    .ZN(_03395_)
  );
  AND2_X1 _13662_ (
    .A1(_03384_),
    .A2(_03394_),
    .ZN(_03396_)
  );
  INV_X1 _13663_ (
    .A(_03396_),
    .ZN(_03397_)
  );
  AND2_X1 _13664_ (
    .A1(_03385_),
    .A2(_03395_),
    .ZN(_03398_)
  );
  INV_X1 _13665_ (
    .A(_03398_),
    .ZN(_03399_)
  );
  AND2_X1 _13666_ (
    .A1(_03397_),
    .A2(_03399_),
    .ZN(_03400_)
  );
  INV_X1 _13667_ (
    .A(_03400_),
    .ZN(_03401_)
  );
  AND2_X1 _13668_ (
    .A1(_03383_),
    .A2(_03400_),
    .ZN(_03402_)
  );
  INV_X1 _13669_ (
    .A(_03402_),
    .ZN(_03403_)
  );
  AND2_X1 _13670_ (
    .A1(_03382_),
    .A2(_03401_),
    .ZN(_03404_)
  );
  INV_X1 _13671_ (
    .A(_03404_),
    .ZN(_03405_)
  );
  AND2_X1 _13672_ (
    .A1(_03403_),
    .A2(_03405_),
    .ZN(_03406_)
  );
  INV_X1 _13673_ (
    .A(_03406_),
    .ZN(_03407_)
  );
  AND2_X1 _13674_ (
    .A1(_03046_),
    .A2(_03406_),
    .ZN(_03408_)
  );
  INV_X1 _13675_ (
    .A(_03408_),
    .ZN(_03409_)
  );
  AND2_X1 _13676_ (
    .A1(_03047_),
    .A2(_03407_),
    .ZN(_03410_)
  );
  INV_X1 _13677_ (
    .A(_03410_),
    .ZN(_03411_)
  );
  AND2_X1 _13678_ (
    .A1(_03409_),
    .A2(_03411_),
    .ZN(_03412_)
  );
  INV_X1 _13679_ (
    .A(_03412_),
    .ZN(_03413_)
  );
  AND2_X1 _13680_ (
    .A1(_03281_),
    .A2(_03412_),
    .ZN(_03414_)
  );
  INV_X1 _13681_ (
    .A(_03414_),
    .ZN(_03415_)
  );
  AND2_X1 _13682_ (
    .A1(_03282_),
    .A2(_03413_),
    .ZN(_03416_)
  );
  INV_X1 _13683_ (
    .A(_03416_),
    .ZN(_03417_)
  );
  AND2_X1 _13684_ (
    .A1(_03415_),
    .A2(_03417_),
    .ZN(_03418_)
  );
  INV_X1 _13685_ (
    .A(_03418_),
    .ZN(_03419_)
  );
  AND2_X1 _13686_ (
    .A1(_03381_),
    .A2(_03418_),
    .ZN(_03420_)
  );
  INV_X1 _13687_ (
    .A(_03420_),
    .ZN(_03421_)
  );
  AND2_X1 _13688_ (
    .A1(_03380_),
    .A2(_03419_),
    .ZN(_03422_)
  );
  INV_X1 _13689_ (
    .A(_03422_),
    .ZN(_03423_)
  );
  AND2_X1 _13690_ (
    .A1(_03421_),
    .A2(_03423_),
    .ZN(_03424_)
  );
  INV_X1 _13691_ (
    .A(_03424_),
    .ZN(_03425_)
  );
  AND2_X1 _13692_ (
    .A1(_03287_),
    .A2(_03424_),
    .ZN(_03426_)
  );
  INV_X1 _13693_ (
    .A(_03426_),
    .ZN(_03427_)
  );
  AND2_X1 _13694_ (
    .A1(_03288_),
    .A2(_03425_),
    .ZN(_03428_)
  );
  INV_X1 _13695_ (
    .A(_03428_),
    .ZN(_03429_)
  );
  AND2_X1 _13696_ (
    .A1(_03427_),
    .A2(_03429_),
    .ZN(_03430_)
  );
  INV_X1 _13697_ (
    .A(_03430_),
    .ZN(_03431_)
  );
  AND2_X1 _13698_ (
    .A1(_03379_),
    .A2(_03430_),
    .ZN(_03432_)
  );
  INV_X1 _13699_ (
    .A(_03432_),
    .ZN(_03433_)
  );
  AND2_X1 _13700_ (
    .A1(_03378_),
    .A2(_03431_),
    .ZN(_03434_)
  );
  INV_X1 _13701_ (
    .A(_03434_),
    .ZN(_03435_)
  );
  AND2_X1 _13702_ (
    .A1(_03433_),
    .A2(_03435_),
    .ZN(_03436_)
  );
  INV_X1 _13703_ (
    .A(_03436_),
    .ZN(_03437_)
  );
  AND2_X1 _13704_ (
    .A1(_03377_),
    .A2(_03436_),
    .ZN(_03438_)
  );
  INV_X1 _13705_ (
    .A(_03438_),
    .ZN(_03439_)
  );
  AND2_X1 _13706_ (
    .A1(_03376_),
    .A2(_03437_),
    .ZN(_03440_)
  );
  INV_X1 _13707_ (
    .A(_03440_),
    .ZN(_03441_)
  );
  AND2_X1 _13708_ (
    .A1(_03439_),
    .A2(_03441_),
    .ZN(_03442_)
  );
  INV_X1 _13709_ (
    .A(_03442_),
    .ZN(_03443_)
  );
  AND2_X1 _13710_ (
    .A1(_03170_),
    .A2(_03442_),
    .ZN(_03444_)
  );
  INV_X1 _13711_ (
    .A(_03444_),
    .ZN(_03445_)
  );
  AND2_X1 _13712_ (
    .A1(_03169_),
    .A2(_03443_),
    .ZN(_03446_)
  );
  INV_X1 _13713_ (
    .A(_03446_),
    .ZN(_03447_)
  );
  AND2_X1 _13714_ (
    .A1(_03445_),
    .A2(_03447_),
    .ZN(_03448_)
  );
  INV_X1 _13715_ (
    .A(_03448_),
    .ZN(_03449_)
  );
  AND2_X1 _13716_ (
    .A1(_03375_),
    .A2(_03448_),
    .ZN(_03450_)
  );
  INV_X1 _13717_ (
    .A(_03450_),
    .ZN(_03451_)
  );
  AND2_X1 _13718_ (
    .A1(_03374_),
    .A2(_03449_),
    .ZN(_03452_)
  );
  INV_X1 _13719_ (
    .A(_03452_),
    .ZN(_03453_)
  );
  AND2_X1 _13720_ (
    .A1(_03451_),
    .A2(_03453_),
    .ZN(_03454_)
  );
  INV_X1 _13721_ (
    .A(_03454_),
    .ZN(_03455_)
  );
  AND2_X1 _13722_ (
    .A1(divisor[10]),
    .A2(remainder[2]),
    .ZN(_03456_)
  );
  INV_X1 _13723_ (
    .A(_03456_),
    .ZN(_03457_)
  );
  AND2_X1 _13724_ (
    .A1(divisor[12]),
    .A2(remainder[0]),
    .ZN(_03458_)
  );
  INV_X1 _13725_ (
    .A(_03458_),
    .ZN(_03459_)
  );
  AND2_X1 _13726_ (
    .A1(divisor[12]),
    .A2(remainder[1]),
    .ZN(_03460_)
  );
  INV_X1 _13727_ (
    .A(_03460_),
    .ZN(_03461_)
  );
  AND2_X1 _13728_ (
    .A1(_03251_),
    .A2(_03460_),
    .ZN(_03462_)
  );
  INV_X1 _13729_ (
    .A(_03462_),
    .ZN(_03463_)
  );
  AND2_X1 _13730_ (
    .A1(_03256_),
    .A2(_03459_),
    .ZN(_03464_)
  );
  INV_X1 _13731_ (
    .A(_03464_),
    .ZN(_03465_)
  );
  AND2_X1 _13732_ (
    .A1(_03463_),
    .A2(_03465_),
    .ZN(_03466_)
  );
  INV_X1 _13733_ (
    .A(_03466_),
    .ZN(_03467_)
  );
  AND2_X1 _13734_ (
    .A1(_03456_),
    .A2(_03466_),
    .ZN(_03468_)
  );
  INV_X1 _13735_ (
    .A(_03468_),
    .ZN(_03469_)
  );
  AND2_X1 _13736_ (
    .A1(_03457_),
    .A2(_03467_),
    .ZN(_03470_)
  );
  INV_X1 _13737_ (
    .A(_03470_),
    .ZN(_03471_)
  );
  AND2_X1 _13738_ (
    .A1(_03469_),
    .A2(_03471_),
    .ZN(_03472_)
  );
  INV_X1 _13739_ (
    .A(_03472_),
    .ZN(_03473_)
  );
  AND2_X1 _13740_ (
    .A1(_03270_),
    .A2(_03276_),
    .ZN(_03474_)
  );
  INV_X1 _13741_ (
    .A(_03474_),
    .ZN(_03475_)
  );
  AND2_X1 _13742_ (
    .A1(divisor[7]),
    .A2(remainder[5]),
    .ZN(_03476_)
  );
  INV_X1 _13743_ (
    .A(_03476_),
    .ZN(_03477_)
  );
  AND2_X1 _13744_ (
    .A1(divisor[8]),
    .A2(remainder[4]),
    .ZN(_03478_)
  );
  INV_X1 _13745_ (
    .A(_03478_),
    .ZN(_03479_)
  );
  AND2_X1 _13746_ (
    .A1(divisor[9]),
    .A2(remainder[4]),
    .ZN(_03480_)
  );
  INV_X1 _13747_ (
    .A(_03480_),
    .ZN(_03481_)
  );
  AND2_X1 _13748_ (
    .A1(_03267_),
    .A2(_03478_),
    .ZN(_03482_)
  );
  INV_X1 _13749_ (
    .A(_03482_),
    .ZN(_03483_)
  );
  AND2_X1 _13750_ (
    .A1(_03268_),
    .A2(_03479_),
    .ZN(_03484_)
  );
  INV_X1 _13751_ (
    .A(_03484_),
    .ZN(_03485_)
  );
  AND2_X1 _13752_ (
    .A1(_03483_),
    .A2(_03485_),
    .ZN(_03486_)
  );
  INV_X1 _13753_ (
    .A(_03486_),
    .ZN(_03487_)
  );
  AND2_X1 _13754_ (
    .A1(_03476_),
    .A2(_03486_),
    .ZN(_03488_)
  );
  INV_X1 _13755_ (
    .A(_03488_),
    .ZN(_03489_)
  );
  AND2_X1 _13756_ (
    .A1(_03477_),
    .A2(_03487_),
    .ZN(_03490_)
  );
  INV_X1 _13757_ (
    .A(_03490_),
    .ZN(_03491_)
  );
  AND2_X1 _13758_ (
    .A1(_03489_),
    .A2(_03491_),
    .ZN(_03492_)
  );
  INV_X1 _13759_ (
    .A(_03492_),
    .ZN(_03493_)
  );
  AND2_X1 _13760_ (
    .A1(_03257_),
    .A2(_03492_),
    .ZN(_03494_)
  );
  INV_X1 _13761_ (
    .A(_03494_),
    .ZN(_03495_)
  );
  AND2_X1 _13762_ (
    .A1(_03258_),
    .A2(_03493_),
    .ZN(_03496_)
  );
  INV_X1 _13763_ (
    .A(_03496_),
    .ZN(_03497_)
  );
  AND2_X1 _13764_ (
    .A1(_03495_),
    .A2(_03497_),
    .ZN(_03498_)
  );
  INV_X1 _13765_ (
    .A(_03498_),
    .ZN(_03499_)
  );
  AND2_X1 _13766_ (
    .A1(_03475_),
    .A2(_03498_),
    .ZN(_03500_)
  );
  INV_X1 _13767_ (
    .A(_03500_),
    .ZN(_03501_)
  );
  AND2_X1 _13768_ (
    .A1(_03474_),
    .A2(_03499_),
    .ZN(_03502_)
  );
  INV_X1 _13769_ (
    .A(_03502_),
    .ZN(_03503_)
  );
  AND2_X1 _13770_ (
    .A1(_03501_),
    .A2(_03503_),
    .ZN(_03504_)
  );
  INV_X1 _13771_ (
    .A(_03504_),
    .ZN(_03505_)
  );
  AND2_X1 _13772_ (
    .A1(_03472_),
    .A2(_03504_),
    .ZN(_03506_)
  );
  INV_X1 _13773_ (
    .A(_03506_),
    .ZN(_03507_)
  );
  AND2_X1 _13774_ (
    .A1(_03473_),
    .A2(_03505_),
    .ZN(_03508_)
  );
  INV_X1 _13775_ (
    .A(_03508_),
    .ZN(_03509_)
  );
  AND2_X1 _13776_ (
    .A1(_03507_),
    .A2(_03509_),
    .ZN(_03510_)
  );
  INV_X1 _13777_ (
    .A(_03510_),
    .ZN(_03511_)
  );
  AND2_X1 _13778_ (
    .A1(_03294_),
    .A2(_03511_),
    .ZN(_03512_)
  );
  INV_X1 _13779_ (
    .A(_03512_),
    .ZN(_03513_)
  );
  AND2_X1 _13780_ (
    .A1(_03293_),
    .A2(_03510_),
    .ZN(_03514_)
  );
  INV_X1 _13781_ (
    .A(_03514_),
    .ZN(_03515_)
  );
  AND2_X1 _13782_ (
    .A1(_03293_),
    .A2(_03511_),
    .ZN(_03516_)
  );
  INV_X1 _13783_ (
    .A(_03516_),
    .ZN(_03517_)
  );
  AND2_X1 _13784_ (
    .A1(_03294_),
    .A2(_03510_),
    .ZN(_03518_)
  );
  INV_X1 _13785_ (
    .A(_03518_),
    .ZN(_03519_)
  );
  AND2_X1 _13786_ (
    .A1(_03513_),
    .A2(_03515_),
    .ZN(_03520_)
  );
  AND2_X1 _13787_ (
    .A1(_03517_),
    .A2(_03519_),
    .ZN(_03521_)
  );
  AND2_X1 _13788_ (
    .A1(_03454_),
    .A2(_03520_),
    .ZN(_03522_)
  );
  INV_X1 _13789_ (
    .A(_03522_),
    .ZN(_03523_)
  );
  AND2_X1 _13790_ (
    .A1(_03455_),
    .A2(_03521_),
    .ZN(_03524_)
  );
  INV_X1 _13791_ (
    .A(_03524_),
    .ZN(_03525_)
  );
  AND2_X1 _13792_ (
    .A1(_03523_),
    .A2(_03525_),
    .ZN(_03526_)
  );
  INV_X1 _13793_ (
    .A(_03526_),
    .ZN(_03527_)
  );
  AND2_X1 _13794_ (
    .A1(_03373_),
    .A2(_03526_),
    .ZN(_03528_)
  );
  INV_X1 _13795_ (
    .A(_03528_),
    .ZN(_03529_)
  );
  AND2_X1 _13796_ (
    .A1(_03372_),
    .A2(_03527_),
    .ZN(_03530_)
  );
  INV_X1 _13797_ (
    .A(_03530_),
    .ZN(_03531_)
  );
  AND2_X1 _13798_ (
    .A1(_03529_),
    .A2(_03531_),
    .ZN(_03532_)
  );
  INV_X1 _13799_ (
    .A(_03532_),
    .ZN(_03533_)
  );
  AND2_X1 _13800_ (
    .A1(_03243_),
    .A2(_03532_),
    .ZN(_03534_)
  );
  INV_X1 _13801_ (
    .A(_03534_),
    .ZN(_03535_)
  );
  AND2_X1 _13802_ (
    .A1(_03244_),
    .A2(_03533_),
    .ZN(_03536_)
  );
  INV_X1 _13803_ (
    .A(_03536_),
    .ZN(_03537_)
  );
  AND2_X1 _13804_ (
    .A1(_03535_),
    .A2(_03537_),
    .ZN(_03538_)
  );
  INV_X1 _13805_ (
    .A(_03538_),
    .ZN(_03539_)
  );
  AND2_X1 _13806_ (
    .A1(_03371_),
    .A2(_03538_),
    .ZN(_03540_)
  );
  INV_X1 _13807_ (
    .A(_03540_),
    .ZN(_03541_)
  );
  AND2_X1 _13808_ (
    .A1(_03370_),
    .A2(_03539_),
    .ZN(_03542_)
  );
  INV_X1 _13809_ (
    .A(_03542_),
    .ZN(_03543_)
  );
  AND2_X1 _13810_ (
    .A1(_03541_),
    .A2(_03543_),
    .ZN(_03544_)
  );
  INV_X1 _13811_ (
    .A(_03544_),
    .ZN(_03545_)
  );
  AND2_X1 _13812_ (
    .A1(_03323_),
    .A2(_03544_),
    .ZN(_03546_)
  );
  INV_X1 _13813_ (
    .A(_03546_),
    .ZN(_03547_)
  );
  AND2_X1 _13814_ (
    .A1(_03324_),
    .A2(_03545_),
    .ZN(_03548_)
  );
  INV_X1 _13815_ (
    .A(_03548_),
    .ZN(_03549_)
  );
  AND2_X1 _13816_ (
    .A1(_03547_),
    .A2(_03549_),
    .ZN(_03550_)
  );
  INV_X1 _13817_ (
    .A(_03550_),
    .ZN(_03551_)
  );
  AND2_X1 _13818_ (
    .A1(_03369_),
    .A2(_03550_),
    .ZN(_03552_)
  );
  INV_X1 _13819_ (
    .A(_03552_),
    .ZN(_03553_)
  );
  AND2_X1 _13820_ (
    .A1(_03368_),
    .A2(_03551_),
    .ZN(_03554_)
  );
  INV_X1 _13821_ (
    .A(_03554_),
    .ZN(_03555_)
  );
  AND2_X1 _13822_ (
    .A1(_03553_),
    .A2(_03555_),
    .ZN(_03556_)
  );
  INV_X1 _13823_ (
    .A(_03556_),
    .ZN(_03557_)
  );
  AND2_X1 _13824_ (
    .A1(remainder[45]),
    .A2(_03556_),
    .ZN(_03558_)
  );
  INV_X1 _13825_ (
    .A(_03558_),
    .ZN(_03559_)
  );
  AND2_X1 _13826_ (
    .A1(_04623_),
    .A2(_03557_),
    .ZN(_03560_)
  );
  INV_X1 _13827_ (
    .A(_03560_),
    .ZN(_03561_)
  );
  AND2_X1 _13828_ (
    .A1(_03559_),
    .A2(_03561_),
    .ZN(_03562_)
  );
  INV_X1 _13829_ (
    .A(_03562_),
    .ZN(_03563_)
  );
  AND2_X1 _13830_ (
    .A1(_03367_),
    .A2(_03562_),
    .ZN(_03564_)
  );
  INV_X1 _13831_ (
    .A(_03564_),
    .ZN(_03565_)
  );
  AND2_X1 _13832_ (
    .A1(_03366_),
    .A2(_03563_),
    .ZN(_03566_)
  );
  INV_X1 _13833_ (
    .A(_03566_),
    .ZN(_03567_)
  );
  AND2_X1 _13834_ (
    .A1(_02082_),
    .A2(_03567_),
    .ZN(_03568_)
  );
  AND2_X1 _13835_ (
    .A1(_03565_),
    .A2(_03568_),
    .ZN(_03569_)
  );
  INV_X1 _13836_ (
    .A(_03569_),
    .ZN(_03570_)
  );
  AND2_X1 _13837_ (
    .A1(_03365_),
    .A2(_03570_),
    .ZN(_03571_)
  );
  AND2_X1 _13838_ (
    .A1(_03363_),
    .A2(_03571_),
    .ZN(_03572_)
  );
  INV_X1 _13839_ (
    .A(_03572_),
    .ZN(_03573_)
  );
  AND2_X1 _13840_ (
    .A1(_06201_),
    .A2(_03573_),
    .ZN(_00058_)
  );
  AND2_X1 _13841_ (
    .A1(_04711_),
    .A2(_10451_),
    .ZN(_03574_)
  );
  INV_X1 _13842_ (
    .A(_03574_),
    .ZN(_03575_)
  );
  AND2_X1 _13843_ (
    .A1(_10462_),
    .A2(_01005_),
    .ZN(_03576_)
  );
  INV_X1 _13844_ (
    .A(_03576_),
    .ZN(_03577_)
  );
  AND2_X1 _13845_ (
    .A1(_05983_),
    .A2(_03577_),
    .ZN(_03578_)
  );
  AND2_X1 _13846_ (
    .A1(_03575_),
    .A2(_03578_),
    .ZN(_03579_)
  );
  INV_X1 _13847_ (
    .A(_03579_),
    .ZN(_03580_)
  );
  AND2_X1 _13848_ (
    .A1(remainder[38]),
    .A2(_02077_),
    .ZN(_03581_)
  );
  INV_X1 _13849_ (
    .A(_03581_),
    .ZN(_03582_)
  );
  AND2_X1 _13850_ (
    .A1(_03559_),
    .A2(_03565_),
    .ZN(_03583_)
  );
  INV_X1 _13851_ (
    .A(_03583_),
    .ZN(_03584_)
  );
  AND2_X1 _13852_ (
    .A1(_03547_),
    .A2(_03553_),
    .ZN(_03585_)
  );
  INV_X1 _13853_ (
    .A(_03585_),
    .ZN(_03586_)
  );
  AND2_X1 _13854_ (
    .A1(_03529_),
    .A2(_03535_),
    .ZN(_03587_)
  );
  INV_X1 _13855_ (
    .A(_03587_),
    .ZN(_03588_)
  );
  AND2_X1 _13856_ (
    .A1(_03249_),
    .A2(_03511_),
    .ZN(_03589_)
  );
  INV_X1 _13857_ (
    .A(_03589_),
    .ZN(_03590_)
  );
  AND2_X1 _13858_ (
    .A1(_03291_),
    .A2(_03589_),
    .ZN(_03591_)
  );
  INV_X1 _13859_ (
    .A(_03591_),
    .ZN(_03592_)
  );
  AND2_X1 _13860_ (
    .A1(_03523_),
    .A2(_03592_),
    .ZN(_03593_)
  );
  INV_X1 _13861_ (
    .A(_03593_),
    .ZN(_03594_)
  );
  AND2_X1 _13862_ (
    .A1(_03439_),
    .A2(_03445_),
    .ZN(_03595_)
  );
  INV_X1 _13863_ (
    .A(_03595_),
    .ZN(_03596_)
  );
  AND2_X1 _13864_ (
    .A1(_03427_),
    .A2(_03433_),
    .ZN(_03597_)
  );
  INV_X1 _13865_ (
    .A(_03597_),
    .ZN(_03598_)
  );
  AND2_X1 _13866_ (
    .A1(_03415_),
    .A2(_03421_),
    .ZN(_03599_)
  );
  INV_X1 _13867_ (
    .A(_03599_),
    .ZN(_03600_)
  );
  AND2_X1 _13868_ (
    .A1(_03403_),
    .A2(_03409_),
    .ZN(_03601_)
  );
  INV_X1 _13869_ (
    .A(_03601_),
    .ZN(_03602_)
  );
  AND2_X1 _13870_ (
    .A1(_03495_),
    .A2(_03501_),
    .ZN(_03603_)
  );
  INV_X1 _13871_ (
    .A(_03603_),
    .ZN(_03604_)
  );
  AND2_X1 _13872_ (
    .A1(_03391_),
    .A2(_03397_),
    .ZN(_03605_)
  );
  INV_X1 _13873_ (
    .A(_03605_),
    .ZN(_03606_)
  );
  AND2_X1 _13874_ (
    .A1(remainder[32]),
    .A2(divisor[6]),
    .ZN(_03607_)
  );
  INV_X1 _13875_ (
    .A(_03607_),
    .ZN(_03608_)
  );
  AND2_X1 _13876_ (
    .A1(remainder[32]),
    .A2(divisor[5]),
    .ZN(_03609_)
  );
  INV_X1 _13877_ (
    .A(_03609_),
    .ZN(_03610_)
  );
  AND2_X1 _13878_ (
    .A1(_03388_),
    .A2(_03609_),
    .ZN(_03611_)
  );
  INV_X1 _13879_ (
    .A(_03611_),
    .ZN(_03612_)
  );
  AND2_X1 _13880_ (
    .A1(_03389_),
    .A2(_03610_),
    .ZN(_03613_)
  );
  INV_X1 _13881_ (
    .A(_03613_),
    .ZN(_03614_)
  );
  AND2_X1 _13882_ (
    .A1(_03612_),
    .A2(_03614_),
    .ZN(_03615_)
  );
  INV_X1 _13883_ (
    .A(_03615_),
    .ZN(_03616_)
  );
  AND2_X1 _13884_ (
    .A1(_03384_),
    .A2(_03615_),
    .ZN(_03617_)
  );
  INV_X1 _13885_ (
    .A(_03617_),
    .ZN(_03618_)
  );
  AND2_X1 _13886_ (
    .A1(_03385_),
    .A2(_03616_),
    .ZN(_03619_)
  );
  INV_X1 _13887_ (
    .A(_03619_),
    .ZN(_03620_)
  );
  AND2_X1 _13888_ (
    .A1(_03618_),
    .A2(_03620_),
    .ZN(_03621_)
  );
  INV_X1 _13889_ (
    .A(_03621_),
    .ZN(_03622_)
  );
  AND2_X1 _13890_ (
    .A1(_03606_),
    .A2(_03621_),
    .ZN(_03623_)
  );
  INV_X1 _13891_ (
    .A(_03623_),
    .ZN(_03624_)
  );
  AND2_X1 _13892_ (
    .A1(_03605_),
    .A2(_03622_),
    .ZN(_03625_)
  );
  INV_X1 _13893_ (
    .A(_03625_),
    .ZN(_03626_)
  );
  AND2_X1 _13894_ (
    .A1(_03624_),
    .A2(_03626_),
    .ZN(_03627_)
  );
  INV_X1 _13895_ (
    .A(_03627_),
    .ZN(_03628_)
  );
  AND2_X1 _13896_ (
    .A1(_03046_),
    .A2(_03627_),
    .ZN(_03629_)
  );
  INV_X1 _13897_ (
    .A(_03629_),
    .ZN(_03630_)
  );
  AND2_X1 _13898_ (
    .A1(_03047_),
    .A2(_03628_),
    .ZN(_03631_)
  );
  INV_X1 _13899_ (
    .A(_03631_),
    .ZN(_03632_)
  );
  AND2_X1 _13900_ (
    .A1(_03630_),
    .A2(_03632_),
    .ZN(_03633_)
  );
  INV_X1 _13901_ (
    .A(_03633_),
    .ZN(_03634_)
  );
  AND2_X1 _13902_ (
    .A1(_03604_),
    .A2(_03633_),
    .ZN(_03635_)
  );
  INV_X1 _13903_ (
    .A(_03635_),
    .ZN(_03636_)
  );
  AND2_X1 _13904_ (
    .A1(_03603_),
    .A2(_03634_),
    .ZN(_03637_)
  );
  INV_X1 _13905_ (
    .A(_03637_),
    .ZN(_03638_)
  );
  AND2_X1 _13906_ (
    .A1(_03636_),
    .A2(_03638_),
    .ZN(_03639_)
  );
  INV_X1 _13907_ (
    .A(_03639_),
    .ZN(_03640_)
  );
  AND2_X1 _13908_ (
    .A1(_03602_),
    .A2(_03639_),
    .ZN(_03641_)
  );
  INV_X1 _13909_ (
    .A(_03641_),
    .ZN(_03642_)
  );
  AND2_X1 _13910_ (
    .A1(_03601_),
    .A2(_03640_),
    .ZN(_03643_)
  );
  INV_X1 _13911_ (
    .A(_03643_),
    .ZN(_03644_)
  );
  AND2_X1 _13912_ (
    .A1(_03642_),
    .A2(_03644_),
    .ZN(_03645_)
  );
  INV_X1 _13913_ (
    .A(_03645_),
    .ZN(_03646_)
  );
  AND2_X1 _13914_ (
    .A1(_03506_),
    .A2(_03645_),
    .ZN(_03647_)
  );
  INV_X1 _13915_ (
    .A(_03647_),
    .ZN(_03648_)
  );
  AND2_X1 _13916_ (
    .A1(_03507_),
    .A2(_03646_),
    .ZN(_03649_)
  );
  INV_X1 _13917_ (
    .A(_03649_),
    .ZN(_03650_)
  );
  AND2_X1 _13918_ (
    .A1(_03648_),
    .A2(_03650_),
    .ZN(_03651_)
  );
  INV_X1 _13919_ (
    .A(_03651_),
    .ZN(_03652_)
  );
  AND2_X1 _13920_ (
    .A1(_03600_),
    .A2(_03651_),
    .ZN(_03653_)
  );
  INV_X1 _13921_ (
    .A(_03653_),
    .ZN(_03654_)
  );
  AND2_X1 _13922_ (
    .A1(_03599_),
    .A2(_03652_),
    .ZN(_03655_)
  );
  INV_X1 _13923_ (
    .A(_03655_),
    .ZN(_03656_)
  );
  AND2_X1 _13924_ (
    .A1(_03654_),
    .A2(_03656_),
    .ZN(_03657_)
  );
  INV_X1 _13925_ (
    .A(_03657_),
    .ZN(_03658_)
  );
  AND2_X1 _13926_ (
    .A1(_03598_),
    .A2(_03657_),
    .ZN(_03659_)
  );
  INV_X1 _13927_ (
    .A(_03659_),
    .ZN(_03660_)
  );
  AND2_X1 _13928_ (
    .A1(_03597_),
    .A2(_03658_),
    .ZN(_03661_)
  );
  INV_X1 _13929_ (
    .A(_03661_),
    .ZN(_03662_)
  );
  AND2_X1 _13930_ (
    .A1(_03660_),
    .A2(_03662_),
    .ZN(_03663_)
  );
  INV_X1 _13931_ (
    .A(_03663_),
    .ZN(_03664_)
  );
  AND2_X1 _13932_ (
    .A1(_03170_),
    .A2(_03663_),
    .ZN(_03665_)
  );
  INV_X1 _13933_ (
    .A(_03665_),
    .ZN(_03666_)
  );
  AND2_X1 _13934_ (
    .A1(_03169_),
    .A2(_03664_),
    .ZN(_03667_)
  );
  INV_X1 _13935_ (
    .A(_03667_),
    .ZN(_03668_)
  );
  AND2_X1 _13936_ (
    .A1(_03666_),
    .A2(_03668_),
    .ZN(_03669_)
  );
  INV_X1 _13937_ (
    .A(_03669_),
    .ZN(_03670_)
  );
  AND2_X1 _13938_ (
    .A1(_03596_),
    .A2(_03669_),
    .ZN(_03671_)
  );
  INV_X1 _13939_ (
    .A(_03671_),
    .ZN(_03672_)
  );
  AND2_X1 _13940_ (
    .A1(_03595_),
    .A2(_03670_),
    .ZN(_03673_)
  );
  INV_X1 _13941_ (
    .A(_03673_),
    .ZN(_03674_)
  );
  AND2_X1 _13942_ (
    .A1(_03672_),
    .A2(_03674_),
    .ZN(_03675_)
  );
  INV_X1 _13943_ (
    .A(_03675_),
    .ZN(_03676_)
  );
  AND2_X1 _13944_ (
    .A1(divisor[13]),
    .A2(remainder[0]),
    .ZN(_03677_)
  );
  INV_X1 _13945_ (
    .A(_03677_),
    .ZN(_03678_)
  );
  AND2_X1 _13946_ (
    .A1(divisor[10]),
    .A2(remainder[3]),
    .ZN(_03679_)
  );
  INV_X1 _13947_ (
    .A(_03679_),
    .ZN(_03680_)
  );
  AND2_X1 _13948_ (
    .A1(divisor[11]),
    .A2(remainder[2]),
    .ZN(_03681_)
  );
  INV_X1 _13949_ (
    .A(_03681_),
    .ZN(_03682_)
  );
  AND2_X1 _13950_ (
    .A1(divisor[12]),
    .A2(remainder[2]),
    .ZN(_03683_)
  );
  INV_X1 _13951_ (
    .A(_03683_),
    .ZN(_03684_)
  );
  AND2_X1 _13952_ (
    .A1(_03255_),
    .A2(_03683_),
    .ZN(_03685_)
  );
  INV_X1 _13953_ (
    .A(_03685_),
    .ZN(_03686_)
  );
  AND2_X1 _13954_ (
    .A1(_03461_),
    .A2(_03682_),
    .ZN(_03687_)
  );
  INV_X1 _13955_ (
    .A(_03687_),
    .ZN(_03688_)
  );
  AND2_X1 _13956_ (
    .A1(_03686_),
    .A2(_03688_),
    .ZN(_03689_)
  );
  INV_X1 _13957_ (
    .A(_03689_),
    .ZN(_03690_)
  );
  AND2_X1 _13958_ (
    .A1(_03679_),
    .A2(_03689_),
    .ZN(_03691_)
  );
  INV_X1 _13959_ (
    .A(_03691_),
    .ZN(_03692_)
  );
  AND2_X1 _13960_ (
    .A1(_03680_),
    .A2(_03690_),
    .ZN(_03693_)
  );
  INV_X1 _13961_ (
    .A(_03693_),
    .ZN(_03694_)
  );
  AND2_X1 _13962_ (
    .A1(_03692_),
    .A2(_03694_),
    .ZN(_03695_)
  );
  INV_X1 _13963_ (
    .A(_03695_),
    .ZN(_03696_)
  );
  AND2_X1 _13964_ (
    .A1(_03677_),
    .A2(_03695_),
    .ZN(_03697_)
  );
  INV_X1 _13965_ (
    .A(_03697_),
    .ZN(_03698_)
  );
  AND2_X1 _13966_ (
    .A1(_03678_),
    .A2(_03696_),
    .ZN(_03699_)
  );
  INV_X1 _13967_ (
    .A(_03699_),
    .ZN(_03700_)
  );
  AND2_X1 _13968_ (
    .A1(_03698_),
    .A2(_03700_),
    .ZN(_03701_)
  );
  INV_X1 _13969_ (
    .A(_03701_),
    .ZN(_03702_)
  );
  AND2_X1 _13970_ (
    .A1(_03483_),
    .A2(_03489_),
    .ZN(_03703_)
  );
  INV_X1 _13971_ (
    .A(_03703_),
    .ZN(_03704_)
  );
  AND2_X1 _13972_ (
    .A1(_03463_),
    .A2(_03469_),
    .ZN(_03705_)
  );
  INV_X1 _13973_ (
    .A(_03705_),
    .ZN(_03706_)
  );
  AND2_X1 _13974_ (
    .A1(divisor[7]),
    .A2(remainder[6]),
    .ZN(_03707_)
  );
  INV_X1 _13975_ (
    .A(_03707_),
    .ZN(_03708_)
  );
  AND2_X1 _13976_ (
    .A1(divisor[8]),
    .A2(remainder[5]),
    .ZN(_03709_)
  );
  INV_X1 _13977_ (
    .A(_03709_),
    .ZN(_03710_)
  );
  AND2_X1 _13978_ (
    .A1(divisor[9]),
    .A2(remainder[5]),
    .ZN(_03711_)
  );
  INV_X1 _13979_ (
    .A(_03711_),
    .ZN(_03712_)
  );
  AND2_X1 _13980_ (
    .A1(_03480_),
    .A2(_03709_),
    .ZN(_03713_)
  );
  INV_X1 _13981_ (
    .A(_03713_),
    .ZN(_03714_)
  );
  AND2_X1 _13982_ (
    .A1(_03481_),
    .A2(_03710_),
    .ZN(_03715_)
  );
  INV_X1 _13983_ (
    .A(_03715_),
    .ZN(_03716_)
  );
  AND2_X1 _13984_ (
    .A1(_03714_),
    .A2(_03716_),
    .ZN(_03717_)
  );
  INV_X1 _13985_ (
    .A(_03717_),
    .ZN(_03718_)
  );
  AND2_X1 _13986_ (
    .A1(_03707_),
    .A2(_03717_),
    .ZN(_03719_)
  );
  INV_X1 _13987_ (
    .A(_03719_),
    .ZN(_03720_)
  );
  AND2_X1 _13988_ (
    .A1(_03708_),
    .A2(_03718_),
    .ZN(_03721_)
  );
  INV_X1 _13989_ (
    .A(_03721_),
    .ZN(_03722_)
  );
  AND2_X1 _13990_ (
    .A1(_03720_),
    .A2(_03722_),
    .ZN(_03723_)
  );
  INV_X1 _13991_ (
    .A(_03723_),
    .ZN(_03724_)
  );
  AND2_X1 _13992_ (
    .A1(_03706_),
    .A2(_03723_),
    .ZN(_03725_)
  );
  INV_X1 _13993_ (
    .A(_03725_),
    .ZN(_03726_)
  );
  AND2_X1 _13994_ (
    .A1(_03705_),
    .A2(_03724_),
    .ZN(_03727_)
  );
  INV_X1 _13995_ (
    .A(_03727_),
    .ZN(_03728_)
  );
  AND2_X1 _13996_ (
    .A1(_03726_),
    .A2(_03728_),
    .ZN(_03729_)
  );
  INV_X1 _13997_ (
    .A(_03729_),
    .ZN(_03730_)
  );
  AND2_X1 _13998_ (
    .A1(_03704_),
    .A2(_03729_),
    .ZN(_03731_)
  );
  INV_X1 _13999_ (
    .A(_03731_),
    .ZN(_03732_)
  );
  AND2_X1 _14000_ (
    .A1(_03703_),
    .A2(_03730_),
    .ZN(_03733_)
  );
  INV_X1 _14001_ (
    .A(_03733_),
    .ZN(_03734_)
  );
  AND2_X1 _14002_ (
    .A1(_03732_),
    .A2(_03734_),
    .ZN(_03735_)
  );
  INV_X1 _14003_ (
    .A(_03735_),
    .ZN(_03736_)
  );
  AND2_X1 _14004_ (
    .A1(_03701_),
    .A2(_03735_),
    .ZN(_03737_)
  );
  INV_X1 _14005_ (
    .A(_03737_),
    .ZN(_03738_)
  );
  AND2_X1 _14006_ (
    .A1(_03702_),
    .A2(_03736_),
    .ZN(_03739_)
  );
  INV_X1 _14007_ (
    .A(_03739_),
    .ZN(_03740_)
  );
  AND2_X1 _14008_ (
    .A1(_03738_),
    .A2(_03740_),
    .ZN(_03741_)
  );
  INV_X1 _14009_ (
    .A(_03741_),
    .ZN(_03742_)
  );
  AND2_X1 _14010_ (
    .A1(_03589_),
    .A2(_03742_),
    .ZN(_03743_)
  );
  INV_X1 _14011_ (
    .A(_03743_),
    .ZN(_03744_)
  );
  AND2_X1 _14012_ (
    .A1(_03590_),
    .A2(_03741_),
    .ZN(_03745_)
  );
  INV_X1 _14013_ (
    .A(_03745_),
    .ZN(_03746_)
  );
  AND2_X1 _14014_ (
    .A1(_03590_),
    .A2(_03742_),
    .ZN(_03747_)
  );
  INV_X1 _14015_ (
    .A(_03747_),
    .ZN(_03748_)
  );
  AND2_X1 _14016_ (
    .A1(_03589_),
    .A2(_03741_),
    .ZN(_03749_)
  );
  INV_X1 _14017_ (
    .A(_03749_),
    .ZN(_03750_)
  );
  AND2_X1 _14018_ (
    .A1(_03744_),
    .A2(_03746_),
    .ZN(_03751_)
  );
  AND2_X1 _14019_ (
    .A1(_03748_),
    .A2(_03750_),
    .ZN(_03752_)
  );
  AND2_X1 _14020_ (
    .A1(_03675_),
    .A2(_03752_),
    .ZN(_03753_)
  );
  INV_X1 _14021_ (
    .A(_03753_),
    .ZN(_03754_)
  );
  AND2_X1 _14022_ (
    .A1(_03676_),
    .A2(_03751_),
    .ZN(_03755_)
  );
  INV_X1 _14023_ (
    .A(_03755_),
    .ZN(_03756_)
  );
  AND2_X1 _14024_ (
    .A1(_03754_),
    .A2(_03756_),
    .ZN(_03757_)
  );
  INV_X1 _14025_ (
    .A(_03757_),
    .ZN(_03758_)
  );
  AND2_X1 _14026_ (
    .A1(_03594_),
    .A2(_03757_),
    .ZN(_03759_)
  );
  INV_X1 _14027_ (
    .A(_03759_),
    .ZN(_03760_)
  );
  AND2_X1 _14028_ (
    .A1(_03593_),
    .A2(_03758_),
    .ZN(_03761_)
  );
  INV_X1 _14029_ (
    .A(_03761_),
    .ZN(_03762_)
  );
  AND2_X1 _14030_ (
    .A1(_03760_),
    .A2(_03762_),
    .ZN(_03763_)
  );
  INV_X1 _14031_ (
    .A(_03763_),
    .ZN(_03764_)
  );
  AND2_X1 _14032_ (
    .A1(_03450_),
    .A2(_03763_),
    .ZN(_03765_)
  );
  INV_X1 _14033_ (
    .A(_03765_),
    .ZN(_03766_)
  );
  AND2_X1 _14034_ (
    .A1(_03451_),
    .A2(_03764_),
    .ZN(_03767_)
  );
  INV_X1 _14035_ (
    .A(_03767_),
    .ZN(_03768_)
  );
  AND2_X1 _14036_ (
    .A1(_03766_),
    .A2(_03768_),
    .ZN(_03769_)
  );
  INV_X1 _14037_ (
    .A(_03769_),
    .ZN(_03770_)
  );
  AND2_X1 _14038_ (
    .A1(_03588_),
    .A2(_03769_),
    .ZN(_03771_)
  );
  INV_X1 _14039_ (
    .A(_03771_),
    .ZN(_03772_)
  );
  AND2_X1 _14040_ (
    .A1(_03587_),
    .A2(_03770_),
    .ZN(_03773_)
  );
  INV_X1 _14041_ (
    .A(_03773_),
    .ZN(_03774_)
  );
  AND2_X1 _14042_ (
    .A1(_03772_),
    .A2(_03774_),
    .ZN(_03775_)
  );
  INV_X1 _14043_ (
    .A(_03775_),
    .ZN(_03776_)
  );
  AND2_X1 _14044_ (
    .A1(_03540_),
    .A2(_03775_),
    .ZN(_03777_)
  );
  INV_X1 _14045_ (
    .A(_03777_),
    .ZN(_03778_)
  );
  AND2_X1 _14046_ (
    .A1(_03541_),
    .A2(_03776_),
    .ZN(_03779_)
  );
  INV_X1 _14047_ (
    .A(_03779_),
    .ZN(_03780_)
  );
  AND2_X1 _14048_ (
    .A1(_03778_),
    .A2(_03780_),
    .ZN(_03781_)
  );
  INV_X1 _14049_ (
    .A(_03781_),
    .ZN(_03782_)
  );
  AND2_X1 _14050_ (
    .A1(_03585_),
    .A2(_03782_),
    .ZN(_03783_)
  );
  INV_X1 _14051_ (
    .A(_03783_),
    .ZN(_03784_)
  );
  AND2_X1 _14052_ (
    .A1(_03586_),
    .A2(_03781_),
    .ZN(_03785_)
  );
  INV_X1 _14053_ (
    .A(_03785_),
    .ZN(_03786_)
  );
  AND2_X1 _14054_ (
    .A1(_03784_),
    .A2(_03786_),
    .ZN(_03787_)
  );
  INV_X1 _14055_ (
    .A(_03787_),
    .ZN(_03788_)
  );
  AND2_X1 _14056_ (
    .A1(remainder[46]),
    .A2(_03787_),
    .ZN(_03789_)
  );
  INV_X1 _14057_ (
    .A(_03789_),
    .ZN(_03790_)
  );
  AND2_X1 _14058_ (
    .A1(_04612_),
    .A2(_03788_),
    .ZN(_03791_)
  );
  INV_X1 _14059_ (
    .A(_03791_),
    .ZN(_03792_)
  );
  AND2_X1 _14060_ (
    .A1(_03790_),
    .A2(_03792_),
    .ZN(_03793_)
  );
  INV_X1 _14061_ (
    .A(_03793_),
    .ZN(_03794_)
  );
  AND2_X1 _14062_ (
    .A1(_03584_),
    .A2(_03793_),
    .ZN(_03795_)
  );
  INV_X1 _14063_ (
    .A(_03795_),
    .ZN(_03796_)
  );
  AND2_X1 _14064_ (
    .A1(_03583_),
    .A2(_03794_),
    .ZN(_03797_)
  );
  INV_X1 _14065_ (
    .A(_03797_),
    .ZN(_03798_)
  );
  AND2_X1 _14066_ (
    .A1(_03796_),
    .A2(_03798_),
    .ZN(_03799_)
  );
  AND2_X1 _14067_ (
    .A1(_02082_),
    .A2(_03799_),
    .ZN(_03800_)
  );
  INV_X1 _14068_ (
    .A(_03800_),
    .ZN(_03801_)
  );
  AND2_X1 _14069_ (
    .A1(_03582_),
    .A2(_03801_),
    .ZN(_03802_)
  );
  AND2_X1 _14070_ (
    .A1(_03580_),
    .A2(_03802_),
    .ZN(_03803_)
  );
  INV_X1 _14071_ (
    .A(_03803_),
    .ZN(_03804_)
  );
  AND2_X1 _14072_ (
    .A1(_06201_),
    .A2(_03804_),
    .ZN(_00059_)
  );
  AND2_X1 _14073_ (
    .A1(_04700_),
    .A2(_10451_),
    .ZN(_03805_)
  );
  INV_X1 _14074_ (
    .A(_03805_),
    .ZN(_03806_)
  );
  AND2_X1 _14075_ (
    .A1(_10462_),
    .A2(_01136_),
    .ZN(_03807_)
  );
  INV_X1 _14076_ (
    .A(_03807_),
    .ZN(_03808_)
  );
  AND2_X1 _14077_ (
    .A1(_05983_),
    .A2(_03808_),
    .ZN(_03809_)
  );
  AND2_X1 _14078_ (
    .A1(_03806_),
    .A2(_03809_),
    .ZN(_03810_)
  );
  INV_X1 _14079_ (
    .A(_03810_),
    .ZN(_03811_)
  );
  AND2_X1 _14080_ (
    .A1(remainder[39]),
    .A2(_02077_),
    .ZN(_03812_)
  );
  INV_X1 _14081_ (
    .A(_03812_),
    .ZN(_03813_)
  );
  AND2_X1 _14082_ (
    .A1(_03760_),
    .A2(_03766_),
    .ZN(_03814_)
  );
  INV_X1 _14083_ (
    .A(_03814_),
    .ZN(_03815_)
  );
  AND2_X1 _14084_ (
    .A1(_03249_),
    .A2(_03742_),
    .ZN(_03816_)
  );
  INV_X1 _14085_ (
    .A(_03816_),
    .ZN(_03817_)
  );
  AND2_X1 _14086_ (
    .A1(_03510_),
    .A2(_03816_),
    .ZN(_03818_)
  );
  INV_X1 _14087_ (
    .A(_03818_),
    .ZN(_03819_)
  );
  AND2_X1 _14088_ (
    .A1(_03754_),
    .A2(_03819_),
    .ZN(_03820_)
  );
  INV_X1 _14089_ (
    .A(_03820_),
    .ZN(_03821_)
  );
  AND2_X1 _14090_ (
    .A1(_03660_),
    .A2(_03666_),
    .ZN(_03822_)
  );
  INV_X1 _14091_ (
    .A(_03822_),
    .ZN(_03823_)
  );
  AND2_X1 _14092_ (
    .A1(_03648_),
    .A2(_03654_),
    .ZN(_03824_)
  );
  INV_X1 _14093_ (
    .A(_03824_),
    .ZN(_03825_)
  );
  AND2_X1 _14094_ (
    .A1(_03636_),
    .A2(_03642_),
    .ZN(_03826_)
  );
  INV_X1 _14095_ (
    .A(_03826_),
    .ZN(_03827_)
  );
  AND2_X1 _14096_ (
    .A1(_03624_),
    .A2(_03630_),
    .ZN(_03828_)
  );
  INV_X1 _14097_ (
    .A(_03828_),
    .ZN(_03829_)
  );
  AND2_X1 _14098_ (
    .A1(_03726_),
    .A2(_03732_),
    .ZN(_03830_)
  );
  INV_X1 _14099_ (
    .A(_03830_),
    .ZN(_03831_)
  );
  AND2_X1 _14100_ (
    .A1(_03612_),
    .A2(_03618_),
    .ZN(_03832_)
  );
  INV_X1 _14101_ (
    .A(_03832_),
    .ZN(_03833_)
  );
  AND2_X1 _14102_ (
    .A1(_03608_),
    .A2(_03610_),
    .ZN(_03834_)
  );
  MUX2_X1 _14103_ (
    .A(_03609_),
    .B(_04886_),
    .S(_03607_),
    .Z(_03835_)
  );
  MUX2_X1 _14104_ (
    .A(_03384_),
    .B(_04875_),
    .S(_03835_),
    .Z(_03836_)
  );
  MUX2_X1 _14105_ (
    .A(_03385_),
    .B(divisor[4]),
    .S(_03835_),
    .Z(_03837_)
  );
  AND2_X1 _14106_ (
    .A1(_03833_),
    .A2(_03836_),
    .ZN(_03838_)
  );
  INV_X1 _14107_ (
    .A(_03838_),
    .ZN(_03839_)
  );
  AND2_X1 _14108_ (
    .A1(_03832_),
    .A2(_03837_),
    .ZN(_03840_)
  );
  INV_X1 _14109_ (
    .A(_03840_),
    .ZN(_03841_)
  );
  AND2_X1 _14110_ (
    .A1(_03839_),
    .A2(_03841_),
    .ZN(_03842_)
  );
  INV_X1 _14111_ (
    .A(_03842_),
    .ZN(_03843_)
  );
  AND2_X1 _14112_ (
    .A1(_03046_),
    .A2(_03842_),
    .ZN(_03844_)
  );
  INV_X1 _14113_ (
    .A(_03844_),
    .ZN(_03845_)
  );
  AND2_X1 _14114_ (
    .A1(_03047_),
    .A2(_03843_),
    .ZN(_03846_)
  );
  INV_X1 _14115_ (
    .A(_03846_),
    .ZN(_03847_)
  );
  AND2_X1 _14116_ (
    .A1(_03845_),
    .A2(_03847_),
    .ZN(_03848_)
  );
  INV_X1 _14117_ (
    .A(_03848_),
    .ZN(_03849_)
  );
  AND2_X1 _14118_ (
    .A1(_03831_),
    .A2(_03848_),
    .ZN(_03850_)
  );
  INV_X1 _14119_ (
    .A(_03850_),
    .ZN(_03851_)
  );
  AND2_X1 _14120_ (
    .A1(_03830_),
    .A2(_03849_),
    .ZN(_03852_)
  );
  INV_X1 _14121_ (
    .A(_03852_),
    .ZN(_03853_)
  );
  AND2_X1 _14122_ (
    .A1(_03851_),
    .A2(_03853_),
    .ZN(_03854_)
  );
  INV_X1 _14123_ (
    .A(_03854_),
    .ZN(_03855_)
  );
  AND2_X1 _14124_ (
    .A1(_03829_),
    .A2(_03854_),
    .ZN(_03856_)
  );
  INV_X1 _14125_ (
    .A(_03856_),
    .ZN(_03857_)
  );
  AND2_X1 _14126_ (
    .A1(_03828_),
    .A2(_03855_),
    .ZN(_03858_)
  );
  INV_X1 _14127_ (
    .A(_03858_),
    .ZN(_03859_)
  );
  AND2_X1 _14128_ (
    .A1(_03857_),
    .A2(_03859_),
    .ZN(_03860_)
  );
  INV_X1 _14129_ (
    .A(_03860_),
    .ZN(_03861_)
  );
  AND2_X1 _14130_ (
    .A1(_03737_),
    .A2(_03860_),
    .ZN(_03862_)
  );
  INV_X1 _14131_ (
    .A(_03862_),
    .ZN(_03863_)
  );
  AND2_X1 _14132_ (
    .A1(_03738_),
    .A2(_03861_),
    .ZN(_03864_)
  );
  INV_X1 _14133_ (
    .A(_03864_),
    .ZN(_03865_)
  );
  AND2_X1 _14134_ (
    .A1(_03863_),
    .A2(_03865_),
    .ZN(_03866_)
  );
  INV_X1 _14135_ (
    .A(_03866_),
    .ZN(_03867_)
  );
  AND2_X1 _14136_ (
    .A1(_03827_),
    .A2(_03866_),
    .ZN(_03868_)
  );
  INV_X1 _14137_ (
    .A(_03868_),
    .ZN(_03869_)
  );
  AND2_X1 _14138_ (
    .A1(_03826_),
    .A2(_03867_),
    .ZN(_03870_)
  );
  INV_X1 _14139_ (
    .A(_03870_),
    .ZN(_03871_)
  );
  AND2_X1 _14140_ (
    .A1(_03869_),
    .A2(_03871_),
    .ZN(_03872_)
  );
  INV_X1 _14141_ (
    .A(_03872_),
    .ZN(_03873_)
  );
  AND2_X1 _14142_ (
    .A1(_03825_),
    .A2(_03872_),
    .ZN(_03874_)
  );
  INV_X1 _14143_ (
    .A(_03874_),
    .ZN(_03875_)
  );
  AND2_X1 _14144_ (
    .A1(_03824_),
    .A2(_03873_),
    .ZN(_03876_)
  );
  INV_X1 _14145_ (
    .A(_03876_),
    .ZN(_03877_)
  );
  AND2_X1 _14146_ (
    .A1(_03875_),
    .A2(_03877_),
    .ZN(_03878_)
  );
  INV_X1 _14147_ (
    .A(_03878_),
    .ZN(_03879_)
  );
  AND2_X1 _14148_ (
    .A1(_03170_),
    .A2(_03878_),
    .ZN(_03880_)
  );
  INV_X1 _14149_ (
    .A(_03880_),
    .ZN(_03881_)
  );
  AND2_X1 _14150_ (
    .A1(_03169_),
    .A2(_03879_),
    .ZN(_03882_)
  );
  INV_X1 _14151_ (
    .A(_03882_),
    .ZN(_03883_)
  );
  AND2_X1 _14152_ (
    .A1(_03881_),
    .A2(_03883_),
    .ZN(_03884_)
  );
  INV_X1 _14153_ (
    .A(_03884_),
    .ZN(_03885_)
  );
  AND2_X1 _14154_ (
    .A1(_03823_),
    .A2(_03884_),
    .ZN(_03886_)
  );
  INV_X1 _14155_ (
    .A(_03886_),
    .ZN(_03887_)
  );
  AND2_X1 _14156_ (
    .A1(_03822_),
    .A2(_03885_),
    .ZN(_03888_)
  );
  INV_X1 _14157_ (
    .A(_03888_),
    .ZN(_03889_)
  );
  AND2_X1 _14158_ (
    .A1(_03887_),
    .A2(_03889_),
    .ZN(_03890_)
  );
  INV_X1 _14159_ (
    .A(_03890_),
    .ZN(_03891_)
  );
  AND2_X1 _14160_ (
    .A1(divisor[14]),
    .A2(remainder[0]),
    .ZN(_03892_)
  );
  INV_X1 _14161_ (
    .A(_03892_),
    .ZN(_03893_)
  );
  AND2_X1 _14162_ (
    .A1(divisor[13]),
    .A2(remainder[1]),
    .ZN(_03894_)
  );
  INV_X1 _14163_ (
    .A(_03894_),
    .ZN(_03895_)
  );
  AND2_X1 _14164_ (
    .A1(divisor[14]),
    .A2(remainder[1]),
    .ZN(_03896_)
  );
  INV_X1 _14165_ (
    .A(_03896_),
    .ZN(_03897_)
  );
  AND2_X1 _14166_ (
    .A1(_03677_),
    .A2(_03896_),
    .ZN(_03898_)
  );
  INV_X1 _14167_ (
    .A(_03898_),
    .ZN(_03899_)
  );
  AND2_X1 _14168_ (
    .A1(_03893_),
    .A2(_03895_),
    .ZN(_03900_)
  );
  INV_X1 _14169_ (
    .A(_03900_),
    .ZN(_03901_)
  );
  AND2_X1 _14170_ (
    .A1(_03899_),
    .A2(_03901_),
    .ZN(_03902_)
  );
  INV_X1 _14171_ (
    .A(_03902_),
    .ZN(_03903_)
  );
  AND2_X1 _14172_ (
    .A1(divisor[10]),
    .A2(remainder[4]),
    .ZN(_03904_)
  );
  INV_X1 _14173_ (
    .A(_03904_),
    .ZN(_03905_)
  );
  AND2_X1 _14174_ (
    .A1(divisor[11]),
    .A2(remainder[3]),
    .ZN(_03906_)
  );
  INV_X1 _14175_ (
    .A(_03906_),
    .ZN(_03907_)
  );
  AND2_X1 _14176_ (
    .A1(divisor[12]),
    .A2(remainder[3]),
    .ZN(_03908_)
  );
  INV_X1 _14177_ (
    .A(_03908_),
    .ZN(_03909_)
  );
  AND2_X1 _14178_ (
    .A1(_03683_),
    .A2(_03906_),
    .ZN(_03910_)
  );
  INV_X1 _14179_ (
    .A(_03910_),
    .ZN(_03911_)
  );
  AND2_X1 _14180_ (
    .A1(_03684_),
    .A2(_03907_),
    .ZN(_03912_)
  );
  INV_X1 _14181_ (
    .A(_03912_),
    .ZN(_03913_)
  );
  AND2_X1 _14182_ (
    .A1(_03911_),
    .A2(_03913_),
    .ZN(_03914_)
  );
  INV_X1 _14183_ (
    .A(_03914_),
    .ZN(_03915_)
  );
  AND2_X1 _14184_ (
    .A1(_03904_),
    .A2(_03914_),
    .ZN(_03916_)
  );
  INV_X1 _14185_ (
    .A(_03916_),
    .ZN(_03917_)
  );
  AND2_X1 _14186_ (
    .A1(_03905_),
    .A2(_03915_),
    .ZN(_03918_)
  );
  INV_X1 _14187_ (
    .A(_03918_),
    .ZN(_03919_)
  );
  AND2_X1 _14188_ (
    .A1(_03917_),
    .A2(_03919_),
    .ZN(_03920_)
  );
  INV_X1 _14189_ (
    .A(_03920_),
    .ZN(_03921_)
  );
  AND2_X1 _14190_ (
    .A1(_03902_),
    .A2(_03920_),
    .ZN(_03922_)
  );
  INV_X1 _14191_ (
    .A(_03922_),
    .ZN(_03923_)
  );
  AND2_X1 _14192_ (
    .A1(_03903_),
    .A2(_03921_),
    .ZN(_03924_)
  );
  INV_X1 _14193_ (
    .A(_03924_),
    .ZN(_03925_)
  );
  AND2_X1 _14194_ (
    .A1(_03923_),
    .A2(_03925_),
    .ZN(_03926_)
  );
  INV_X1 _14195_ (
    .A(_03926_),
    .ZN(_03927_)
  );
  AND2_X1 _14196_ (
    .A1(_03697_),
    .A2(_03926_),
    .ZN(_03928_)
  );
  INV_X1 _14197_ (
    .A(_03928_),
    .ZN(_03929_)
  );
  AND2_X1 _14198_ (
    .A1(_03698_),
    .A2(_03927_),
    .ZN(_03930_)
  );
  INV_X1 _14199_ (
    .A(_03930_),
    .ZN(_03931_)
  );
  AND2_X1 _14200_ (
    .A1(_03929_),
    .A2(_03931_),
    .ZN(_03932_)
  );
  INV_X1 _14201_ (
    .A(_03932_),
    .ZN(_03933_)
  );
  AND2_X1 _14202_ (
    .A1(_03714_),
    .A2(_03720_),
    .ZN(_03934_)
  );
  INV_X1 _14203_ (
    .A(_03934_),
    .ZN(_03935_)
  );
  AND2_X1 _14204_ (
    .A1(_03686_),
    .A2(_03692_),
    .ZN(_03936_)
  );
  INV_X1 _14205_ (
    .A(_03936_),
    .ZN(_03937_)
  );
  AND2_X1 _14206_ (
    .A1(divisor[7]),
    .A2(remainder[7]),
    .ZN(_03938_)
  );
  INV_X1 _14207_ (
    .A(_03938_),
    .ZN(_03939_)
  );
  AND2_X1 _14208_ (
    .A1(divisor[8]),
    .A2(remainder[6]),
    .ZN(_03940_)
  );
  INV_X1 _14209_ (
    .A(_03940_),
    .ZN(_03941_)
  );
  AND2_X1 _14210_ (
    .A1(divisor[9]),
    .A2(remainder[6]),
    .ZN(_03942_)
  );
  INV_X1 _14211_ (
    .A(_03942_),
    .ZN(_03943_)
  );
  AND2_X1 _14212_ (
    .A1(_03711_),
    .A2(_03940_),
    .ZN(_03944_)
  );
  INV_X1 _14213_ (
    .A(_03944_),
    .ZN(_03945_)
  );
  AND2_X1 _14214_ (
    .A1(_03712_),
    .A2(_03941_),
    .ZN(_03946_)
  );
  INV_X1 _14215_ (
    .A(_03946_),
    .ZN(_03947_)
  );
  AND2_X1 _14216_ (
    .A1(_03945_),
    .A2(_03947_),
    .ZN(_03948_)
  );
  INV_X1 _14217_ (
    .A(_03948_),
    .ZN(_03949_)
  );
  AND2_X1 _14218_ (
    .A1(_03938_),
    .A2(_03948_),
    .ZN(_03950_)
  );
  INV_X1 _14219_ (
    .A(_03950_),
    .ZN(_03951_)
  );
  AND2_X1 _14220_ (
    .A1(_03939_),
    .A2(_03949_),
    .ZN(_03952_)
  );
  INV_X1 _14221_ (
    .A(_03952_),
    .ZN(_03953_)
  );
  AND2_X1 _14222_ (
    .A1(_03951_),
    .A2(_03953_),
    .ZN(_03954_)
  );
  INV_X1 _14223_ (
    .A(_03954_),
    .ZN(_03955_)
  );
  AND2_X1 _14224_ (
    .A1(_03937_),
    .A2(_03954_),
    .ZN(_03956_)
  );
  INV_X1 _14225_ (
    .A(_03956_),
    .ZN(_03957_)
  );
  AND2_X1 _14226_ (
    .A1(_03936_),
    .A2(_03955_),
    .ZN(_03958_)
  );
  INV_X1 _14227_ (
    .A(_03958_),
    .ZN(_03959_)
  );
  AND2_X1 _14228_ (
    .A1(_03957_),
    .A2(_03959_),
    .ZN(_03960_)
  );
  INV_X1 _14229_ (
    .A(_03960_),
    .ZN(_03961_)
  );
  AND2_X1 _14230_ (
    .A1(_03935_),
    .A2(_03960_),
    .ZN(_03962_)
  );
  INV_X1 _14231_ (
    .A(_03962_),
    .ZN(_03963_)
  );
  AND2_X1 _14232_ (
    .A1(_03934_),
    .A2(_03961_),
    .ZN(_03964_)
  );
  INV_X1 _14233_ (
    .A(_03964_),
    .ZN(_03965_)
  );
  AND2_X1 _14234_ (
    .A1(_03963_),
    .A2(_03965_),
    .ZN(_03966_)
  );
  INV_X1 _14235_ (
    .A(_03966_),
    .ZN(_03967_)
  );
  AND2_X1 _14236_ (
    .A1(_03932_),
    .A2(_03966_),
    .ZN(_03968_)
  );
  INV_X1 _14237_ (
    .A(_03968_),
    .ZN(_03969_)
  );
  AND2_X1 _14238_ (
    .A1(_03933_),
    .A2(_03967_),
    .ZN(_03970_)
  );
  INV_X1 _14239_ (
    .A(_03970_),
    .ZN(_03971_)
  );
  AND2_X1 _14240_ (
    .A1(_03969_),
    .A2(_03971_),
    .ZN(_03972_)
  );
  INV_X1 _14241_ (
    .A(_03972_),
    .ZN(_03973_)
  );
  AND2_X1 _14242_ (
    .A1(_03816_),
    .A2(_03973_),
    .ZN(_03974_)
  );
  INV_X1 _14243_ (
    .A(_03974_),
    .ZN(_03975_)
  );
  AND2_X1 _14244_ (
    .A1(_03817_),
    .A2(_03972_),
    .ZN(_03976_)
  );
  INV_X1 _14245_ (
    .A(_03976_),
    .ZN(_03977_)
  );
  AND2_X1 _14246_ (
    .A1(_03817_),
    .A2(_03973_),
    .ZN(_03978_)
  );
  INV_X1 _14247_ (
    .A(_03978_),
    .ZN(_03979_)
  );
  AND2_X1 _14248_ (
    .A1(_03816_),
    .A2(_03972_),
    .ZN(_03980_)
  );
  INV_X1 _14249_ (
    .A(_03980_),
    .ZN(_03981_)
  );
  AND2_X1 _14250_ (
    .A1(_03975_),
    .A2(_03977_),
    .ZN(_03982_)
  );
  AND2_X1 _14251_ (
    .A1(_03979_),
    .A2(_03981_),
    .ZN(_03983_)
  );
  AND2_X1 _14252_ (
    .A1(_03890_),
    .A2(_03983_),
    .ZN(_03984_)
  );
  INV_X1 _14253_ (
    .A(_03984_),
    .ZN(_03985_)
  );
  AND2_X1 _14254_ (
    .A1(_03891_),
    .A2(_03982_),
    .ZN(_03986_)
  );
  INV_X1 _14255_ (
    .A(_03986_),
    .ZN(_03987_)
  );
  AND2_X1 _14256_ (
    .A1(_03985_),
    .A2(_03987_),
    .ZN(_03988_)
  );
  INV_X1 _14257_ (
    .A(_03988_),
    .ZN(_03989_)
  );
  AND2_X1 _14258_ (
    .A1(_03821_),
    .A2(_03988_),
    .ZN(_03990_)
  );
  INV_X1 _14259_ (
    .A(_03990_),
    .ZN(_03991_)
  );
  AND2_X1 _14260_ (
    .A1(_03820_),
    .A2(_03989_),
    .ZN(_03992_)
  );
  INV_X1 _14261_ (
    .A(_03992_),
    .ZN(_03993_)
  );
  AND2_X1 _14262_ (
    .A1(_03991_),
    .A2(_03993_),
    .ZN(_03994_)
  );
  INV_X1 _14263_ (
    .A(_03994_),
    .ZN(_03995_)
  );
  AND2_X1 _14264_ (
    .A1(_03671_),
    .A2(_03994_),
    .ZN(_03996_)
  );
  INV_X1 _14265_ (
    .A(_03996_),
    .ZN(_03997_)
  );
  AND2_X1 _14266_ (
    .A1(_03672_),
    .A2(_03995_),
    .ZN(_03998_)
  );
  INV_X1 _14267_ (
    .A(_03998_),
    .ZN(_03999_)
  );
  AND2_X1 _14268_ (
    .A1(_03997_),
    .A2(_03999_),
    .ZN(_04000_)
  );
  INV_X1 _14269_ (
    .A(_04000_),
    .ZN(_04001_)
  );
  AND2_X1 _14270_ (
    .A1(_03815_),
    .A2(_04000_),
    .ZN(_04002_)
  );
  INV_X1 _14271_ (
    .A(_04002_),
    .ZN(_04003_)
  );
  AND2_X1 _14272_ (
    .A1(_03814_),
    .A2(_04001_),
    .ZN(_04004_)
  );
  INV_X1 _14273_ (
    .A(_04004_),
    .ZN(_04005_)
  );
  AND2_X1 _14274_ (
    .A1(_04003_),
    .A2(_04005_),
    .ZN(_04006_)
  );
  INV_X1 _14275_ (
    .A(_04006_),
    .ZN(_04007_)
  );
  AND2_X1 _14276_ (
    .A1(_03771_),
    .A2(_04006_),
    .ZN(_04008_)
  );
  INV_X1 _14277_ (
    .A(_04008_),
    .ZN(_04009_)
  );
  AND2_X1 _14278_ (
    .A1(_03772_),
    .A2(_04007_),
    .ZN(_04010_)
  );
  INV_X1 _14279_ (
    .A(_04010_),
    .ZN(_04011_)
  );
  AND2_X1 _14280_ (
    .A1(_04009_),
    .A2(_04011_),
    .ZN(_04012_)
  );
  INV_X1 _14281_ (
    .A(_04012_),
    .ZN(_04013_)
  );
  AND2_X1 _14282_ (
    .A1(_03585_),
    .A2(_03778_),
    .ZN(_04014_)
  );
  INV_X1 _14283_ (
    .A(_04014_),
    .ZN(_04015_)
  );
  AND2_X1 _14284_ (
    .A1(_03778_),
    .A2(_03786_),
    .ZN(_04016_)
  );
  AND2_X1 _14285_ (
    .A1(_03780_),
    .A2(_04015_),
    .ZN(_04017_)
  );
  AND2_X1 _14286_ (
    .A1(_04012_),
    .A2(_04017_),
    .ZN(_04018_)
  );
  INV_X1 _14287_ (
    .A(_04018_),
    .ZN(_04019_)
  );
  AND2_X1 _14288_ (
    .A1(_04013_),
    .A2(_04016_),
    .ZN(_04020_)
  );
  INV_X1 _14289_ (
    .A(_04020_),
    .ZN(_04021_)
  );
  AND2_X1 _14290_ (
    .A1(_04019_),
    .A2(_04021_),
    .ZN(_04022_)
  );
  INV_X1 _14291_ (
    .A(_04022_),
    .ZN(_04023_)
  );
  AND2_X1 _14292_ (
    .A1(remainder[47]),
    .A2(_04022_),
    .ZN(_04024_)
  );
  INV_X1 _14293_ (
    .A(_04024_),
    .ZN(_04025_)
  );
  AND2_X1 _14294_ (
    .A1(_04601_),
    .A2(_04023_),
    .ZN(_04026_)
  );
  INV_X1 _14295_ (
    .A(_04026_),
    .ZN(_04027_)
  );
  AND2_X1 _14296_ (
    .A1(_04025_),
    .A2(_04027_),
    .ZN(_04028_)
  );
  INV_X1 _14297_ (
    .A(_04028_),
    .ZN(_04029_)
  );
  AND2_X1 _14298_ (
    .A1(_03583_),
    .A2(_03790_),
    .ZN(_04030_)
  );
  INV_X1 _14299_ (
    .A(_04030_),
    .ZN(_04031_)
  );
  AND2_X1 _14300_ (
    .A1(_03584_),
    .A2(_03792_),
    .ZN(_04032_)
  );
  INV_X1 _14301_ (
    .A(_04032_),
    .ZN(_04033_)
  );
  AND2_X1 _14302_ (
    .A1(_03792_),
    .A2(_04031_),
    .ZN(_04034_)
  );
  AND2_X1 _14303_ (
    .A1(_03790_),
    .A2(_04033_),
    .ZN(_04035_)
  );
  AND2_X1 _14304_ (
    .A1(_04028_),
    .A2(_04034_),
    .ZN(_04036_)
  );
  INV_X1 _14305_ (
    .A(_04036_),
    .ZN(_04037_)
  );
  AND2_X1 _14306_ (
    .A1(_04029_),
    .A2(_04035_),
    .ZN(_04038_)
  );
  INV_X1 _14307_ (
    .A(_04038_),
    .ZN(_04039_)
  );
  AND2_X1 _14308_ (
    .A1(_02082_),
    .A2(_04037_),
    .ZN(_04040_)
  );
  AND2_X1 _14309_ (
    .A1(_04039_),
    .A2(_04040_),
    .ZN(_04041_)
  );
  INV_X1 _14310_ (
    .A(_04041_),
    .ZN(_04042_)
  );
  AND2_X1 _14311_ (
    .A1(_03813_),
    .A2(_04042_),
    .ZN(_04043_)
  );
  AND2_X1 _14312_ (
    .A1(_03811_),
    .A2(_04043_),
    .ZN(_04044_)
  );
  INV_X1 _14313_ (
    .A(_04044_),
    .ZN(_04045_)
  );
  AND2_X1 _14314_ (
    .A1(_06201_),
    .A2(_04045_),
    .ZN(_00060_)
  );
  AND2_X1 _14315_ (
    .A1(_04689_),
    .A2(_10451_),
    .ZN(_04046_)
  );
  INV_X1 _14316_ (
    .A(_04046_),
    .ZN(_04047_)
  );
  AND2_X1 _14317_ (
    .A1(_10462_),
    .A2(_01298_),
    .ZN(_04048_)
  );
  INV_X1 _14318_ (
    .A(_04048_),
    .ZN(_04049_)
  );
  AND2_X1 _14319_ (
    .A1(_05983_),
    .A2(_04049_),
    .ZN(_04050_)
  );
  AND2_X1 _14320_ (
    .A1(_04047_),
    .A2(_04050_),
    .ZN(_04051_)
  );
  INV_X1 _14321_ (
    .A(_04051_),
    .ZN(_04052_)
  );
  AND2_X1 _14322_ (
    .A1(remainder[40]),
    .A2(_02077_),
    .ZN(_04053_)
  );
  INV_X1 _14323_ (
    .A(_04053_),
    .ZN(_04054_)
  );
  AND2_X1 _14324_ (
    .A1(_04025_),
    .A2(_04037_),
    .ZN(_04055_)
  );
  INV_X1 _14325_ (
    .A(_04055_),
    .ZN(_04056_)
  );
  AND2_X1 _14326_ (
    .A1(_04009_),
    .A2(_04019_),
    .ZN(_04057_)
  );
  INV_X1 _14327_ (
    .A(_04057_),
    .ZN(_04058_)
  );
  AND2_X1 _14328_ (
    .A1(_03991_),
    .A2(_03997_),
    .ZN(_04059_)
  );
  INV_X1 _14329_ (
    .A(_04059_),
    .ZN(_04060_)
  );
  AND2_X1 _14330_ (
    .A1(_03249_),
    .A2(_03973_),
    .ZN(_04061_)
  );
  INV_X1 _14331_ (
    .A(_04061_),
    .ZN(_04062_)
  );
  AND2_X1 _14332_ (
    .A1(_03741_),
    .A2(_04061_),
    .ZN(_04063_)
  );
  INV_X1 _14333_ (
    .A(_04063_),
    .ZN(_04064_)
  );
  AND2_X1 _14334_ (
    .A1(_03985_),
    .A2(_04064_),
    .ZN(_04065_)
  );
  INV_X1 _14335_ (
    .A(_04065_),
    .ZN(_04066_)
  );
  AND2_X1 _14336_ (
    .A1(_03875_),
    .A2(_03881_),
    .ZN(_04067_)
  );
  INV_X1 _14337_ (
    .A(_04067_),
    .ZN(_04068_)
  );
  AND2_X1 _14338_ (
    .A1(_03863_),
    .A2(_03869_),
    .ZN(_04069_)
  );
  INV_X1 _14339_ (
    .A(_04069_),
    .ZN(_04070_)
  );
  AND2_X1 _14340_ (
    .A1(_03851_),
    .A2(_03857_),
    .ZN(_04071_)
  );
  INV_X1 _14341_ (
    .A(_04071_),
    .ZN(_04072_)
  );
  AND2_X1 _14342_ (
    .A1(_03929_),
    .A2(_03969_),
    .ZN(_04073_)
  );
  INV_X1 _14343_ (
    .A(_04073_),
    .ZN(_04074_)
  );
  AND2_X1 _14344_ (
    .A1(_03839_),
    .A2(_03845_),
    .ZN(_04075_)
  );
  INV_X1 _14345_ (
    .A(_04075_),
    .ZN(_04076_)
  );
  AND2_X1 _14346_ (
    .A1(_03957_),
    .A2(_03963_),
    .ZN(_04077_)
  );
  INV_X1 _14347_ (
    .A(_04077_),
    .ZN(_04078_)
  );
  AND2_X1 _14348_ (
    .A1(_03385_),
    .A2(_03834_),
    .ZN(_04079_)
  );
  INV_X1 _14349_ (
    .A(_04079_),
    .ZN(_04080_)
  );
  AND2_X1 _14350_ (
    .A1(_03839_),
    .A2(_04080_),
    .ZN(_04081_)
  );
  INV_X1 _14351_ (
    .A(_04081_),
    .ZN(_04082_)
  );
  AND2_X1 _14352_ (
    .A1(_03046_),
    .A2(_04081_),
    .ZN(_04083_)
  );
  INV_X1 _14353_ (
    .A(_04083_),
    .ZN(_04084_)
  );
  AND2_X1 _14354_ (
    .A1(_03047_),
    .A2(_04082_),
    .ZN(_04085_)
  );
  INV_X1 _14355_ (
    .A(_04085_),
    .ZN(_04086_)
  );
  AND2_X1 _14356_ (
    .A1(_04084_),
    .A2(_04086_),
    .ZN(_04087_)
  );
  INV_X1 _14357_ (
    .A(_04087_),
    .ZN(_04088_)
  );
  AND2_X1 _14358_ (
    .A1(_04078_),
    .A2(_04087_),
    .ZN(_04089_)
  );
  INV_X1 _14359_ (
    .A(_04089_),
    .ZN(_04090_)
  );
  AND2_X1 _14360_ (
    .A1(_04077_),
    .A2(_04088_),
    .ZN(_04091_)
  );
  INV_X1 _14361_ (
    .A(_04091_),
    .ZN(_04092_)
  );
  AND2_X1 _14362_ (
    .A1(_04090_),
    .A2(_04092_),
    .ZN(_04093_)
  );
  INV_X1 _14363_ (
    .A(_04093_),
    .ZN(_04094_)
  );
  AND2_X1 _14364_ (
    .A1(_04076_),
    .A2(_04093_),
    .ZN(_04095_)
  );
  INV_X1 _14365_ (
    .A(_04095_),
    .ZN(_04096_)
  );
  AND2_X1 _14366_ (
    .A1(_04075_),
    .A2(_04094_),
    .ZN(_04097_)
  );
  INV_X1 _14367_ (
    .A(_04097_),
    .ZN(_04098_)
  );
  AND2_X1 _14368_ (
    .A1(_04096_),
    .A2(_04098_),
    .ZN(_04099_)
  );
  INV_X1 _14369_ (
    .A(_04099_),
    .ZN(_04100_)
  );
  AND2_X1 _14370_ (
    .A1(_04074_),
    .A2(_04099_),
    .ZN(_04101_)
  );
  INV_X1 _14371_ (
    .A(_04101_),
    .ZN(_04102_)
  );
  AND2_X1 _14372_ (
    .A1(_04073_),
    .A2(_04100_),
    .ZN(_04103_)
  );
  INV_X1 _14373_ (
    .A(_04103_),
    .ZN(_04104_)
  );
  AND2_X1 _14374_ (
    .A1(_04102_),
    .A2(_04104_),
    .ZN(_04105_)
  );
  INV_X1 _14375_ (
    .A(_04105_),
    .ZN(_04106_)
  );
  AND2_X1 _14376_ (
    .A1(_04072_),
    .A2(_04105_),
    .ZN(_04107_)
  );
  INV_X1 _14377_ (
    .A(_04107_),
    .ZN(_04108_)
  );
  AND2_X1 _14378_ (
    .A1(_04071_),
    .A2(_04106_),
    .ZN(_04109_)
  );
  INV_X1 _14379_ (
    .A(_04109_),
    .ZN(_04110_)
  );
  AND2_X1 _14380_ (
    .A1(_04108_),
    .A2(_04110_),
    .ZN(_04111_)
  );
  INV_X1 _14381_ (
    .A(_04111_),
    .ZN(_04112_)
  );
  AND2_X1 _14382_ (
    .A1(_04070_),
    .A2(_04111_),
    .ZN(_04113_)
  );
  INV_X1 _14383_ (
    .A(_04113_),
    .ZN(_04114_)
  );
  AND2_X1 _14384_ (
    .A1(_04069_),
    .A2(_04112_),
    .ZN(_04115_)
  );
  INV_X1 _14385_ (
    .A(_04115_),
    .ZN(_04116_)
  );
  AND2_X1 _14386_ (
    .A1(_04114_),
    .A2(_04116_),
    .ZN(_04117_)
  );
  INV_X1 _14387_ (
    .A(_04117_),
    .ZN(_04118_)
  );
  AND2_X1 _14388_ (
    .A1(_03170_),
    .A2(_04117_),
    .ZN(_04119_)
  );
  INV_X1 _14389_ (
    .A(_04119_),
    .ZN(_04120_)
  );
  AND2_X1 _14390_ (
    .A1(_03169_),
    .A2(_04118_),
    .ZN(_04121_)
  );
  INV_X1 _14391_ (
    .A(_04121_),
    .ZN(_04122_)
  );
  AND2_X1 _14392_ (
    .A1(_04120_),
    .A2(_04122_),
    .ZN(_04123_)
  );
  INV_X1 _14393_ (
    .A(_04123_),
    .ZN(_04124_)
  );
  AND2_X1 _14394_ (
    .A1(_04068_),
    .A2(_04123_),
    .ZN(_04125_)
  );
  INV_X1 _14395_ (
    .A(_04125_),
    .ZN(_04126_)
  );
  AND2_X1 _14396_ (
    .A1(_04067_),
    .A2(_04124_),
    .ZN(_04127_)
  );
  INV_X1 _14397_ (
    .A(_04127_),
    .ZN(_04128_)
  );
  AND2_X1 _14398_ (
    .A1(_04126_),
    .A2(_04128_),
    .ZN(_04129_)
  );
  INV_X1 _14399_ (
    .A(_04129_),
    .ZN(_04130_)
  );
  AND2_X1 _14400_ (
    .A1(divisor[13]),
    .A2(remainder[2]),
    .ZN(_04131_)
  );
  INV_X1 _14401_ (
    .A(_04131_),
    .ZN(_04132_)
  );
  AND2_X1 _14402_ (
    .A1(divisor[15]),
    .A2(remainder[0]),
    .ZN(_04133_)
  );
  INV_X1 _14403_ (
    .A(_04133_),
    .ZN(_04134_)
  );
  AND2_X1 _14404_ (
    .A1(divisor[15]),
    .A2(remainder[1]),
    .ZN(_04135_)
  );
  INV_X1 _14405_ (
    .A(_04135_),
    .ZN(_04136_)
  );
  AND2_X1 _14406_ (
    .A1(_03892_),
    .A2(_04135_),
    .ZN(_04137_)
  );
  INV_X1 _14407_ (
    .A(_04137_),
    .ZN(_04138_)
  );
  AND2_X1 _14408_ (
    .A1(_03897_),
    .A2(_04134_),
    .ZN(_04139_)
  );
  INV_X1 _14409_ (
    .A(_04139_),
    .ZN(_04140_)
  );
  AND2_X1 _14410_ (
    .A1(_04138_),
    .A2(_04140_),
    .ZN(_04141_)
  );
  INV_X1 _14411_ (
    .A(_04141_),
    .ZN(_04142_)
  );
  AND2_X1 _14412_ (
    .A1(_04131_),
    .A2(_04141_),
    .ZN(_04143_)
  );
  INV_X1 _14413_ (
    .A(_04143_),
    .ZN(_04144_)
  );
  AND2_X1 _14414_ (
    .A1(_04132_),
    .A2(_04142_),
    .ZN(_04145_)
  );
  INV_X1 _14415_ (
    .A(_04145_),
    .ZN(_04146_)
  );
  AND2_X1 _14416_ (
    .A1(_04144_),
    .A2(_04146_),
    .ZN(_04147_)
  );
  INV_X1 _14417_ (
    .A(_04147_),
    .ZN(_04148_)
  );
  AND2_X1 _14418_ (
    .A1(_03898_),
    .A2(_04147_),
    .ZN(_04149_)
  );
  INV_X1 _14419_ (
    .A(_04149_),
    .ZN(_04150_)
  );
  AND2_X1 _14420_ (
    .A1(_03899_),
    .A2(_04148_),
    .ZN(_04151_)
  );
  INV_X1 _14421_ (
    .A(_04151_),
    .ZN(_04152_)
  );
  AND2_X1 _14422_ (
    .A1(_04150_),
    .A2(_04152_),
    .ZN(_04153_)
  );
  INV_X1 _14423_ (
    .A(_04153_),
    .ZN(_04154_)
  );
  AND2_X1 _14424_ (
    .A1(divisor[10]),
    .A2(remainder[5]),
    .ZN(_04155_)
  );
  INV_X1 _14425_ (
    .A(_04155_),
    .ZN(_04156_)
  );
  AND2_X1 _14426_ (
    .A1(divisor[11]),
    .A2(remainder[4]),
    .ZN(_04157_)
  );
  INV_X1 _14427_ (
    .A(_04157_),
    .ZN(_04158_)
  );
  AND2_X1 _14428_ (
    .A1(divisor[12]),
    .A2(remainder[4]),
    .ZN(_04159_)
  );
  INV_X1 _14429_ (
    .A(_04159_),
    .ZN(_04160_)
  );
  AND2_X1 _14430_ (
    .A1(_03908_),
    .A2(_04157_),
    .ZN(_04161_)
  );
  INV_X1 _14431_ (
    .A(_04161_),
    .ZN(_04162_)
  );
  AND2_X1 _14432_ (
    .A1(_03909_),
    .A2(_04158_),
    .ZN(_04163_)
  );
  INV_X1 _14433_ (
    .A(_04163_),
    .ZN(_04164_)
  );
  AND2_X1 _14434_ (
    .A1(_04162_),
    .A2(_04164_),
    .ZN(_04165_)
  );
  INV_X1 _14435_ (
    .A(_04165_),
    .ZN(_04166_)
  );
  AND2_X1 _14436_ (
    .A1(_04155_),
    .A2(_04165_),
    .ZN(_04167_)
  );
  INV_X1 _14437_ (
    .A(_04167_),
    .ZN(_04168_)
  );
  AND2_X1 _14438_ (
    .A1(_04156_),
    .A2(_04166_),
    .ZN(_04169_)
  );
  INV_X1 _14439_ (
    .A(_04169_),
    .ZN(_04170_)
  );
  AND2_X1 _14440_ (
    .A1(_04168_),
    .A2(_04170_),
    .ZN(_04171_)
  );
  INV_X1 _14441_ (
    .A(_04171_),
    .ZN(_04172_)
  );
  AND2_X1 _14442_ (
    .A1(_04153_),
    .A2(_04171_),
    .ZN(_04173_)
  );
  INV_X1 _14443_ (
    .A(_04173_),
    .ZN(_04174_)
  );
  AND2_X1 _14444_ (
    .A1(_04154_),
    .A2(_04172_),
    .ZN(_04175_)
  );
  INV_X1 _14445_ (
    .A(_04175_),
    .ZN(_04176_)
  );
  AND2_X1 _14446_ (
    .A1(_04174_),
    .A2(_04176_),
    .ZN(_04177_)
  );
  INV_X1 _14447_ (
    .A(_04177_),
    .ZN(_04178_)
  );
  AND2_X1 _14448_ (
    .A1(_03922_),
    .A2(_04177_),
    .ZN(_04179_)
  );
  INV_X1 _14449_ (
    .A(_04179_),
    .ZN(_04180_)
  );
  AND2_X1 _14450_ (
    .A1(_03923_),
    .A2(_04178_),
    .ZN(_04181_)
  );
  INV_X1 _14451_ (
    .A(_04181_),
    .ZN(_04182_)
  );
  AND2_X1 _14452_ (
    .A1(_04180_),
    .A2(_04182_),
    .ZN(_04183_)
  );
  INV_X1 _14453_ (
    .A(_04183_),
    .ZN(_04184_)
  );
  AND2_X1 _14454_ (
    .A1(_03945_),
    .A2(_03951_),
    .ZN(_04185_)
  );
  INV_X1 _14455_ (
    .A(_04185_),
    .ZN(_04186_)
  );
  AND2_X1 _14456_ (
    .A1(_03911_),
    .A2(_03917_),
    .ZN(_04187_)
  );
  INV_X1 _14457_ (
    .A(_04187_),
    .ZN(_04188_)
  );
  AND2_X1 _14458_ (
    .A1(remainder[32]),
    .A2(divisor[7]),
    .ZN(_04189_)
  );
  INV_X1 _14459_ (
    .A(_04189_),
    .ZN(_04190_)
  );
  AND2_X1 _14460_ (
    .A1(divisor[8]),
    .A2(remainder[7]),
    .ZN(_04191_)
  );
  INV_X1 _14461_ (
    .A(_04191_),
    .ZN(_04192_)
  );
  AND2_X1 _14462_ (
    .A1(divisor[9]),
    .A2(remainder[7]),
    .ZN(_04193_)
  );
  INV_X1 _14463_ (
    .A(_04193_),
    .ZN(_04194_)
  );
  AND2_X1 _14464_ (
    .A1(_03940_),
    .A2(_04193_),
    .ZN(_04195_)
  );
  INV_X1 _14465_ (
    .A(_04195_),
    .ZN(_04196_)
  );
  AND2_X1 _14466_ (
    .A1(_03943_),
    .A2(_04192_),
    .ZN(_04197_)
  );
  INV_X1 _14467_ (
    .A(_04197_),
    .ZN(_04198_)
  );
  AND2_X1 _14468_ (
    .A1(_04196_),
    .A2(_04198_),
    .ZN(_04199_)
  );
  INV_X1 _14469_ (
    .A(_04199_),
    .ZN(_04200_)
  );
  AND2_X1 _14470_ (
    .A1(_04189_),
    .A2(_04199_),
    .ZN(_04201_)
  );
  INV_X1 _14471_ (
    .A(_04201_),
    .ZN(_04202_)
  );
  AND2_X1 _14472_ (
    .A1(_04190_),
    .A2(_04200_),
    .ZN(_04203_)
  );
  INV_X1 _14473_ (
    .A(_04203_),
    .ZN(_04204_)
  );
  AND2_X1 _14474_ (
    .A1(_04202_),
    .A2(_04204_),
    .ZN(_04205_)
  );
  INV_X1 _14475_ (
    .A(_04205_),
    .ZN(_04206_)
  );
  AND2_X1 _14476_ (
    .A1(_04188_),
    .A2(_04205_),
    .ZN(_04207_)
  );
  INV_X1 _14477_ (
    .A(_04207_),
    .ZN(_04208_)
  );
  AND2_X1 _14478_ (
    .A1(_04187_),
    .A2(_04206_),
    .ZN(_04209_)
  );
  INV_X1 _14479_ (
    .A(_04209_),
    .ZN(_04210_)
  );
  AND2_X1 _14480_ (
    .A1(_04208_),
    .A2(_04210_),
    .ZN(_04211_)
  );
  INV_X1 _14481_ (
    .A(_04211_),
    .ZN(_04212_)
  );
  AND2_X1 _14482_ (
    .A1(_04186_),
    .A2(_04211_),
    .ZN(_04213_)
  );
  INV_X1 _14483_ (
    .A(_04213_),
    .ZN(_04214_)
  );
  AND2_X1 _14484_ (
    .A1(_04185_),
    .A2(_04212_),
    .ZN(_04215_)
  );
  INV_X1 _14485_ (
    .A(_04215_),
    .ZN(_04216_)
  );
  AND2_X1 _14486_ (
    .A1(_04214_),
    .A2(_04216_),
    .ZN(_04217_)
  );
  INV_X1 _14487_ (
    .A(_04217_),
    .ZN(_04218_)
  );
  AND2_X1 _14488_ (
    .A1(_04183_),
    .A2(_04217_),
    .ZN(_04219_)
  );
  INV_X1 _14489_ (
    .A(_04219_),
    .ZN(_04220_)
  );
  AND2_X1 _14490_ (
    .A1(_04184_),
    .A2(_04218_),
    .ZN(_04221_)
  );
  INV_X1 _14491_ (
    .A(_04221_),
    .ZN(_04222_)
  );
  AND2_X1 _14492_ (
    .A1(_04220_),
    .A2(_04222_),
    .ZN(_04223_)
  );
  INV_X1 _14493_ (
    .A(_04223_),
    .ZN(_04224_)
  );
  AND2_X1 _14494_ (
    .A1(_04062_),
    .A2(_04224_),
    .ZN(_04225_)
  );
  INV_X1 _14495_ (
    .A(_04225_),
    .ZN(_04226_)
  );
  AND2_X1 _14496_ (
    .A1(_04061_),
    .A2(_04223_),
    .ZN(_04227_)
  );
  INV_X1 _14497_ (
    .A(_04227_),
    .ZN(_04228_)
  );
  AND2_X1 _14498_ (
    .A1(_04062_),
    .A2(_04223_),
    .ZN(_04229_)
  );
  INV_X1 _14499_ (
    .A(_04229_),
    .ZN(_04230_)
  );
  AND2_X1 _14500_ (
    .A1(_04061_),
    .A2(_04224_),
    .ZN(_04231_)
  );
  INV_X1 _14501_ (
    .A(_04231_),
    .ZN(_04232_)
  );
  AND2_X1 _14502_ (
    .A1(_04226_),
    .A2(_04228_),
    .ZN(_04233_)
  );
  AND2_X1 _14503_ (
    .A1(_04230_),
    .A2(_04232_),
    .ZN(_04234_)
  );
  AND2_X1 _14504_ (
    .A1(_04129_),
    .A2(_04233_),
    .ZN(_04235_)
  );
  INV_X1 _14505_ (
    .A(_04235_),
    .ZN(_04236_)
  );
  AND2_X1 _14506_ (
    .A1(_04130_),
    .A2(_04234_),
    .ZN(_04237_)
  );
  INV_X1 _14507_ (
    .A(_04237_),
    .ZN(_04238_)
  );
  AND2_X1 _14508_ (
    .A1(_04236_),
    .A2(_04238_),
    .ZN(_04239_)
  );
  INV_X1 _14509_ (
    .A(_04239_),
    .ZN(_04240_)
  );
  AND2_X1 _14510_ (
    .A1(_04066_),
    .A2(_04239_),
    .ZN(_04241_)
  );
  INV_X1 _14511_ (
    .A(_04241_),
    .ZN(_04242_)
  );
  AND2_X1 _14512_ (
    .A1(_04065_),
    .A2(_04240_),
    .ZN(_04243_)
  );
  INV_X1 _14513_ (
    .A(_04243_),
    .ZN(_04244_)
  );
  AND2_X1 _14514_ (
    .A1(_04242_),
    .A2(_04244_),
    .ZN(_04245_)
  );
  INV_X1 _14515_ (
    .A(_04245_),
    .ZN(_04246_)
  );
  AND2_X1 _14516_ (
    .A1(_03886_),
    .A2(_04245_),
    .ZN(_04247_)
  );
  INV_X1 _14517_ (
    .A(_04247_),
    .ZN(_04248_)
  );
  AND2_X1 _14518_ (
    .A1(_03887_),
    .A2(_04246_),
    .ZN(_04249_)
  );
  INV_X1 _14519_ (
    .A(_04249_),
    .ZN(_04250_)
  );
  AND2_X1 _14520_ (
    .A1(_04248_),
    .A2(_04250_),
    .ZN(_04251_)
  );
  INV_X1 _14521_ (
    .A(_04251_),
    .ZN(_04252_)
  );
  AND2_X1 _14522_ (
    .A1(_04060_),
    .A2(_04251_),
    .ZN(_04253_)
  );
  INV_X1 _14523_ (
    .A(_04253_),
    .ZN(_04254_)
  );
  AND2_X1 _14524_ (
    .A1(_04059_),
    .A2(_04252_),
    .ZN(_04255_)
  );
  INV_X1 _14525_ (
    .A(_04255_),
    .ZN(_04256_)
  );
  AND2_X1 _14526_ (
    .A1(_04254_),
    .A2(_04256_),
    .ZN(_04257_)
  );
  INV_X1 _14527_ (
    .A(_04257_),
    .ZN(_04258_)
  );
  AND2_X1 _14528_ (
    .A1(_04002_),
    .A2(_04257_),
    .ZN(_04259_)
  );
  INV_X1 _14529_ (
    .A(_04259_),
    .ZN(_04260_)
  );
  AND2_X1 _14530_ (
    .A1(_04003_),
    .A2(_04258_),
    .ZN(_04261_)
  );
  INV_X1 _14531_ (
    .A(_04261_),
    .ZN(_04262_)
  );
  AND2_X1 _14532_ (
    .A1(_04260_),
    .A2(_04262_),
    .ZN(_04263_)
  );
  INV_X1 _14533_ (
    .A(_04263_),
    .ZN(_04264_)
  );
  AND2_X1 _14534_ (
    .A1(_04058_),
    .A2(_04263_),
    .ZN(_04265_)
  );
  INV_X1 _14535_ (
    .A(_04265_),
    .ZN(_04266_)
  );
  AND2_X1 _14536_ (
    .A1(_04057_),
    .A2(_04264_),
    .ZN(_04267_)
  );
  INV_X1 _14537_ (
    .A(_04267_),
    .ZN(_04268_)
  );
  AND2_X1 _14538_ (
    .A1(_04266_),
    .A2(_04268_),
    .ZN(_04269_)
  );
  INV_X1 _14539_ (
    .A(_04269_),
    .ZN(_04270_)
  );
  AND2_X1 _14540_ (
    .A1(remainder[48]),
    .A2(_04269_),
    .ZN(_04271_)
  );
  INV_X1 _14541_ (
    .A(_04271_),
    .ZN(_04272_)
  );
  AND2_X1 _14542_ (
    .A1(_04590_),
    .A2(_04270_),
    .ZN(_04273_)
  );
  INV_X1 _14543_ (
    .A(_04273_),
    .ZN(_04274_)
  );
  AND2_X1 _14544_ (
    .A1(_04272_),
    .A2(_04274_),
    .ZN(_04275_)
  );
  INV_X1 _14545_ (
    .A(_04275_),
    .ZN(_04276_)
  );
  AND2_X1 _14546_ (
    .A1(_04056_),
    .A2(_04275_),
    .ZN(_04277_)
  );
  INV_X1 _14547_ (
    .A(_04277_),
    .ZN(_04278_)
  );
  AND2_X1 _14548_ (
    .A1(_04055_),
    .A2(_04276_),
    .ZN(_04279_)
  );
  INV_X1 _14549_ (
    .A(_04279_),
    .ZN(_04280_)
  );
  AND2_X1 _14550_ (
    .A1(_02082_),
    .A2(_04280_),
    .ZN(_04281_)
  );
  AND2_X1 _14551_ (
    .A1(_04278_),
    .A2(_04281_),
    .ZN(_04282_)
  );
  INV_X1 _14552_ (
    .A(_04282_),
    .ZN(_04283_)
  );
  AND2_X1 _14553_ (
    .A1(_04054_),
    .A2(_04283_),
    .ZN(_04284_)
  );
  AND2_X1 _14554_ (
    .A1(_04052_),
    .A2(_04284_),
    .ZN(_04285_)
  );
  INV_X1 _14555_ (
    .A(_04285_),
    .ZN(_04286_)
  );
  AND2_X1 _14556_ (
    .A1(_06201_),
    .A2(_04286_),
    .ZN(_00061_)
  );
  AND2_X1 _14557_ (
    .A1(_04678_),
    .A2(_10451_),
    .ZN(_04287_)
  );
  INV_X1 _14558_ (
    .A(_04287_),
    .ZN(_04288_)
  );
  AND2_X1 _14559_ (
    .A1(_10462_),
    .A2(_01441_),
    .ZN(_04289_)
  );
  INV_X1 _14560_ (
    .A(_04289_),
    .ZN(_04290_)
  );
  AND2_X1 _14561_ (
    .A1(_05983_),
    .A2(_04290_),
    .ZN(_04291_)
  );
  AND2_X1 _14562_ (
    .A1(_04288_),
    .A2(_04291_),
    .ZN(_04292_)
  );
  INV_X1 _14563_ (
    .A(_04292_),
    .ZN(_04293_)
  );
  AND2_X1 _14564_ (
    .A1(remainder[41]),
    .A2(_02077_),
    .ZN(_04294_)
  );
  INV_X1 _14565_ (
    .A(_04294_),
    .ZN(_04295_)
  );
  AND2_X1 _14566_ (
    .A1(_04272_),
    .A2(_04278_),
    .ZN(_04296_)
  );
  INV_X1 _14567_ (
    .A(_04296_),
    .ZN(_04297_)
  );
  AND2_X1 _14568_ (
    .A1(_04260_),
    .A2(_04266_),
    .ZN(_04298_)
  );
  INV_X1 _14569_ (
    .A(_04298_),
    .ZN(_04299_)
  );
  AND2_X1 _14570_ (
    .A1(_04242_),
    .A2(_04248_),
    .ZN(_04300_)
  );
  INV_X1 _14571_ (
    .A(_04300_),
    .ZN(_04301_)
  );
  AND2_X1 _14572_ (
    .A1(_03249_),
    .A2(_04224_),
    .ZN(_04302_)
  );
  INV_X1 _14573_ (
    .A(_04302_),
    .ZN(_04303_)
  );
  AND2_X1 _14574_ (
    .A1(_03972_),
    .A2(_04302_),
    .ZN(_04304_)
  );
  INV_X1 _14575_ (
    .A(_04304_),
    .ZN(_04305_)
  );
  AND2_X1 _14576_ (
    .A1(_04236_),
    .A2(_04305_),
    .ZN(_04306_)
  );
  INV_X1 _14577_ (
    .A(_04306_),
    .ZN(_04307_)
  );
  AND2_X1 _14578_ (
    .A1(_04114_),
    .A2(_04120_),
    .ZN(_04308_)
  );
  INV_X1 _14579_ (
    .A(_04308_),
    .ZN(_04309_)
  );
  AND2_X1 _14580_ (
    .A1(_04102_),
    .A2(_04108_),
    .ZN(_04310_)
  );
  INV_X1 _14581_ (
    .A(_04310_),
    .ZN(_04311_)
  );
  AND2_X1 _14582_ (
    .A1(_04090_),
    .A2(_04096_),
    .ZN(_04312_)
  );
  INV_X1 _14583_ (
    .A(_04312_),
    .ZN(_04313_)
  );
  AND2_X1 _14584_ (
    .A1(_04180_),
    .A2(_04220_),
    .ZN(_04314_)
  );
  INV_X1 _14585_ (
    .A(_04314_),
    .ZN(_04315_)
  );
  AND2_X1 _14586_ (
    .A1(_03839_),
    .A2(_04084_),
    .ZN(_04316_)
  );
  INV_X1 _14587_ (
    .A(_04316_),
    .ZN(_04317_)
  );
  AND2_X1 _14588_ (
    .A1(_04208_),
    .A2(_04214_),
    .ZN(_04318_)
  );
  INV_X1 _14589_ (
    .A(_04318_),
    .ZN(_04319_)
  );
  AND2_X1 _14590_ (
    .A1(_04087_),
    .A2(_04319_),
    .ZN(_04320_)
  );
  INV_X1 _14591_ (
    .A(_04320_),
    .ZN(_04321_)
  );
  AND2_X1 _14592_ (
    .A1(_04088_),
    .A2(_04318_),
    .ZN(_04322_)
  );
  INV_X1 _14593_ (
    .A(_04322_),
    .ZN(_04323_)
  );
  AND2_X1 _14594_ (
    .A1(_04321_),
    .A2(_04323_),
    .ZN(_04324_)
  );
  INV_X1 _14595_ (
    .A(_04324_),
    .ZN(_04325_)
  );
  AND2_X1 _14596_ (
    .A1(_04317_),
    .A2(_04324_),
    .ZN(_04326_)
  );
  INV_X1 _14597_ (
    .A(_04326_),
    .ZN(_04327_)
  );
  AND2_X1 _14598_ (
    .A1(_04316_),
    .A2(_04325_),
    .ZN(_04328_)
  );
  INV_X1 _14599_ (
    .A(_04328_),
    .ZN(_04329_)
  );
  AND2_X1 _14600_ (
    .A1(_04327_),
    .A2(_04329_),
    .ZN(_04330_)
  );
  INV_X1 _14601_ (
    .A(_04330_),
    .ZN(_04331_)
  );
  AND2_X1 _14602_ (
    .A1(_04315_),
    .A2(_04330_),
    .ZN(_04332_)
  );
  INV_X1 _14603_ (
    .A(_04332_),
    .ZN(_04333_)
  );
  AND2_X1 _14604_ (
    .A1(_04314_),
    .A2(_04331_),
    .ZN(_04334_)
  );
  INV_X1 _14605_ (
    .A(_04334_),
    .ZN(_04335_)
  );
  AND2_X1 _14606_ (
    .A1(_04333_),
    .A2(_04335_),
    .ZN(_04336_)
  );
  INV_X1 _14607_ (
    .A(_04336_),
    .ZN(_04337_)
  );
  AND2_X1 _14608_ (
    .A1(_04313_),
    .A2(_04336_),
    .ZN(_04338_)
  );
  INV_X1 _14609_ (
    .A(_04338_),
    .ZN(_04339_)
  );
  AND2_X1 _14610_ (
    .A1(_04312_),
    .A2(_04337_),
    .ZN(_04340_)
  );
  INV_X1 _14611_ (
    .A(_04340_),
    .ZN(_04341_)
  );
  AND2_X1 _14612_ (
    .A1(_04339_),
    .A2(_04341_),
    .ZN(_04342_)
  );
  INV_X1 _14613_ (
    .A(_04342_),
    .ZN(_04343_)
  );
  AND2_X1 _14614_ (
    .A1(_04311_),
    .A2(_04342_),
    .ZN(_04344_)
  );
  INV_X1 _14615_ (
    .A(_04344_),
    .ZN(_04345_)
  );
  AND2_X1 _14616_ (
    .A1(_04310_),
    .A2(_04343_),
    .ZN(_04346_)
  );
  INV_X1 _14617_ (
    .A(_04346_),
    .ZN(_04347_)
  );
  AND2_X1 _14618_ (
    .A1(_04345_),
    .A2(_04347_),
    .ZN(_04348_)
  );
  INV_X1 _14619_ (
    .A(_04348_),
    .ZN(_04349_)
  );
  AND2_X1 _14620_ (
    .A1(_03170_),
    .A2(_04348_),
    .ZN(_04350_)
  );
  INV_X1 _14621_ (
    .A(_04350_),
    .ZN(_04351_)
  );
  AND2_X1 _14622_ (
    .A1(_03169_),
    .A2(_04349_),
    .ZN(_04352_)
  );
  INV_X1 _14623_ (
    .A(_04352_),
    .ZN(_04353_)
  );
  AND2_X1 _14624_ (
    .A1(_04351_),
    .A2(_04353_),
    .ZN(_04354_)
  );
  INV_X1 _14625_ (
    .A(_04354_),
    .ZN(_04355_)
  );
  AND2_X1 _14626_ (
    .A1(_04309_),
    .A2(_04354_),
    .ZN(_04356_)
  );
  INV_X1 _14627_ (
    .A(_04356_),
    .ZN(_04357_)
  );
  AND2_X1 _14628_ (
    .A1(_04308_),
    .A2(_04355_),
    .ZN(_04358_)
  );
  INV_X1 _14629_ (
    .A(_04358_),
    .ZN(_04359_)
  );
  AND2_X1 _14630_ (
    .A1(_04357_),
    .A2(_04359_),
    .ZN(_04360_)
  );
  INV_X1 _14631_ (
    .A(_04360_),
    .ZN(_04361_)
  );
  AND2_X1 _14632_ (
    .A1(divisor[16]),
    .A2(remainder[0]),
    .ZN(_04362_)
  );
  INV_X1 _14633_ (
    .A(_04362_),
    .ZN(_04363_)
  );
  AND2_X1 _14634_ (
    .A1(_04150_),
    .A2(_04174_),
    .ZN(_04364_)
  );
  INV_X1 _14635_ (
    .A(_04364_),
    .ZN(_04365_)
  );
  AND2_X1 _14636_ (
    .A1(_04138_),
    .A2(_04144_),
    .ZN(_04366_)
  );
  INV_X1 _14637_ (
    .A(_04366_),
    .ZN(_04367_)
  );
  AND2_X1 _14638_ (
    .A1(divisor[13]),
    .A2(remainder[3]),
    .ZN(_04368_)
  );
  INV_X1 _14639_ (
    .A(_04368_),
    .ZN(_04369_)
  );
  AND2_X1 _14640_ (
    .A1(divisor[14]),
    .A2(remainder[2]),
    .ZN(_04370_)
  );
  INV_X1 _14641_ (
    .A(_04370_),
    .ZN(_04371_)
  );
  AND2_X1 _14642_ (
    .A1(divisor[15]),
    .A2(remainder[2]),
    .ZN(_04372_)
  );
  INV_X1 _14643_ (
    .A(_04372_),
    .ZN(_04373_)
  );
  AND2_X1 _14644_ (
    .A1(_03896_),
    .A2(_04372_),
    .ZN(_04374_)
  );
  INV_X1 _14645_ (
    .A(_04374_),
    .ZN(_04375_)
  );
  AND2_X1 _14646_ (
    .A1(_04136_),
    .A2(_04371_),
    .ZN(_04376_)
  );
  INV_X1 _14647_ (
    .A(_04376_),
    .ZN(_04377_)
  );
  AND2_X1 _14648_ (
    .A1(_04375_),
    .A2(_04377_),
    .ZN(_04378_)
  );
  INV_X1 _14649_ (
    .A(_04378_),
    .ZN(_04379_)
  );
  AND2_X1 _14650_ (
    .A1(_04368_),
    .A2(_04378_),
    .ZN(_04380_)
  );
  INV_X1 _14651_ (
    .A(_04380_),
    .ZN(_04381_)
  );
  AND2_X1 _14652_ (
    .A1(_04369_),
    .A2(_04379_),
    .ZN(_04382_)
  );
  INV_X1 _14653_ (
    .A(_04382_),
    .ZN(_04383_)
  );
  AND2_X1 _14654_ (
    .A1(_04381_),
    .A2(_04383_),
    .ZN(_04384_)
  );
  INV_X1 _14655_ (
    .A(_04384_),
    .ZN(_04385_)
  );
  AND2_X1 _14656_ (
    .A1(_04367_),
    .A2(_04384_),
    .ZN(_04386_)
  );
  INV_X1 _14657_ (
    .A(_04386_),
    .ZN(_04387_)
  );
  AND2_X1 _14658_ (
    .A1(_04366_),
    .A2(_04385_),
    .ZN(_04388_)
  );
  INV_X1 _14659_ (
    .A(_04388_),
    .ZN(_04389_)
  );
  AND2_X1 _14660_ (
    .A1(_04387_),
    .A2(_04389_),
    .ZN(_04390_)
  );
  INV_X1 _14661_ (
    .A(_04390_),
    .ZN(_04391_)
  );
  AND2_X1 _14662_ (
    .A1(divisor[10]),
    .A2(remainder[6]),
    .ZN(_04392_)
  );
  INV_X1 _14663_ (
    .A(_04392_),
    .ZN(_04393_)
  );
  AND2_X1 _14664_ (
    .A1(divisor[11]),
    .A2(remainder[5]),
    .ZN(_04394_)
  );
  INV_X1 _14665_ (
    .A(_04394_),
    .ZN(_04395_)
  );
  AND2_X1 _14666_ (
    .A1(divisor[12]),
    .A2(remainder[5]),
    .ZN(_04396_)
  );
  INV_X1 _14667_ (
    .A(_04396_),
    .ZN(_04397_)
  );
  AND2_X1 _14668_ (
    .A1(_04159_),
    .A2(_04394_),
    .ZN(_04398_)
  );
  INV_X1 _14669_ (
    .A(_04398_),
    .ZN(_04399_)
  );
  AND2_X1 _14670_ (
    .A1(_04160_),
    .A2(_04395_),
    .ZN(_04400_)
  );
  INV_X1 _14671_ (
    .A(_04400_),
    .ZN(_04401_)
  );
  AND2_X1 _14672_ (
    .A1(_04399_),
    .A2(_04401_),
    .ZN(_04402_)
  );
  INV_X1 _14673_ (
    .A(_04402_),
    .ZN(_04403_)
  );
  AND2_X1 _14674_ (
    .A1(_04392_),
    .A2(_04402_),
    .ZN(_04405_)
  );
  INV_X1 _14675_ (
    .A(_04405_),
    .ZN(_04406_)
  );
  AND2_X1 _14676_ (
    .A1(_04393_),
    .A2(_04403_),
    .ZN(_04407_)
  );
  INV_X1 _14677_ (
    .A(_04407_),
    .ZN(_04408_)
  );
  AND2_X1 _14678_ (
    .A1(_04406_),
    .A2(_04408_),
    .ZN(_04409_)
  );
  INV_X1 _14679_ (
    .A(_04409_),
    .ZN(_04410_)
  );
  AND2_X1 _14680_ (
    .A1(_04390_),
    .A2(_04409_),
    .ZN(_04411_)
  );
  INV_X1 _14681_ (
    .A(_04411_),
    .ZN(_04412_)
  );
  AND2_X1 _14682_ (
    .A1(_04391_),
    .A2(_04410_),
    .ZN(_04413_)
  );
  INV_X1 _14683_ (
    .A(_04413_),
    .ZN(_04414_)
  );
  AND2_X1 _14684_ (
    .A1(_04412_),
    .A2(_04414_),
    .ZN(_04416_)
  );
  INV_X1 _14685_ (
    .A(_04416_),
    .ZN(_04417_)
  );
  AND2_X1 _14686_ (
    .A1(_04365_),
    .A2(_04416_),
    .ZN(_04418_)
  );
  INV_X1 _14687_ (
    .A(_04418_),
    .ZN(_04419_)
  );
  AND2_X1 _14688_ (
    .A1(_04364_),
    .A2(_04417_),
    .ZN(_04420_)
  );
  INV_X1 _14689_ (
    .A(_04420_),
    .ZN(_04421_)
  );
  AND2_X1 _14690_ (
    .A1(_04419_),
    .A2(_04421_),
    .ZN(_04422_)
  );
  INV_X1 _14691_ (
    .A(_04422_),
    .ZN(_04423_)
  );
  AND2_X1 _14692_ (
    .A1(_04196_),
    .A2(_04202_),
    .ZN(_04424_)
  );
  INV_X1 _14693_ (
    .A(_04424_),
    .ZN(_04425_)
  );
  AND2_X1 _14694_ (
    .A1(_04162_),
    .A2(_04168_),
    .ZN(_04427_)
  );
  INV_X1 _14695_ (
    .A(_04427_),
    .ZN(_04428_)
  );
  AND2_X1 _14696_ (
    .A1(remainder[32]),
    .A2(divisor[9]),
    .ZN(_04429_)
  );
  AND2_X1 _14697_ (
    .A1(remainder[32]),
    .A2(divisor[8]),
    .ZN(_04430_)
  );
  INV_X1 _14698_ (
    .A(_04430_),
    .ZN(_04431_)
  );
  AND2_X1 _14699_ (
    .A1(divisor[9]),
    .A2(_04430_),
    .ZN(_04432_)
  );
  INV_X1 _14700_ (
    .A(_04432_),
    .ZN(_04433_)
  );
  AND2_X1 _14701_ (
    .A1(_04193_),
    .A2(_04430_),
    .ZN(_04434_)
  );
  INV_X1 _14702_ (
    .A(_04434_),
    .ZN(_04435_)
  );
  AND2_X1 _14703_ (
    .A1(_04194_),
    .A2(_04431_),
    .ZN(_04436_)
  );
  INV_X1 _14704_ (
    .A(_04436_),
    .ZN(_04438_)
  );
  AND2_X1 _14705_ (
    .A1(_04435_),
    .A2(_04438_),
    .ZN(_04439_)
  );
  INV_X1 _14706_ (
    .A(_04439_),
    .ZN(_04440_)
  );
  AND2_X1 _14707_ (
    .A1(_04189_),
    .A2(_04439_),
    .ZN(_04441_)
  );
  INV_X1 _14708_ (
    .A(_04441_),
    .ZN(_04442_)
  );
  AND2_X1 _14709_ (
    .A1(_04190_),
    .A2(_04440_),
    .ZN(_04443_)
  );
  INV_X1 _14710_ (
    .A(_04443_),
    .ZN(_04444_)
  );
  AND2_X1 _14711_ (
    .A1(_04442_),
    .A2(_04444_),
    .ZN(_04445_)
  );
  INV_X1 _14712_ (
    .A(_04445_),
    .ZN(_04446_)
  );
  AND2_X1 _14713_ (
    .A1(_04428_),
    .A2(_04445_),
    .ZN(_04447_)
  );
  INV_X1 _14714_ (
    .A(_04447_),
    .ZN(_04449_)
  );
  AND2_X1 _14715_ (
    .A1(_04427_),
    .A2(_04446_),
    .ZN(_04450_)
  );
  INV_X1 _14716_ (
    .A(_04450_),
    .ZN(_04451_)
  );
  AND2_X1 _14717_ (
    .A1(_04449_),
    .A2(_04451_),
    .ZN(_04452_)
  );
  INV_X1 _14718_ (
    .A(_04452_),
    .ZN(_04453_)
  );
  AND2_X1 _14719_ (
    .A1(_04425_),
    .A2(_04452_),
    .ZN(_04454_)
  );
  INV_X1 _14720_ (
    .A(_04454_),
    .ZN(_04455_)
  );
  AND2_X1 _14721_ (
    .A1(_04424_),
    .A2(_04453_),
    .ZN(_04456_)
  );
  INV_X1 _14722_ (
    .A(_04456_),
    .ZN(_04457_)
  );
  AND2_X1 _14723_ (
    .A1(_04455_),
    .A2(_04457_),
    .ZN(_04458_)
  );
  INV_X1 _14724_ (
    .A(_04458_),
    .ZN(_04460_)
  );
  AND2_X1 _14725_ (
    .A1(_04422_),
    .A2(_04458_),
    .ZN(_04461_)
  );
  INV_X1 _14726_ (
    .A(_04461_),
    .ZN(_04462_)
  );
  AND2_X1 _14727_ (
    .A1(_04423_),
    .A2(_04460_),
    .ZN(_04463_)
  );
  INV_X1 _14728_ (
    .A(_04463_),
    .ZN(_04464_)
  );
  AND2_X1 _14729_ (
    .A1(_04462_),
    .A2(_04464_),
    .ZN(_04465_)
  );
  INV_X1 _14730_ (
    .A(_04465_),
    .ZN(_04466_)
  );
  AND2_X1 _14731_ (
    .A1(_04362_),
    .A2(_04465_),
    .ZN(_04467_)
  );
  INV_X1 _14732_ (
    .A(_04467_),
    .ZN(_04468_)
  );
  AND2_X1 _14733_ (
    .A1(_04363_),
    .A2(_04466_),
    .ZN(_04469_)
  );
  INV_X1 _14734_ (
    .A(_04469_),
    .ZN(_04471_)
  );
  AND2_X1 _14735_ (
    .A1(_04468_),
    .A2(_04471_),
    .ZN(_04472_)
  );
  INV_X1 _14736_ (
    .A(_04472_),
    .ZN(_04473_)
  );
  AND2_X1 _14737_ (
    .A1(_04303_),
    .A2(_04473_),
    .ZN(_04474_)
  );
  INV_X1 _14738_ (
    .A(_04474_),
    .ZN(_04475_)
  );
  AND2_X1 _14739_ (
    .A1(_04302_),
    .A2(_04472_),
    .ZN(_04476_)
  );
  INV_X1 _14740_ (
    .A(_04476_),
    .ZN(_04477_)
  );
  AND2_X1 _14741_ (
    .A1(_04303_),
    .A2(_04472_),
    .ZN(_04478_)
  );
  INV_X1 _14742_ (
    .A(_04478_),
    .ZN(_04479_)
  );
  AND2_X1 _14743_ (
    .A1(_04302_),
    .A2(_04473_),
    .ZN(_04480_)
  );
  INV_X1 _14744_ (
    .A(_04480_),
    .ZN(_04482_)
  );
  AND2_X1 _14745_ (
    .A1(_04475_),
    .A2(_04477_),
    .ZN(_04483_)
  );
  AND2_X1 _14746_ (
    .A1(_04479_),
    .A2(_04482_),
    .ZN(_04484_)
  );
  AND2_X1 _14747_ (
    .A1(_04360_),
    .A2(_04483_),
    .ZN(_04485_)
  );
  INV_X1 _14748_ (
    .A(_04485_),
    .ZN(_04486_)
  );
  AND2_X1 _14749_ (
    .A1(_04361_),
    .A2(_04484_),
    .ZN(_04487_)
  );
  INV_X1 _14750_ (
    .A(_04487_),
    .ZN(_04488_)
  );
  AND2_X1 _14751_ (
    .A1(_04486_),
    .A2(_04488_),
    .ZN(_04489_)
  );
  INV_X1 _14752_ (
    .A(_04489_),
    .ZN(_04490_)
  );
  AND2_X1 _14753_ (
    .A1(_04307_),
    .A2(_04489_),
    .ZN(_04491_)
  );
  INV_X1 _14754_ (
    .A(_04491_),
    .ZN(_04493_)
  );
  AND2_X1 _14755_ (
    .A1(_04306_),
    .A2(_04490_),
    .ZN(_04494_)
  );
  INV_X1 _14756_ (
    .A(_04494_),
    .ZN(_04495_)
  );
  AND2_X1 _14757_ (
    .A1(_04493_),
    .A2(_04495_),
    .ZN(_04496_)
  );
  INV_X1 _14758_ (
    .A(_04496_),
    .ZN(_04497_)
  );
  AND2_X1 _14759_ (
    .A1(_04125_),
    .A2(_04496_),
    .ZN(_04498_)
  );
  INV_X1 _14760_ (
    .A(_04498_),
    .ZN(_04499_)
  );
  AND2_X1 _14761_ (
    .A1(_04126_),
    .A2(_04497_),
    .ZN(_04500_)
  );
  INV_X1 _14762_ (
    .A(_04500_),
    .ZN(_04501_)
  );
  AND2_X1 _14763_ (
    .A1(_04499_),
    .A2(_04501_),
    .ZN(_04502_)
  );
  INV_X1 _14764_ (
    .A(_04502_),
    .ZN(_04504_)
  );
  AND2_X1 _14765_ (
    .A1(_04301_),
    .A2(_04502_),
    .ZN(_04505_)
  );
  INV_X1 _14766_ (
    .A(_04505_),
    .ZN(_04506_)
  );
  AND2_X1 _14767_ (
    .A1(_04300_),
    .A2(_04504_),
    .ZN(_04507_)
  );
  INV_X1 _14768_ (
    .A(_04507_),
    .ZN(_04508_)
  );
  AND2_X1 _14769_ (
    .A1(_04506_),
    .A2(_04508_),
    .ZN(_04509_)
  );
  INV_X1 _14770_ (
    .A(_04509_),
    .ZN(_04510_)
  );
  AND2_X1 _14771_ (
    .A1(_04253_),
    .A2(_04509_),
    .ZN(_04511_)
  );
  INV_X1 _14772_ (
    .A(_04511_),
    .ZN(_04512_)
  );
  AND2_X1 _14773_ (
    .A1(_04254_),
    .A2(_04510_),
    .ZN(_04513_)
  );
  INV_X1 _14774_ (
    .A(_04513_),
    .ZN(_04515_)
  );
  AND2_X1 _14775_ (
    .A1(_04512_),
    .A2(_04515_),
    .ZN(_04516_)
  );
  INV_X1 _14776_ (
    .A(_04516_),
    .ZN(_04517_)
  );
  AND2_X1 _14777_ (
    .A1(_04299_),
    .A2(_04516_),
    .ZN(_04518_)
  );
  INV_X1 _14778_ (
    .A(_04518_),
    .ZN(_04519_)
  );
  AND2_X1 _14779_ (
    .A1(_04298_),
    .A2(_04517_),
    .ZN(_04520_)
  );
  INV_X1 _14780_ (
    .A(_04520_),
    .ZN(_04521_)
  );
  AND2_X1 _14781_ (
    .A1(_04519_),
    .A2(_04521_),
    .ZN(_04522_)
  );
  INV_X1 _14782_ (
    .A(_04522_),
    .ZN(_04523_)
  );
  AND2_X1 _14783_ (
    .A1(remainder[49]),
    .A2(_04522_),
    .ZN(_04524_)
  );
  INV_X1 _14784_ (
    .A(_04524_),
    .ZN(_04526_)
  );
  AND2_X1 _14785_ (
    .A1(_04579_),
    .A2(_04523_),
    .ZN(_04527_)
  );
  INV_X1 _14786_ (
    .A(_04527_),
    .ZN(_04528_)
  );
  AND2_X1 _14787_ (
    .A1(_04526_),
    .A2(_04528_),
    .ZN(_04529_)
  );
  INV_X1 _14788_ (
    .A(_04529_),
    .ZN(_04530_)
  );
  AND2_X1 _14789_ (
    .A1(_04297_),
    .A2(_04529_),
    .ZN(_04531_)
  );
  INV_X1 _14790_ (
    .A(_04531_),
    .ZN(_04532_)
  );
  AND2_X1 _14791_ (
    .A1(_04296_),
    .A2(_04530_),
    .ZN(_04533_)
  );
  INV_X1 _14792_ (
    .A(_04533_),
    .ZN(_04534_)
  );
  AND2_X1 _14793_ (
    .A1(_02082_),
    .A2(_04534_),
    .ZN(_04535_)
  );
  AND2_X1 _14794_ (
    .A1(_04532_),
    .A2(_04535_),
    .ZN(_04537_)
  );
  INV_X1 _14795_ (
    .A(_04537_),
    .ZN(_04538_)
  );
  AND2_X1 _14796_ (
    .A1(_04295_),
    .A2(_04538_),
    .ZN(_04539_)
  );
  AND2_X1 _14797_ (
    .A1(_04293_),
    .A2(_04539_),
    .ZN(_04540_)
  );
  INV_X1 _14798_ (
    .A(_04540_),
    .ZN(_04541_)
  );
  AND2_X1 _14799_ (
    .A1(_06201_),
    .A2(_04541_),
    .ZN(_00062_)
  );
  AND2_X1 _14800_ (
    .A1(_04667_),
    .A2(_10451_),
    .ZN(_04542_)
  );
  INV_X1 _14801_ (
    .A(_04542_),
    .ZN(_04543_)
  );
  AND2_X1 _14802_ (
    .A1(_10462_),
    .A2(_01604_),
    .ZN(_04544_)
  );
  INV_X1 _14803_ (
    .A(_04544_),
    .ZN(_04545_)
  );
  AND2_X1 _14804_ (
    .A1(_05983_),
    .A2(_04545_),
    .ZN(_04547_)
  );
  AND2_X1 _14805_ (
    .A1(_04543_),
    .A2(_04547_),
    .ZN(_04548_)
  );
  INV_X1 _14806_ (
    .A(_04548_),
    .ZN(_04549_)
  );
  AND2_X1 _14807_ (
    .A1(remainder[42]),
    .A2(_02077_),
    .ZN(_04550_)
  );
  INV_X1 _14808_ (
    .A(_04550_),
    .ZN(_04551_)
  );
  AND2_X1 _14809_ (
    .A1(_04526_),
    .A2(_04532_),
    .ZN(_04552_)
  );
  INV_X1 _14810_ (
    .A(_04552_),
    .ZN(_04553_)
  );
  AND2_X1 _14811_ (
    .A1(_04512_),
    .A2(_04519_),
    .ZN(_04554_)
  );
  INV_X1 _14812_ (
    .A(_04554_),
    .ZN(_04555_)
  );
  AND2_X1 _14813_ (
    .A1(_04493_),
    .A2(_04499_),
    .ZN(_04556_)
  );
  INV_X1 _14814_ (
    .A(_04556_),
    .ZN(_04558_)
  );
  AND2_X1 _14815_ (
    .A1(_03249_),
    .A2(_04473_),
    .ZN(_04559_)
  );
  INV_X1 _14816_ (
    .A(_04559_),
    .ZN(_04560_)
  );
  AND2_X1 _14817_ (
    .A1(_04223_),
    .A2(_04559_),
    .ZN(_04561_)
  );
  INV_X1 _14818_ (
    .A(_04561_),
    .ZN(_04562_)
  );
  AND2_X1 _14819_ (
    .A1(_04486_),
    .A2(_04562_),
    .ZN(_04563_)
  );
  INV_X1 _14820_ (
    .A(_04563_),
    .ZN(_04564_)
  );
  AND2_X1 _14821_ (
    .A1(_04345_),
    .A2(_04351_),
    .ZN(_04565_)
  );
  INV_X1 _14822_ (
    .A(_04565_),
    .ZN(_04566_)
  );
  AND2_X1 _14823_ (
    .A1(_04333_),
    .A2(_04339_),
    .ZN(_04567_)
  );
  INV_X1 _14824_ (
    .A(_04567_),
    .ZN(_04569_)
  );
  AND2_X1 _14825_ (
    .A1(_04321_),
    .A2(_04327_),
    .ZN(_04570_)
  );
  INV_X1 _14826_ (
    .A(_04570_),
    .ZN(_04571_)
  );
  AND2_X1 _14827_ (
    .A1(_04419_),
    .A2(_04462_),
    .ZN(_04572_)
  );
  INV_X1 _14828_ (
    .A(_04572_),
    .ZN(_04573_)
  );
  AND2_X1 _14829_ (
    .A1(_04449_),
    .A2(_04455_),
    .ZN(_04574_)
  );
  INV_X1 _14830_ (
    .A(_04574_),
    .ZN(_04575_)
  );
  AND2_X1 _14831_ (
    .A1(_04087_),
    .A2(_04575_),
    .ZN(_04576_)
  );
  INV_X1 _14832_ (
    .A(_04576_),
    .ZN(_04577_)
  );
  AND2_X1 _14833_ (
    .A1(_04088_),
    .A2(_04574_),
    .ZN(_04578_)
  );
  INV_X1 _14834_ (
    .A(_04578_),
    .ZN(_04580_)
  );
  AND2_X1 _14835_ (
    .A1(_04577_),
    .A2(_04580_),
    .ZN(_04581_)
  );
  INV_X1 _14836_ (
    .A(_04581_),
    .ZN(_04582_)
  );
  AND2_X1 _14837_ (
    .A1(_04317_),
    .A2(_04581_),
    .ZN(_04583_)
  );
  INV_X1 _14838_ (
    .A(_04583_),
    .ZN(_04584_)
  );
  AND2_X1 _14839_ (
    .A1(_04316_),
    .A2(_04582_),
    .ZN(_04585_)
  );
  INV_X1 _14840_ (
    .A(_04585_),
    .ZN(_04586_)
  );
  AND2_X1 _14841_ (
    .A1(_04584_),
    .A2(_04586_),
    .ZN(_04587_)
  );
  INV_X1 _14842_ (
    .A(_04587_),
    .ZN(_04588_)
  );
  AND2_X1 _14843_ (
    .A1(_04573_),
    .A2(_04587_),
    .ZN(_04589_)
  );
  INV_X1 _14844_ (
    .A(_04589_),
    .ZN(_04591_)
  );
  AND2_X1 _14845_ (
    .A1(_04572_),
    .A2(_04588_),
    .ZN(_04592_)
  );
  INV_X1 _14846_ (
    .A(_04592_),
    .ZN(_04593_)
  );
  AND2_X1 _14847_ (
    .A1(_04591_),
    .A2(_04593_),
    .ZN(_04594_)
  );
  INV_X1 _14848_ (
    .A(_04594_),
    .ZN(_04595_)
  );
  AND2_X1 _14849_ (
    .A1(_04571_),
    .A2(_04594_),
    .ZN(_04596_)
  );
  INV_X1 _14850_ (
    .A(_04596_),
    .ZN(_04597_)
  );
  AND2_X1 _14851_ (
    .A1(_04570_),
    .A2(_04595_),
    .ZN(_04598_)
  );
  INV_X1 _14852_ (
    .A(_04598_),
    .ZN(_04599_)
  );
  AND2_X1 _14853_ (
    .A1(_04597_),
    .A2(_04599_),
    .ZN(_04600_)
  );
  INV_X1 _14854_ (
    .A(_04600_),
    .ZN(_04602_)
  );
  AND2_X1 _14855_ (
    .A1(_04569_),
    .A2(_04600_),
    .ZN(_04603_)
  );
  INV_X1 _14856_ (
    .A(_04603_),
    .ZN(_04604_)
  );
  AND2_X1 _14857_ (
    .A1(_04567_),
    .A2(_04602_),
    .ZN(_04605_)
  );
  INV_X1 _14858_ (
    .A(_04605_),
    .ZN(_04606_)
  );
  AND2_X1 _14859_ (
    .A1(_04604_),
    .A2(_04606_),
    .ZN(_04607_)
  );
  INV_X1 _14860_ (
    .A(_04607_),
    .ZN(_04608_)
  );
  AND2_X1 _14861_ (
    .A1(_03170_),
    .A2(_04607_),
    .ZN(_04609_)
  );
  INV_X1 _14862_ (
    .A(_04609_),
    .ZN(_04610_)
  );
  AND2_X1 _14863_ (
    .A1(_03169_),
    .A2(_04608_),
    .ZN(_04611_)
  );
  INV_X1 _14864_ (
    .A(_04611_),
    .ZN(_04613_)
  );
  AND2_X1 _14865_ (
    .A1(_04610_),
    .A2(_04613_),
    .ZN(_04614_)
  );
  INV_X1 _14866_ (
    .A(_04614_),
    .ZN(_04615_)
  );
  AND2_X1 _14867_ (
    .A1(_04566_),
    .A2(_04614_),
    .ZN(_04616_)
  );
  INV_X1 _14868_ (
    .A(_04616_),
    .ZN(_04617_)
  );
  AND2_X1 _14869_ (
    .A1(_04565_),
    .A2(_04615_),
    .ZN(_04618_)
  );
  INV_X1 _14870_ (
    .A(_04618_),
    .ZN(_04619_)
  );
  AND2_X1 _14871_ (
    .A1(_04617_),
    .A2(_04619_),
    .ZN(_04620_)
  );
  INV_X1 _14872_ (
    .A(_04620_),
    .ZN(_04621_)
  );
  AND2_X1 _14873_ (
    .A1(divisor[17]),
    .A2(remainder[0]),
    .ZN(_04622_)
  );
  INV_X1 _14874_ (
    .A(_04622_),
    .ZN(_04624_)
  );
  AND2_X1 _14875_ (
    .A1(divisor[16]),
    .A2(remainder[1]),
    .ZN(_04625_)
  );
  INV_X1 _14876_ (
    .A(_04625_),
    .ZN(_04626_)
  );
  AND2_X1 _14877_ (
    .A1(divisor[17]),
    .A2(remainder[1]),
    .ZN(_04627_)
  );
  INV_X1 _14878_ (
    .A(_04627_),
    .ZN(_04628_)
  );
  AND2_X1 _14879_ (
    .A1(_04362_),
    .A2(_04627_),
    .ZN(_04629_)
  );
  INV_X1 _14880_ (
    .A(_04629_),
    .ZN(_04630_)
  );
  AND2_X1 _14881_ (
    .A1(_04624_),
    .A2(_04626_),
    .ZN(_04631_)
  );
  INV_X1 _14882_ (
    .A(_04631_),
    .ZN(_04632_)
  );
  AND2_X1 _14883_ (
    .A1(_04630_),
    .A2(_04632_),
    .ZN(_04633_)
  );
  INV_X1 _14884_ (
    .A(_04633_),
    .ZN(_04635_)
  );
  AND2_X1 _14885_ (
    .A1(_04387_),
    .A2(_04412_),
    .ZN(_04636_)
  );
  INV_X1 _14886_ (
    .A(_04636_),
    .ZN(_04637_)
  );
  AND2_X1 _14887_ (
    .A1(_04375_),
    .A2(_04381_),
    .ZN(_04638_)
  );
  INV_X1 _14888_ (
    .A(_04638_),
    .ZN(_04639_)
  );
  AND2_X1 _14889_ (
    .A1(divisor[13]),
    .A2(remainder[4]),
    .ZN(_04640_)
  );
  INV_X1 _14890_ (
    .A(_04640_),
    .ZN(_04641_)
  );
  AND2_X1 _14891_ (
    .A1(divisor[14]),
    .A2(remainder[3]),
    .ZN(_04642_)
  );
  INV_X1 _14892_ (
    .A(_04642_),
    .ZN(_04643_)
  );
  AND2_X1 _14893_ (
    .A1(divisor[15]),
    .A2(remainder[3]),
    .ZN(_04644_)
  );
  INV_X1 _14894_ (
    .A(_04644_),
    .ZN(_04646_)
  );
  AND2_X1 _14895_ (
    .A1(_04372_),
    .A2(_04642_),
    .ZN(_04647_)
  );
  INV_X1 _14896_ (
    .A(_04647_),
    .ZN(_04648_)
  );
  AND2_X1 _14897_ (
    .A1(_04373_),
    .A2(_04643_),
    .ZN(_04649_)
  );
  INV_X1 _14898_ (
    .A(_04649_),
    .ZN(_04650_)
  );
  AND2_X1 _14899_ (
    .A1(_04648_),
    .A2(_04650_),
    .ZN(_04651_)
  );
  INV_X1 _14900_ (
    .A(_04651_),
    .ZN(_04652_)
  );
  AND2_X1 _14901_ (
    .A1(_04640_),
    .A2(_04651_),
    .ZN(_04653_)
  );
  INV_X1 _14902_ (
    .A(_04653_),
    .ZN(_04654_)
  );
  AND2_X1 _14903_ (
    .A1(_04641_),
    .A2(_04652_),
    .ZN(_04655_)
  );
  INV_X1 _14904_ (
    .A(_04655_),
    .ZN(_04657_)
  );
  AND2_X1 _14905_ (
    .A1(_04654_),
    .A2(_04657_),
    .ZN(_04658_)
  );
  INV_X1 _14906_ (
    .A(_04658_),
    .ZN(_04659_)
  );
  AND2_X1 _14907_ (
    .A1(_04639_),
    .A2(_04658_),
    .ZN(_04660_)
  );
  INV_X1 _14908_ (
    .A(_04660_),
    .ZN(_04661_)
  );
  AND2_X1 _14909_ (
    .A1(_04638_),
    .A2(_04659_),
    .ZN(_04662_)
  );
  INV_X1 _14910_ (
    .A(_04662_),
    .ZN(_04663_)
  );
  AND2_X1 _14911_ (
    .A1(_04661_),
    .A2(_04663_),
    .ZN(_04664_)
  );
  INV_X1 _14912_ (
    .A(_04664_),
    .ZN(_04665_)
  );
  AND2_X1 _14913_ (
    .A1(divisor[10]),
    .A2(remainder[7]),
    .ZN(_04666_)
  );
  INV_X1 _14914_ (
    .A(_04666_),
    .ZN(_04668_)
  );
  AND2_X1 _14915_ (
    .A1(divisor[11]),
    .A2(remainder[6]),
    .ZN(_04669_)
  );
  INV_X1 _14916_ (
    .A(_04669_),
    .ZN(_04670_)
  );
  AND2_X1 _14917_ (
    .A1(divisor[12]),
    .A2(remainder[6]),
    .ZN(_04671_)
  );
  INV_X1 _14918_ (
    .A(_04671_),
    .ZN(_04672_)
  );
  AND2_X1 _14919_ (
    .A1(_04396_),
    .A2(_04669_),
    .ZN(_04673_)
  );
  INV_X1 _14920_ (
    .A(_04673_),
    .ZN(_04674_)
  );
  AND2_X1 _14921_ (
    .A1(_04397_),
    .A2(_04670_),
    .ZN(_04675_)
  );
  INV_X1 _14922_ (
    .A(_04675_),
    .ZN(_04676_)
  );
  AND2_X1 _14923_ (
    .A1(_04674_),
    .A2(_04676_),
    .ZN(_04677_)
  );
  INV_X1 _14924_ (
    .A(_04677_),
    .ZN(_04679_)
  );
  AND2_X1 _14925_ (
    .A1(_04666_),
    .A2(_04677_),
    .ZN(_04680_)
  );
  INV_X1 _14926_ (
    .A(_04680_),
    .ZN(_04681_)
  );
  AND2_X1 _14927_ (
    .A1(_04668_),
    .A2(_04679_),
    .ZN(_04682_)
  );
  INV_X1 _14928_ (
    .A(_04682_),
    .ZN(_04683_)
  );
  AND2_X1 _14929_ (
    .A1(_04681_),
    .A2(_04683_),
    .ZN(_04684_)
  );
  INV_X1 _14930_ (
    .A(_04684_),
    .ZN(_04685_)
  );
  AND2_X1 _14931_ (
    .A1(_04664_),
    .A2(_04684_),
    .ZN(_04686_)
  );
  INV_X1 _14932_ (
    .A(_04686_),
    .ZN(_04687_)
  );
  AND2_X1 _14933_ (
    .A1(_04665_),
    .A2(_04685_),
    .ZN(_04688_)
  );
  INV_X1 _14934_ (
    .A(_04688_),
    .ZN(_04690_)
  );
  AND2_X1 _14935_ (
    .A1(_04687_),
    .A2(_04690_),
    .ZN(_04691_)
  );
  INV_X1 _14936_ (
    .A(_04691_),
    .ZN(_04692_)
  );
  AND2_X1 _14937_ (
    .A1(_04637_),
    .A2(_04691_),
    .ZN(_04693_)
  );
  INV_X1 _14938_ (
    .A(_04693_),
    .ZN(_04694_)
  );
  AND2_X1 _14939_ (
    .A1(_04636_),
    .A2(_04692_),
    .ZN(_04695_)
  );
  INV_X1 _14940_ (
    .A(_04695_),
    .ZN(_04696_)
  );
  AND2_X1 _14941_ (
    .A1(_04694_),
    .A2(_04696_),
    .ZN(_04697_)
  );
  INV_X1 _14942_ (
    .A(_04697_),
    .ZN(_04698_)
  );
  AND2_X1 _14943_ (
    .A1(_04435_),
    .A2(_04442_),
    .ZN(_04699_)
  );
  INV_X1 _14944_ (
    .A(_04699_),
    .ZN(_04701_)
  );
  AND2_X1 _14945_ (
    .A1(_04399_),
    .A2(_04406_),
    .ZN(_04702_)
  );
  INV_X1 _14946_ (
    .A(_04702_),
    .ZN(_04703_)
  );
  MUX2_X1 _14947_ (
    .A(_04430_),
    .B(_04908_),
    .S(_04429_),
    .Z(_04704_)
  );
  AND2_X1 _14948_ (
    .A1(divisor[7]),
    .A2(_04704_),
    .ZN(_04705_)
  );
  INV_X1 _14949_ (
    .A(_04705_),
    .ZN(_04706_)
  );
  MUX2_X1 _14950_ (
    .A(_04189_),
    .B(_04897_),
    .S(_04704_),
    .Z(_04707_)
  );
  MUX2_X1 _14951_ (
    .A(_04190_),
    .B(divisor[7]),
    .S(_04704_),
    .Z(_04708_)
  );
  AND2_X1 _14952_ (
    .A1(_04703_),
    .A2(_04707_),
    .ZN(_04709_)
  );
  INV_X1 _14953_ (
    .A(_04709_),
    .ZN(_04710_)
  );
  AND2_X1 _14954_ (
    .A1(_04702_),
    .A2(_04708_),
    .ZN(_04712_)
  );
  INV_X1 _14955_ (
    .A(_04712_),
    .ZN(_04713_)
  );
  AND2_X1 _14956_ (
    .A1(_04710_),
    .A2(_04713_),
    .ZN(_04714_)
  );
  INV_X1 _14957_ (
    .A(_04714_),
    .ZN(_04715_)
  );
  AND2_X1 _14958_ (
    .A1(_04701_),
    .A2(_04714_),
    .ZN(_04716_)
  );
  INV_X1 _14959_ (
    .A(_04716_),
    .ZN(_04717_)
  );
  AND2_X1 _14960_ (
    .A1(_04699_),
    .A2(_04715_),
    .ZN(_04718_)
  );
  INV_X1 _14961_ (
    .A(_04718_),
    .ZN(_04719_)
  );
  AND2_X1 _14962_ (
    .A1(_04717_),
    .A2(_04719_),
    .ZN(_04720_)
  );
  INV_X1 _14963_ (
    .A(_04720_),
    .ZN(_04721_)
  );
  AND2_X1 _14964_ (
    .A1(_04697_),
    .A2(_04720_),
    .ZN(_04723_)
  );
  INV_X1 _14965_ (
    .A(_04723_),
    .ZN(_04724_)
  );
  AND2_X1 _14966_ (
    .A1(_04698_),
    .A2(_04721_),
    .ZN(_04725_)
  );
  INV_X1 _14967_ (
    .A(_04725_),
    .ZN(_04726_)
  );
  AND2_X1 _14968_ (
    .A1(_04724_),
    .A2(_04726_),
    .ZN(_04727_)
  );
  INV_X1 _14969_ (
    .A(_04727_),
    .ZN(_04728_)
  );
  AND2_X1 _14970_ (
    .A1(_04633_),
    .A2(_04727_),
    .ZN(_04729_)
  );
  INV_X1 _14971_ (
    .A(_04729_),
    .ZN(_04730_)
  );
  AND2_X1 _14972_ (
    .A1(_04635_),
    .A2(_04728_),
    .ZN(_04731_)
  );
  INV_X1 _14973_ (
    .A(_04731_),
    .ZN(_04732_)
  );
  AND2_X1 _14974_ (
    .A1(_04730_),
    .A2(_04732_),
    .ZN(_04734_)
  );
  INV_X1 _14975_ (
    .A(_04734_),
    .ZN(_04735_)
  );
  AND2_X1 _14976_ (
    .A1(_04467_),
    .A2(_04734_),
    .ZN(_04736_)
  );
  INV_X1 _14977_ (
    .A(_04736_),
    .ZN(_04737_)
  );
  AND2_X1 _14978_ (
    .A1(_04468_),
    .A2(_04735_),
    .ZN(_04738_)
  );
  INV_X1 _14979_ (
    .A(_04738_),
    .ZN(_04739_)
  );
  AND2_X1 _14980_ (
    .A1(_04737_),
    .A2(_04739_),
    .ZN(_04740_)
  );
  INV_X1 _14981_ (
    .A(_04740_),
    .ZN(_04741_)
  );
  AND2_X1 _14982_ (
    .A1(_04559_),
    .A2(_04741_),
    .ZN(_04742_)
  );
  INV_X1 _14983_ (
    .A(_04742_),
    .ZN(_04743_)
  );
  AND2_X1 _14984_ (
    .A1(_04560_),
    .A2(_04740_),
    .ZN(_04745_)
  );
  INV_X1 _14985_ (
    .A(_04745_),
    .ZN(_04746_)
  );
  AND2_X1 _14986_ (
    .A1(_04743_),
    .A2(_04746_),
    .ZN(_04747_)
  );
  INV_X1 _14987_ (
    .A(_04747_),
    .ZN(_04748_)
  );
  AND2_X1 _14988_ (
    .A1(_04620_),
    .A2(_04748_),
    .ZN(_04749_)
  );
  INV_X1 _14989_ (
    .A(_04749_),
    .ZN(_04750_)
  );
  AND2_X1 _14990_ (
    .A1(_04621_),
    .A2(_04747_),
    .ZN(_04751_)
  );
  INV_X1 _14991_ (
    .A(_04751_),
    .ZN(_04752_)
  );
  AND2_X1 _14992_ (
    .A1(_04750_),
    .A2(_04752_),
    .ZN(_04753_)
  );
  INV_X1 _14993_ (
    .A(_04753_),
    .ZN(_04754_)
  );
  AND2_X1 _14994_ (
    .A1(_04564_),
    .A2(_04753_),
    .ZN(_04756_)
  );
  INV_X1 _14995_ (
    .A(_04756_),
    .ZN(_04757_)
  );
  AND2_X1 _14996_ (
    .A1(_04563_),
    .A2(_04754_),
    .ZN(_04758_)
  );
  INV_X1 _14997_ (
    .A(_04758_),
    .ZN(_04759_)
  );
  AND2_X1 _14998_ (
    .A1(_04757_),
    .A2(_04759_),
    .ZN(_04760_)
  );
  INV_X1 _14999_ (
    .A(_04760_),
    .ZN(_04761_)
  );
  AND2_X1 _15000_ (
    .A1(_04356_),
    .A2(_04760_),
    .ZN(_04762_)
  );
  INV_X1 _15001_ (
    .A(_04762_),
    .ZN(_04763_)
  );
  AND2_X1 _15002_ (
    .A1(_04357_),
    .A2(_04761_),
    .ZN(_04764_)
  );
  INV_X1 _15003_ (
    .A(_04764_),
    .ZN(_04765_)
  );
  AND2_X1 _15004_ (
    .A1(_04763_),
    .A2(_04765_),
    .ZN(_04767_)
  );
  INV_X1 _15005_ (
    .A(_04767_),
    .ZN(_04768_)
  );
  AND2_X1 _15006_ (
    .A1(_04558_),
    .A2(_04767_),
    .ZN(_04769_)
  );
  INV_X1 _15007_ (
    .A(_04769_),
    .ZN(_04770_)
  );
  AND2_X1 _15008_ (
    .A1(_04556_),
    .A2(_04768_),
    .ZN(_04771_)
  );
  INV_X1 _15009_ (
    .A(_04771_),
    .ZN(_04772_)
  );
  AND2_X1 _15010_ (
    .A1(_04770_),
    .A2(_04772_),
    .ZN(_04773_)
  );
  INV_X1 _15011_ (
    .A(_04773_),
    .ZN(_04774_)
  );
  AND2_X1 _15012_ (
    .A1(_04505_),
    .A2(_04773_),
    .ZN(_04775_)
  );
  INV_X1 _15013_ (
    .A(_04775_),
    .ZN(_04776_)
  );
  AND2_X1 _15014_ (
    .A1(_04506_),
    .A2(_04774_),
    .ZN(_04778_)
  );
  INV_X1 _15015_ (
    .A(_04778_),
    .ZN(_04779_)
  );
  AND2_X1 _15016_ (
    .A1(_04776_),
    .A2(_04779_),
    .ZN(_04780_)
  );
  INV_X1 _15017_ (
    .A(_04780_),
    .ZN(_04781_)
  );
  AND2_X1 _15018_ (
    .A1(_04555_),
    .A2(_04781_),
    .ZN(_04782_)
  );
  INV_X1 _15019_ (
    .A(_04782_),
    .ZN(_04783_)
  );
  AND2_X1 _15020_ (
    .A1(_04554_),
    .A2(_04780_),
    .ZN(_04784_)
  );
  INV_X1 _15021_ (
    .A(_04784_),
    .ZN(_04785_)
  );
  AND2_X1 _15022_ (
    .A1(_04555_),
    .A2(_04780_),
    .ZN(_04786_)
  );
  INV_X1 _15023_ (
    .A(_04786_),
    .ZN(_04787_)
  );
  AND2_X1 _15024_ (
    .A1(_04554_),
    .A2(_04781_),
    .ZN(_04789_)
  );
  INV_X1 _15025_ (
    .A(_04789_),
    .ZN(_04790_)
  );
  AND2_X1 _15026_ (
    .A1(_04783_),
    .A2(_04785_),
    .ZN(_04791_)
  );
  AND2_X1 _15027_ (
    .A1(_04787_),
    .A2(_04790_),
    .ZN(_04792_)
  );
  AND2_X1 _15028_ (
    .A1(remainder[50]),
    .A2(_04792_),
    .ZN(_04793_)
  );
  INV_X1 _15029_ (
    .A(_04793_),
    .ZN(_04794_)
  );
  AND2_X1 _15030_ (
    .A1(_04568_),
    .A2(_04791_),
    .ZN(_04795_)
  );
  INV_X1 _15031_ (
    .A(_04795_),
    .ZN(_04796_)
  );
  AND2_X1 _15032_ (
    .A1(_04794_),
    .A2(_04796_),
    .ZN(_04797_)
  );
  INV_X1 _15033_ (
    .A(_04797_),
    .ZN(_04798_)
  );
  AND2_X1 _15034_ (
    .A1(_04553_),
    .A2(_04797_),
    .ZN(_04800_)
  );
  INV_X1 _15035_ (
    .A(_04800_),
    .ZN(_04801_)
  );
  AND2_X1 _15036_ (
    .A1(_04552_),
    .A2(_04798_),
    .ZN(_04802_)
  );
  INV_X1 _15037_ (
    .A(_04802_),
    .ZN(_04803_)
  );
  AND2_X1 _15038_ (
    .A1(_02082_),
    .A2(_04803_),
    .ZN(_04804_)
  );
  AND2_X1 _15039_ (
    .A1(_04801_),
    .A2(_04804_),
    .ZN(_04805_)
  );
  INV_X1 _15040_ (
    .A(_04805_),
    .ZN(_04806_)
  );
  AND2_X1 _15041_ (
    .A1(_04551_),
    .A2(_04806_),
    .ZN(_04807_)
  );
  AND2_X1 _15042_ (
    .A1(_04549_),
    .A2(_04807_),
    .ZN(_04808_)
  );
  INV_X1 _15043_ (
    .A(_04808_),
    .ZN(_04809_)
  );
  AND2_X1 _15044_ (
    .A1(_06201_),
    .A2(_04809_),
    .ZN(_00063_)
  );
  AND2_X1 _15045_ (
    .A1(_04656_),
    .A2(_10451_),
    .ZN(_04811_)
  );
  INV_X1 _15046_ (
    .A(_04811_),
    .ZN(_04812_)
  );
  AND2_X1 _15047_ (
    .A1(_10462_),
    .A2(_01748_),
    .ZN(_04813_)
  );
  INV_X1 _15048_ (
    .A(_04813_),
    .ZN(_04814_)
  );
  AND2_X1 _15049_ (
    .A1(_05983_),
    .A2(_04814_),
    .ZN(_04815_)
  );
  AND2_X1 _15050_ (
    .A1(_04812_),
    .A2(_04815_),
    .ZN(_04816_)
  );
  INV_X1 _15051_ (
    .A(_04816_),
    .ZN(_04817_)
  );
  AND2_X1 _15052_ (
    .A1(remainder[43]),
    .A2(_02077_),
    .ZN(_04818_)
  );
  INV_X1 _15053_ (
    .A(_04818_),
    .ZN(_04819_)
  );
  AND2_X1 _15054_ (
    .A1(_04518_),
    .A2(_04780_),
    .ZN(_04821_)
  );
  INV_X1 _15055_ (
    .A(_04821_),
    .ZN(_04822_)
  );
  AND2_X1 _15056_ (
    .A1(_04511_),
    .A2(_04779_),
    .ZN(_04823_)
  );
  INV_X1 _15057_ (
    .A(_04823_),
    .ZN(_04824_)
  );
  AND2_X1 _15058_ (
    .A1(_04776_),
    .A2(_04824_),
    .ZN(_04825_)
  );
  AND2_X1 _15059_ (
    .A1(_04822_),
    .A2(_04825_),
    .ZN(_04826_)
  );
  INV_X1 _15060_ (
    .A(_04826_),
    .ZN(_04827_)
  );
  AND2_X1 _15061_ (
    .A1(_04757_),
    .A2(_04763_),
    .ZN(_04828_)
  );
  INV_X1 _15062_ (
    .A(_04828_),
    .ZN(_04829_)
  );
  AND2_X1 _15063_ (
    .A1(_03249_),
    .A2(_04741_),
    .ZN(_04830_)
  );
  INV_X1 _15064_ (
    .A(_04830_),
    .ZN(_04832_)
  );
  AND2_X1 _15065_ (
    .A1(_04472_),
    .A2(_04830_),
    .ZN(_04833_)
  );
  INV_X1 _15066_ (
    .A(_04833_),
    .ZN(_04834_)
  );
  AND2_X1 _15067_ (
    .A1(_04750_),
    .A2(_04834_),
    .ZN(_04835_)
  );
  INV_X1 _15068_ (
    .A(_04835_),
    .ZN(_04836_)
  );
  AND2_X1 _15069_ (
    .A1(_04604_),
    .A2(_04610_),
    .ZN(_04837_)
  );
  INV_X1 _15070_ (
    .A(_04837_),
    .ZN(_04838_)
  );
  AND2_X1 _15071_ (
    .A1(_04591_),
    .A2(_04597_),
    .ZN(_04839_)
  );
  INV_X1 _15072_ (
    .A(_04839_),
    .ZN(_04840_)
  );
  AND2_X1 _15073_ (
    .A1(_04577_),
    .A2(_04584_),
    .ZN(_04841_)
  );
  INV_X1 _15074_ (
    .A(_04841_),
    .ZN(_04843_)
  );
  AND2_X1 _15075_ (
    .A1(_04694_),
    .A2(_04724_),
    .ZN(_04844_)
  );
  INV_X1 _15076_ (
    .A(_04844_),
    .ZN(_04845_)
  );
  AND2_X1 _15077_ (
    .A1(_04710_),
    .A2(_04717_),
    .ZN(_04846_)
  );
  INV_X1 _15078_ (
    .A(_04846_),
    .ZN(_04847_)
  );
  AND2_X1 _15079_ (
    .A1(_04087_),
    .A2(_04847_),
    .ZN(_04848_)
  );
  INV_X1 _15080_ (
    .A(_04848_),
    .ZN(_04849_)
  );
  AND2_X1 _15081_ (
    .A1(_04088_),
    .A2(_04846_),
    .ZN(_04850_)
  );
  INV_X1 _15082_ (
    .A(_04850_),
    .ZN(_04851_)
  );
  AND2_X1 _15083_ (
    .A1(_04849_),
    .A2(_04851_),
    .ZN(_04852_)
  );
  INV_X1 _15084_ (
    .A(_04852_),
    .ZN(_04854_)
  );
  AND2_X1 _15085_ (
    .A1(_04317_),
    .A2(_04852_),
    .ZN(_04855_)
  );
  INV_X1 _15086_ (
    .A(_04855_),
    .ZN(_04856_)
  );
  AND2_X1 _15087_ (
    .A1(_04316_),
    .A2(_04854_),
    .ZN(_04857_)
  );
  INV_X1 _15088_ (
    .A(_04857_),
    .ZN(_04858_)
  );
  AND2_X1 _15089_ (
    .A1(_04856_),
    .A2(_04858_),
    .ZN(_04859_)
  );
  INV_X1 _15090_ (
    .A(_04859_),
    .ZN(_04860_)
  );
  AND2_X1 _15091_ (
    .A1(_04845_),
    .A2(_04859_),
    .ZN(_04861_)
  );
  INV_X1 _15092_ (
    .A(_04861_),
    .ZN(_04862_)
  );
  AND2_X1 _15093_ (
    .A1(_04844_),
    .A2(_04860_),
    .ZN(_04863_)
  );
  INV_X1 _15094_ (
    .A(_04863_),
    .ZN(_04865_)
  );
  AND2_X1 _15095_ (
    .A1(_04862_),
    .A2(_04865_),
    .ZN(_04866_)
  );
  INV_X1 _15096_ (
    .A(_04866_),
    .ZN(_04867_)
  );
  AND2_X1 _15097_ (
    .A1(_04843_),
    .A2(_04866_),
    .ZN(_04868_)
  );
  INV_X1 _15098_ (
    .A(_04868_),
    .ZN(_04869_)
  );
  AND2_X1 _15099_ (
    .A1(_04841_),
    .A2(_04867_),
    .ZN(_04870_)
  );
  INV_X1 _15100_ (
    .A(_04870_),
    .ZN(_04871_)
  );
  AND2_X1 _15101_ (
    .A1(_04869_),
    .A2(_04871_),
    .ZN(_04872_)
  );
  INV_X1 _15102_ (
    .A(_04872_),
    .ZN(_04873_)
  );
  AND2_X1 _15103_ (
    .A1(_04840_),
    .A2(_04872_),
    .ZN(_04874_)
  );
  INV_X1 _15104_ (
    .A(_04874_),
    .ZN(_04876_)
  );
  AND2_X1 _15105_ (
    .A1(_04839_),
    .A2(_04873_),
    .ZN(_04877_)
  );
  INV_X1 _15106_ (
    .A(_04877_),
    .ZN(_04878_)
  );
  AND2_X1 _15107_ (
    .A1(_04876_),
    .A2(_04878_),
    .ZN(_04879_)
  );
  INV_X1 _15108_ (
    .A(_04879_),
    .ZN(_04880_)
  );
  AND2_X1 _15109_ (
    .A1(_03170_),
    .A2(_04879_),
    .ZN(_04881_)
  );
  INV_X1 _15110_ (
    .A(_04881_),
    .ZN(_04882_)
  );
  AND2_X1 _15111_ (
    .A1(_03169_),
    .A2(_04880_),
    .ZN(_04883_)
  );
  INV_X1 _15112_ (
    .A(_04883_),
    .ZN(_04884_)
  );
  AND2_X1 _15113_ (
    .A1(_04882_),
    .A2(_04884_),
    .ZN(_04885_)
  );
  INV_X1 _15114_ (
    .A(_04885_),
    .ZN(_04887_)
  );
  AND2_X1 _15115_ (
    .A1(_04736_),
    .A2(_04885_),
    .ZN(_04888_)
  );
  INV_X1 _15116_ (
    .A(_04888_),
    .ZN(_04889_)
  );
  AND2_X1 _15117_ (
    .A1(_04737_),
    .A2(_04887_),
    .ZN(_04890_)
  );
  INV_X1 _15118_ (
    .A(_04890_),
    .ZN(_04891_)
  );
  AND2_X1 _15119_ (
    .A1(_04889_),
    .A2(_04891_),
    .ZN(_04892_)
  );
  INV_X1 _15120_ (
    .A(_04892_),
    .ZN(_04893_)
  );
  AND2_X1 _15121_ (
    .A1(_04838_),
    .A2(_04892_),
    .ZN(_04894_)
  );
  INV_X1 _15122_ (
    .A(_04894_),
    .ZN(_04895_)
  );
  AND2_X1 _15123_ (
    .A1(_04837_),
    .A2(_04893_),
    .ZN(_04896_)
  );
  INV_X1 _15124_ (
    .A(_04896_),
    .ZN(_04898_)
  );
  AND2_X1 _15125_ (
    .A1(_04895_),
    .A2(_04898_),
    .ZN(_04899_)
  );
  INV_X1 _15126_ (
    .A(_04899_),
    .ZN(_04900_)
  );
  AND2_X1 _15127_ (
    .A1(divisor[16]),
    .A2(remainder[2]),
    .ZN(_04901_)
  );
  INV_X1 _15128_ (
    .A(_04901_),
    .ZN(_04902_)
  );
  AND2_X1 _15129_ (
    .A1(divisor[18]),
    .A2(remainder[0]),
    .ZN(_04903_)
  );
  INV_X1 _15130_ (
    .A(_04903_),
    .ZN(_04904_)
  );
  AND2_X1 _15131_ (
    .A1(divisor[18]),
    .A2(remainder[1]),
    .ZN(_04905_)
  );
  INV_X1 _15132_ (
    .A(_04905_),
    .ZN(_04906_)
  );
  AND2_X1 _15133_ (
    .A1(_04622_),
    .A2(_04905_),
    .ZN(_04907_)
  );
  INV_X1 _15134_ (
    .A(_04907_),
    .ZN(_04909_)
  );
  AND2_X1 _15135_ (
    .A1(_04628_),
    .A2(_04904_),
    .ZN(_04910_)
  );
  INV_X1 _15136_ (
    .A(_04910_),
    .ZN(_04911_)
  );
  AND2_X1 _15137_ (
    .A1(_04909_),
    .A2(_04911_),
    .ZN(_04912_)
  );
  INV_X1 _15138_ (
    .A(_04912_),
    .ZN(_04913_)
  );
  AND2_X1 _15139_ (
    .A1(_04901_),
    .A2(_04912_),
    .ZN(_04914_)
  );
  INV_X1 _15140_ (
    .A(_04914_),
    .ZN(_04915_)
  );
  AND2_X1 _15141_ (
    .A1(_04902_),
    .A2(_04913_),
    .ZN(_04916_)
  );
  INV_X1 _15142_ (
    .A(_04916_),
    .ZN(_04917_)
  );
  AND2_X1 _15143_ (
    .A1(_04915_),
    .A2(_04917_),
    .ZN(_04918_)
  );
  INV_X1 _15144_ (
    .A(_04918_),
    .ZN(_04920_)
  );
  AND2_X1 _15145_ (
    .A1(_04629_),
    .A2(_04918_),
    .ZN(_04921_)
  );
  INV_X1 _15146_ (
    .A(_04921_),
    .ZN(_04922_)
  );
  AND2_X1 _15147_ (
    .A1(_04630_),
    .A2(_04920_),
    .ZN(_04923_)
  );
  INV_X1 _15148_ (
    .A(_04923_),
    .ZN(_04924_)
  );
  AND2_X1 _15149_ (
    .A1(_04922_),
    .A2(_04924_),
    .ZN(_04925_)
  );
  INV_X1 _15150_ (
    .A(_04925_),
    .ZN(_04926_)
  );
  AND2_X1 _15151_ (
    .A1(_04661_),
    .A2(_04687_),
    .ZN(_04927_)
  );
  INV_X1 _15152_ (
    .A(_04927_),
    .ZN(_04928_)
  );
  AND2_X1 _15153_ (
    .A1(_04648_),
    .A2(_04654_),
    .ZN(_04929_)
  );
  INV_X1 _15154_ (
    .A(_04929_),
    .ZN(_04931_)
  );
  AND2_X1 _15155_ (
    .A1(divisor[13]),
    .A2(remainder[5]),
    .ZN(_04932_)
  );
  INV_X1 _15156_ (
    .A(_04932_),
    .ZN(_04933_)
  );
  AND2_X1 _15157_ (
    .A1(divisor[14]),
    .A2(remainder[4]),
    .ZN(_04934_)
  );
  INV_X1 _15158_ (
    .A(_04934_),
    .ZN(_04935_)
  );
  AND2_X1 _15159_ (
    .A1(divisor[15]),
    .A2(remainder[4]),
    .ZN(_04936_)
  );
  INV_X1 _15160_ (
    .A(_04936_),
    .ZN(_04937_)
  );
  AND2_X1 _15161_ (
    .A1(_04644_),
    .A2(_04934_),
    .ZN(_04938_)
  );
  INV_X1 _15162_ (
    .A(_04938_),
    .ZN(_04939_)
  );
  AND2_X1 _15163_ (
    .A1(_04646_),
    .A2(_04935_),
    .ZN(_04940_)
  );
  INV_X1 _15164_ (
    .A(_04940_),
    .ZN(_04942_)
  );
  AND2_X1 _15165_ (
    .A1(_04939_),
    .A2(_04942_),
    .ZN(_04943_)
  );
  INV_X1 _15166_ (
    .A(_04943_),
    .ZN(_04944_)
  );
  AND2_X1 _15167_ (
    .A1(_04932_),
    .A2(_04943_),
    .ZN(_04945_)
  );
  INV_X1 _15168_ (
    .A(_04945_),
    .ZN(_04946_)
  );
  AND2_X1 _15169_ (
    .A1(_04933_),
    .A2(_04944_),
    .ZN(_04947_)
  );
  INV_X1 _15170_ (
    .A(_04947_),
    .ZN(_04948_)
  );
  AND2_X1 _15171_ (
    .A1(_04946_),
    .A2(_04948_),
    .ZN(_04949_)
  );
  INV_X1 _15172_ (
    .A(_04949_),
    .ZN(_04950_)
  );
  AND2_X1 _15173_ (
    .A1(_04931_),
    .A2(_04949_),
    .ZN(_04951_)
  );
  INV_X1 _15174_ (
    .A(_04951_),
    .ZN(_04953_)
  );
  AND2_X1 _15175_ (
    .A1(_04929_),
    .A2(_04950_),
    .ZN(_04954_)
  );
  INV_X1 _15176_ (
    .A(_04954_),
    .ZN(_04955_)
  );
  AND2_X1 _15177_ (
    .A1(_04953_),
    .A2(_04955_),
    .ZN(_04956_)
  );
  INV_X1 _15178_ (
    .A(_04956_),
    .ZN(_04957_)
  );
  AND2_X1 _15179_ (
    .A1(remainder[32]),
    .A2(divisor[10]),
    .ZN(_04958_)
  );
  INV_X1 _15180_ (
    .A(_04958_),
    .ZN(_04959_)
  );
  AND2_X1 _15181_ (
    .A1(divisor[11]),
    .A2(remainder[7]),
    .ZN(_04960_)
  );
  INV_X1 _15182_ (
    .A(_04960_),
    .ZN(_04961_)
  );
  AND2_X1 _15183_ (
    .A1(divisor[12]),
    .A2(remainder[7]),
    .ZN(_04962_)
  );
  INV_X1 _15184_ (
    .A(_04962_),
    .ZN(_04964_)
  );
  AND2_X1 _15185_ (
    .A1(_04669_),
    .A2(_04962_),
    .ZN(_04965_)
  );
  INV_X1 _15186_ (
    .A(_04965_),
    .ZN(_04966_)
  );
  AND2_X1 _15187_ (
    .A1(_04672_),
    .A2(_04961_),
    .ZN(_04967_)
  );
  INV_X1 _15188_ (
    .A(_04967_),
    .ZN(_04968_)
  );
  AND2_X1 _15189_ (
    .A1(_04966_),
    .A2(_04968_),
    .ZN(_04969_)
  );
  INV_X1 _15190_ (
    .A(_04969_),
    .ZN(_04970_)
  );
  AND2_X1 _15191_ (
    .A1(_04958_),
    .A2(_04969_),
    .ZN(_04971_)
  );
  INV_X1 _15192_ (
    .A(_04971_),
    .ZN(_04972_)
  );
  AND2_X1 _15193_ (
    .A1(_04959_),
    .A2(_04970_),
    .ZN(_04973_)
  );
  INV_X1 _15194_ (
    .A(_04973_),
    .ZN(_04975_)
  );
  AND2_X1 _15195_ (
    .A1(_04972_),
    .A2(_04975_),
    .ZN(_04976_)
  );
  INV_X1 _15196_ (
    .A(_04976_),
    .ZN(_04977_)
  );
  AND2_X1 _15197_ (
    .A1(_04956_),
    .A2(_04976_),
    .ZN(_04978_)
  );
  INV_X1 _15198_ (
    .A(_04978_),
    .ZN(_04979_)
  );
  AND2_X1 _15199_ (
    .A1(_04957_),
    .A2(_04977_),
    .ZN(_04980_)
  );
  INV_X1 _15200_ (
    .A(_04980_),
    .ZN(_04981_)
  );
  AND2_X1 _15201_ (
    .A1(_04979_),
    .A2(_04981_),
    .ZN(_04982_)
  );
  INV_X1 _15202_ (
    .A(_04982_),
    .ZN(_04983_)
  );
  AND2_X1 _15203_ (
    .A1(_04928_),
    .A2(_04982_),
    .ZN(_04984_)
  );
  INV_X1 _15204_ (
    .A(_04984_),
    .ZN(_04986_)
  );
  AND2_X1 _15205_ (
    .A1(_04927_),
    .A2(_04983_),
    .ZN(_04987_)
  );
  INV_X1 _15206_ (
    .A(_04987_),
    .ZN(_04988_)
  );
  AND2_X1 _15207_ (
    .A1(_04986_),
    .A2(_04988_),
    .ZN(_04989_)
  );
  INV_X1 _15208_ (
    .A(_04989_),
    .ZN(_04990_)
  );
  AND2_X1 _15209_ (
    .A1(_04433_),
    .A2(_04706_),
    .ZN(_04991_)
  );
  INV_X1 _15210_ (
    .A(_04991_),
    .ZN(_04992_)
  );
  AND2_X1 _15211_ (
    .A1(_04674_),
    .A2(_04681_),
    .ZN(_04993_)
  );
  INV_X1 _15212_ (
    .A(_04993_),
    .ZN(_04994_)
  );
  AND2_X1 _15213_ (
    .A1(_04707_),
    .A2(_04994_),
    .ZN(_04995_)
  );
  INV_X1 _15214_ (
    .A(_04995_),
    .ZN(_04997_)
  );
  AND2_X1 _15215_ (
    .A1(_04708_),
    .A2(_04993_),
    .ZN(_04998_)
  );
  INV_X1 _15216_ (
    .A(_04998_),
    .ZN(_04999_)
  );
  AND2_X1 _15217_ (
    .A1(_04997_),
    .A2(_04999_),
    .ZN(_05000_)
  );
  INV_X1 _15218_ (
    .A(_05000_),
    .ZN(_05001_)
  );
  AND2_X1 _15219_ (
    .A1(_04992_),
    .A2(_05000_),
    .ZN(_05002_)
  );
  INV_X1 _15220_ (
    .A(_05002_),
    .ZN(_05003_)
  );
  AND2_X1 _15221_ (
    .A1(_04991_),
    .A2(_05001_),
    .ZN(_05004_)
  );
  INV_X1 _15222_ (
    .A(_05004_),
    .ZN(_05005_)
  );
  AND2_X1 _15223_ (
    .A1(_05003_),
    .A2(_05005_),
    .ZN(_05006_)
  );
  INV_X1 _15224_ (
    .A(_05006_),
    .ZN(_05008_)
  );
  AND2_X1 _15225_ (
    .A1(_04989_),
    .A2(_05006_),
    .ZN(_05009_)
  );
  INV_X1 _15226_ (
    .A(_05009_),
    .ZN(_05010_)
  );
  AND2_X1 _15227_ (
    .A1(_04990_),
    .A2(_05008_),
    .ZN(_05011_)
  );
  INV_X1 _15228_ (
    .A(_05011_),
    .ZN(_05012_)
  );
  AND2_X1 _15229_ (
    .A1(_05010_),
    .A2(_05012_),
    .ZN(_05013_)
  );
  INV_X1 _15230_ (
    .A(_05013_),
    .ZN(_05014_)
  );
  AND2_X1 _15231_ (
    .A1(_04925_),
    .A2(_05013_),
    .ZN(_05015_)
  );
  INV_X1 _15232_ (
    .A(_05015_),
    .ZN(_05016_)
  );
  AND2_X1 _15233_ (
    .A1(_04926_),
    .A2(_05014_),
    .ZN(_05017_)
  );
  INV_X1 _15234_ (
    .A(_05017_),
    .ZN(_05019_)
  );
  AND2_X1 _15235_ (
    .A1(_05016_),
    .A2(_05019_),
    .ZN(_05020_)
  );
  INV_X1 _15236_ (
    .A(_05020_),
    .ZN(_05021_)
  );
  AND2_X1 _15237_ (
    .A1(_04729_),
    .A2(_05020_),
    .ZN(_05022_)
  );
  INV_X1 _15238_ (
    .A(_05022_),
    .ZN(_05023_)
  );
  AND2_X1 _15239_ (
    .A1(_04730_),
    .A2(_05021_),
    .ZN(_05024_)
  );
  INV_X1 _15240_ (
    .A(_05024_),
    .ZN(_05025_)
  );
  AND2_X1 _15241_ (
    .A1(_05023_),
    .A2(_05025_),
    .ZN(_05026_)
  );
  INV_X1 _15242_ (
    .A(_05026_),
    .ZN(_05027_)
  );
  AND2_X1 _15243_ (
    .A1(_04832_),
    .A2(_05027_),
    .ZN(_05028_)
  );
  INV_X1 _15244_ (
    .A(_05028_),
    .ZN(_05030_)
  );
  AND2_X1 _15245_ (
    .A1(_04830_),
    .A2(_05026_),
    .ZN(_05031_)
  );
  INV_X1 _15246_ (
    .A(_05031_),
    .ZN(_05032_)
  );
  AND2_X1 _15247_ (
    .A1(_04832_),
    .A2(_05026_),
    .ZN(_05033_)
  );
  INV_X1 _15248_ (
    .A(_05033_),
    .ZN(_05034_)
  );
  AND2_X1 _15249_ (
    .A1(_04830_),
    .A2(_05027_),
    .ZN(_05035_)
  );
  INV_X1 _15250_ (
    .A(_05035_),
    .ZN(_05036_)
  );
  AND2_X1 _15251_ (
    .A1(_05030_),
    .A2(_05032_),
    .ZN(_05037_)
  );
  AND2_X1 _15252_ (
    .A1(_05034_),
    .A2(_05036_),
    .ZN(_05038_)
  );
  AND2_X1 _15253_ (
    .A1(_04899_),
    .A2(_05037_),
    .ZN(_05039_)
  );
  INV_X1 _15254_ (
    .A(_05039_),
    .ZN(_05041_)
  );
  AND2_X1 _15255_ (
    .A1(_04900_),
    .A2(_05038_),
    .ZN(_05042_)
  );
  INV_X1 _15256_ (
    .A(_05042_),
    .ZN(_05043_)
  );
  AND2_X1 _15257_ (
    .A1(_05041_),
    .A2(_05043_),
    .ZN(_05044_)
  );
  INV_X1 _15258_ (
    .A(_05044_),
    .ZN(_05045_)
  );
  AND2_X1 _15259_ (
    .A1(_04836_),
    .A2(_05044_),
    .ZN(_05046_)
  );
  INV_X1 _15260_ (
    .A(_05046_),
    .ZN(_05047_)
  );
  AND2_X1 _15261_ (
    .A1(_04835_),
    .A2(_05045_),
    .ZN(_05048_)
  );
  INV_X1 _15262_ (
    .A(_05048_),
    .ZN(_05049_)
  );
  AND2_X1 _15263_ (
    .A1(_05047_),
    .A2(_05049_),
    .ZN(_05050_)
  );
  INV_X1 _15264_ (
    .A(_05050_),
    .ZN(_05052_)
  );
  AND2_X1 _15265_ (
    .A1(_04616_),
    .A2(_05050_),
    .ZN(_05053_)
  );
  INV_X1 _15266_ (
    .A(_05053_),
    .ZN(_05054_)
  );
  AND2_X1 _15267_ (
    .A1(_04617_),
    .A2(_05052_),
    .ZN(_05055_)
  );
  INV_X1 _15268_ (
    .A(_05055_),
    .ZN(_05056_)
  );
  AND2_X1 _15269_ (
    .A1(_05054_),
    .A2(_05056_),
    .ZN(_05057_)
  );
  INV_X1 _15270_ (
    .A(_05057_),
    .ZN(_05058_)
  );
  AND2_X1 _15271_ (
    .A1(_04829_),
    .A2(_05057_),
    .ZN(_05059_)
  );
  INV_X1 _15272_ (
    .A(_05059_),
    .ZN(_05060_)
  );
  AND2_X1 _15273_ (
    .A1(_04828_),
    .A2(_05058_),
    .ZN(_05061_)
  );
  INV_X1 _15274_ (
    .A(_05061_),
    .ZN(_05063_)
  );
  AND2_X1 _15275_ (
    .A1(_05060_),
    .A2(_05063_),
    .ZN(_05064_)
  );
  INV_X1 _15276_ (
    .A(_05064_),
    .ZN(_05065_)
  );
  AND2_X1 _15277_ (
    .A1(_04769_),
    .A2(_05064_),
    .ZN(_05066_)
  );
  INV_X1 _15278_ (
    .A(_05066_),
    .ZN(_05067_)
  );
  AND2_X1 _15279_ (
    .A1(_04770_),
    .A2(_05065_),
    .ZN(_05068_)
  );
  INV_X1 _15280_ (
    .A(_05068_),
    .ZN(_05069_)
  );
  AND2_X1 _15281_ (
    .A1(_05067_),
    .A2(_05069_),
    .ZN(_05070_)
  );
  INV_X1 _15282_ (
    .A(_05070_),
    .ZN(_05071_)
  );
  AND2_X1 _15283_ (
    .A1(_04827_),
    .A2(_05070_),
    .ZN(_05072_)
  );
  INV_X1 _15284_ (
    .A(_05072_),
    .ZN(_05074_)
  );
  AND2_X1 _15285_ (
    .A1(_04826_),
    .A2(_05071_),
    .ZN(_05075_)
  );
  INV_X1 _15286_ (
    .A(_05075_),
    .ZN(_05076_)
  );
  AND2_X1 _15287_ (
    .A1(_05074_),
    .A2(_05076_),
    .ZN(_05077_)
  );
  INV_X1 _15288_ (
    .A(_05077_),
    .ZN(_05078_)
  );
  AND2_X1 _15289_ (
    .A1(remainder[51]),
    .A2(_05077_),
    .ZN(_05079_)
  );
  INV_X1 _15290_ (
    .A(_05079_),
    .ZN(_05080_)
  );
  AND2_X1 _15291_ (
    .A1(_04557_),
    .A2(_05078_),
    .ZN(_05081_)
  );
  INV_X1 _15292_ (
    .A(_05081_),
    .ZN(_05082_)
  );
  AND2_X1 _15293_ (
    .A1(_05080_),
    .A2(_05082_),
    .ZN(_05083_)
  );
  INV_X1 _15294_ (
    .A(_05083_),
    .ZN(_05085_)
  );
  AND2_X1 _15295_ (
    .A1(_04552_),
    .A2(_04794_),
    .ZN(_05086_)
  );
  INV_X1 _15296_ (
    .A(_05086_),
    .ZN(_05087_)
  );
  AND2_X1 _15297_ (
    .A1(_04553_),
    .A2(_04796_),
    .ZN(_05088_)
  );
  INV_X1 _15298_ (
    .A(_05088_),
    .ZN(_05089_)
  );
  AND2_X1 _15299_ (
    .A1(_04796_),
    .A2(_05087_),
    .ZN(_05090_)
  );
  AND2_X1 _15300_ (
    .A1(_04794_),
    .A2(_05089_),
    .ZN(_05091_)
  );
  AND2_X1 _15301_ (
    .A1(_05083_),
    .A2(_05090_),
    .ZN(_05092_)
  );
  INV_X1 _15302_ (
    .A(_05092_),
    .ZN(_05093_)
  );
  AND2_X1 _15303_ (
    .A1(_05085_),
    .A2(_05091_),
    .ZN(_05094_)
  );
  INV_X1 _15304_ (
    .A(_05094_),
    .ZN(_05096_)
  );
  AND2_X1 _15305_ (
    .A1(_02082_),
    .A2(_05093_),
    .ZN(_05097_)
  );
  AND2_X1 _15306_ (
    .A1(_05096_),
    .A2(_05097_),
    .ZN(_05098_)
  );
  INV_X1 _15307_ (
    .A(_05098_),
    .ZN(_05099_)
  );
  AND2_X1 _15308_ (
    .A1(_04819_),
    .A2(_05099_),
    .ZN(_05100_)
  );
  AND2_X1 _15309_ (
    .A1(_04817_),
    .A2(_05100_),
    .ZN(_05101_)
  );
  INV_X1 _15310_ (
    .A(_05101_),
    .ZN(_05102_)
  );
  AND2_X1 _15311_ (
    .A1(_06201_),
    .A2(_05102_),
    .ZN(_00064_)
  );
  AND2_X1 _15312_ (
    .A1(_10462_),
    .A2(_01770_),
    .ZN(_05103_)
  );
  INV_X1 _15313_ (
    .A(_05103_),
    .ZN(_05104_)
  );
  AND2_X1 _15314_ (
    .A1(_04645_),
    .A2(_10451_),
    .ZN(_05106_)
  );
  INV_X1 _15315_ (
    .A(_05106_),
    .ZN(_05107_)
  );
  AND2_X1 _15316_ (
    .A1(_05983_),
    .A2(_05104_),
    .ZN(_05108_)
  );
  AND2_X1 _15317_ (
    .A1(_05107_),
    .A2(_05108_),
    .ZN(_05109_)
  );
  INV_X1 _15318_ (
    .A(_05109_),
    .ZN(_05110_)
  );
  AND2_X1 _15319_ (
    .A1(remainder[44]),
    .A2(_02077_),
    .ZN(_05111_)
  );
  INV_X1 _15320_ (
    .A(_05111_),
    .ZN(_05112_)
  );
  AND2_X1 _15321_ (
    .A1(_05080_),
    .A2(_05093_),
    .ZN(_05113_)
  );
  INV_X1 _15322_ (
    .A(_05113_),
    .ZN(_05114_)
  );
  AND2_X1 _15323_ (
    .A1(_05067_),
    .A2(_05074_),
    .ZN(_05115_)
  );
  INV_X1 _15324_ (
    .A(_05115_),
    .ZN(_05117_)
  );
  AND2_X1 _15325_ (
    .A1(_05047_),
    .A2(_05054_),
    .ZN(_05118_)
  );
  INV_X1 _15326_ (
    .A(_05118_),
    .ZN(_05119_)
  );
  AND2_X1 _15327_ (
    .A1(_04889_),
    .A2(_04895_),
    .ZN(_05120_)
  );
  INV_X1 _15328_ (
    .A(_05120_),
    .ZN(_05121_)
  );
  AND2_X1 _15329_ (
    .A1(_03249_),
    .A2(_04740_),
    .ZN(_05122_)
  );
  AND2_X1 _15330_ (
    .A1(_05027_),
    .A2(_05122_),
    .ZN(_05123_)
  );
  INV_X1 _15331_ (
    .A(_05123_),
    .ZN(_05124_)
  );
  AND2_X1 _15332_ (
    .A1(_05041_),
    .A2(_05124_),
    .ZN(_05125_)
  );
  INV_X1 _15333_ (
    .A(_05125_),
    .ZN(_05126_)
  );
  AND2_X1 _15334_ (
    .A1(_03249_),
    .A2(_05026_),
    .ZN(_05128_)
  );
  INV_X1 _15335_ (
    .A(_05128_),
    .ZN(_05129_)
  );
  AND2_X1 _15336_ (
    .A1(_04909_),
    .A2(_04915_),
    .ZN(_05130_)
  );
  INV_X1 _15337_ (
    .A(_05130_),
    .ZN(_05131_)
  );
  AND2_X1 _15338_ (
    .A1(divisor[16]),
    .A2(remainder[3]),
    .ZN(_05132_)
  );
  INV_X1 _15339_ (
    .A(_05132_),
    .ZN(_05133_)
  );
  AND2_X1 _15340_ (
    .A1(divisor[17]),
    .A2(remainder[2]),
    .ZN(_05134_)
  );
  INV_X1 _15341_ (
    .A(_05134_),
    .ZN(_05135_)
  );
  AND2_X1 _15342_ (
    .A1(divisor[18]),
    .A2(remainder[2]),
    .ZN(_05136_)
  );
  INV_X1 _15343_ (
    .A(_05136_),
    .ZN(_05137_)
  );
  AND2_X1 _15344_ (
    .A1(_04627_),
    .A2(_05136_),
    .ZN(_05139_)
  );
  INV_X1 _15345_ (
    .A(_05139_),
    .ZN(_05140_)
  );
  AND2_X1 _15346_ (
    .A1(_04906_),
    .A2(_05135_),
    .ZN(_05141_)
  );
  INV_X1 _15347_ (
    .A(_05141_),
    .ZN(_05142_)
  );
  AND2_X1 _15348_ (
    .A1(_05140_),
    .A2(_05142_),
    .ZN(_05143_)
  );
  INV_X1 _15349_ (
    .A(_05143_),
    .ZN(_05144_)
  );
  AND2_X1 _15350_ (
    .A1(_05132_),
    .A2(_05143_),
    .ZN(_05145_)
  );
  INV_X1 _15351_ (
    .A(_05145_),
    .ZN(_05146_)
  );
  AND2_X1 _15352_ (
    .A1(_05133_),
    .A2(_05144_),
    .ZN(_05147_)
  );
  INV_X1 _15353_ (
    .A(_05147_),
    .ZN(_05148_)
  );
  AND2_X1 _15354_ (
    .A1(_05146_),
    .A2(_05148_),
    .ZN(_05150_)
  );
  INV_X1 _15355_ (
    .A(_05150_),
    .ZN(_05151_)
  );
  AND2_X1 _15356_ (
    .A1(_05131_),
    .A2(_05150_),
    .ZN(_05152_)
  );
  INV_X1 _15357_ (
    .A(_05152_),
    .ZN(_05153_)
  );
  AND2_X1 _15358_ (
    .A1(_05130_),
    .A2(_05151_),
    .ZN(_05154_)
  );
  INV_X1 _15359_ (
    .A(_05154_),
    .ZN(_05155_)
  );
  AND2_X1 _15360_ (
    .A1(_05153_),
    .A2(_05155_),
    .ZN(_05156_)
  );
  INV_X1 _15361_ (
    .A(_05156_),
    .ZN(_05157_)
  );
  AND2_X1 _15362_ (
    .A1(_04921_),
    .A2(_05156_),
    .ZN(_05158_)
  );
  INV_X1 _15363_ (
    .A(_05158_),
    .ZN(_05159_)
  );
  AND2_X1 _15364_ (
    .A1(_04922_),
    .A2(_05157_),
    .ZN(_05161_)
  );
  INV_X1 _15365_ (
    .A(_05161_),
    .ZN(_05162_)
  );
  AND2_X1 _15366_ (
    .A1(_05159_),
    .A2(_05162_),
    .ZN(_05163_)
  );
  INV_X1 _15367_ (
    .A(_05163_),
    .ZN(_05164_)
  );
  AND2_X1 _15368_ (
    .A1(_04953_),
    .A2(_04979_),
    .ZN(_05165_)
  );
  INV_X1 _15369_ (
    .A(_05165_),
    .ZN(_05166_)
  );
  AND2_X1 _15370_ (
    .A1(_04939_),
    .A2(_04946_),
    .ZN(_05167_)
  );
  INV_X1 _15371_ (
    .A(_05167_),
    .ZN(_05168_)
  );
  AND2_X1 _15372_ (
    .A1(divisor[13]),
    .A2(remainder[6]),
    .ZN(_05169_)
  );
  INV_X1 _15373_ (
    .A(_05169_),
    .ZN(_05170_)
  );
  AND2_X1 _15374_ (
    .A1(divisor[14]),
    .A2(remainder[5]),
    .ZN(_05172_)
  );
  INV_X1 _15375_ (
    .A(_05172_),
    .ZN(_05173_)
  );
  AND2_X1 _15376_ (
    .A1(divisor[15]),
    .A2(remainder[5]),
    .ZN(_05174_)
  );
  INV_X1 _15377_ (
    .A(_05174_),
    .ZN(_05175_)
  );
  AND2_X1 _15378_ (
    .A1(_04936_),
    .A2(_05172_),
    .ZN(_05176_)
  );
  INV_X1 _15379_ (
    .A(_05176_),
    .ZN(_05177_)
  );
  AND2_X1 _15380_ (
    .A1(_04937_),
    .A2(_05173_),
    .ZN(_05178_)
  );
  INV_X1 _15381_ (
    .A(_05178_),
    .ZN(_05179_)
  );
  AND2_X1 _15382_ (
    .A1(_05177_),
    .A2(_05179_),
    .ZN(_05180_)
  );
  INV_X1 _15383_ (
    .A(_05180_),
    .ZN(_05181_)
  );
  AND2_X1 _15384_ (
    .A1(_05169_),
    .A2(_05180_),
    .ZN(_05183_)
  );
  INV_X1 _15385_ (
    .A(_05183_),
    .ZN(_05184_)
  );
  AND2_X1 _15386_ (
    .A1(_05170_),
    .A2(_05181_),
    .ZN(_05185_)
  );
  INV_X1 _15387_ (
    .A(_05185_),
    .ZN(_05186_)
  );
  AND2_X1 _15388_ (
    .A1(_05184_),
    .A2(_05186_),
    .ZN(_05187_)
  );
  INV_X1 _15389_ (
    .A(_05187_),
    .ZN(_05188_)
  );
  AND2_X1 _15390_ (
    .A1(_05168_),
    .A2(_05187_),
    .ZN(_05189_)
  );
  INV_X1 _15391_ (
    .A(_05189_),
    .ZN(_05190_)
  );
  AND2_X1 _15392_ (
    .A1(_05167_),
    .A2(_05188_),
    .ZN(_05191_)
  );
  INV_X1 _15393_ (
    .A(_05191_),
    .ZN(_05192_)
  );
  AND2_X1 _15394_ (
    .A1(_05190_),
    .A2(_05192_),
    .ZN(_05194_)
  );
  INV_X1 _15395_ (
    .A(_05194_),
    .ZN(_05195_)
  );
  AND2_X1 _15396_ (
    .A1(remainder[32]),
    .A2(divisor[12]),
    .ZN(_05196_)
  );
  AND2_X1 _15397_ (
    .A1(remainder[32]),
    .A2(divisor[11]),
    .ZN(_05197_)
  );
  INV_X1 _15398_ (
    .A(_05197_),
    .ZN(_05198_)
  );
  AND2_X1 _15399_ (
    .A1(divisor[12]),
    .A2(_05197_),
    .ZN(_05199_)
  );
  INV_X1 _15400_ (
    .A(_05199_),
    .ZN(_05200_)
  );
  AND2_X1 _15401_ (
    .A1(_04962_),
    .A2(_05197_),
    .ZN(_05201_)
  );
  INV_X1 _15402_ (
    .A(_05201_),
    .ZN(_05202_)
  );
  AND2_X1 _15403_ (
    .A1(_04964_),
    .A2(_05198_),
    .ZN(_05203_)
  );
  INV_X1 _15404_ (
    .A(_05203_),
    .ZN(_05205_)
  );
  AND2_X1 _15405_ (
    .A1(_05202_),
    .A2(_05205_),
    .ZN(_05206_)
  );
  INV_X1 _15406_ (
    .A(_05206_),
    .ZN(_05207_)
  );
  AND2_X1 _15407_ (
    .A1(_04958_),
    .A2(_05206_),
    .ZN(_05208_)
  );
  INV_X1 _15408_ (
    .A(_05208_),
    .ZN(_05209_)
  );
  AND2_X1 _15409_ (
    .A1(_04959_),
    .A2(_05207_),
    .ZN(_05210_)
  );
  INV_X1 _15410_ (
    .A(_05210_),
    .ZN(_05211_)
  );
  AND2_X1 _15411_ (
    .A1(_05209_),
    .A2(_05211_),
    .ZN(_05212_)
  );
  INV_X1 _15412_ (
    .A(_05212_),
    .ZN(_05213_)
  );
  AND2_X1 _15413_ (
    .A1(_05194_),
    .A2(_05212_),
    .ZN(_05214_)
  );
  INV_X1 _15414_ (
    .A(_05214_),
    .ZN(_05216_)
  );
  AND2_X1 _15415_ (
    .A1(_05195_),
    .A2(_05213_),
    .ZN(_05217_)
  );
  INV_X1 _15416_ (
    .A(_05217_),
    .ZN(_05218_)
  );
  AND2_X1 _15417_ (
    .A1(_05216_),
    .A2(_05218_),
    .ZN(_05219_)
  );
  INV_X1 _15418_ (
    .A(_05219_),
    .ZN(_05220_)
  );
  AND2_X1 _15419_ (
    .A1(_05166_),
    .A2(_05219_),
    .ZN(_05221_)
  );
  INV_X1 _15420_ (
    .A(_05221_),
    .ZN(_05222_)
  );
  AND2_X1 _15421_ (
    .A1(_05165_),
    .A2(_05220_),
    .ZN(_05223_)
  );
  INV_X1 _15422_ (
    .A(_05223_),
    .ZN(_05224_)
  );
  AND2_X1 _15423_ (
    .A1(_05222_),
    .A2(_05224_),
    .ZN(_05225_)
  );
  INV_X1 _15424_ (
    .A(_05225_),
    .ZN(_05227_)
  );
  AND2_X1 _15425_ (
    .A1(_04966_),
    .A2(_04972_),
    .ZN(_05228_)
  );
  INV_X1 _15426_ (
    .A(_05228_),
    .ZN(_05229_)
  );
  AND2_X1 _15427_ (
    .A1(_04707_),
    .A2(_05229_),
    .ZN(_05230_)
  );
  INV_X1 _15428_ (
    .A(_05230_),
    .ZN(_05231_)
  );
  AND2_X1 _15429_ (
    .A1(_04708_),
    .A2(_05228_),
    .ZN(_05232_)
  );
  INV_X1 _15430_ (
    .A(_05232_),
    .ZN(_05233_)
  );
  AND2_X1 _15431_ (
    .A1(_05231_),
    .A2(_05233_),
    .ZN(_05234_)
  );
  INV_X1 _15432_ (
    .A(_05234_),
    .ZN(_05235_)
  );
  AND2_X1 _15433_ (
    .A1(_04992_),
    .A2(_05234_),
    .ZN(_05236_)
  );
  INV_X1 _15434_ (
    .A(_05236_),
    .ZN(_05238_)
  );
  AND2_X1 _15435_ (
    .A1(_04991_),
    .A2(_05235_),
    .ZN(_05239_)
  );
  INV_X1 _15436_ (
    .A(_05239_),
    .ZN(_05240_)
  );
  AND2_X1 _15437_ (
    .A1(_05238_),
    .A2(_05240_),
    .ZN(_05241_)
  );
  INV_X1 _15438_ (
    .A(_05241_),
    .ZN(_05242_)
  );
  AND2_X1 _15439_ (
    .A1(_05225_),
    .A2(_05241_),
    .ZN(_05243_)
  );
  INV_X1 _15440_ (
    .A(_05243_),
    .ZN(_05244_)
  );
  AND2_X1 _15441_ (
    .A1(_05227_),
    .A2(_05242_),
    .ZN(_05245_)
  );
  INV_X1 _15442_ (
    .A(_05245_),
    .ZN(_05246_)
  );
  AND2_X1 _15443_ (
    .A1(_05244_),
    .A2(_05246_),
    .ZN(_05247_)
  );
  INV_X1 _15444_ (
    .A(_05247_),
    .ZN(_05249_)
  );
  AND2_X1 _15445_ (
    .A1(_05163_),
    .A2(_05247_),
    .ZN(_05250_)
  );
  INV_X1 _15446_ (
    .A(_05250_),
    .ZN(_05251_)
  );
  AND2_X1 _15447_ (
    .A1(_05164_),
    .A2(_05249_),
    .ZN(_05252_)
  );
  INV_X1 _15448_ (
    .A(_05252_),
    .ZN(_05253_)
  );
  AND2_X1 _15449_ (
    .A1(_05251_),
    .A2(_05253_),
    .ZN(_05254_)
  );
  INV_X1 _15450_ (
    .A(_05254_),
    .ZN(_05255_)
  );
  AND2_X1 _15451_ (
    .A1(_05015_),
    .A2(_05254_),
    .ZN(_05256_)
  );
  INV_X1 _15452_ (
    .A(_05256_),
    .ZN(_05257_)
  );
  AND2_X1 _15453_ (
    .A1(_05016_),
    .A2(_05255_),
    .ZN(_05258_)
  );
  INV_X1 _15454_ (
    .A(_05258_),
    .ZN(_05260_)
  );
  AND2_X1 _15455_ (
    .A1(_05257_),
    .A2(_05260_),
    .ZN(_05261_)
  );
  INV_X1 _15456_ (
    .A(_05261_),
    .ZN(_05262_)
  );
  AND2_X1 _15457_ (
    .A1(divisor[19]),
    .A2(remainder[0]),
    .ZN(_05263_)
  );
  INV_X1 _15458_ (
    .A(_05263_),
    .ZN(_05264_)
  );
  AND2_X1 _15459_ (
    .A1(_03249_),
    .A2(_05264_),
    .ZN(_05265_)
  );
  INV_X1 _15460_ (
    .A(_05265_),
    .ZN(_05266_)
  );
  AND2_X1 _15461_ (
    .A1(_03250_),
    .A2(_05263_),
    .ZN(_05267_)
  );
  INV_X1 _15462_ (
    .A(_05267_),
    .ZN(_05268_)
  );
  AND2_X1 _15463_ (
    .A1(remainder[32]),
    .A2(divisor[19]),
    .ZN(_05269_)
  );
  INV_X1 _15464_ (
    .A(_05269_),
    .ZN(_05271_)
  );
  AND2_X1 _15465_ (
    .A1(_05266_),
    .A2(_05268_),
    .ZN(_05272_)
  );
  INV_X1 _15466_ (
    .A(_05272_),
    .ZN(_05273_)
  );
  AND2_X1 _15467_ (
    .A1(_05261_),
    .A2(_05273_),
    .ZN(_05274_)
  );
  INV_X1 _15468_ (
    .A(_05274_),
    .ZN(_05275_)
  );
  AND2_X1 _15469_ (
    .A1(_05262_),
    .A2(_05272_),
    .ZN(_05276_)
  );
  INV_X1 _15470_ (
    .A(_05276_),
    .ZN(_05277_)
  );
  AND2_X1 _15471_ (
    .A1(_05275_),
    .A2(_05277_),
    .ZN(_05278_)
  );
  INV_X1 _15472_ (
    .A(_05278_),
    .ZN(_05279_)
  );
  AND2_X1 _15473_ (
    .A1(_05128_),
    .A2(_05278_),
    .ZN(_05280_)
  );
  INV_X1 _15474_ (
    .A(_05280_),
    .ZN(_05282_)
  );
  AND2_X1 _15475_ (
    .A1(_05129_),
    .A2(_05279_),
    .ZN(_05283_)
  );
  INV_X1 _15476_ (
    .A(_05283_),
    .ZN(_05284_)
  );
  AND2_X1 _15477_ (
    .A1(_05282_),
    .A2(_05284_),
    .ZN(_05285_)
  );
  INV_X1 _15478_ (
    .A(_05285_),
    .ZN(_05286_)
  );
  AND2_X1 _15479_ (
    .A1(_04876_),
    .A2(_04882_),
    .ZN(_05287_)
  );
  INV_X1 _15480_ (
    .A(_05287_),
    .ZN(_05288_)
  );
  AND2_X1 _15481_ (
    .A1(_04862_),
    .A2(_04869_),
    .ZN(_05289_)
  );
  INV_X1 _15482_ (
    .A(_05289_),
    .ZN(_05290_)
  );
  AND2_X1 _15483_ (
    .A1(_04849_),
    .A2(_04856_),
    .ZN(_05291_)
  );
  INV_X1 _15484_ (
    .A(_05291_),
    .ZN(_05293_)
  );
  AND2_X1 _15485_ (
    .A1(_04986_),
    .A2(_05010_),
    .ZN(_05294_)
  );
  INV_X1 _15486_ (
    .A(_05294_),
    .ZN(_05295_)
  );
  AND2_X1 _15487_ (
    .A1(_04997_),
    .A2(_05003_),
    .ZN(_05296_)
  );
  INV_X1 _15488_ (
    .A(_05296_),
    .ZN(_05297_)
  );
  AND2_X1 _15489_ (
    .A1(_04087_),
    .A2(_05297_),
    .ZN(_05298_)
  );
  INV_X1 _15490_ (
    .A(_05298_),
    .ZN(_05299_)
  );
  AND2_X1 _15491_ (
    .A1(_04088_),
    .A2(_05296_),
    .ZN(_05300_)
  );
  INV_X1 _15492_ (
    .A(_05300_),
    .ZN(_05301_)
  );
  AND2_X1 _15493_ (
    .A1(_05299_),
    .A2(_05301_),
    .ZN(_05302_)
  );
  INV_X1 _15494_ (
    .A(_05302_),
    .ZN(_05304_)
  );
  AND2_X1 _15495_ (
    .A1(_04317_),
    .A2(_05302_),
    .ZN(_05305_)
  );
  INV_X1 _15496_ (
    .A(_05305_),
    .ZN(_05306_)
  );
  AND2_X1 _15497_ (
    .A1(_04316_),
    .A2(_05304_),
    .ZN(_05307_)
  );
  INV_X1 _15498_ (
    .A(_05307_),
    .ZN(_05308_)
  );
  AND2_X1 _15499_ (
    .A1(_05306_),
    .A2(_05308_),
    .ZN(_05309_)
  );
  INV_X1 _15500_ (
    .A(_05309_),
    .ZN(_05310_)
  );
  AND2_X1 _15501_ (
    .A1(_05295_),
    .A2(_05309_),
    .ZN(_05311_)
  );
  INV_X1 _15502_ (
    .A(_05311_),
    .ZN(_05312_)
  );
  AND2_X1 _15503_ (
    .A1(_05294_),
    .A2(_05310_),
    .ZN(_05313_)
  );
  INV_X1 _15504_ (
    .A(_05313_),
    .ZN(_05315_)
  );
  AND2_X1 _15505_ (
    .A1(_05312_),
    .A2(_05315_),
    .ZN(_05316_)
  );
  INV_X1 _15506_ (
    .A(_05316_),
    .ZN(_05317_)
  );
  AND2_X1 _15507_ (
    .A1(_05293_),
    .A2(_05316_),
    .ZN(_05318_)
  );
  INV_X1 _15508_ (
    .A(_05318_),
    .ZN(_05319_)
  );
  AND2_X1 _15509_ (
    .A1(_05291_),
    .A2(_05317_),
    .ZN(_05320_)
  );
  INV_X1 _15510_ (
    .A(_05320_),
    .ZN(_05321_)
  );
  AND2_X1 _15511_ (
    .A1(_05319_),
    .A2(_05321_),
    .ZN(_05322_)
  );
  INV_X1 _15512_ (
    .A(_05322_),
    .ZN(_05323_)
  );
  AND2_X1 _15513_ (
    .A1(_05290_),
    .A2(_05322_),
    .ZN(_05324_)
  );
  INV_X1 _15514_ (
    .A(_05324_),
    .ZN(_05326_)
  );
  AND2_X1 _15515_ (
    .A1(_05289_),
    .A2(_05323_),
    .ZN(_05327_)
  );
  INV_X1 _15516_ (
    .A(_05327_),
    .ZN(_05328_)
  );
  AND2_X1 _15517_ (
    .A1(_05326_),
    .A2(_05328_),
    .ZN(_05329_)
  );
  INV_X1 _15518_ (
    .A(_05329_),
    .ZN(_05330_)
  );
  AND2_X1 _15519_ (
    .A1(_03170_),
    .A2(_05329_),
    .ZN(_05331_)
  );
  INV_X1 _15520_ (
    .A(_05331_),
    .ZN(_05332_)
  );
  AND2_X1 _15521_ (
    .A1(_03169_),
    .A2(_05330_),
    .ZN(_05333_)
  );
  INV_X1 _15522_ (
    .A(_05333_),
    .ZN(_05334_)
  );
  AND2_X1 _15523_ (
    .A1(_05332_),
    .A2(_05334_),
    .ZN(_05335_)
  );
  INV_X1 _15524_ (
    .A(_05335_),
    .ZN(_05337_)
  );
  AND2_X1 _15525_ (
    .A1(_05022_),
    .A2(_05335_),
    .ZN(_05338_)
  );
  INV_X1 _15526_ (
    .A(_05338_),
    .ZN(_05339_)
  );
  AND2_X1 _15527_ (
    .A1(_05023_),
    .A2(_05337_),
    .ZN(_05340_)
  );
  INV_X1 _15528_ (
    .A(_05340_),
    .ZN(_05341_)
  );
  AND2_X1 _15529_ (
    .A1(_05339_),
    .A2(_05341_),
    .ZN(_05342_)
  );
  INV_X1 _15530_ (
    .A(_05342_),
    .ZN(_05343_)
  );
  AND2_X1 _15531_ (
    .A1(_05288_),
    .A2(_05342_),
    .ZN(_05344_)
  );
  INV_X1 _15532_ (
    .A(_05344_),
    .ZN(_05345_)
  );
  AND2_X1 _15533_ (
    .A1(_05287_),
    .A2(_05343_),
    .ZN(_05346_)
  );
  INV_X1 _15534_ (
    .A(_05346_),
    .ZN(_05348_)
  );
  AND2_X1 _15535_ (
    .A1(_05345_),
    .A2(_05348_),
    .ZN(_05349_)
  );
  INV_X1 _15536_ (
    .A(_05349_),
    .ZN(_05350_)
  );
  AND2_X1 _15537_ (
    .A1(_05285_),
    .A2(_05349_),
    .ZN(_05351_)
  );
  INV_X1 _15538_ (
    .A(_05351_),
    .ZN(_05352_)
  );
  AND2_X1 _15539_ (
    .A1(_05286_),
    .A2(_05350_),
    .ZN(_05353_)
  );
  INV_X1 _15540_ (
    .A(_05353_),
    .ZN(_05354_)
  );
  AND2_X1 _15541_ (
    .A1(_05352_),
    .A2(_05354_),
    .ZN(_05355_)
  );
  INV_X1 _15542_ (
    .A(_05355_),
    .ZN(_05356_)
  );
  AND2_X1 _15543_ (
    .A1(_05126_),
    .A2(_05355_),
    .ZN(_05357_)
  );
  INV_X1 _15544_ (
    .A(_05357_),
    .ZN(_05359_)
  );
  AND2_X1 _15545_ (
    .A1(_05125_),
    .A2(_05356_),
    .ZN(_05360_)
  );
  INV_X1 _15546_ (
    .A(_05360_),
    .ZN(_05361_)
  );
  AND2_X1 _15547_ (
    .A1(_05359_),
    .A2(_05361_),
    .ZN(_05362_)
  );
  INV_X1 _15548_ (
    .A(_05362_),
    .ZN(_05363_)
  );
  AND2_X1 _15549_ (
    .A1(_05121_),
    .A2(_05362_),
    .ZN(_05364_)
  );
  INV_X1 _15550_ (
    .A(_05364_),
    .ZN(_05365_)
  );
  AND2_X1 _15551_ (
    .A1(_05120_),
    .A2(_05363_),
    .ZN(_05366_)
  );
  INV_X1 _15552_ (
    .A(_05366_),
    .ZN(_05367_)
  );
  AND2_X1 _15553_ (
    .A1(_05365_),
    .A2(_05367_),
    .ZN(_05368_)
  );
  INV_X1 _15554_ (
    .A(_05368_),
    .ZN(_05370_)
  );
  AND2_X1 _15555_ (
    .A1(_05119_),
    .A2(_05368_),
    .ZN(_05371_)
  );
  INV_X1 _15556_ (
    .A(_05371_),
    .ZN(_05372_)
  );
  AND2_X1 _15557_ (
    .A1(_05118_),
    .A2(_05370_),
    .ZN(_05373_)
  );
  INV_X1 _15558_ (
    .A(_05373_),
    .ZN(_05374_)
  );
  AND2_X1 _15559_ (
    .A1(_05372_),
    .A2(_05374_),
    .ZN(_05375_)
  );
  INV_X1 _15560_ (
    .A(_05375_),
    .ZN(_05376_)
  );
  AND2_X1 _15561_ (
    .A1(_05059_),
    .A2(_05375_),
    .ZN(_05377_)
  );
  INV_X1 _15562_ (
    .A(_05377_),
    .ZN(_05378_)
  );
  AND2_X1 _15563_ (
    .A1(_05060_),
    .A2(_05376_),
    .ZN(_05379_)
  );
  INV_X1 _15564_ (
    .A(_05379_),
    .ZN(_05381_)
  );
  AND2_X1 _15565_ (
    .A1(_05378_),
    .A2(_05381_),
    .ZN(_05382_)
  );
  INV_X1 _15566_ (
    .A(_05382_),
    .ZN(_05383_)
  );
  AND2_X1 _15567_ (
    .A1(_05115_),
    .A2(_05382_),
    .ZN(_05384_)
  );
  INV_X1 _15568_ (
    .A(_05384_),
    .ZN(_05385_)
  );
  AND2_X1 _15569_ (
    .A1(_05117_),
    .A2(_05383_),
    .ZN(_05386_)
  );
  INV_X1 _15570_ (
    .A(_05386_),
    .ZN(_05387_)
  );
  AND2_X1 _15571_ (
    .A1(_05117_),
    .A2(_05382_),
    .ZN(_05388_)
  );
  INV_X1 _15572_ (
    .A(_05388_),
    .ZN(_05389_)
  );
  AND2_X1 _15573_ (
    .A1(_05115_),
    .A2(_05383_),
    .ZN(_05390_)
  );
  INV_X1 _15574_ (
    .A(_05390_),
    .ZN(_05392_)
  );
  AND2_X1 _15575_ (
    .A1(_05385_),
    .A2(_05387_),
    .ZN(_05393_)
  );
  AND2_X1 _15576_ (
    .A1(_05389_),
    .A2(_05392_),
    .ZN(_05394_)
  );
  AND2_X1 _15577_ (
    .A1(remainder[52]),
    .A2(_05394_),
    .ZN(_05395_)
  );
  INV_X1 _15578_ (
    .A(_05395_),
    .ZN(_05396_)
  );
  AND2_X1 _15579_ (
    .A1(_04546_),
    .A2(_05393_),
    .ZN(_05397_)
  );
  INV_X1 _15580_ (
    .A(_05397_),
    .ZN(_05398_)
  );
  AND2_X1 _15581_ (
    .A1(_05396_),
    .A2(_05398_),
    .ZN(_05399_)
  );
  INV_X1 _15582_ (
    .A(_05399_),
    .ZN(_05400_)
  );
  AND2_X1 _15583_ (
    .A1(_05113_),
    .A2(_05400_),
    .ZN(_05401_)
  );
  INV_X1 _15584_ (
    .A(_05401_),
    .ZN(_05403_)
  );
  AND2_X1 _15585_ (
    .A1(_05114_),
    .A2(_05399_),
    .ZN(_05404_)
  );
  INV_X1 _15586_ (
    .A(_05404_),
    .ZN(_05405_)
  );
  AND2_X1 _15587_ (
    .A1(_05403_),
    .A2(_05405_),
    .ZN(_05406_)
  );
  AND2_X1 _15588_ (
    .A1(_02082_),
    .A2(_05406_),
    .ZN(_05407_)
  );
  INV_X1 _15589_ (
    .A(_05407_),
    .ZN(_05408_)
  );
  AND2_X1 _15590_ (
    .A1(_05112_),
    .A2(_05408_),
    .ZN(_05409_)
  );
  AND2_X1 _15591_ (
    .A1(_05110_),
    .A2(_05409_),
    .ZN(_05410_)
  );
  INV_X1 _15592_ (
    .A(_05410_),
    .ZN(_05411_)
  );
  AND2_X1 _15593_ (
    .A1(_06201_),
    .A2(_05411_),
    .ZN(_00065_)
  );
  AND2_X1 _15594_ (
    .A1(_04634_),
    .A2(_10451_),
    .ZN(_05413_)
  );
  INV_X1 _15595_ (
    .A(_05413_),
    .ZN(_05414_)
  );
  AND2_X1 _15596_ (
    .A1(_10462_),
    .A2(_01783_),
    .ZN(_05415_)
  );
  INV_X1 _15597_ (
    .A(_05415_),
    .ZN(_05416_)
  );
  AND2_X1 _15598_ (
    .A1(_05983_),
    .A2(_05416_),
    .ZN(_05417_)
  );
  AND2_X1 _15599_ (
    .A1(_05414_),
    .A2(_05417_),
    .ZN(_05418_)
  );
  INV_X1 _15600_ (
    .A(_05418_),
    .ZN(_05419_)
  );
  AND2_X1 _15601_ (
    .A1(_05359_),
    .A2(_05365_),
    .ZN(_05420_)
  );
  INV_X1 _15602_ (
    .A(_05420_),
    .ZN(_05421_)
  );
  AND2_X1 _15603_ (
    .A1(_05339_),
    .A2(_05345_),
    .ZN(_05422_)
  );
  INV_X1 _15604_ (
    .A(_05422_),
    .ZN(_05424_)
  );
  AND2_X1 _15605_ (
    .A1(_05282_),
    .A2(_05352_),
    .ZN(_05425_)
  );
  INV_X1 _15606_ (
    .A(_05425_),
    .ZN(_05426_)
  );
  AND2_X1 _15607_ (
    .A1(_05140_),
    .A2(_05146_),
    .ZN(_05427_)
  );
  INV_X1 _15608_ (
    .A(_05427_),
    .ZN(_05428_)
  );
  AND2_X1 _15609_ (
    .A1(divisor[16]),
    .A2(remainder[4]),
    .ZN(_05429_)
  );
  INV_X1 _15610_ (
    .A(_05429_),
    .ZN(_05430_)
  );
  AND2_X1 _15611_ (
    .A1(divisor[17]),
    .A2(remainder[3]),
    .ZN(_05431_)
  );
  INV_X1 _15612_ (
    .A(_05431_),
    .ZN(_05432_)
  );
  AND2_X1 _15613_ (
    .A1(divisor[18]),
    .A2(remainder[3]),
    .ZN(_05433_)
  );
  INV_X1 _15614_ (
    .A(_05433_),
    .ZN(_05435_)
  );
  AND2_X1 _15615_ (
    .A1(_05136_),
    .A2(_05431_),
    .ZN(_05436_)
  );
  INV_X1 _15616_ (
    .A(_05436_),
    .ZN(_05437_)
  );
  AND2_X1 _15617_ (
    .A1(_05137_),
    .A2(_05432_),
    .ZN(_05438_)
  );
  INV_X1 _15618_ (
    .A(_05438_),
    .ZN(_05439_)
  );
  AND2_X1 _15619_ (
    .A1(_05437_),
    .A2(_05439_),
    .ZN(_05440_)
  );
  INV_X1 _15620_ (
    .A(_05440_),
    .ZN(_05441_)
  );
  AND2_X1 _15621_ (
    .A1(_05429_),
    .A2(_05440_),
    .ZN(_05442_)
  );
  INV_X1 _15622_ (
    .A(_05442_),
    .ZN(_05443_)
  );
  AND2_X1 _15623_ (
    .A1(_05430_),
    .A2(_05441_),
    .ZN(_05444_)
  );
  INV_X1 _15624_ (
    .A(_05444_),
    .ZN(_05446_)
  );
  AND2_X1 _15625_ (
    .A1(_05443_),
    .A2(_05446_),
    .ZN(_05447_)
  );
  INV_X1 _15626_ (
    .A(_05447_),
    .ZN(_05448_)
  );
  AND2_X1 _15627_ (
    .A1(_05428_),
    .A2(_05447_),
    .ZN(_05449_)
  );
  INV_X1 _15628_ (
    .A(_05449_),
    .ZN(_05450_)
  );
  AND2_X1 _15629_ (
    .A1(_05427_),
    .A2(_05448_),
    .ZN(_05451_)
  );
  INV_X1 _15630_ (
    .A(_05451_),
    .ZN(_05452_)
  );
  AND2_X1 _15631_ (
    .A1(_05450_),
    .A2(_05452_),
    .ZN(_05453_)
  );
  INV_X1 _15632_ (
    .A(_05453_),
    .ZN(_05454_)
  );
  AND2_X1 _15633_ (
    .A1(_05152_),
    .A2(_05453_),
    .ZN(_05455_)
  );
  INV_X1 _15634_ (
    .A(_05455_),
    .ZN(_05457_)
  );
  AND2_X1 _15635_ (
    .A1(_05158_),
    .A2(_05453_),
    .ZN(_05458_)
  );
  INV_X1 _15636_ (
    .A(_05458_),
    .ZN(_05459_)
  );
  AND2_X1 _15637_ (
    .A1(_05159_),
    .A2(_05454_),
    .ZN(_05460_)
  );
  INV_X1 _15638_ (
    .A(_05460_),
    .ZN(_05461_)
  );
  AND2_X1 _15639_ (
    .A1(_05459_),
    .A2(_05461_),
    .ZN(_05462_)
  );
  MUX2_X1 _15640_ (
    .A(_05454_),
    .B(_05462_),
    .S(_05153_),
    .Z(_05463_)
  );
  INV_X1 _15641_ (
    .A(_05463_),
    .ZN(_05464_)
  );
  AND2_X1 _15642_ (
    .A1(_05190_),
    .A2(_05216_),
    .ZN(_05465_)
  );
  INV_X1 _15643_ (
    .A(_05465_),
    .ZN(_05466_)
  );
  AND2_X1 _15644_ (
    .A1(_05177_),
    .A2(_05184_),
    .ZN(_05468_)
  );
  INV_X1 _15645_ (
    .A(_05468_),
    .ZN(_05469_)
  );
  AND2_X1 _15646_ (
    .A1(divisor[13]),
    .A2(remainder[7]),
    .ZN(_05470_)
  );
  INV_X1 _15647_ (
    .A(_05470_),
    .ZN(_05471_)
  );
  AND2_X1 _15648_ (
    .A1(divisor[14]),
    .A2(remainder[6]),
    .ZN(_05472_)
  );
  INV_X1 _15649_ (
    .A(_05472_),
    .ZN(_05473_)
  );
  AND2_X1 _15650_ (
    .A1(divisor[15]),
    .A2(remainder[6]),
    .ZN(_05474_)
  );
  INV_X1 _15651_ (
    .A(_05474_),
    .ZN(_05475_)
  );
  AND2_X1 _15652_ (
    .A1(_05174_),
    .A2(_05472_),
    .ZN(_05476_)
  );
  INV_X1 _15653_ (
    .A(_05476_),
    .ZN(_05477_)
  );
  AND2_X1 _15654_ (
    .A1(_05175_),
    .A2(_05473_),
    .ZN(_05479_)
  );
  INV_X1 _15655_ (
    .A(_05479_),
    .ZN(_05480_)
  );
  AND2_X1 _15656_ (
    .A1(_05477_),
    .A2(_05480_),
    .ZN(_05481_)
  );
  INV_X1 _15657_ (
    .A(_05481_),
    .ZN(_05482_)
  );
  AND2_X1 _15658_ (
    .A1(_05470_),
    .A2(_05481_),
    .ZN(_05483_)
  );
  INV_X1 _15659_ (
    .A(_05483_),
    .ZN(_05484_)
  );
  AND2_X1 _15660_ (
    .A1(_05471_),
    .A2(_05482_),
    .ZN(_05485_)
  );
  INV_X1 _15661_ (
    .A(_05485_),
    .ZN(_05486_)
  );
  AND2_X1 _15662_ (
    .A1(_05484_),
    .A2(_05486_),
    .ZN(_05487_)
  );
  INV_X1 _15663_ (
    .A(_05487_),
    .ZN(_05488_)
  );
  AND2_X1 _15664_ (
    .A1(_05469_),
    .A2(_05487_),
    .ZN(_05490_)
  );
  INV_X1 _15665_ (
    .A(_05490_),
    .ZN(_05491_)
  );
  AND2_X1 _15666_ (
    .A1(_05468_),
    .A2(_05488_),
    .ZN(_05492_)
  );
  INV_X1 _15667_ (
    .A(_05492_),
    .ZN(_05493_)
  );
  AND2_X1 _15668_ (
    .A1(_05491_),
    .A2(_05493_),
    .ZN(_05494_)
  );
  INV_X1 _15669_ (
    .A(_05494_),
    .ZN(_05495_)
  );
  MUX2_X1 _15670_ (
    .A(_05197_),
    .B(_04930_),
    .S(_05196_),
    .Z(_05496_)
  );
  AND2_X1 _15671_ (
    .A1(divisor[10]),
    .A2(_05496_),
    .ZN(_05497_)
  );
  INV_X1 _15672_ (
    .A(_05497_),
    .ZN(_05498_)
  );
  MUX2_X1 _15673_ (
    .A(_04958_),
    .B(_04919_),
    .S(_05496_),
    .Z(_05499_)
  );
  MUX2_X1 _15674_ (
    .A(_04959_),
    .B(divisor[10]),
    .S(_05496_),
    .Z(_05501_)
  );
  AND2_X1 _15675_ (
    .A1(_05494_),
    .A2(_05499_),
    .ZN(_05502_)
  );
  INV_X1 _15676_ (
    .A(_05502_),
    .ZN(_05503_)
  );
  AND2_X1 _15677_ (
    .A1(_05495_),
    .A2(_05501_),
    .ZN(_05504_)
  );
  INV_X1 _15678_ (
    .A(_05504_),
    .ZN(_05505_)
  );
  AND2_X1 _15679_ (
    .A1(_05503_),
    .A2(_05505_),
    .ZN(_05506_)
  );
  INV_X1 _15680_ (
    .A(_05506_),
    .ZN(_05507_)
  );
  AND2_X1 _15681_ (
    .A1(_05466_),
    .A2(_05506_),
    .ZN(_05508_)
  );
  INV_X1 _15682_ (
    .A(_05508_),
    .ZN(_05509_)
  );
  AND2_X1 _15683_ (
    .A1(_05465_),
    .A2(_05507_),
    .ZN(_05510_)
  );
  INV_X1 _15684_ (
    .A(_05510_),
    .ZN(_05512_)
  );
  AND2_X1 _15685_ (
    .A1(_05509_),
    .A2(_05512_),
    .ZN(_05513_)
  );
  INV_X1 _15686_ (
    .A(_05513_),
    .ZN(_05514_)
  );
  AND2_X1 _15687_ (
    .A1(_05202_),
    .A2(_05209_),
    .ZN(_05515_)
  );
  INV_X1 _15688_ (
    .A(_05515_),
    .ZN(_05516_)
  );
  AND2_X1 _15689_ (
    .A1(_04707_),
    .A2(_05516_),
    .ZN(_05517_)
  );
  INV_X1 _15690_ (
    .A(_05517_),
    .ZN(_05518_)
  );
  AND2_X1 _15691_ (
    .A1(_04708_),
    .A2(_05515_),
    .ZN(_05519_)
  );
  INV_X1 _15692_ (
    .A(_05519_),
    .ZN(_05520_)
  );
  AND2_X1 _15693_ (
    .A1(_05518_),
    .A2(_05520_),
    .ZN(_05521_)
  );
  INV_X1 _15694_ (
    .A(_05521_),
    .ZN(_05523_)
  );
  AND2_X1 _15695_ (
    .A1(_04992_),
    .A2(_05521_),
    .ZN(_05524_)
  );
  INV_X1 _15696_ (
    .A(_05524_),
    .ZN(_05525_)
  );
  AND2_X1 _15697_ (
    .A1(_04991_),
    .A2(_05523_),
    .ZN(_05526_)
  );
  INV_X1 _15698_ (
    .A(_05526_),
    .ZN(_05527_)
  );
  AND2_X1 _15699_ (
    .A1(_05525_),
    .A2(_05527_),
    .ZN(_05528_)
  );
  INV_X1 _15700_ (
    .A(_05528_),
    .ZN(_05529_)
  );
  AND2_X1 _15701_ (
    .A1(_05513_),
    .A2(_05528_),
    .ZN(_05530_)
  );
  INV_X1 _15702_ (
    .A(_05530_),
    .ZN(_05531_)
  );
  AND2_X1 _15703_ (
    .A1(_05514_),
    .A2(_05529_),
    .ZN(_05532_)
  );
  INV_X1 _15704_ (
    .A(_05532_),
    .ZN(_05534_)
  );
  AND2_X1 _15705_ (
    .A1(_05531_),
    .A2(_05534_),
    .ZN(_05535_)
  );
  INV_X1 _15706_ (
    .A(_05535_),
    .ZN(_05536_)
  );
  AND2_X1 _15707_ (
    .A1(_05463_),
    .A2(_05535_),
    .ZN(_05537_)
  );
  INV_X1 _15708_ (
    .A(_05537_),
    .ZN(_05538_)
  );
  AND2_X1 _15709_ (
    .A1(_05464_),
    .A2(_05536_),
    .ZN(_05539_)
  );
  INV_X1 _15710_ (
    .A(_05539_),
    .ZN(_05540_)
  );
  AND2_X1 _15711_ (
    .A1(_05538_),
    .A2(_05540_),
    .ZN(_05541_)
  );
  INV_X1 _15712_ (
    .A(_05541_),
    .ZN(_05542_)
  );
  AND2_X1 _15713_ (
    .A1(_05250_),
    .A2(_05541_),
    .ZN(_05543_)
  );
  INV_X1 _15714_ (
    .A(_05543_),
    .ZN(_05545_)
  );
  AND2_X1 _15715_ (
    .A1(_05251_),
    .A2(_05542_),
    .ZN(_05546_)
  );
  INV_X1 _15716_ (
    .A(_05546_),
    .ZN(_05547_)
  );
  AND2_X1 _15717_ (
    .A1(_05545_),
    .A2(_05547_),
    .ZN(_05548_)
  );
  INV_X1 _15718_ (
    .A(_05548_),
    .ZN(_05549_)
  );
  AND2_X1 _15719_ (
    .A1(divisor[20]),
    .A2(remainder[0]),
    .ZN(_05550_)
  );
  INV_X1 _15720_ (
    .A(_05550_),
    .ZN(_05551_)
  );
  AND2_X1 _15721_ (
    .A1(divisor[19]),
    .A2(remainder[1]),
    .ZN(_05552_)
  );
  INV_X1 _15722_ (
    .A(_05552_),
    .ZN(_05553_)
  );
  AND2_X1 _15723_ (
    .A1(divisor[20]),
    .A2(remainder[1]),
    .ZN(_05554_)
  );
  INV_X1 _15724_ (
    .A(_05554_),
    .ZN(_05556_)
  );
  AND2_X1 _15725_ (
    .A1(_05263_),
    .A2(_05554_),
    .ZN(_05557_)
  );
  INV_X1 _15726_ (
    .A(_05557_),
    .ZN(_05558_)
  );
  AND2_X1 _15727_ (
    .A1(_05551_),
    .A2(_05553_),
    .ZN(_05559_)
  );
  INV_X1 _15728_ (
    .A(_05559_),
    .ZN(_05560_)
  );
  AND2_X1 _15729_ (
    .A1(_05558_),
    .A2(_05560_),
    .ZN(_05561_)
  );
  INV_X1 _15730_ (
    .A(_05561_),
    .ZN(_05562_)
  );
  AND2_X1 _15731_ (
    .A1(_05266_),
    .A2(_05562_),
    .ZN(_05563_)
  );
  INV_X1 _15732_ (
    .A(_05563_),
    .ZN(_05564_)
  );
  AND2_X1 _15733_ (
    .A1(_05265_),
    .A2(_05561_),
    .ZN(_05565_)
  );
  INV_X1 _15734_ (
    .A(_05565_),
    .ZN(_05567_)
  );
  AND2_X1 _15735_ (
    .A1(_05266_),
    .A2(_05561_),
    .ZN(_05568_)
  );
  INV_X1 _15736_ (
    .A(_05568_),
    .ZN(_05569_)
  );
  AND2_X1 _15737_ (
    .A1(_05265_),
    .A2(_05562_),
    .ZN(_05570_)
  );
  INV_X1 _15738_ (
    .A(_05570_),
    .ZN(_05571_)
  );
  AND2_X1 _15739_ (
    .A1(_05564_),
    .A2(_05567_),
    .ZN(_05572_)
  );
  AND2_X1 _15740_ (
    .A1(_05569_),
    .A2(_05571_),
    .ZN(_05573_)
  );
  AND2_X1 _15741_ (
    .A1(_05548_),
    .A2(_05572_),
    .ZN(_05574_)
  );
  INV_X1 _15742_ (
    .A(_05574_),
    .ZN(_05575_)
  );
  AND2_X1 _15743_ (
    .A1(_05549_),
    .A2(_05573_),
    .ZN(_05576_)
  );
  INV_X1 _15744_ (
    .A(_05576_),
    .ZN(_05578_)
  );
  AND2_X1 _15745_ (
    .A1(_05575_),
    .A2(_05578_),
    .ZN(_05579_)
  );
  INV_X1 _15746_ (
    .A(_05579_),
    .ZN(_05580_)
  );
  AND2_X1 _15747_ (
    .A1(_05274_),
    .A2(_05579_),
    .ZN(_05581_)
  );
  INV_X1 _15748_ (
    .A(_05581_),
    .ZN(_05582_)
  );
  AND2_X1 _15749_ (
    .A1(_05275_),
    .A2(_05580_),
    .ZN(_05583_)
  );
  INV_X1 _15750_ (
    .A(_05583_),
    .ZN(_05584_)
  );
  AND2_X1 _15751_ (
    .A1(_05582_),
    .A2(_05584_),
    .ZN(_05585_)
  );
  INV_X1 _15752_ (
    .A(_05585_),
    .ZN(_05586_)
  );
  AND2_X1 _15753_ (
    .A1(_05326_),
    .A2(_05332_),
    .ZN(_05587_)
  );
  INV_X1 _15754_ (
    .A(_05587_),
    .ZN(_05589_)
  );
  AND2_X1 _15755_ (
    .A1(_05312_),
    .A2(_05319_),
    .ZN(_05590_)
  );
  INV_X1 _15756_ (
    .A(_05590_),
    .ZN(_05591_)
  );
  AND2_X1 _15757_ (
    .A1(_05299_),
    .A2(_05306_),
    .ZN(_05592_)
  );
  INV_X1 _15758_ (
    .A(_05592_),
    .ZN(_05593_)
  );
  AND2_X1 _15759_ (
    .A1(_05222_),
    .A2(_05244_),
    .ZN(_05594_)
  );
  INV_X1 _15760_ (
    .A(_05594_),
    .ZN(_05595_)
  );
  AND2_X1 _15761_ (
    .A1(_05231_),
    .A2(_05238_),
    .ZN(_05596_)
  );
  INV_X1 _15762_ (
    .A(_05596_),
    .ZN(_05597_)
  );
  AND2_X1 _15763_ (
    .A1(_04087_),
    .A2(_05597_),
    .ZN(_05598_)
  );
  INV_X1 _15764_ (
    .A(_05598_),
    .ZN(_05600_)
  );
  AND2_X1 _15765_ (
    .A1(_04088_),
    .A2(_05596_),
    .ZN(_05601_)
  );
  INV_X1 _15766_ (
    .A(_05601_),
    .ZN(_05602_)
  );
  AND2_X1 _15767_ (
    .A1(_05600_),
    .A2(_05602_),
    .ZN(_05603_)
  );
  INV_X1 _15768_ (
    .A(_05603_),
    .ZN(_05604_)
  );
  AND2_X1 _15769_ (
    .A1(_04317_),
    .A2(_05603_),
    .ZN(_05605_)
  );
  INV_X1 _15770_ (
    .A(_05605_),
    .ZN(_05606_)
  );
  AND2_X1 _15771_ (
    .A1(_04316_),
    .A2(_05604_),
    .ZN(_05607_)
  );
  INV_X1 _15772_ (
    .A(_05607_),
    .ZN(_05608_)
  );
  AND2_X1 _15773_ (
    .A1(_05606_),
    .A2(_05608_),
    .ZN(_05609_)
  );
  INV_X1 _15774_ (
    .A(_05609_),
    .ZN(_05611_)
  );
  AND2_X1 _15775_ (
    .A1(_05595_),
    .A2(_05609_),
    .ZN(_05612_)
  );
  INV_X1 _15776_ (
    .A(_05612_),
    .ZN(_05613_)
  );
  AND2_X1 _15777_ (
    .A1(_05594_),
    .A2(_05611_),
    .ZN(_05614_)
  );
  INV_X1 _15778_ (
    .A(_05614_),
    .ZN(_05615_)
  );
  AND2_X1 _15779_ (
    .A1(_05613_),
    .A2(_05615_),
    .ZN(_05616_)
  );
  INV_X1 _15780_ (
    .A(_05616_),
    .ZN(_05617_)
  );
  AND2_X1 _15781_ (
    .A1(_05593_),
    .A2(_05616_),
    .ZN(_05618_)
  );
  INV_X1 _15782_ (
    .A(_05618_),
    .ZN(_05619_)
  );
  AND2_X1 _15783_ (
    .A1(_05592_),
    .A2(_05617_),
    .ZN(_05620_)
  );
  INV_X1 _15784_ (
    .A(_05620_),
    .ZN(_05622_)
  );
  AND2_X1 _15785_ (
    .A1(_05619_),
    .A2(_05622_),
    .ZN(_05623_)
  );
  INV_X1 _15786_ (
    .A(_05623_),
    .ZN(_05624_)
  );
  AND2_X1 _15787_ (
    .A1(_05591_),
    .A2(_05623_),
    .ZN(_05625_)
  );
  INV_X1 _15788_ (
    .A(_05625_),
    .ZN(_05626_)
  );
  AND2_X1 _15789_ (
    .A1(_05590_),
    .A2(_05624_),
    .ZN(_05627_)
  );
  INV_X1 _15790_ (
    .A(_05627_),
    .ZN(_05628_)
  );
  AND2_X1 _15791_ (
    .A1(_05626_),
    .A2(_05628_),
    .ZN(_05629_)
  );
  INV_X1 _15792_ (
    .A(_05629_),
    .ZN(_05630_)
  );
  AND2_X1 _15793_ (
    .A1(_03170_),
    .A2(_05629_),
    .ZN(_05631_)
  );
  INV_X1 _15794_ (
    .A(_05631_),
    .ZN(_05633_)
  );
  AND2_X1 _15795_ (
    .A1(_03169_),
    .A2(_05630_),
    .ZN(_05634_)
  );
  INV_X1 _15796_ (
    .A(_05634_),
    .ZN(_05635_)
  );
  AND2_X1 _15797_ (
    .A1(_05633_),
    .A2(_05635_),
    .ZN(_05636_)
  );
  INV_X1 _15798_ (
    .A(_05636_),
    .ZN(_05637_)
  );
  AND2_X1 _15799_ (
    .A1(_05256_),
    .A2(_05636_),
    .ZN(_05638_)
  );
  INV_X1 _15800_ (
    .A(_05638_),
    .ZN(_05639_)
  );
  AND2_X1 _15801_ (
    .A1(_05257_),
    .A2(_05637_),
    .ZN(_05640_)
  );
  INV_X1 _15802_ (
    .A(_05640_),
    .ZN(_05641_)
  );
  AND2_X1 _15803_ (
    .A1(_05639_),
    .A2(_05641_),
    .ZN(_05642_)
  );
  INV_X1 _15804_ (
    .A(_05642_),
    .ZN(_05644_)
  );
  AND2_X1 _15805_ (
    .A1(_05589_),
    .A2(_05642_),
    .ZN(_05645_)
  );
  INV_X1 _15806_ (
    .A(_05645_),
    .ZN(_05646_)
  );
  AND2_X1 _15807_ (
    .A1(_05587_),
    .A2(_05644_),
    .ZN(_05647_)
  );
  INV_X1 _15808_ (
    .A(_05647_),
    .ZN(_05648_)
  );
  AND2_X1 _15809_ (
    .A1(_05646_),
    .A2(_05648_),
    .ZN(_05649_)
  );
  INV_X1 _15810_ (
    .A(_05649_),
    .ZN(_05650_)
  );
  AND2_X1 _15811_ (
    .A1(_05585_),
    .A2(_05649_),
    .ZN(_05651_)
  );
  INV_X1 _15812_ (
    .A(_05651_),
    .ZN(_05652_)
  );
  AND2_X1 _15813_ (
    .A1(_05586_),
    .A2(_05650_),
    .ZN(_05653_)
  );
  INV_X1 _15814_ (
    .A(_05653_),
    .ZN(_05655_)
  );
  AND2_X1 _15815_ (
    .A1(_05652_),
    .A2(_05655_),
    .ZN(_05656_)
  );
  INV_X1 _15816_ (
    .A(_05656_),
    .ZN(_05657_)
  );
  AND2_X1 _15817_ (
    .A1(_05426_),
    .A2(_05656_),
    .ZN(_05658_)
  );
  INV_X1 _15818_ (
    .A(_05658_),
    .ZN(_05659_)
  );
  AND2_X1 _15819_ (
    .A1(_05425_),
    .A2(_05657_),
    .ZN(_05660_)
  );
  INV_X1 _15820_ (
    .A(_05660_),
    .ZN(_05661_)
  );
  AND2_X1 _15821_ (
    .A1(_05659_),
    .A2(_05661_),
    .ZN(_05662_)
  );
  INV_X1 _15822_ (
    .A(_05662_),
    .ZN(_05663_)
  );
  AND2_X1 _15823_ (
    .A1(_05424_),
    .A2(_05662_),
    .ZN(_05664_)
  );
  INV_X1 _15824_ (
    .A(_05664_),
    .ZN(_05666_)
  );
  AND2_X1 _15825_ (
    .A1(_05422_),
    .A2(_05663_),
    .ZN(_05667_)
  );
  INV_X1 _15826_ (
    .A(_05667_),
    .ZN(_05668_)
  );
  AND2_X1 _15827_ (
    .A1(_05666_),
    .A2(_05668_),
    .ZN(_05669_)
  );
  INV_X1 _15828_ (
    .A(_05669_),
    .ZN(_05670_)
  );
  AND2_X1 _15829_ (
    .A1(_05421_),
    .A2(_05669_),
    .ZN(_05671_)
  );
  INV_X1 _15830_ (
    .A(_05671_),
    .ZN(_05672_)
  );
  AND2_X1 _15831_ (
    .A1(_05420_),
    .A2(_05670_),
    .ZN(_05673_)
  );
  INV_X1 _15832_ (
    .A(_05673_),
    .ZN(_05674_)
  );
  AND2_X1 _15833_ (
    .A1(_05672_),
    .A2(_05674_),
    .ZN(_05675_)
  );
  INV_X1 _15834_ (
    .A(_05675_),
    .ZN(_05677_)
  );
  AND2_X1 _15835_ (
    .A1(_05371_),
    .A2(_05675_),
    .ZN(_05678_)
  );
  INV_X1 _15836_ (
    .A(_05678_),
    .ZN(_05679_)
  );
  AND2_X1 _15837_ (
    .A1(_05372_),
    .A2(_05677_),
    .ZN(_05680_)
  );
  INV_X1 _15838_ (
    .A(_05680_),
    .ZN(_05681_)
  );
  AND2_X1 _15839_ (
    .A1(_05679_),
    .A2(_05681_),
    .ZN(_05682_)
  );
  INV_X1 _15840_ (
    .A(_05682_),
    .ZN(_05683_)
  );
  AND2_X1 _15841_ (
    .A1(_05067_),
    .A2(_05378_),
    .ZN(_05684_)
  );
  INV_X1 _15842_ (
    .A(_05684_),
    .ZN(_05685_)
  );
  AND2_X1 _15843_ (
    .A1(_05072_),
    .A2(_05382_),
    .ZN(_05686_)
  );
  INV_X1 _15844_ (
    .A(_05686_),
    .ZN(_05688_)
  );
  AND2_X1 _15845_ (
    .A1(_05381_),
    .A2(_05685_),
    .ZN(_05689_)
  );
  INV_X1 _15846_ (
    .A(_05689_),
    .ZN(_05690_)
  );
  AND2_X1 _15847_ (
    .A1(_05688_),
    .A2(_05690_),
    .ZN(_05691_)
  );
  INV_X1 _15848_ (
    .A(_05691_),
    .ZN(_05692_)
  );
  AND2_X1 _15849_ (
    .A1(_05682_),
    .A2(_05692_),
    .ZN(_05693_)
  );
  INV_X1 _15850_ (
    .A(_05693_),
    .ZN(_05694_)
  );
  AND2_X1 _15851_ (
    .A1(_05683_),
    .A2(_05691_),
    .ZN(_05695_)
  );
  INV_X1 _15852_ (
    .A(_05695_),
    .ZN(_05696_)
  );
  AND2_X1 _15853_ (
    .A1(_05694_),
    .A2(_05696_),
    .ZN(_05697_)
  );
  INV_X1 _15854_ (
    .A(_05697_),
    .ZN(_05699_)
  );
  AND2_X1 _15855_ (
    .A1(remainder[53]),
    .A2(_05697_),
    .ZN(_05700_)
  );
  INV_X1 _15856_ (
    .A(_05700_),
    .ZN(_05701_)
  );
  AND2_X1 _15857_ (
    .A1(_04536_),
    .A2(_05699_),
    .ZN(_05702_)
  );
  INV_X1 _15858_ (
    .A(_05702_),
    .ZN(_05703_)
  );
  AND2_X1 _15859_ (
    .A1(_05701_),
    .A2(_05703_),
    .ZN(_05704_)
  );
  INV_X1 _15860_ (
    .A(_05704_),
    .ZN(_05705_)
  );
  AND2_X1 _15861_ (
    .A1(_05114_),
    .A2(_05398_),
    .ZN(_05706_)
  );
  INV_X1 _15862_ (
    .A(_05706_),
    .ZN(_05707_)
  );
  AND2_X1 _15863_ (
    .A1(_05113_),
    .A2(_05396_),
    .ZN(_05708_)
  );
  INV_X1 _15864_ (
    .A(_05708_),
    .ZN(_05710_)
  );
  AND2_X1 _15865_ (
    .A1(_05396_),
    .A2(_05707_),
    .ZN(_05711_)
  );
  AND2_X1 _15866_ (
    .A1(_05398_),
    .A2(_05710_),
    .ZN(_05712_)
  );
  AND2_X1 _15867_ (
    .A1(_05704_),
    .A2(_05712_),
    .ZN(_05713_)
  );
  INV_X1 _15868_ (
    .A(_05713_),
    .ZN(_05714_)
  );
  AND2_X1 _15869_ (
    .A1(_05705_),
    .A2(_05711_),
    .ZN(_05715_)
  );
  INV_X1 _15870_ (
    .A(_05715_),
    .ZN(_05716_)
  );
  AND2_X1 _15871_ (
    .A1(_02082_),
    .A2(_05714_),
    .ZN(_05717_)
  );
  AND2_X1 _15872_ (
    .A1(_05716_),
    .A2(_05717_),
    .ZN(_05718_)
  );
  INV_X1 _15873_ (
    .A(_05718_),
    .ZN(_05719_)
  );
  AND2_X1 _15874_ (
    .A1(remainder[45]),
    .A2(_02077_),
    .ZN(_05721_)
  );
  INV_X1 _15875_ (
    .A(_05721_),
    .ZN(_05722_)
  );
  AND2_X1 _15876_ (
    .A1(_05719_),
    .A2(_05722_),
    .ZN(_05723_)
  );
  AND2_X1 _15877_ (
    .A1(_05419_),
    .A2(_05723_),
    .ZN(_05724_)
  );
  INV_X1 _15878_ (
    .A(_05724_),
    .ZN(_05725_)
  );
  AND2_X1 _15879_ (
    .A1(_06201_),
    .A2(_05725_),
    .ZN(_00066_)
  );
  AND2_X1 _15880_ (
    .A1(_04623_),
    .A2(_10451_),
    .ZN(_05726_)
  );
  INV_X1 _15881_ (
    .A(_05726_),
    .ZN(_05727_)
  );
  AND2_X1 _15882_ (
    .A1(_10462_),
    .A2(_01802_),
    .ZN(_05728_)
  );
  INV_X1 _15883_ (
    .A(_05728_),
    .ZN(_05729_)
  );
  AND2_X1 _15884_ (
    .A1(_05983_),
    .A2(_05729_),
    .ZN(_05731_)
  );
  AND2_X1 _15885_ (
    .A1(_05727_),
    .A2(_05731_),
    .ZN(_05732_)
  );
  INV_X1 _15886_ (
    .A(_05732_),
    .ZN(_05733_)
  );
  AND2_X1 _15887_ (
    .A1(remainder[46]),
    .A2(_02077_),
    .ZN(_05734_)
  );
  INV_X1 _15888_ (
    .A(_05734_),
    .ZN(_05735_)
  );
  AND2_X1 _15889_ (
    .A1(_05701_),
    .A2(_05714_),
    .ZN(_05736_)
  );
  INV_X1 _15890_ (
    .A(_05736_),
    .ZN(_05737_)
  );
  AND2_X1 _15891_ (
    .A1(_05679_),
    .A2(_05694_),
    .ZN(_05738_)
  );
  INV_X1 _15892_ (
    .A(_05738_),
    .ZN(_05739_)
  );
  AND2_X1 _15893_ (
    .A1(_05659_),
    .A2(_05666_),
    .ZN(_05740_)
  );
  INV_X1 _15894_ (
    .A(_05740_),
    .ZN(_05742_)
  );
  AND2_X1 _15895_ (
    .A1(_05639_),
    .A2(_05646_),
    .ZN(_05743_)
  );
  INV_X1 _15896_ (
    .A(_05743_),
    .ZN(_05744_)
  );
  AND2_X1 _15897_ (
    .A1(_05582_),
    .A2(_05652_),
    .ZN(_05745_)
  );
  INV_X1 _15898_ (
    .A(_05745_),
    .ZN(_05746_)
  );
  AND2_X1 _15899_ (
    .A1(_03249_),
    .A2(_05562_),
    .ZN(_05747_)
  );
  INV_X1 _15900_ (
    .A(_05747_),
    .ZN(_05748_)
  );
  AND2_X1 _15901_ (
    .A1(_05263_),
    .A2(_05747_),
    .ZN(_05749_)
  );
  INV_X1 _15902_ (
    .A(_05749_),
    .ZN(_05750_)
  );
  AND2_X1 _15903_ (
    .A1(_05575_),
    .A2(_05750_),
    .ZN(_05751_)
  );
  INV_X1 _15904_ (
    .A(_05751_),
    .ZN(_05753_)
  );
  AND2_X1 _15905_ (
    .A1(_05459_),
    .A2(_05538_),
    .ZN(_05754_)
  );
  INV_X1 _15906_ (
    .A(_05754_),
    .ZN(_05755_)
  );
  AND2_X1 _15907_ (
    .A1(_05491_),
    .A2(_05503_),
    .ZN(_05756_)
  );
  INV_X1 _15908_ (
    .A(_05756_),
    .ZN(_05757_)
  );
  AND2_X1 _15909_ (
    .A1(_05477_),
    .A2(_05484_),
    .ZN(_05758_)
  );
  INV_X1 _15910_ (
    .A(_05758_),
    .ZN(_05759_)
  );
  AND2_X1 _15911_ (
    .A1(remainder[32]),
    .A2(divisor[13]),
    .ZN(_05760_)
  );
  INV_X1 _15912_ (
    .A(_05760_),
    .ZN(_05761_)
  );
  AND2_X1 _15913_ (
    .A1(divisor[14]),
    .A2(remainder[7]),
    .ZN(_05762_)
  );
  INV_X1 _15914_ (
    .A(_05762_),
    .ZN(_05764_)
  );
  AND2_X1 _15915_ (
    .A1(divisor[15]),
    .A2(remainder[7]),
    .ZN(_05765_)
  );
  INV_X1 _15916_ (
    .A(_05765_),
    .ZN(_05766_)
  );
  AND2_X1 _15917_ (
    .A1(_05472_),
    .A2(_05765_),
    .ZN(_05767_)
  );
  INV_X1 _15918_ (
    .A(_05767_),
    .ZN(_05768_)
  );
  AND2_X1 _15919_ (
    .A1(_05475_),
    .A2(_05764_),
    .ZN(_05769_)
  );
  INV_X1 _15920_ (
    .A(_05769_),
    .ZN(_05770_)
  );
  AND2_X1 _15921_ (
    .A1(_05768_),
    .A2(_05770_),
    .ZN(_05771_)
  );
  INV_X1 _15922_ (
    .A(_05771_),
    .ZN(_05772_)
  );
  AND2_X1 _15923_ (
    .A1(_05760_),
    .A2(_05771_),
    .ZN(_05773_)
  );
  INV_X1 _15924_ (
    .A(_05773_),
    .ZN(_05775_)
  );
  AND2_X1 _15925_ (
    .A1(_05761_),
    .A2(_05772_),
    .ZN(_05776_)
  );
  INV_X1 _15926_ (
    .A(_05776_),
    .ZN(_05777_)
  );
  AND2_X1 _15927_ (
    .A1(_05775_),
    .A2(_05777_),
    .ZN(_05778_)
  );
  INV_X1 _15928_ (
    .A(_05778_),
    .ZN(_05779_)
  );
  AND2_X1 _15929_ (
    .A1(_05759_),
    .A2(_05778_),
    .ZN(_05780_)
  );
  INV_X1 _15930_ (
    .A(_05780_),
    .ZN(_05781_)
  );
  AND2_X1 _15931_ (
    .A1(_05758_),
    .A2(_05779_),
    .ZN(_05782_)
  );
  INV_X1 _15932_ (
    .A(_05782_),
    .ZN(_05783_)
  );
  AND2_X1 _15933_ (
    .A1(_05781_),
    .A2(_05783_),
    .ZN(_05784_)
  );
  INV_X1 _15934_ (
    .A(_05784_),
    .ZN(_05786_)
  );
  AND2_X1 _15935_ (
    .A1(_05499_),
    .A2(_05784_),
    .ZN(_05787_)
  );
  INV_X1 _15936_ (
    .A(_05787_),
    .ZN(_05788_)
  );
  AND2_X1 _15937_ (
    .A1(_05501_),
    .A2(_05786_),
    .ZN(_05789_)
  );
  INV_X1 _15938_ (
    .A(_05789_),
    .ZN(_05790_)
  );
  AND2_X1 _15939_ (
    .A1(_05788_),
    .A2(_05790_),
    .ZN(_05791_)
  );
  INV_X1 _15940_ (
    .A(_05791_),
    .ZN(_05792_)
  );
  AND2_X1 _15941_ (
    .A1(_05757_),
    .A2(_05791_),
    .ZN(_05793_)
  );
  INV_X1 _15942_ (
    .A(_05793_),
    .ZN(_05794_)
  );
  AND2_X1 _15943_ (
    .A1(_05756_),
    .A2(_05792_),
    .ZN(_05795_)
  );
  INV_X1 _15944_ (
    .A(_05795_),
    .ZN(_05797_)
  );
  AND2_X1 _15945_ (
    .A1(_05794_),
    .A2(_05797_),
    .ZN(_05798_)
  );
  INV_X1 _15946_ (
    .A(_05798_),
    .ZN(_05799_)
  );
  AND2_X1 _15947_ (
    .A1(_05200_),
    .A2(_05498_),
    .ZN(_05800_)
  );
  INV_X1 _15948_ (
    .A(_05800_),
    .ZN(_05801_)
  );
  AND2_X1 _15949_ (
    .A1(_04707_),
    .A2(_05801_),
    .ZN(_05802_)
  );
  INV_X1 _15950_ (
    .A(_05802_),
    .ZN(_05803_)
  );
  AND2_X1 _15951_ (
    .A1(_04708_),
    .A2(_05800_),
    .ZN(_05804_)
  );
  INV_X1 _15952_ (
    .A(_05804_),
    .ZN(_05805_)
  );
  AND2_X1 _15953_ (
    .A1(_05803_),
    .A2(_05805_),
    .ZN(_05806_)
  );
  INV_X1 _15954_ (
    .A(_05806_),
    .ZN(_05808_)
  );
  AND2_X1 _15955_ (
    .A1(_04992_),
    .A2(_05806_),
    .ZN(_05809_)
  );
  INV_X1 _15956_ (
    .A(_05809_),
    .ZN(_05810_)
  );
  AND2_X1 _15957_ (
    .A1(_04991_),
    .A2(_05808_),
    .ZN(_05811_)
  );
  INV_X1 _15958_ (
    .A(_05811_),
    .ZN(_05812_)
  );
  AND2_X1 _15959_ (
    .A1(_05810_),
    .A2(_05812_),
    .ZN(_05813_)
  );
  INV_X1 _15960_ (
    .A(_05813_),
    .ZN(_05814_)
  );
  AND2_X1 _15961_ (
    .A1(_05798_),
    .A2(_05813_),
    .ZN(_05815_)
  );
  INV_X1 _15962_ (
    .A(_05815_),
    .ZN(_05816_)
  );
  AND2_X1 _15963_ (
    .A1(_05799_),
    .A2(_05814_),
    .ZN(_05817_)
  );
  INV_X1 _15964_ (
    .A(_05817_),
    .ZN(_05819_)
  );
  AND2_X1 _15965_ (
    .A1(_05816_),
    .A2(_05819_),
    .ZN(_05820_)
  );
  INV_X1 _15966_ (
    .A(_05820_),
    .ZN(_05821_)
  );
  AND2_X1 _15967_ (
    .A1(_05437_),
    .A2(_05443_),
    .ZN(_05822_)
  );
  INV_X1 _15968_ (
    .A(_05822_),
    .ZN(_05823_)
  );
  AND2_X1 _15969_ (
    .A1(divisor[16]),
    .A2(remainder[5]),
    .ZN(_05824_)
  );
  INV_X1 _15970_ (
    .A(_05824_),
    .ZN(_05825_)
  );
  AND2_X1 _15971_ (
    .A1(divisor[17]),
    .A2(remainder[4]),
    .ZN(_05826_)
  );
  INV_X1 _15972_ (
    .A(_05826_),
    .ZN(_05827_)
  );
  AND2_X1 _15973_ (
    .A1(divisor[18]),
    .A2(remainder[4]),
    .ZN(_05828_)
  );
  INV_X1 _15974_ (
    .A(_05828_),
    .ZN(_05830_)
  );
  AND2_X1 _15975_ (
    .A1(_05433_),
    .A2(_05826_),
    .ZN(_05831_)
  );
  INV_X1 _15976_ (
    .A(_05831_),
    .ZN(_05832_)
  );
  AND2_X1 _15977_ (
    .A1(_05435_),
    .A2(_05827_),
    .ZN(_05833_)
  );
  INV_X1 _15978_ (
    .A(_05833_),
    .ZN(_05834_)
  );
  AND2_X1 _15979_ (
    .A1(_05832_),
    .A2(_05834_),
    .ZN(_05835_)
  );
  INV_X1 _15980_ (
    .A(_05835_),
    .ZN(_05836_)
  );
  AND2_X1 _15981_ (
    .A1(_05824_),
    .A2(_05835_),
    .ZN(_05837_)
  );
  INV_X1 _15982_ (
    .A(_05837_),
    .ZN(_05838_)
  );
  AND2_X1 _15983_ (
    .A1(_05825_),
    .A2(_05836_),
    .ZN(_05839_)
  );
  INV_X1 _15984_ (
    .A(_05839_),
    .ZN(_05841_)
  );
  AND2_X1 _15985_ (
    .A1(_05838_),
    .A2(_05841_),
    .ZN(_05842_)
  );
  INV_X1 _15986_ (
    .A(_05842_),
    .ZN(_05843_)
  );
  AND2_X1 _15987_ (
    .A1(_05557_),
    .A2(_05842_),
    .ZN(_05844_)
  );
  INV_X1 _15988_ (
    .A(_05844_),
    .ZN(_05845_)
  );
  AND2_X1 _15989_ (
    .A1(_05558_),
    .A2(_05843_),
    .ZN(_05846_)
  );
  INV_X1 _15990_ (
    .A(_05846_),
    .ZN(_05847_)
  );
  AND2_X1 _15991_ (
    .A1(_05845_),
    .A2(_05847_),
    .ZN(_05848_)
  );
  INV_X1 _15992_ (
    .A(_05848_),
    .ZN(_05849_)
  );
  AND2_X1 _15993_ (
    .A1(_05823_),
    .A2(_05848_),
    .ZN(_05850_)
  );
  INV_X1 _15994_ (
    .A(_05850_),
    .ZN(_05852_)
  );
  AND2_X1 _15995_ (
    .A1(_05822_),
    .A2(_05849_),
    .ZN(_05853_)
  );
  INV_X1 _15996_ (
    .A(_05853_),
    .ZN(_05854_)
  );
  AND2_X1 _15997_ (
    .A1(_05852_),
    .A2(_05854_),
    .ZN(_05855_)
  );
  INV_X1 _15998_ (
    .A(_05855_),
    .ZN(_05856_)
  );
  AND2_X1 _15999_ (
    .A1(_05450_),
    .A2(_05457_),
    .ZN(_05857_)
  );
  INV_X1 _16000_ (
    .A(_05857_),
    .ZN(_05858_)
  );
  AND2_X1 _16001_ (
    .A1(_05855_),
    .A2(_05857_),
    .ZN(_05859_)
  );
  INV_X1 _16002_ (
    .A(_05859_),
    .ZN(_05860_)
  );
  AND2_X1 _16003_ (
    .A1(_05856_),
    .A2(_05858_),
    .ZN(_05861_)
  );
  INV_X1 _16004_ (
    .A(_05861_),
    .ZN(_05863_)
  );
  AND2_X1 _16005_ (
    .A1(_05856_),
    .A2(_05857_),
    .ZN(_05864_)
  );
  INV_X1 _16006_ (
    .A(_05864_),
    .ZN(_05865_)
  );
  AND2_X1 _16007_ (
    .A1(_05855_),
    .A2(_05858_),
    .ZN(_05866_)
  );
  INV_X1 _16008_ (
    .A(_05866_),
    .ZN(_05867_)
  );
  AND2_X1 _16009_ (
    .A1(_05860_),
    .A2(_05863_),
    .ZN(_05868_)
  );
  AND2_X1 _16010_ (
    .A1(_05865_),
    .A2(_05867_),
    .ZN(_05869_)
  );
  AND2_X1 _16011_ (
    .A1(_05820_),
    .A2(_05869_),
    .ZN(_05870_)
  );
  INV_X1 _16012_ (
    .A(_05870_),
    .ZN(_05871_)
  );
  AND2_X1 _16013_ (
    .A1(_05821_),
    .A2(_05868_),
    .ZN(_05872_)
  );
  INV_X1 _16014_ (
    .A(_05872_),
    .ZN(_05874_)
  );
  AND2_X1 _16015_ (
    .A1(_05871_),
    .A2(_05874_),
    .ZN(_05875_)
  );
  INV_X1 _16016_ (
    .A(_05875_),
    .ZN(_05876_)
  );
  AND2_X1 _16017_ (
    .A1(_05755_),
    .A2(_05875_),
    .ZN(_05877_)
  );
  INV_X1 _16018_ (
    .A(_05877_),
    .ZN(_05878_)
  );
  AND2_X1 _16019_ (
    .A1(_05754_),
    .A2(_05876_),
    .ZN(_05879_)
  );
  INV_X1 _16020_ (
    .A(_05879_),
    .ZN(_05880_)
  );
  AND2_X1 _16021_ (
    .A1(_05878_),
    .A2(_05880_),
    .ZN(_05881_)
  );
  INV_X1 _16022_ (
    .A(_05881_),
    .ZN(_05882_)
  );
  AND2_X1 _16023_ (
    .A1(divisor[19]),
    .A2(remainder[2]),
    .ZN(_05883_)
  );
  INV_X1 _16024_ (
    .A(_05883_),
    .ZN(_05885_)
  );
  AND2_X1 _16025_ (
    .A1(divisor[21]),
    .A2(remainder[0]),
    .ZN(_05886_)
  );
  INV_X1 _16026_ (
    .A(_05886_),
    .ZN(_05887_)
  );
  AND2_X1 _16027_ (
    .A1(divisor[21]),
    .A2(remainder[1]),
    .ZN(_05888_)
  );
  INV_X1 _16028_ (
    .A(_05888_),
    .ZN(_05889_)
  );
  AND2_X1 _16029_ (
    .A1(_05550_),
    .A2(_05888_),
    .ZN(_05890_)
  );
  INV_X1 _16030_ (
    .A(_05890_),
    .ZN(_05891_)
  );
  AND2_X1 _16031_ (
    .A1(_05556_),
    .A2(_05887_),
    .ZN(_05892_)
  );
  INV_X1 _16032_ (
    .A(_05892_),
    .ZN(_05893_)
  );
  AND2_X1 _16033_ (
    .A1(_05891_),
    .A2(_05893_),
    .ZN(_05894_)
  );
  INV_X1 _16034_ (
    .A(_05894_),
    .ZN(_05896_)
  );
  AND2_X1 _16035_ (
    .A1(_05883_),
    .A2(_05894_),
    .ZN(_05897_)
  );
  INV_X1 _16036_ (
    .A(_05897_),
    .ZN(_05898_)
  );
  AND2_X1 _16037_ (
    .A1(_05885_),
    .A2(_05896_),
    .ZN(_05899_)
  );
  INV_X1 _16038_ (
    .A(_05899_),
    .ZN(_05900_)
  );
  AND2_X1 _16039_ (
    .A1(_05898_),
    .A2(_05900_),
    .ZN(_05901_)
  );
  INV_X1 _16040_ (
    .A(_05901_),
    .ZN(_05902_)
  );
  AND2_X1 _16041_ (
    .A1(_05747_),
    .A2(_05902_),
    .ZN(_05903_)
  );
  INV_X1 _16042_ (
    .A(_05903_),
    .ZN(_05904_)
  );
  AND2_X1 _16043_ (
    .A1(_05748_),
    .A2(_05901_),
    .ZN(_05905_)
  );
  INV_X1 _16044_ (
    .A(_05905_),
    .ZN(_05907_)
  );
  AND2_X1 _16045_ (
    .A1(_05748_),
    .A2(_05902_),
    .ZN(_05908_)
  );
  INV_X1 _16046_ (
    .A(_05908_),
    .ZN(_05909_)
  );
  AND2_X1 _16047_ (
    .A1(_05747_),
    .A2(_05901_),
    .ZN(_05910_)
  );
  INV_X1 _16048_ (
    .A(_05910_),
    .ZN(_05911_)
  );
  AND2_X1 _16049_ (
    .A1(_05904_),
    .A2(_05907_),
    .ZN(_05912_)
  );
  AND2_X1 _16050_ (
    .A1(_05909_),
    .A2(_05911_),
    .ZN(_05913_)
  );
  AND2_X1 _16051_ (
    .A1(_05881_),
    .A2(_05913_),
    .ZN(_05914_)
  );
  INV_X1 _16052_ (
    .A(_05914_),
    .ZN(_05915_)
  );
  AND2_X1 _16053_ (
    .A1(_05882_),
    .A2(_05912_),
    .ZN(_05916_)
  );
  INV_X1 _16054_ (
    .A(_05916_),
    .ZN(_05918_)
  );
  AND2_X1 _16055_ (
    .A1(_05915_),
    .A2(_05918_),
    .ZN(_05919_)
  );
  INV_X1 _16056_ (
    .A(_05919_),
    .ZN(_05920_)
  );
  AND2_X1 _16057_ (
    .A1(_05753_),
    .A2(_05919_),
    .ZN(_05921_)
  );
  INV_X1 _16058_ (
    .A(_05921_),
    .ZN(_05922_)
  );
  AND2_X1 _16059_ (
    .A1(_05751_),
    .A2(_05920_),
    .ZN(_05923_)
  );
  INV_X1 _16060_ (
    .A(_05923_),
    .ZN(_05924_)
  );
  AND2_X1 _16061_ (
    .A1(_05922_),
    .A2(_05924_),
    .ZN(_05925_)
  );
  INV_X1 _16062_ (
    .A(_05925_),
    .ZN(_05926_)
  );
  AND2_X1 _16063_ (
    .A1(_05626_),
    .A2(_05633_),
    .ZN(_05927_)
  );
  INV_X1 _16064_ (
    .A(_05927_),
    .ZN(_05929_)
  );
  AND2_X1 _16065_ (
    .A1(_05613_),
    .A2(_05619_),
    .ZN(_05930_)
  );
  INV_X1 _16066_ (
    .A(_05930_),
    .ZN(_05931_)
  );
  AND2_X1 _16067_ (
    .A1(_05600_),
    .A2(_05606_),
    .ZN(_05932_)
  );
  INV_X1 _16068_ (
    .A(_05932_),
    .ZN(_05933_)
  );
  AND2_X1 _16069_ (
    .A1(_05509_),
    .A2(_05531_),
    .ZN(_05934_)
  );
  INV_X1 _16070_ (
    .A(_05934_),
    .ZN(_05935_)
  );
  AND2_X1 _16071_ (
    .A1(_05518_),
    .A2(_05525_),
    .ZN(_05936_)
  );
  INV_X1 _16072_ (
    .A(_05936_),
    .ZN(_05937_)
  );
  AND2_X1 _16073_ (
    .A1(_04087_),
    .A2(_05937_),
    .ZN(_05938_)
  );
  INV_X1 _16074_ (
    .A(_05938_),
    .ZN(_05940_)
  );
  AND2_X1 _16075_ (
    .A1(_04088_),
    .A2(_05936_),
    .ZN(_05941_)
  );
  INV_X1 _16076_ (
    .A(_05941_),
    .ZN(_05942_)
  );
  AND2_X1 _16077_ (
    .A1(_05940_),
    .A2(_05942_),
    .ZN(_05943_)
  );
  INV_X1 _16078_ (
    .A(_05943_),
    .ZN(_05944_)
  );
  AND2_X1 _16079_ (
    .A1(_04317_),
    .A2(_05943_),
    .ZN(_05945_)
  );
  INV_X1 _16080_ (
    .A(_05945_),
    .ZN(_05946_)
  );
  AND2_X1 _16081_ (
    .A1(_04316_),
    .A2(_05944_),
    .ZN(_05947_)
  );
  INV_X1 _16082_ (
    .A(_05947_),
    .ZN(_05948_)
  );
  AND2_X1 _16083_ (
    .A1(_05946_),
    .A2(_05948_),
    .ZN(_05949_)
  );
  INV_X1 _16084_ (
    .A(_05949_),
    .ZN(_05951_)
  );
  AND2_X1 _16085_ (
    .A1(_05935_),
    .A2(_05949_),
    .ZN(_05952_)
  );
  INV_X1 _16086_ (
    .A(_05952_),
    .ZN(_05953_)
  );
  AND2_X1 _16087_ (
    .A1(_05934_),
    .A2(_05951_),
    .ZN(_05954_)
  );
  INV_X1 _16088_ (
    .A(_05954_),
    .ZN(_05955_)
  );
  AND2_X1 _16089_ (
    .A1(_05953_),
    .A2(_05955_),
    .ZN(_05956_)
  );
  INV_X1 _16090_ (
    .A(_05956_),
    .ZN(_05957_)
  );
  AND2_X1 _16091_ (
    .A1(_05933_),
    .A2(_05956_),
    .ZN(_05958_)
  );
  INV_X1 _16092_ (
    .A(_05958_),
    .ZN(_05959_)
  );
  AND2_X1 _16093_ (
    .A1(_05932_),
    .A2(_05957_),
    .ZN(_05960_)
  );
  INV_X1 _16094_ (
    .A(_05960_),
    .ZN(_05962_)
  );
  AND2_X1 _16095_ (
    .A1(_05959_),
    .A2(_05962_),
    .ZN(_05963_)
  );
  INV_X1 _16096_ (
    .A(_05963_),
    .ZN(_05964_)
  );
  AND2_X1 _16097_ (
    .A1(_05931_),
    .A2(_05963_),
    .ZN(_05965_)
  );
  INV_X1 _16098_ (
    .A(_05965_),
    .ZN(_05966_)
  );
  AND2_X1 _16099_ (
    .A1(_05930_),
    .A2(_05964_),
    .ZN(_05967_)
  );
  INV_X1 _16100_ (
    .A(_05967_),
    .ZN(_05968_)
  );
  AND2_X1 _16101_ (
    .A1(_05966_),
    .A2(_05968_),
    .ZN(_05969_)
  );
  INV_X1 _16102_ (
    .A(_05969_),
    .ZN(_05970_)
  );
  AND2_X1 _16103_ (
    .A1(_03170_),
    .A2(_05969_),
    .ZN(_05971_)
  );
  INV_X1 _16104_ (
    .A(_05971_),
    .ZN(_05973_)
  );
  AND2_X1 _16105_ (
    .A1(_03169_),
    .A2(_05970_),
    .ZN(_05974_)
  );
  INV_X1 _16106_ (
    .A(_05974_),
    .ZN(_05975_)
  );
  AND2_X1 _16107_ (
    .A1(_05973_),
    .A2(_05975_),
    .ZN(_05976_)
  );
  INV_X1 _16108_ (
    .A(_05976_),
    .ZN(_05977_)
  );
  AND2_X1 _16109_ (
    .A1(_05543_),
    .A2(_05976_),
    .ZN(_05978_)
  );
  INV_X1 _16110_ (
    .A(_05978_),
    .ZN(_05979_)
  );
  AND2_X1 _16111_ (
    .A1(_05545_),
    .A2(_05977_),
    .ZN(_05980_)
  );
  INV_X1 _16112_ (
    .A(_05980_),
    .ZN(_05981_)
  );
  AND2_X1 _16113_ (
    .A1(_05979_),
    .A2(_05981_),
    .ZN(_05982_)
  );
  INV_X1 _16114_ (
    .A(_05982_),
    .ZN(_05984_)
  );
  AND2_X1 _16115_ (
    .A1(_05929_),
    .A2(_05982_),
    .ZN(_05985_)
  );
  INV_X1 _16116_ (
    .A(_05985_),
    .ZN(_05986_)
  );
  AND2_X1 _16117_ (
    .A1(_05927_),
    .A2(_05984_),
    .ZN(_05987_)
  );
  INV_X1 _16118_ (
    .A(_05987_),
    .ZN(_05988_)
  );
  AND2_X1 _16119_ (
    .A1(_05986_),
    .A2(_05988_),
    .ZN(_05989_)
  );
  INV_X1 _16120_ (
    .A(_05989_),
    .ZN(_05990_)
  );
  AND2_X1 _16121_ (
    .A1(_05925_),
    .A2(_05989_),
    .ZN(_05991_)
  );
  INV_X1 _16122_ (
    .A(_05991_),
    .ZN(_05992_)
  );
  AND2_X1 _16123_ (
    .A1(_05926_),
    .A2(_05990_),
    .ZN(_05993_)
  );
  INV_X1 _16124_ (
    .A(_05993_),
    .ZN(_05995_)
  );
  AND2_X1 _16125_ (
    .A1(_05992_),
    .A2(_05995_),
    .ZN(_05996_)
  );
  INV_X1 _16126_ (
    .A(_05996_),
    .ZN(_05997_)
  );
  AND2_X1 _16127_ (
    .A1(_05746_),
    .A2(_05996_),
    .ZN(_05998_)
  );
  INV_X1 _16128_ (
    .A(_05998_),
    .ZN(_05999_)
  );
  AND2_X1 _16129_ (
    .A1(_05745_),
    .A2(_05997_),
    .ZN(_06000_)
  );
  INV_X1 _16130_ (
    .A(_06000_),
    .ZN(_06001_)
  );
  AND2_X1 _16131_ (
    .A1(_05999_),
    .A2(_06001_),
    .ZN(_06002_)
  );
  INV_X1 _16132_ (
    .A(_06002_),
    .ZN(_06003_)
  );
  AND2_X1 _16133_ (
    .A1(_05744_),
    .A2(_06002_),
    .ZN(_06004_)
  );
  INV_X1 _16134_ (
    .A(_06004_),
    .ZN(_06006_)
  );
  AND2_X1 _16135_ (
    .A1(_05743_),
    .A2(_06003_),
    .ZN(_06007_)
  );
  INV_X1 _16136_ (
    .A(_06007_),
    .ZN(_06008_)
  );
  AND2_X1 _16137_ (
    .A1(_06006_),
    .A2(_06008_),
    .ZN(_06009_)
  );
  INV_X1 _16138_ (
    .A(_06009_),
    .ZN(_06010_)
  );
  AND2_X1 _16139_ (
    .A1(_05742_),
    .A2(_06009_),
    .ZN(_06011_)
  );
  INV_X1 _16140_ (
    .A(_06011_),
    .ZN(_06012_)
  );
  AND2_X1 _16141_ (
    .A1(_05740_),
    .A2(_06010_),
    .ZN(_06013_)
  );
  INV_X1 _16142_ (
    .A(_06013_),
    .ZN(_06014_)
  );
  AND2_X1 _16143_ (
    .A1(_06012_),
    .A2(_06014_),
    .ZN(_06015_)
  );
  INV_X1 _16144_ (
    .A(_06015_),
    .ZN(_06017_)
  );
  AND2_X1 _16145_ (
    .A1(_05671_),
    .A2(_06015_),
    .ZN(_06018_)
  );
  INV_X1 _16146_ (
    .A(_06018_),
    .ZN(_06019_)
  );
  AND2_X1 _16147_ (
    .A1(_05672_),
    .A2(_06017_),
    .ZN(_06020_)
  );
  INV_X1 _16148_ (
    .A(_06020_),
    .ZN(_06021_)
  );
  AND2_X1 _16149_ (
    .A1(_06019_),
    .A2(_06021_),
    .ZN(_06022_)
  );
  INV_X1 _16150_ (
    .A(_06022_),
    .ZN(_06023_)
  );
  AND2_X1 _16151_ (
    .A1(_05738_),
    .A2(_06023_),
    .ZN(_06024_)
  );
  INV_X1 _16152_ (
    .A(_06024_),
    .ZN(_06025_)
  );
  AND2_X1 _16153_ (
    .A1(_05739_),
    .A2(_06022_),
    .ZN(_06026_)
  );
  INV_X1 _16154_ (
    .A(_06026_),
    .ZN(_06028_)
  );
  AND2_X1 _16155_ (
    .A1(_06025_),
    .A2(_06028_),
    .ZN(_06029_)
  );
  INV_X1 _16156_ (
    .A(_06029_),
    .ZN(_06030_)
  );
  AND2_X1 _16157_ (
    .A1(remainder[54]),
    .A2(_06029_),
    .ZN(_06031_)
  );
  INV_X1 _16158_ (
    .A(_06031_),
    .ZN(_06032_)
  );
  AND2_X1 _16159_ (
    .A1(_04525_),
    .A2(_06030_),
    .ZN(_06033_)
  );
  INV_X1 _16160_ (
    .A(_06033_),
    .ZN(_06034_)
  );
  AND2_X1 _16161_ (
    .A1(_06032_),
    .A2(_06034_),
    .ZN(_06035_)
  );
  INV_X1 _16162_ (
    .A(_06035_),
    .ZN(_06036_)
  );
  AND2_X1 _16163_ (
    .A1(_05737_),
    .A2(_06035_),
    .ZN(_06037_)
  );
  INV_X1 _16164_ (
    .A(_06037_),
    .ZN(_06039_)
  );
  AND2_X1 _16165_ (
    .A1(_05736_),
    .A2(_06036_),
    .ZN(_06040_)
  );
  INV_X1 _16166_ (
    .A(_06040_),
    .ZN(_06041_)
  );
  AND2_X1 _16167_ (
    .A1(_02082_),
    .A2(_06041_),
    .ZN(_06042_)
  );
  AND2_X1 _16168_ (
    .A1(_06039_),
    .A2(_06042_),
    .ZN(_06043_)
  );
  INV_X1 _16169_ (
    .A(_06043_),
    .ZN(_06044_)
  );
  AND2_X1 _16170_ (
    .A1(_05733_),
    .A2(_06044_),
    .ZN(_06045_)
  );
  AND2_X1 _16171_ (
    .A1(_05735_),
    .A2(_06045_),
    .ZN(_06046_)
  );
  INV_X1 _16172_ (
    .A(_06046_),
    .ZN(_06047_)
  );
  AND2_X1 _16173_ (
    .A1(_06201_),
    .A2(_06047_),
    .ZN(_00067_)
  );
  AND2_X1 _16174_ (
    .A1(_10462_),
    .A2(_01815_),
    .ZN(_06049_)
  );
  INV_X1 _16175_ (
    .A(_06049_),
    .ZN(_06050_)
  );
  AND2_X1 _16176_ (
    .A1(_04612_),
    .A2(_10451_),
    .ZN(_06051_)
  );
  INV_X1 _16177_ (
    .A(_06051_),
    .ZN(_06052_)
  );
  AND2_X1 _16178_ (
    .A1(_05983_),
    .A2(_06050_),
    .ZN(_06053_)
  );
  AND2_X1 _16179_ (
    .A1(_06052_),
    .A2(_06053_),
    .ZN(_06054_)
  );
  INV_X1 _16180_ (
    .A(_06054_),
    .ZN(_06055_)
  );
  AND2_X1 _16181_ (
    .A1(remainder[47]),
    .A2(_02077_),
    .ZN(_06056_)
  );
  INV_X1 _16182_ (
    .A(_06056_),
    .ZN(_06057_)
  );
  AND2_X1 _16183_ (
    .A1(_05999_),
    .A2(_06006_),
    .ZN(_06058_)
  );
  INV_X1 _16184_ (
    .A(_06058_),
    .ZN(_06060_)
  );
  AND2_X1 _16185_ (
    .A1(_05979_),
    .A2(_05986_),
    .ZN(_06061_)
  );
  INV_X1 _16186_ (
    .A(_06061_),
    .ZN(_06062_)
  );
  AND2_X1 _16187_ (
    .A1(_05922_),
    .A2(_05992_),
    .ZN(_06063_)
  );
  INV_X1 _16188_ (
    .A(_06063_),
    .ZN(_06064_)
  );
  AND2_X1 _16189_ (
    .A1(_03249_),
    .A2(_05902_),
    .ZN(_06065_)
  );
  INV_X1 _16190_ (
    .A(_06065_),
    .ZN(_06066_)
  );
  AND2_X1 _16191_ (
    .A1(_05561_),
    .A2(_06065_),
    .ZN(_06067_)
  );
  INV_X1 _16192_ (
    .A(_06067_),
    .ZN(_06068_)
  );
  AND2_X1 _16193_ (
    .A1(_05915_),
    .A2(_06068_),
    .ZN(_06069_)
  );
  INV_X1 _16194_ (
    .A(_06069_),
    .ZN(_06071_)
  );
  AND2_X1 _16195_ (
    .A1(_05455_),
    .A2(_05855_),
    .ZN(_06072_)
  );
  INV_X1 _16196_ (
    .A(_06072_),
    .ZN(_06073_)
  );
  AND2_X1 _16197_ (
    .A1(_05871_),
    .A2(_06073_),
    .ZN(_06074_)
  );
  INV_X1 _16198_ (
    .A(_06074_),
    .ZN(_06075_)
  );
  AND2_X1 _16199_ (
    .A1(_05449_),
    .A2(_05855_),
    .ZN(_06076_)
  );
  INV_X1 _16200_ (
    .A(_06076_),
    .ZN(_06077_)
  );
  AND2_X1 _16201_ (
    .A1(_05845_),
    .A2(_05852_),
    .ZN(_06078_)
  );
  INV_X1 _16202_ (
    .A(_06078_),
    .ZN(_06079_)
  );
  AND2_X1 _16203_ (
    .A1(_05832_),
    .A2(_05838_),
    .ZN(_06080_)
  );
  INV_X1 _16204_ (
    .A(_06080_),
    .ZN(_06082_)
  );
  AND2_X1 _16205_ (
    .A1(_05891_),
    .A2(_05898_),
    .ZN(_06083_)
  );
  INV_X1 _16206_ (
    .A(_06083_),
    .ZN(_06084_)
  );
  AND2_X1 _16207_ (
    .A1(divisor[16]),
    .A2(remainder[6]),
    .ZN(_06085_)
  );
  INV_X1 _16208_ (
    .A(_06085_),
    .ZN(_06086_)
  );
  AND2_X1 _16209_ (
    .A1(divisor[17]),
    .A2(remainder[5]),
    .ZN(_06087_)
  );
  INV_X1 _16210_ (
    .A(_06087_),
    .ZN(_06088_)
  );
  AND2_X1 _16211_ (
    .A1(divisor[18]),
    .A2(remainder[5]),
    .ZN(_06089_)
  );
  INV_X1 _16212_ (
    .A(_06089_),
    .ZN(_06090_)
  );
  AND2_X1 _16213_ (
    .A1(_05828_),
    .A2(_06087_),
    .ZN(_06091_)
  );
  INV_X1 _16214_ (
    .A(_06091_),
    .ZN(_06093_)
  );
  AND2_X1 _16215_ (
    .A1(_05830_),
    .A2(_06088_),
    .ZN(_06094_)
  );
  INV_X1 _16216_ (
    .A(_06094_),
    .ZN(_06095_)
  );
  AND2_X1 _16217_ (
    .A1(_06093_),
    .A2(_06095_),
    .ZN(_06096_)
  );
  INV_X1 _16218_ (
    .A(_06096_),
    .ZN(_06097_)
  );
  AND2_X1 _16219_ (
    .A1(_06085_),
    .A2(_06096_),
    .ZN(_06098_)
  );
  INV_X1 _16220_ (
    .A(_06098_),
    .ZN(_06099_)
  );
  AND2_X1 _16221_ (
    .A1(_06086_),
    .A2(_06097_),
    .ZN(_06100_)
  );
  INV_X1 _16222_ (
    .A(_06100_),
    .ZN(_06101_)
  );
  AND2_X1 _16223_ (
    .A1(_06099_),
    .A2(_06101_),
    .ZN(_06102_)
  );
  INV_X1 _16224_ (
    .A(_06102_),
    .ZN(_06104_)
  );
  AND2_X1 _16225_ (
    .A1(_06084_),
    .A2(_06102_),
    .ZN(_06105_)
  );
  INV_X1 _16226_ (
    .A(_06105_),
    .ZN(_06106_)
  );
  AND2_X1 _16227_ (
    .A1(_06083_),
    .A2(_06104_),
    .ZN(_06107_)
  );
  INV_X1 _16228_ (
    .A(_06107_),
    .ZN(_06108_)
  );
  AND2_X1 _16229_ (
    .A1(_06106_),
    .A2(_06108_),
    .ZN(_06109_)
  );
  INV_X1 _16230_ (
    .A(_06109_),
    .ZN(_06110_)
  );
  AND2_X1 _16231_ (
    .A1(_06082_),
    .A2(_06109_),
    .ZN(_06111_)
  );
  INV_X1 _16232_ (
    .A(_06111_),
    .ZN(_06112_)
  );
  AND2_X1 _16233_ (
    .A1(_06080_),
    .A2(_06110_),
    .ZN(_06113_)
  );
  INV_X1 _16234_ (
    .A(_06113_),
    .ZN(_06115_)
  );
  AND2_X1 _16235_ (
    .A1(_06112_),
    .A2(_06115_),
    .ZN(_06116_)
  );
  INV_X1 _16236_ (
    .A(_06116_),
    .ZN(_06117_)
  );
  AND2_X1 _16237_ (
    .A1(_06079_),
    .A2(_06116_),
    .ZN(_06118_)
  );
  INV_X1 _16238_ (
    .A(_06118_),
    .ZN(_06119_)
  );
  AND2_X1 _16239_ (
    .A1(_06078_),
    .A2(_06117_),
    .ZN(_06120_)
  );
  INV_X1 _16240_ (
    .A(_06120_),
    .ZN(_06121_)
  );
  AND2_X1 _16241_ (
    .A1(_06119_),
    .A2(_06121_),
    .ZN(_06122_)
  );
  INV_X1 _16242_ (
    .A(_06122_),
    .ZN(_06123_)
  );
  AND2_X1 _16243_ (
    .A1(_06076_),
    .A2(_06122_),
    .ZN(_06124_)
  );
  INV_X1 _16244_ (
    .A(_06124_),
    .ZN(_06126_)
  );
  AND2_X1 _16245_ (
    .A1(_06077_),
    .A2(_06123_),
    .ZN(_06127_)
  );
  INV_X1 _16246_ (
    .A(_06127_),
    .ZN(_06128_)
  );
  AND2_X1 _16247_ (
    .A1(_06126_),
    .A2(_06128_),
    .ZN(_06129_)
  );
  INV_X1 _16248_ (
    .A(_06129_),
    .ZN(_06130_)
  );
  AND2_X1 _16249_ (
    .A1(_05781_),
    .A2(_05788_),
    .ZN(_06131_)
  );
  INV_X1 _16250_ (
    .A(_06131_),
    .ZN(_06132_)
  );
  AND2_X1 _16251_ (
    .A1(_05768_),
    .A2(_05775_),
    .ZN(_06133_)
  );
  INV_X1 _16252_ (
    .A(_06133_),
    .ZN(_06134_)
  );
  AND2_X1 _16253_ (
    .A1(remainder[32]),
    .A2(divisor[15]),
    .ZN(_06135_)
  );
  INV_X1 _16254_ (
    .A(_06135_),
    .ZN(_06137_)
  );
  AND2_X1 _16255_ (
    .A1(remainder[32]),
    .A2(divisor[14]),
    .ZN(_06138_)
  );
  INV_X1 _16256_ (
    .A(_06138_),
    .ZN(_06139_)
  );
  AND2_X1 _16257_ (
    .A1(_05765_),
    .A2(_06138_),
    .ZN(_06140_)
  );
  INV_X1 _16258_ (
    .A(_06140_),
    .ZN(_06141_)
  );
  AND2_X1 _16259_ (
    .A1(_05766_),
    .A2(_06139_),
    .ZN(_06142_)
  );
  INV_X1 _16260_ (
    .A(_06142_),
    .ZN(_06143_)
  );
  AND2_X1 _16261_ (
    .A1(_06141_),
    .A2(_06143_),
    .ZN(_06144_)
  );
  INV_X1 _16262_ (
    .A(_06144_),
    .ZN(_06145_)
  );
  AND2_X1 _16263_ (
    .A1(_05760_),
    .A2(_06144_),
    .ZN(_06146_)
  );
  INV_X1 _16264_ (
    .A(_06146_),
    .ZN(_06148_)
  );
  AND2_X1 _16265_ (
    .A1(_05761_),
    .A2(_06145_),
    .ZN(_06149_)
  );
  INV_X1 _16266_ (
    .A(_06149_),
    .ZN(_06150_)
  );
  AND2_X1 _16267_ (
    .A1(_06148_),
    .A2(_06150_),
    .ZN(_06151_)
  );
  INV_X1 _16268_ (
    .A(_06151_),
    .ZN(_06152_)
  );
  AND2_X1 _16269_ (
    .A1(_06134_),
    .A2(_06151_),
    .ZN(_06153_)
  );
  INV_X1 _16270_ (
    .A(_06153_),
    .ZN(_06154_)
  );
  AND2_X1 _16271_ (
    .A1(_06133_),
    .A2(_06152_),
    .ZN(_06155_)
  );
  INV_X1 _16272_ (
    .A(_06155_),
    .ZN(_06156_)
  );
  AND2_X1 _16273_ (
    .A1(_06154_),
    .A2(_06156_),
    .ZN(_06157_)
  );
  INV_X1 _16274_ (
    .A(_06157_),
    .ZN(_06159_)
  );
  AND2_X1 _16275_ (
    .A1(_05499_),
    .A2(_06157_),
    .ZN(_06160_)
  );
  INV_X1 _16276_ (
    .A(_06160_),
    .ZN(_06161_)
  );
  AND2_X1 _16277_ (
    .A1(_05501_),
    .A2(_06159_),
    .ZN(_06162_)
  );
  INV_X1 _16278_ (
    .A(_06162_),
    .ZN(_06163_)
  );
  AND2_X1 _16279_ (
    .A1(_06161_),
    .A2(_06163_),
    .ZN(_06164_)
  );
  INV_X1 _16280_ (
    .A(_06164_),
    .ZN(_06165_)
  );
  AND2_X1 _16281_ (
    .A1(_06132_),
    .A2(_06164_),
    .ZN(_06166_)
  );
  INV_X1 _16282_ (
    .A(_06166_),
    .ZN(_06167_)
  );
  AND2_X1 _16283_ (
    .A1(_06131_),
    .A2(_06165_),
    .ZN(_06168_)
  );
  INV_X1 _16284_ (
    .A(_06168_),
    .ZN(_06170_)
  );
  AND2_X1 _16285_ (
    .A1(_06167_),
    .A2(_06170_),
    .ZN(_06171_)
  );
  INV_X1 _16286_ (
    .A(_06171_),
    .ZN(_06172_)
  );
  AND2_X1 _16287_ (
    .A1(_05813_),
    .A2(_06171_),
    .ZN(_06173_)
  );
  INV_X1 _16288_ (
    .A(_06173_),
    .ZN(_06174_)
  );
  AND2_X1 _16289_ (
    .A1(_05814_),
    .A2(_06172_),
    .ZN(_06175_)
  );
  INV_X1 _16290_ (
    .A(_06175_),
    .ZN(_06176_)
  );
  AND2_X1 _16291_ (
    .A1(_06174_),
    .A2(_06176_),
    .ZN(_06177_)
  );
  INV_X1 _16292_ (
    .A(_06177_),
    .ZN(_06178_)
  );
  AND2_X1 _16293_ (
    .A1(_06129_),
    .A2(_06177_),
    .ZN(_06179_)
  );
  INV_X1 _16294_ (
    .A(_06179_),
    .ZN(_06180_)
  );
  AND2_X1 _16295_ (
    .A1(_06130_),
    .A2(_06178_),
    .ZN(_06181_)
  );
  INV_X1 _16296_ (
    .A(_06181_),
    .ZN(_06182_)
  );
  AND2_X1 _16297_ (
    .A1(_06180_),
    .A2(_06182_),
    .ZN(_06183_)
  );
  INV_X1 _16298_ (
    .A(_06183_),
    .ZN(_06184_)
  );
  AND2_X1 _16299_ (
    .A1(_06075_),
    .A2(_06183_),
    .ZN(_06185_)
  );
  INV_X1 _16300_ (
    .A(_06185_),
    .ZN(_06186_)
  );
  AND2_X1 _16301_ (
    .A1(_06074_),
    .A2(_06184_),
    .ZN(_06187_)
  );
  INV_X1 _16302_ (
    .A(_06187_),
    .ZN(_06188_)
  );
  AND2_X1 _16303_ (
    .A1(_06186_),
    .A2(_06188_),
    .ZN(_06189_)
  );
  INV_X1 _16304_ (
    .A(_06189_),
    .ZN(_06191_)
  );
  AND2_X1 _16305_ (
    .A1(divisor[22]),
    .A2(remainder[0]),
    .ZN(_06192_)
  );
  INV_X1 _16306_ (
    .A(_06192_),
    .ZN(_06193_)
  );
  AND2_X1 _16307_ (
    .A1(divisor[19]),
    .A2(remainder[3]),
    .ZN(_06194_)
  );
  INV_X1 _16308_ (
    .A(_06194_),
    .ZN(_06195_)
  );
  AND2_X1 _16309_ (
    .A1(divisor[20]),
    .A2(remainder[2]),
    .ZN(_06196_)
  );
  INV_X1 _16310_ (
    .A(_06196_),
    .ZN(_06197_)
  );
  AND2_X1 _16311_ (
    .A1(divisor[21]),
    .A2(remainder[2]),
    .ZN(_06198_)
  );
  INV_X1 _16312_ (
    .A(_06198_),
    .ZN(_06199_)
  );
  AND2_X1 _16313_ (
    .A1(_05554_),
    .A2(_06198_),
    .ZN(_06200_)
  );
  INV_X1 _16314_ (
    .A(_06200_),
    .ZN(_06202_)
  );
  AND2_X1 _16315_ (
    .A1(_05889_),
    .A2(_06197_),
    .ZN(_06203_)
  );
  INV_X1 _16316_ (
    .A(_06203_),
    .ZN(_06204_)
  );
  AND2_X1 _16317_ (
    .A1(_06202_),
    .A2(_06204_),
    .ZN(_06205_)
  );
  INV_X1 _16318_ (
    .A(_06205_),
    .ZN(_06206_)
  );
  AND2_X1 _16319_ (
    .A1(_06194_),
    .A2(_06205_),
    .ZN(_06207_)
  );
  INV_X1 _16320_ (
    .A(_06207_),
    .ZN(_06208_)
  );
  AND2_X1 _16321_ (
    .A1(_06195_),
    .A2(_06206_),
    .ZN(_06209_)
  );
  INV_X1 _16322_ (
    .A(_06209_),
    .ZN(_06210_)
  );
  AND2_X1 _16323_ (
    .A1(_06208_),
    .A2(_06210_),
    .ZN(_06211_)
  );
  INV_X1 _16324_ (
    .A(_06211_),
    .ZN(_06213_)
  );
  AND2_X1 _16325_ (
    .A1(_06192_),
    .A2(_06211_),
    .ZN(_06214_)
  );
  INV_X1 _16326_ (
    .A(_06214_),
    .ZN(_06215_)
  );
  AND2_X1 _16327_ (
    .A1(_06193_),
    .A2(_06213_),
    .ZN(_06216_)
  );
  INV_X1 _16328_ (
    .A(_06216_),
    .ZN(_06217_)
  );
  AND2_X1 _16329_ (
    .A1(_06215_),
    .A2(_06217_),
    .ZN(_06218_)
  );
  INV_X1 _16330_ (
    .A(_06218_),
    .ZN(_06219_)
  );
  AND2_X1 _16331_ (
    .A1(_06066_),
    .A2(_06219_),
    .ZN(_06220_)
  );
  INV_X1 _16332_ (
    .A(_06220_),
    .ZN(_06221_)
  );
  AND2_X1 _16333_ (
    .A1(_06065_),
    .A2(_06218_),
    .ZN(_06222_)
  );
  INV_X1 _16334_ (
    .A(_06222_),
    .ZN(_06224_)
  );
  AND2_X1 _16335_ (
    .A1(_06065_),
    .A2(_06219_),
    .ZN(_06225_)
  );
  INV_X1 _16336_ (
    .A(_06225_),
    .ZN(_06226_)
  );
  AND2_X1 _16337_ (
    .A1(_06066_),
    .A2(_06218_),
    .ZN(_06227_)
  );
  INV_X1 _16338_ (
    .A(_06227_),
    .ZN(_06228_)
  );
  AND2_X1 _16339_ (
    .A1(_06221_),
    .A2(_06224_),
    .ZN(_06229_)
  );
  AND2_X1 _16340_ (
    .A1(_06226_),
    .A2(_06228_),
    .ZN(_06230_)
  );
  AND2_X1 _16341_ (
    .A1(_06189_),
    .A2(_06229_),
    .ZN(_06231_)
  );
  INV_X1 _16342_ (
    .A(_06231_),
    .ZN(_06232_)
  );
  AND2_X1 _16343_ (
    .A1(_06191_),
    .A2(_06230_),
    .ZN(_06233_)
  );
  INV_X1 _16344_ (
    .A(_06233_),
    .ZN(_06235_)
  );
  AND2_X1 _16345_ (
    .A1(_06232_),
    .A2(_06235_),
    .ZN(_06236_)
  );
  INV_X1 _16346_ (
    .A(_06236_),
    .ZN(_06237_)
  );
  AND2_X1 _16347_ (
    .A1(_06071_),
    .A2(_06236_),
    .ZN(_06238_)
  );
  INV_X1 _16348_ (
    .A(_06238_),
    .ZN(_06239_)
  );
  AND2_X1 _16349_ (
    .A1(_06069_),
    .A2(_06237_),
    .ZN(_06240_)
  );
  INV_X1 _16350_ (
    .A(_06240_),
    .ZN(_06241_)
  );
  AND2_X1 _16351_ (
    .A1(_06239_),
    .A2(_06241_),
    .ZN(_06242_)
  );
  INV_X1 _16352_ (
    .A(_06242_),
    .ZN(_06243_)
  );
  AND2_X1 _16353_ (
    .A1(_05966_),
    .A2(_05973_),
    .ZN(_06244_)
  );
  INV_X1 _16354_ (
    .A(_06244_),
    .ZN(_06246_)
  );
  AND2_X1 _16355_ (
    .A1(_05953_),
    .A2(_05959_),
    .ZN(_06247_)
  );
  INV_X1 _16356_ (
    .A(_06247_),
    .ZN(_06248_)
  );
  AND2_X1 _16357_ (
    .A1(_05940_),
    .A2(_05946_),
    .ZN(_06249_)
  );
  INV_X1 _16358_ (
    .A(_06249_),
    .ZN(_06250_)
  );
  AND2_X1 _16359_ (
    .A1(_05794_),
    .A2(_05816_),
    .ZN(_06251_)
  );
  INV_X1 _16360_ (
    .A(_06251_),
    .ZN(_06252_)
  );
  AND2_X1 _16361_ (
    .A1(_05803_),
    .A2(_05810_),
    .ZN(_06253_)
  );
  INV_X1 _16362_ (
    .A(_06253_),
    .ZN(_06254_)
  );
  AND2_X1 _16363_ (
    .A1(_04087_),
    .A2(_06254_),
    .ZN(_06255_)
  );
  INV_X1 _16364_ (
    .A(_06255_),
    .ZN(_06257_)
  );
  AND2_X1 _16365_ (
    .A1(_04088_),
    .A2(_06253_),
    .ZN(_06258_)
  );
  INV_X1 _16366_ (
    .A(_06258_),
    .ZN(_06259_)
  );
  AND2_X1 _16367_ (
    .A1(_06257_),
    .A2(_06259_),
    .ZN(_06260_)
  );
  INV_X1 _16368_ (
    .A(_06260_),
    .ZN(_06261_)
  );
  AND2_X1 _16369_ (
    .A1(_04317_),
    .A2(_06260_),
    .ZN(_06262_)
  );
  INV_X1 _16370_ (
    .A(_06262_),
    .ZN(_06263_)
  );
  AND2_X1 _16371_ (
    .A1(_04316_),
    .A2(_06261_),
    .ZN(_06264_)
  );
  INV_X1 _16372_ (
    .A(_06264_),
    .ZN(_06265_)
  );
  AND2_X1 _16373_ (
    .A1(_06263_),
    .A2(_06265_),
    .ZN(_06266_)
  );
  INV_X1 _16374_ (
    .A(_06266_),
    .ZN(_06268_)
  );
  AND2_X1 _16375_ (
    .A1(_06252_),
    .A2(_06266_),
    .ZN(_06269_)
  );
  INV_X1 _16376_ (
    .A(_06269_),
    .ZN(_06270_)
  );
  AND2_X1 _16377_ (
    .A1(_06251_),
    .A2(_06268_),
    .ZN(_06271_)
  );
  INV_X1 _16378_ (
    .A(_06271_),
    .ZN(_06272_)
  );
  AND2_X1 _16379_ (
    .A1(_06270_),
    .A2(_06272_),
    .ZN(_06273_)
  );
  INV_X1 _16380_ (
    .A(_06273_),
    .ZN(_06274_)
  );
  AND2_X1 _16381_ (
    .A1(_06250_),
    .A2(_06273_),
    .ZN(_06275_)
  );
  INV_X1 _16382_ (
    .A(_06275_),
    .ZN(_06276_)
  );
  AND2_X1 _16383_ (
    .A1(_06249_),
    .A2(_06274_),
    .ZN(_06277_)
  );
  INV_X1 _16384_ (
    .A(_06277_),
    .ZN(_06279_)
  );
  AND2_X1 _16385_ (
    .A1(_06276_),
    .A2(_06279_),
    .ZN(_06280_)
  );
  INV_X1 _16386_ (
    .A(_06280_),
    .ZN(_06281_)
  );
  AND2_X1 _16387_ (
    .A1(_06248_),
    .A2(_06280_),
    .ZN(_06282_)
  );
  INV_X1 _16388_ (
    .A(_06282_),
    .ZN(_06283_)
  );
  AND2_X1 _16389_ (
    .A1(_06247_),
    .A2(_06281_),
    .ZN(_06284_)
  );
  INV_X1 _16390_ (
    .A(_06284_),
    .ZN(_06285_)
  );
  AND2_X1 _16391_ (
    .A1(_06283_),
    .A2(_06285_),
    .ZN(_06286_)
  );
  INV_X1 _16392_ (
    .A(_06286_),
    .ZN(_06287_)
  );
  AND2_X1 _16393_ (
    .A1(_03170_),
    .A2(_06286_),
    .ZN(_06288_)
  );
  INV_X1 _16394_ (
    .A(_06288_),
    .ZN(_06289_)
  );
  AND2_X1 _16395_ (
    .A1(_03169_),
    .A2(_06287_),
    .ZN(_06290_)
  );
  INV_X1 _16396_ (
    .A(_06290_),
    .ZN(_06291_)
  );
  AND2_X1 _16397_ (
    .A1(_06289_),
    .A2(_06291_),
    .ZN(_06292_)
  );
  INV_X1 _16398_ (
    .A(_06292_),
    .ZN(_06293_)
  );
  AND2_X1 _16399_ (
    .A1(_05877_),
    .A2(_06292_),
    .ZN(_06294_)
  );
  INV_X1 _16400_ (
    .A(_06294_),
    .ZN(_06295_)
  );
  AND2_X1 _16401_ (
    .A1(_05878_),
    .A2(_06293_),
    .ZN(_06296_)
  );
  INV_X1 _16402_ (
    .A(_06296_),
    .ZN(_06297_)
  );
  AND2_X1 _16403_ (
    .A1(_06295_),
    .A2(_06297_),
    .ZN(_06298_)
  );
  INV_X1 _16404_ (
    .A(_06298_),
    .ZN(_06300_)
  );
  AND2_X1 _16405_ (
    .A1(_06246_),
    .A2(_06298_),
    .ZN(_06301_)
  );
  INV_X1 _16406_ (
    .A(_06301_),
    .ZN(_06302_)
  );
  AND2_X1 _16407_ (
    .A1(_06244_),
    .A2(_06300_),
    .ZN(_06303_)
  );
  INV_X1 _16408_ (
    .A(_06303_),
    .ZN(_06304_)
  );
  AND2_X1 _16409_ (
    .A1(_06302_),
    .A2(_06304_),
    .ZN(_06305_)
  );
  INV_X1 _16410_ (
    .A(_06305_),
    .ZN(_06306_)
  );
  AND2_X1 _16411_ (
    .A1(_06242_),
    .A2(_06305_),
    .ZN(_06307_)
  );
  INV_X1 _16412_ (
    .A(_06307_),
    .ZN(_06308_)
  );
  AND2_X1 _16413_ (
    .A1(_06243_),
    .A2(_06306_),
    .ZN(_06309_)
  );
  INV_X1 _16414_ (
    .A(_06309_),
    .ZN(_06311_)
  );
  AND2_X1 _16415_ (
    .A1(_06308_),
    .A2(_06311_),
    .ZN(_06312_)
  );
  INV_X1 _16416_ (
    .A(_06312_),
    .ZN(_06313_)
  );
  AND2_X1 _16417_ (
    .A1(_06064_),
    .A2(_06312_),
    .ZN(_06314_)
  );
  INV_X1 _16418_ (
    .A(_06314_),
    .ZN(_06315_)
  );
  AND2_X1 _16419_ (
    .A1(_06063_),
    .A2(_06313_),
    .ZN(_06316_)
  );
  INV_X1 _16420_ (
    .A(_06316_),
    .ZN(_06317_)
  );
  AND2_X1 _16421_ (
    .A1(_06315_),
    .A2(_06317_),
    .ZN(_06318_)
  );
  INV_X1 _16422_ (
    .A(_06318_),
    .ZN(_06319_)
  );
  AND2_X1 _16423_ (
    .A1(_06062_),
    .A2(_06318_),
    .ZN(_06320_)
  );
  INV_X1 _16424_ (
    .A(_06320_),
    .ZN(_06322_)
  );
  AND2_X1 _16425_ (
    .A1(_06061_),
    .A2(_06319_),
    .ZN(_06323_)
  );
  INV_X1 _16426_ (
    .A(_06323_),
    .ZN(_06324_)
  );
  AND2_X1 _16427_ (
    .A1(_06322_),
    .A2(_06324_),
    .ZN(_06325_)
  );
  INV_X1 _16428_ (
    .A(_06325_),
    .ZN(_06326_)
  );
  AND2_X1 _16429_ (
    .A1(_06060_),
    .A2(_06325_),
    .ZN(_06327_)
  );
  INV_X1 _16430_ (
    .A(_06327_),
    .ZN(_06328_)
  );
  AND2_X1 _16431_ (
    .A1(_06058_),
    .A2(_06326_),
    .ZN(_06329_)
  );
  INV_X1 _16432_ (
    .A(_06329_),
    .ZN(_06330_)
  );
  AND2_X1 _16433_ (
    .A1(_06328_),
    .A2(_06330_),
    .ZN(_06331_)
  );
  INV_X1 _16434_ (
    .A(_06331_),
    .ZN(_06333_)
  );
  AND2_X1 _16435_ (
    .A1(_06011_),
    .A2(_06331_),
    .ZN(_06334_)
  );
  INV_X1 _16436_ (
    .A(_06334_),
    .ZN(_06335_)
  );
  AND2_X1 _16437_ (
    .A1(_06012_),
    .A2(_06333_),
    .ZN(_06336_)
  );
  INV_X1 _16438_ (
    .A(_06336_),
    .ZN(_06337_)
  );
  AND2_X1 _16439_ (
    .A1(_06335_),
    .A2(_06337_),
    .ZN(_06338_)
  );
  INV_X1 _16440_ (
    .A(_06338_),
    .ZN(_06339_)
  );
  AND2_X1 _16441_ (
    .A1(_05738_),
    .A2(_06019_),
    .ZN(_06340_)
  );
  INV_X1 _16442_ (
    .A(_06340_),
    .ZN(_06341_)
  );
  AND2_X1 _16443_ (
    .A1(_06019_),
    .A2(_06028_),
    .ZN(_06342_)
  );
  AND2_X1 _16444_ (
    .A1(_06021_),
    .A2(_06341_),
    .ZN(_06344_)
  );
  AND2_X1 _16445_ (
    .A1(_06338_),
    .A2(_06344_),
    .ZN(_06345_)
  );
  INV_X1 _16446_ (
    .A(_06345_),
    .ZN(_06346_)
  );
  AND2_X1 _16447_ (
    .A1(_06339_),
    .A2(_06342_),
    .ZN(_06347_)
  );
  INV_X1 _16448_ (
    .A(_06347_),
    .ZN(_06348_)
  );
  AND2_X1 _16449_ (
    .A1(_06346_),
    .A2(_06348_),
    .ZN(_06349_)
  );
  INV_X1 _16450_ (
    .A(_06349_),
    .ZN(_06350_)
  );
  AND2_X1 _16451_ (
    .A1(remainder[55]),
    .A2(_06349_),
    .ZN(_06351_)
  );
  INV_X1 _16452_ (
    .A(_06351_),
    .ZN(_06352_)
  );
  AND2_X1 _16453_ (
    .A1(_04514_),
    .A2(_06350_),
    .ZN(_06353_)
  );
  INV_X1 _16454_ (
    .A(_06353_),
    .ZN(_06355_)
  );
  AND2_X1 _16455_ (
    .A1(_06352_),
    .A2(_06355_),
    .ZN(_06356_)
  );
  INV_X1 _16456_ (
    .A(_06356_),
    .ZN(_06357_)
  );
  AND2_X1 _16457_ (
    .A1(_05736_),
    .A2(_06032_),
    .ZN(_06358_)
  );
  INV_X1 _16458_ (
    .A(_06358_),
    .ZN(_06359_)
  );
  AND2_X1 _16459_ (
    .A1(_05737_),
    .A2(_06034_),
    .ZN(_06360_)
  );
  INV_X1 _16460_ (
    .A(_06360_),
    .ZN(_06361_)
  );
  AND2_X1 _16461_ (
    .A1(_06034_),
    .A2(_06359_),
    .ZN(_06362_)
  );
  AND2_X1 _16462_ (
    .A1(_06032_),
    .A2(_06361_),
    .ZN(_06363_)
  );
  AND2_X1 _16463_ (
    .A1(_06357_),
    .A2(_06363_),
    .ZN(_06364_)
  );
  INV_X1 _16464_ (
    .A(_06364_),
    .ZN(_06366_)
  );
  AND2_X1 _16465_ (
    .A1(_06356_),
    .A2(_06362_),
    .ZN(_06367_)
  );
  INV_X1 _16466_ (
    .A(_06367_),
    .ZN(_06368_)
  );
  AND2_X1 _16467_ (
    .A1(_02082_),
    .A2(_06368_),
    .ZN(_06369_)
  );
  AND2_X1 _16468_ (
    .A1(_06366_),
    .A2(_06369_),
    .ZN(_06370_)
  );
  INV_X1 _16469_ (
    .A(_06370_),
    .ZN(_06371_)
  );
  AND2_X1 _16470_ (
    .A1(_06055_),
    .A2(_06371_),
    .ZN(_06372_)
  );
  AND2_X1 _16471_ (
    .A1(_06057_),
    .A2(_06372_),
    .ZN(_06373_)
  );
  INV_X1 _16472_ (
    .A(_06373_),
    .ZN(_06374_)
  );
  AND2_X1 _16473_ (
    .A1(_06201_),
    .A2(_06374_),
    .ZN(_00068_)
  );
  AND2_X1 _16474_ (
    .A1(_04601_),
    .A2(_10451_),
    .ZN(_06376_)
  );
  INV_X1 _16475_ (
    .A(_06376_),
    .ZN(_06377_)
  );
  AND2_X1 _16476_ (
    .A1(_10462_),
    .A2(_01834_),
    .ZN(_06378_)
  );
  INV_X1 _16477_ (
    .A(_06378_),
    .ZN(_06379_)
  );
  AND2_X1 _16478_ (
    .A1(_05983_),
    .A2(_06379_),
    .ZN(_06380_)
  );
  AND2_X1 _16479_ (
    .A1(_06377_),
    .A2(_06380_),
    .ZN(_06381_)
  );
  INV_X1 _16480_ (
    .A(_06381_),
    .ZN(_06382_)
  );
  AND2_X1 _16481_ (
    .A1(remainder[48]),
    .A2(_02077_),
    .ZN(_06383_)
  );
  INV_X1 _16482_ (
    .A(_06383_),
    .ZN(_06384_)
  );
  AND2_X1 _16483_ (
    .A1(_06352_),
    .A2(_06368_),
    .ZN(_06385_)
  );
  INV_X1 _16484_ (
    .A(_06385_),
    .ZN(_06387_)
  );
  AND2_X1 _16485_ (
    .A1(_06335_),
    .A2(_06346_),
    .ZN(_06388_)
  );
  INV_X1 _16486_ (
    .A(_06388_),
    .ZN(_06389_)
  );
  AND2_X1 _16487_ (
    .A1(_06315_),
    .A2(_06322_),
    .ZN(_06390_)
  );
  INV_X1 _16488_ (
    .A(_06390_),
    .ZN(_06391_)
  );
  AND2_X1 _16489_ (
    .A1(_06295_),
    .A2(_06302_),
    .ZN(_06392_)
  );
  INV_X1 _16490_ (
    .A(_06392_),
    .ZN(_06393_)
  );
  AND2_X1 _16491_ (
    .A1(_06239_),
    .A2(_06308_),
    .ZN(_06394_)
  );
  INV_X1 _16492_ (
    .A(_06394_),
    .ZN(_06395_)
  );
  AND2_X1 _16493_ (
    .A1(_03249_),
    .A2(_06219_),
    .ZN(_06396_)
  );
  INV_X1 _16494_ (
    .A(_06396_),
    .ZN(_06398_)
  );
  AND2_X1 _16495_ (
    .A1(_05901_),
    .A2(_06396_),
    .ZN(_06399_)
  );
  INV_X1 _16496_ (
    .A(_06399_),
    .ZN(_06400_)
  );
  AND2_X1 _16497_ (
    .A1(_06232_),
    .A2(_06400_),
    .ZN(_06401_)
  );
  INV_X1 _16498_ (
    .A(_06401_),
    .ZN(_06402_)
  );
  AND2_X1 _16499_ (
    .A1(_06126_),
    .A2(_06180_),
    .ZN(_06403_)
  );
  INV_X1 _16500_ (
    .A(_06403_),
    .ZN(_06404_)
  );
  AND2_X1 _16501_ (
    .A1(_06154_),
    .A2(_06161_),
    .ZN(_06405_)
  );
  INV_X1 _16502_ (
    .A(_06405_),
    .ZN(_06406_)
  );
  AND2_X1 _16503_ (
    .A1(_06141_),
    .A2(_06148_),
    .ZN(_06407_)
  );
  INV_X1 _16504_ (
    .A(_06407_),
    .ZN(_06409_)
  );
  AND2_X1 _16505_ (
    .A1(_06137_),
    .A2(_06139_),
    .ZN(_06410_)
  );
  MUX2_X1 _16506_ (
    .A(_06138_),
    .B(_04952_),
    .S(_06135_),
    .Z(_06411_)
  );
  MUX2_X1 _16507_ (
    .A(_05760_),
    .B(_04941_),
    .S(_06411_),
    .Z(_06412_)
  );
  MUX2_X1 _16508_ (
    .A(_05761_),
    .B(divisor[13]),
    .S(_06411_),
    .Z(_06413_)
  );
  AND2_X1 _16509_ (
    .A1(_06409_),
    .A2(_06412_),
    .ZN(_06414_)
  );
  INV_X1 _16510_ (
    .A(_06414_),
    .ZN(_06415_)
  );
  AND2_X1 _16511_ (
    .A1(_06407_),
    .A2(_06413_),
    .ZN(_06416_)
  );
  INV_X1 _16512_ (
    .A(_06416_),
    .ZN(_06417_)
  );
  AND2_X1 _16513_ (
    .A1(_06415_),
    .A2(_06417_),
    .ZN(_06418_)
  );
  INV_X1 _16514_ (
    .A(_06418_),
    .ZN(_06419_)
  );
  AND2_X1 _16515_ (
    .A1(_05499_),
    .A2(_06419_),
    .ZN(_06420_)
  );
  INV_X1 _16516_ (
    .A(_06420_),
    .ZN(_06421_)
  );
  AND2_X1 _16517_ (
    .A1(_05501_),
    .A2(_06418_),
    .ZN(_06422_)
  );
  INV_X1 _16518_ (
    .A(_06422_),
    .ZN(_06423_)
  );
  AND2_X1 _16519_ (
    .A1(_05499_),
    .A2(_06417_),
    .ZN(_06424_)
  );
  AND2_X1 _16520_ (
    .A1(_06421_),
    .A2(_06423_),
    .ZN(_06425_)
  );
  INV_X1 _16521_ (
    .A(_06425_),
    .ZN(_06426_)
  );
  AND2_X1 _16522_ (
    .A1(_06406_),
    .A2(_06426_),
    .ZN(_06427_)
  );
  INV_X1 _16523_ (
    .A(_06427_),
    .ZN(_06428_)
  );
  AND2_X1 _16524_ (
    .A1(_06405_),
    .A2(_06425_),
    .ZN(_06430_)
  );
  INV_X1 _16525_ (
    .A(_06430_),
    .ZN(_06431_)
  );
  AND2_X1 _16526_ (
    .A1(_06428_),
    .A2(_06431_),
    .ZN(_06432_)
  );
  INV_X1 _16527_ (
    .A(_06432_),
    .ZN(_06433_)
  );
  AND2_X1 _16528_ (
    .A1(_05813_),
    .A2(_06432_),
    .ZN(_06434_)
  );
  INV_X1 _16529_ (
    .A(_06434_),
    .ZN(_06435_)
  );
  AND2_X1 _16530_ (
    .A1(_05814_),
    .A2(_06433_),
    .ZN(_06436_)
  );
  INV_X1 _16531_ (
    .A(_06436_),
    .ZN(_06437_)
  );
  AND2_X1 _16532_ (
    .A1(_06435_),
    .A2(_06437_),
    .ZN(_06438_)
  );
  INV_X1 _16533_ (
    .A(_06438_),
    .ZN(_06439_)
  );
  AND2_X1 _16534_ (
    .A1(_06106_),
    .A2(_06112_),
    .ZN(_06441_)
  );
  INV_X1 _16535_ (
    .A(_06441_),
    .ZN(_06442_)
  );
  AND2_X1 _16536_ (
    .A1(_06093_),
    .A2(_06099_),
    .ZN(_06443_)
  );
  INV_X1 _16537_ (
    .A(_06443_),
    .ZN(_06444_)
  );
  AND2_X1 _16538_ (
    .A1(_06202_),
    .A2(_06208_),
    .ZN(_06445_)
  );
  INV_X1 _16539_ (
    .A(_06445_),
    .ZN(_06446_)
  );
  AND2_X1 _16540_ (
    .A1(divisor[16]),
    .A2(remainder[7]),
    .ZN(_06447_)
  );
  INV_X1 _16541_ (
    .A(_06447_),
    .ZN(_06448_)
  );
  AND2_X1 _16542_ (
    .A1(divisor[17]),
    .A2(remainder[6]),
    .ZN(_06449_)
  );
  INV_X1 _16543_ (
    .A(_06449_),
    .ZN(_06450_)
  );
  AND2_X1 _16544_ (
    .A1(divisor[18]),
    .A2(remainder[6]),
    .ZN(_06452_)
  );
  INV_X1 _16545_ (
    .A(_06452_),
    .ZN(_06453_)
  );
  AND2_X1 _16546_ (
    .A1(_06089_),
    .A2(_06449_),
    .ZN(_06454_)
  );
  INV_X1 _16547_ (
    .A(_06454_),
    .ZN(_06455_)
  );
  AND2_X1 _16548_ (
    .A1(_06090_),
    .A2(_06450_),
    .ZN(_06456_)
  );
  INV_X1 _16549_ (
    .A(_06456_),
    .ZN(_06457_)
  );
  AND2_X1 _16550_ (
    .A1(_06455_),
    .A2(_06457_),
    .ZN(_06458_)
  );
  INV_X1 _16551_ (
    .A(_06458_),
    .ZN(_06459_)
  );
  AND2_X1 _16552_ (
    .A1(_06447_),
    .A2(_06458_),
    .ZN(_06460_)
  );
  INV_X1 _16553_ (
    .A(_06460_),
    .ZN(_06461_)
  );
  AND2_X1 _16554_ (
    .A1(_06448_),
    .A2(_06459_),
    .ZN(_06463_)
  );
  INV_X1 _16555_ (
    .A(_06463_),
    .ZN(_06464_)
  );
  AND2_X1 _16556_ (
    .A1(_06461_),
    .A2(_06464_),
    .ZN(_06465_)
  );
  INV_X1 _16557_ (
    .A(_06465_),
    .ZN(_06466_)
  );
  AND2_X1 _16558_ (
    .A1(_06446_),
    .A2(_06465_),
    .ZN(_06467_)
  );
  INV_X1 _16559_ (
    .A(_06467_),
    .ZN(_06468_)
  );
  AND2_X1 _16560_ (
    .A1(_06445_),
    .A2(_06466_),
    .ZN(_06469_)
  );
  INV_X1 _16561_ (
    .A(_06469_),
    .ZN(_06470_)
  );
  AND2_X1 _16562_ (
    .A1(_06468_),
    .A2(_06470_),
    .ZN(_06471_)
  );
  INV_X1 _16563_ (
    .A(_06471_),
    .ZN(_06472_)
  );
  AND2_X1 _16564_ (
    .A1(_06444_),
    .A2(_06471_),
    .ZN(_06474_)
  );
  INV_X1 _16565_ (
    .A(_06474_),
    .ZN(_06475_)
  );
  AND2_X1 _16566_ (
    .A1(_06443_),
    .A2(_06472_),
    .ZN(_06476_)
  );
  INV_X1 _16567_ (
    .A(_06476_),
    .ZN(_06477_)
  );
  AND2_X1 _16568_ (
    .A1(_06475_),
    .A2(_06477_),
    .ZN(_06478_)
  );
  INV_X1 _16569_ (
    .A(_06478_),
    .ZN(_06479_)
  );
  AND2_X1 _16570_ (
    .A1(_06214_),
    .A2(_06478_),
    .ZN(_06480_)
  );
  INV_X1 _16571_ (
    .A(_06480_),
    .ZN(_06481_)
  );
  AND2_X1 _16572_ (
    .A1(_06215_),
    .A2(_06479_),
    .ZN(_06482_)
  );
  INV_X1 _16573_ (
    .A(_06482_),
    .ZN(_06483_)
  );
  AND2_X1 _16574_ (
    .A1(_06481_),
    .A2(_06483_),
    .ZN(_06485_)
  );
  INV_X1 _16575_ (
    .A(_06485_),
    .ZN(_06486_)
  );
  AND2_X1 _16576_ (
    .A1(_06442_),
    .A2(_06485_),
    .ZN(_06487_)
  );
  INV_X1 _16577_ (
    .A(_06487_),
    .ZN(_06488_)
  );
  AND2_X1 _16578_ (
    .A1(_06441_),
    .A2(_06486_),
    .ZN(_06489_)
  );
  INV_X1 _16579_ (
    .A(_06489_),
    .ZN(_06490_)
  );
  AND2_X1 _16580_ (
    .A1(_06488_),
    .A2(_06490_),
    .ZN(_06491_)
  );
  INV_X1 _16581_ (
    .A(_06491_),
    .ZN(_06492_)
  );
  AND2_X1 _16582_ (
    .A1(_06118_),
    .A2(_06491_),
    .ZN(_06493_)
  );
  INV_X1 _16583_ (
    .A(_06493_),
    .ZN(_06494_)
  );
  AND2_X1 _16584_ (
    .A1(_06119_),
    .A2(_06492_),
    .ZN(_06496_)
  );
  INV_X1 _16585_ (
    .A(_06496_),
    .ZN(_06497_)
  );
  AND2_X1 _16586_ (
    .A1(_06494_),
    .A2(_06497_),
    .ZN(_06498_)
  );
  INV_X1 _16587_ (
    .A(_06498_),
    .ZN(_06499_)
  );
  AND2_X1 _16588_ (
    .A1(_06438_),
    .A2(_06498_),
    .ZN(_06500_)
  );
  INV_X1 _16589_ (
    .A(_06500_),
    .ZN(_06501_)
  );
  AND2_X1 _16590_ (
    .A1(_06439_),
    .A2(_06499_),
    .ZN(_06502_)
  );
  INV_X1 _16591_ (
    .A(_06502_),
    .ZN(_06503_)
  );
  AND2_X1 _16592_ (
    .A1(_06501_),
    .A2(_06503_),
    .ZN(_06504_)
  );
  INV_X1 _16593_ (
    .A(_06504_),
    .ZN(_06505_)
  );
  AND2_X1 _16594_ (
    .A1(_06404_),
    .A2(_06504_),
    .ZN(_06507_)
  );
  INV_X1 _16595_ (
    .A(_06507_),
    .ZN(_06508_)
  );
  AND2_X1 _16596_ (
    .A1(_06403_),
    .A2(_06505_),
    .ZN(_06509_)
  );
  INV_X1 _16597_ (
    .A(_06509_),
    .ZN(_06510_)
  );
  AND2_X1 _16598_ (
    .A1(_06508_),
    .A2(_06510_),
    .ZN(_06511_)
  );
  INV_X1 _16599_ (
    .A(_06511_),
    .ZN(_06512_)
  );
  AND2_X1 _16600_ (
    .A1(divisor[23]),
    .A2(remainder[0]),
    .ZN(_06513_)
  );
  INV_X1 _16601_ (
    .A(_06513_),
    .ZN(_06514_)
  );
  AND2_X1 _16602_ (
    .A1(divisor[22]),
    .A2(remainder[1]),
    .ZN(_06515_)
  );
  INV_X1 _16603_ (
    .A(_06515_),
    .ZN(_06516_)
  );
  AND2_X1 _16604_ (
    .A1(divisor[23]),
    .A2(remainder[1]),
    .ZN(_06518_)
  );
  INV_X1 _16605_ (
    .A(_06518_),
    .ZN(_06519_)
  );
  AND2_X1 _16606_ (
    .A1(_06192_),
    .A2(_06518_),
    .ZN(_06520_)
  );
  INV_X1 _16607_ (
    .A(_06520_),
    .ZN(_06521_)
  );
  AND2_X1 _16608_ (
    .A1(_06514_),
    .A2(_06516_),
    .ZN(_06522_)
  );
  INV_X1 _16609_ (
    .A(_06522_),
    .ZN(_06523_)
  );
  AND2_X1 _16610_ (
    .A1(_06521_),
    .A2(_06523_),
    .ZN(_06524_)
  );
  INV_X1 _16611_ (
    .A(_06524_),
    .ZN(_06525_)
  );
  AND2_X1 _16612_ (
    .A1(divisor[19]),
    .A2(remainder[4]),
    .ZN(_06526_)
  );
  INV_X1 _16613_ (
    .A(_06526_),
    .ZN(_06527_)
  );
  AND2_X1 _16614_ (
    .A1(divisor[20]),
    .A2(remainder[3]),
    .ZN(_06529_)
  );
  INV_X1 _16615_ (
    .A(_06529_),
    .ZN(_06530_)
  );
  AND2_X1 _16616_ (
    .A1(divisor[21]),
    .A2(remainder[3]),
    .ZN(_06531_)
  );
  INV_X1 _16617_ (
    .A(_06531_),
    .ZN(_06532_)
  );
  AND2_X1 _16618_ (
    .A1(_06198_),
    .A2(_06529_),
    .ZN(_06533_)
  );
  INV_X1 _16619_ (
    .A(_06533_),
    .ZN(_06534_)
  );
  AND2_X1 _16620_ (
    .A1(_06199_),
    .A2(_06530_),
    .ZN(_06535_)
  );
  INV_X1 _16621_ (
    .A(_06535_),
    .ZN(_06536_)
  );
  AND2_X1 _16622_ (
    .A1(_06534_),
    .A2(_06536_),
    .ZN(_06537_)
  );
  INV_X1 _16623_ (
    .A(_06537_),
    .ZN(_06538_)
  );
  AND2_X1 _16624_ (
    .A1(_06526_),
    .A2(_06537_),
    .ZN(_06539_)
  );
  INV_X1 _16625_ (
    .A(_06539_),
    .ZN(_06540_)
  );
  AND2_X1 _16626_ (
    .A1(_06527_),
    .A2(_06538_),
    .ZN(_06541_)
  );
  INV_X1 _16627_ (
    .A(_06541_),
    .ZN(_06542_)
  );
  AND2_X1 _16628_ (
    .A1(_06540_),
    .A2(_06542_),
    .ZN(_06543_)
  );
  INV_X1 _16629_ (
    .A(_06543_),
    .ZN(_06544_)
  );
  AND2_X1 _16630_ (
    .A1(_06524_),
    .A2(_06543_),
    .ZN(_06545_)
  );
  INV_X1 _16631_ (
    .A(_06545_),
    .ZN(_06546_)
  );
  AND2_X1 _16632_ (
    .A1(_06525_),
    .A2(_06544_),
    .ZN(_06547_)
  );
  INV_X1 _16633_ (
    .A(_06547_),
    .ZN(_06548_)
  );
  AND2_X1 _16634_ (
    .A1(_06546_),
    .A2(_06548_),
    .ZN(_06550_)
  );
  INV_X1 _16635_ (
    .A(_06550_),
    .ZN(_06551_)
  );
  AND2_X1 _16636_ (
    .A1(_06396_),
    .A2(_06551_),
    .ZN(_06552_)
  );
  INV_X1 _16637_ (
    .A(_06552_),
    .ZN(_06553_)
  );
  AND2_X1 _16638_ (
    .A1(_06398_),
    .A2(_06550_),
    .ZN(_06554_)
  );
  INV_X1 _16639_ (
    .A(_06554_),
    .ZN(_06555_)
  );
  AND2_X1 _16640_ (
    .A1(_06398_),
    .A2(_06551_),
    .ZN(_06556_)
  );
  INV_X1 _16641_ (
    .A(_06556_),
    .ZN(_06557_)
  );
  AND2_X1 _16642_ (
    .A1(_06396_),
    .A2(_06550_),
    .ZN(_06558_)
  );
  INV_X1 _16643_ (
    .A(_06558_),
    .ZN(_06559_)
  );
  AND2_X1 _16644_ (
    .A1(_06553_),
    .A2(_06555_),
    .ZN(_06561_)
  );
  AND2_X1 _16645_ (
    .A1(_06557_),
    .A2(_06559_),
    .ZN(_06562_)
  );
  AND2_X1 _16646_ (
    .A1(_06511_),
    .A2(_06562_),
    .ZN(_06563_)
  );
  INV_X1 _16647_ (
    .A(_06563_),
    .ZN(_06564_)
  );
  AND2_X1 _16648_ (
    .A1(_06512_),
    .A2(_06561_),
    .ZN(_06565_)
  );
  INV_X1 _16649_ (
    .A(_06565_),
    .ZN(_06566_)
  );
  AND2_X1 _16650_ (
    .A1(_06564_),
    .A2(_06566_),
    .ZN(_06567_)
  );
  INV_X1 _16651_ (
    .A(_06567_),
    .ZN(_06568_)
  );
  AND2_X1 _16652_ (
    .A1(_06402_),
    .A2(_06567_),
    .ZN(_06569_)
  );
  INV_X1 _16653_ (
    .A(_06569_),
    .ZN(_06570_)
  );
  AND2_X1 _16654_ (
    .A1(_06401_),
    .A2(_06568_),
    .ZN(_06572_)
  );
  INV_X1 _16655_ (
    .A(_06572_),
    .ZN(_06573_)
  );
  AND2_X1 _16656_ (
    .A1(_06570_),
    .A2(_06573_),
    .ZN(_06574_)
  );
  INV_X1 _16657_ (
    .A(_06574_),
    .ZN(_06575_)
  );
  AND2_X1 _16658_ (
    .A1(_06283_),
    .A2(_06289_),
    .ZN(_06576_)
  );
  INV_X1 _16659_ (
    .A(_06576_),
    .ZN(_06577_)
  );
  AND2_X1 _16660_ (
    .A1(_06270_),
    .A2(_06276_),
    .ZN(_06578_)
  );
  INV_X1 _16661_ (
    .A(_06578_),
    .ZN(_06579_)
  );
  AND2_X1 _16662_ (
    .A1(_06257_),
    .A2(_06263_),
    .ZN(_06580_)
  );
  INV_X1 _16663_ (
    .A(_06580_),
    .ZN(_06581_)
  );
  AND2_X1 _16664_ (
    .A1(_06167_),
    .A2(_06174_),
    .ZN(_06583_)
  );
  INV_X1 _16665_ (
    .A(_06583_),
    .ZN(_06584_)
  );
  AND2_X1 _16666_ (
    .A1(_06266_),
    .A2(_06584_),
    .ZN(_06585_)
  );
  INV_X1 _16667_ (
    .A(_06585_),
    .ZN(_06586_)
  );
  AND2_X1 _16668_ (
    .A1(_06268_),
    .A2(_06583_),
    .ZN(_06587_)
  );
  INV_X1 _16669_ (
    .A(_06587_),
    .ZN(_06588_)
  );
  AND2_X1 _16670_ (
    .A1(_06586_),
    .A2(_06588_),
    .ZN(_06589_)
  );
  INV_X1 _16671_ (
    .A(_06589_),
    .ZN(_06590_)
  );
  AND2_X1 _16672_ (
    .A1(_06581_),
    .A2(_06589_),
    .ZN(_06591_)
  );
  INV_X1 _16673_ (
    .A(_06591_),
    .ZN(_06592_)
  );
  AND2_X1 _16674_ (
    .A1(_06580_),
    .A2(_06590_),
    .ZN(_06594_)
  );
  INV_X1 _16675_ (
    .A(_06594_),
    .ZN(_06595_)
  );
  AND2_X1 _16676_ (
    .A1(_06592_),
    .A2(_06595_),
    .ZN(_06596_)
  );
  INV_X1 _16677_ (
    .A(_06596_),
    .ZN(_06597_)
  );
  AND2_X1 _16678_ (
    .A1(_06579_),
    .A2(_06596_),
    .ZN(_06598_)
  );
  INV_X1 _16679_ (
    .A(_06598_),
    .ZN(_06599_)
  );
  AND2_X1 _16680_ (
    .A1(_06578_),
    .A2(_06597_),
    .ZN(_06600_)
  );
  INV_X1 _16681_ (
    .A(_06600_),
    .ZN(_06601_)
  );
  AND2_X1 _16682_ (
    .A1(_06599_),
    .A2(_06601_),
    .ZN(_06602_)
  );
  INV_X1 _16683_ (
    .A(_06602_),
    .ZN(_06603_)
  );
  AND2_X1 _16684_ (
    .A1(_03170_),
    .A2(_06602_),
    .ZN(_06605_)
  );
  INV_X1 _16685_ (
    .A(_06605_),
    .ZN(_06606_)
  );
  AND2_X1 _16686_ (
    .A1(_03169_),
    .A2(_06603_),
    .ZN(_06607_)
  );
  INV_X1 _16687_ (
    .A(_06607_),
    .ZN(_06608_)
  );
  AND2_X1 _16688_ (
    .A1(_06606_),
    .A2(_06608_),
    .ZN(_06609_)
  );
  INV_X1 _16689_ (
    .A(_06609_),
    .ZN(_06610_)
  );
  AND2_X1 _16690_ (
    .A1(_06185_),
    .A2(_06609_),
    .ZN(_06611_)
  );
  INV_X1 _16691_ (
    .A(_06611_),
    .ZN(_06612_)
  );
  AND2_X1 _16692_ (
    .A1(_06186_),
    .A2(_06610_),
    .ZN(_06613_)
  );
  INV_X1 _16693_ (
    .A(_06613_),
    .ZN(_06614_)
  );
  AND2_X1 _16694_ (
    .A1(_06612_),
    .A2(_06614_),
    .ZN(_06616_)
  );
  INV_X1 _16695_ (
    .A(_06616_),
    .ZN(_06617_)
  );
  AND2_X1 _16696_ (
    .A1(_06577_),
    .A2(_06616_),
    .ZN(_06618_)
  );
  INV_X1 _16697_ (
    .A(_06618_),
    .ZN(_06619_)
  );
  AND2_X1 _16698_ (
    .A1(_06576_),
    .A2(_06617_),
    .ZN(_06620_)
  );
  INV_X1 _16699_ (
    .A(_06620_),
    .ZN(_06621_)
  );
  AND2_X1 _16700_ (
    .A1(_06619_),
    .A2(_06621_),
    .ZN(_06622_)
  );
  INV_X1 _16701_ (
    .A(_06622_),
    .ZN(_06623_)
  );
  AND2_X1 _16702_ (
    .A1(_06574_),
    .A2(_06622_),
    .ZN(_06624_)
  );
  INV_X1 _16703_ (
    .A(_06624_),
    .ZN(_06625_)
  );
  AND2_X1 _16704_ (
    .A1(_06575_),
    .A2(_06623_),
    .ZN(_06627_)
  );
  INV_X1 _16705_ (
    .A(_06627_),
    .ZN(_06628_)
  );
  AND2_X1 _16706_ (
    .A1(_06625_),
    .A2(_06628_),
    .ZN(_06629_)
  );
  INV_X1 _16707_ (
    .A(_06629_),
    .ZN(_06630_)
  );
  AND2_X1 _16708_ (
    .A1(_06395_),
    .A2(_06629_),
    .ZN(_06631_)
  );
  INV_X1 _16709_ (
    .A(_06631_),
    .ZN(_06632_)
  );
  AND2_X1 _16710_ (
    .A1(_06394_),
    .A2(_06630_),
    .ZN(_06633_)
  );
  INV_X1 _16711_ (
    .A(_06633_),
    .ZN(_06634_)
  );
  AND2_X1 _16712_ (
    .A1(_06632_),
    .A2(_06634_),
    .ZN(_06635_)
  );
  INV_X1 _16713_ (
    .A(_06635_),
    .ZN(_06636_)
  );
  AND2_X1 _16714_ (
    .A1(_06393_),
    .A2(_06635_),
    .ZN(_06638_)
  );
  INV_X1 _16715_ (
    .A(_06638_),
    .ZN(_06639_)
  );
  AND2_X1 _16716_ (
    .A1(_06392_),
    .A2(_06636_),
    .ZN(_06640_)
  );
  INV_X1 _16717_ (
    .A(_06640_),
    .ZN(_06641_)
  );
  AND2_X1 _16718_ (
    .A1(_06639_),
    .A2(_06641_),
    .ZN(_06642_)
  );
  INV_X1 _16719_ (
    .A(_06642_),
    .ZN(_06643_)
  );
  AND2_X1 _16720_ (
    .A1(_06391_),
    .A2(_06642_),
    .ZN(_06644_)
  );
  INV_X1 _16721_ (
    .A(_06644_),
    .ZN(_06645_)
  );
  AND2_X1 _16722_ (
    .A1(_06390_),
    .A2(_06643_),
    .ZN(_06646_)
  );
  INV_X1 _16723_ (
    .A(_06646_),
    .ZN(_06647_)
  );
  AND2_X1 _16724_ (
    .A1(_06645_),
    .A2(_06647_),
    .ZN(_06649_)
  );
  INV_X1 _16725_ (
    .A(_06649_),
    .ZN(_06650_)
  );
  AND2_X1 _16726_ (
    .A1(_06327_),
    .A2(_06649_),
    .ZN(_06651_)
  );
  INV_X1 _16727_ (
    .A(_06651_),
    .ZN(_06652_)
  );
  AND2_X1 _16728_ (
    .A1(_06328_),
    .A2(_06650_),
    .ZN(_06653_)
  );
  INV_X1 _16729_ (
    .A(_06653_),
    .ZN(_06654_)
  );
  AND2_X1 _16730_ (
    .A1(_06652_),
    .A2(_06654_),
    .ZN(_06655_)
  );
  INV_X1 _16731_ (
    .A(_06655_),
    .ZN(_06656_)
  );
  AND2_X1 _16732_ (
    .A1(_06388_),
    .A2(_06656_),
    .ZN(_06657_)
  );
  INV_X1 _16733_ (
    .A(_06657_),
    .ZN(_06658_)
  );
  AND2_X1 _16734_ (
    .A1(_06389_),
    .A2(_06655_),
    .ZN(_06660_)
  );
  INV_X1 _16735_ (
    .A(_06660_),
    .ZN(_06661_)
  );
  AND2_X1 _16736_ (
    .A1(_06658_),
    .A2(_06661_),
    .ZN(_06662_)
  );
  INV_X1 _16737_ (
    .A(_06662_),
    .ZN(_06663_)
  );
  AND2_X1 _16738_ (
    .A1(remainder[56]),
    .A2(_06662_),
    .ZN(_06664_)
  );
  INV_X1 _16739_ (
    .A(_06664_),
    .ZN(_06665_)
  );
  AND2_X1 _16740_ (
    .A1(_04503_),
    .A2(_06663_),
    .ZN(_06666_)
  );
  INV_X1 _16741_ (
    .A(_06666_),
    .ZN(_06667_)
  );
  AND2_X1 _16742_ (
    .A1(_06665_),
    .A2(_06667_),
    .ZN(_06668_)
  );
  INV_X1 _16743_ (
    .A(_06668_),
    .ZN(_06669_)
  );
  AND2_X1 _16744_ (
    .A1(_06387_),
    .A2(_06668_),
    .ZN(_06671_)
  );
  INV_X1 _16745_ (
    .A(_06671_),
    .ZN(_06672_)
  );
  AND2_X1 _16746_ (
    .A1(_06385_),
    .A2(_06669_),
    .ZN(_06673_)
  );
  INV_X1 _16747_ (
    .A(_06673_),
    .ZN(_06674_)
  );
  AND2_X1 _16748_ (
    .A1(_02082_),
    .A2(_06674_),
    .ZN(_06675_)
  );
  AND2_X1 _16749_ (
    .A1(_06672_),
    .A2(_06675_),
    .ZN(_06676_)
  );
  INV_X1 _16750_ (
    .A(_06676_),
    .ZN(_06677_)
  );
  AND2_X1 _16751_ (
    .A1(_06382_),
    .A2(_06677_),
    .ZN(_06678_)
  );
  AND2_X1 _16752_ (
    .A1(_06384_),
    .A2(_06678_),
    .ZN(_06679_)
  );
  INV_X1 _16753_ (
    .A(_06679_),
    .ZN(_06680_)
  );
  AND2_X1 _16754_ (
    .A1(_06201_),
    .A2(_06680_),
    .ZN(_00069_)
  );
  AND2_X1 _16755_ (
    .A1(_04590_),
    .A2(_10451_),
    .ZN(_06682_)
  );
  INV_X1 _16756_ (
    .A(_06682_),
    .ZN(_06683_)
  );
  AND2_X1 _16757_ (
    .A1(_10462_),
    .A2(_01847_),
    .ZN(_06684_)
  );
  INV_X1 _16758_ (
    .A(_06684_),
    .ZN(_06685_)
  );
  AND2_X1 _16759_ (
    .A1(_05983_),
    .A2(_06685_),
    .ZN(_06686_)
  );
  AND2_X1 _16760_ (
    .A1(_06683_),
    .A2(_06686_),
    .ZN(_06687_)
  );
  INV_X1 _16761_ (
    .A(_06687_),
    .ZN(_06688_)
  );
  AND2_X1 _16762_ (
    .A1(_06665_),
    .A2(_06672_),
    .ZN(_06689_)
  );
  INV_X1 _16763_ (
    .A(_06689_),
    .ZN(_06690_)
  );
  AND2_X1 _16764_ (
    .A1(_06632_),
    .A2(_06639_),
    .ZN(_06692_)
  );
  INV_X1 _16765_ (
    .A(_06692_),
    .ZN(_06693_)
  );
  AND2_X1 _16766_ (
    .A1(_06612_),
    .A2(_06619_),
    .ZN(_06694_)
  );
  INV_X1 _16767_ (
    .A(_06694_),
    .ZN(_06695_)
  );
  AND2_X1 _16768_ (
    .A1(_06570_),
    .A2(_06625_),
    .ZN(_06696_)
  );
  INV_X1 _16769_ (
    .A(_06696_),
    .ZN(_06697_)
  );
  AND2_X1 _16770_ (
    .A1(_03249_),
    .A2(_06551_),
    .ZN(_06698_)
  );
  INV_X1 _16771_ (
    .A(_06698_),
    .ZN(_06699_)
  );
  AND2_X1 _16772_ (
    .A1(_06218_),
    .A2(_06698_),
    .ZN(_06700_)
  );
  INV_X1 _16773_ (
    .A(_06700_),
    .ZN(_06701_)
  );
  AND2_X1 _16774_ (
    .A1(_06564_),
    .A2(_06701_),
    .ZN(_06703_)
  );
  INV_X1 _16775_ (
    .A(_06703_),
    .ZN(_06704_)
  );
  AND2_X1 _16776_ (
    .A1(_06494_),
    .A2(_06501_),
    .ZN(_06705_)
  );
  INV_X1 _16777_ (
    .A(_06705_),
    .ZN(_06706_)
  );
  AND2_X1 _16778_ (
    .A1(_06481_),
    .A2(_06488_),
    .ZN(_06707_)
  );
  INV_X1 _16779_ (
    .A(_06707_),
    .ZN(_06708_)
  );
  AND2_X1 _16780_ (
    .A1(_06468_),
    .A2(_06475_),
    .ZN(_06709_)
  );
  INV_X1 _16781_ (
    .A(_06709_),
    .ZN(_06710_)
  );
  AND2_X1 _16782_ (
    .A1(_06455_),
    .A2(_06461_),
    .ZN(_06711_)
  );
  INV_X1 _16783_ (
    .A(_06711_),
    .ZN(_06712_)
  );
  AND2_X1 _16784_ (
    .A1(_06534_),
    .A2(_06540_),
    .ZN(_06714_)
  );
  INV_X1 _16785_ (
    .A(_06714_),
    .ZN(_06715_)
  );
  AND2_X1 _16786_ (
    .A1(remainder[32]),
    .A2(divisor[16]),
    .ZN(_06716_)
  );
  INV_X1 _16787_ (
    .A(_06716_),
    .ZN(_06717_)
  );
  AND2_X1 _16788_ (
    .A1(divisor[17]),
    .A2(remainder[7]),
    .ZN(_06718_)
  );
  INV_X1 _16789_ (
    .A(_06718_),
    .ZN(_06719_)
  );
  AND2_X1 _16790_ (
    .A1(divisor[18]),
    .A2(remainder[7]),
    .ZN(_06720_)
  );
  INV_X1 _16791_ (
    .A(_06720_),
    .ZN(_06721_)
  );
  AND2_X1 _16792_ (
    .A1(_06449_),
    .A2(_06720_),
    .ZN(_06722_)
  );
  INV_X1 _16793_ (
    .A(_06722_),
    .ZN(_06723_)
  );
  AND2_X1 _16794_ (
    .A1(_06453_),
    .A2(_06719_),
    .ZN(_06725_)
  );
  INV_X1 _16795_ (
    .A(_06725_),
    .ZN(_06726_)
  );
  AND2_X1 _16796_ (
    .A1(_06723_),
    .A2(_06726_),
    .ZN(_06727_)
  );
  INV_X1 _16797_ (
    .A(_06727_),
    .ZN(_06728_)
  );
  AND2_X1 _16798_ (
    .A1(_06716_),
    .A2(_06727_),
    .ZN(_06729_)
  );
  INV_X1 _16799_ (
    .A(_06729_),
    .ZN(_06730_)
  );
  AND2_X1 _16800_ (
    .A1(_06717_),
    .A2(_06728_),
    .ZN(_06731_)
  );
  INV_X1 _16801_ (
    .A(_06731_),
    .ZN(_06732_)
  );
  AND2_X1 _16802_ (
    .A1(_06730_),
    .A2(_06732_),
    .ZN(_06733_)
  );
  INV_X1 _16803_ (
    .A(_06733_),
    .ZN(_06734_)
  );
  AND2_X1 _16804_ (
    .A1(_06715_),
    .A2(_06733_),
    .ZN(_06736_)
  );
  INV_X1 _16805_ (
    .A(_06736_),
    .ZN(_06737_)
  );
  AND2_X1 _16806_ (
    .A1(_06714_),
    .A2(_06734_),
    .ZN(_06738_)
  );
  INV_X1 _16807_ (
    .A(_06738_),
    .ZN(_06739_)
  );
  AND2_X1 _16808_ (
    .A1(_06737_),
    .A2(_06739_),
    .ZN(_06740_)
  );
  INV_X1 _16809_ (
    .A(_06740_),
    .ZN(_06741_)
  );
  AND2_X1 _16810_ (
    .A1(_06712_),
    .A2(_06740_),
    .ZN(_06742_)
  );
  INV_X1 _16811_ (
    .A(_06742_),
    .ZN(_06743_)
  );
  AND2_X1 _16812_ (
    .A1(_06711_),
    .A2(_06741_),
    .ZN(_06744_)
  );
  INV_X1 _16813_ (
    .A(_06744_),
    .ZN(_06745_)
  );
  AND2_X1 _16814_ (
    .A1(_06743_),
    .A2(_06745_),
    .ZN(_06747_)
  );
  INV_X1 _16815_ (
    .A(_06747_),
    .ZN(_06748_)
  );
  AND2_X1 _16816_ (
    .A1(_06545_),
    .A2(_06747_),
    .ZN(_06749_)
  );
  INV_X1 _16817_ (
    .A(_06749_),
    .ZN(_06750_)
  );
  AND2_X1 _16818_ (
    .A1(_06546_),
    .A2(_06748_),
    .ZN(_06751_)
  );
  INV_X1 _16819_ (
    .A(_06751_),
    .ZN(_06752_)
  );
  AND2_X1 _16820_ (
    .A1(_06750_),
    .A2(_06752_),
    .ZN(_06753_)
  );
  INV_X1 _16821_ (
    .A(_06753_),
    .ZN(_06754_)
  );
  AND2_X1 _16822_ (
    .A1(_06710_),
    .A2(_06753_),
    .ZN(_06755_)
  );
  INV_X1 _16823_ (
    .A(_06755_),
    .ZN(_06756_)
  );
  AND2_X1 _16824_ (
    .A1(_06709_),
    .A2(_06754_),
    .ZN(_06758_)
  );
  INV_X1 _16825_ (
    .A(_06758_),
    .ZN(_06759_)
  );
  AND2_X1 _16826_ (
    .A1(_06756_),
    .A2(_06759_),
    .ZN(_06760_)
  );
  INV_X1 _16827_ (
    .A(_06760_),
    .ZN(_06761_)
  );
  AND2_X1 _16828_ (
    .A1(_06708_),
    .A2(_06760_),
    .ZN(_06762_)
  );
  INV_X1 _16829_ (
    .A(_06762_),
    .ZN(_06763_)
  );
  AND2_X1 _16830_ (
    .A1(_06707_),
    .A2(_06761_),
    .ZN(_06764_)
  );
  INV_X1 _16831_ (
    .A(_06764_),
    .ZN(_06765_)
  );
  AND2_X1 _16832_ (
    .A1(_06763_),
    .A2(_06765_),
    .ZN(_06766_)
  );
  INV_X1 _16833_ (
    .A(_06766_),
    .ZN(_06767_)
  );
  AND2_X1 _16834_ (
    .A1(_05761_),
    .A2(_06410_),
    .ZN(_06769_)
  );
  INV_X1 _16835_ (
    .A(_06769_),
    .ZN(_06770_)
  );
  AND2_X1 _16836_ (
    .A1(_05501_),
    .A2(_06769_),
    .ZN(_06771_)
  );
  INV_X1 _16837_ (
    .A(_06771_),
    .ZN(_06772_)
  );
  AND2_X1 _16838_ (
    .A1(_06420_),
    .A2(_06770_),
    .ZN(_06773_)
  );
  INV_X1 _16839_ (
    .A(_06773_),
    .ZN(_06774_)
  );
  AND2_X1 _16840_ (
    .A1(_06415_),
    .A2(_06770_),
    .ZN(_06775_)
  );
  INV_X1 _16841_ (
    .A(_06775_),
    .ZN(_06776_)
  );
  AND2_X1 _16842_ (
    .A1(_06424_),
    .A2(_06776_),
    .ZN(_06777_)
  );
  INV_X1 _16843_ (
    .A(_06777_),
    .ZN(_06778_)
  );
  AND2_X1 _16844_ (
    .A1(_06772_),
    .A2(_06774_),
    .ZN(_06780_)
  );
  INV_X1 _16845_ (
    .A(_06780_),
    .ZN(_06781_)
  );
  AND2_X1 _16846_ (
    .A1(_05813_),
    .A2(_06780_),
    .ZN(_06782_)
  );
  INV_X1 _16847_ (
    .A(_06782_),
    .ZN(_06783_)
  );
  AND2_X1 _16848_ (
    .A1(_05814_),
    .A2(_06781_),
    .ZN(_06784_)
  );
  INV_X1 _16849_ (
    .A(_06784_),
    .ZN(_06785_)
  );
  AND2_X1 _16850_ (
    .A1(_06783_),
    .A2(_06785_),
    .ZN(_06786_)
  );
  INV_X1 _16851_ (
    .A(_06786_),
    .ZN(_06787_)
  );
  AND2_X1 _16852_ (
    .A1(_06766_),
    .A2(_06786_),
    .ZN(_06788_)
  );
  INV_X1 _16853_ (
    .A(_06788_),
    .ZN(_06789_)
  );
  AND2_X1 _16854_ (
    .A1(_06767_),
    .A2(_06787_),
    .ZN(_06791_)
  );
  INV_X1 _16855_ (
    .A(_06791_),
    .ZN(_06792_)
  );
  AND2_X1 _16856_ (
    .A1(_06789_),
    .A2(_06792_),
    .ZN(_06793_)
  );
  INV_X1 _16857_ (
    .A(_06793_),
    .ZN(_06794_)
  );
  AND2_X1 _16858_ (
    .A1(_06706_),
    .A2(_06793_),
    .ZN(_06795_)
  );
  INV_X1 _16859_ (
    .A(_06795_),
    .ZN(_06796_)
  );
  AND2_X1 _16860_ (
    .A1(_06705_),
    .A2(_06794_),
    .ZN(_06797_)
  );
  INV_X1 _16861_ (
    .A(_06797_),
    .ZN(_06798_)
  );
  AND2_X1 _16862_ (
    .A1(_06796_),
    .A2(_06798_),
    .ZN(_06799_)
  );
  INV_X1 _16863_ (
    .A(_06799_),
    .ZN(_06800_)
  );
  AND2_X1 _16864_ (
    .A1(divisor[22]),
    .A2(remainder[2]),
    .ZN(_06802_)
  );
  INV_X1 _16865_ (
    .A(_06802_),
    .ZN(_06803_)
  );
  AND2_X1 _16866_ (
    .A1(divisor[24]),
    .A2(remainder[0]),
    .ZN(_06804_)
  );
  INV_X1 _16867_ (
    .A(_06804_),
    .ZN(_06805_)
  );
  AND2_X1 _16868_ (
    .A1(divisor[24]),
    .A2(remainder[1]),
    .ZN(_06806_)
  );
  INV_X1 _16869_ (
    .A(_06806_),
    .ZN(_06807_)
  );
  AND2_X1 _16870_ (
    .A1(_06513_),
    .A2(_06806_),
    .ZN(_06808_)
  );
  INV_X1 _16871_ (
    .A(_06808_),
    .ZN(_06809_)
  );
  AND2_X1 _16872_ (
    .A1(_06519_),
    .A2(_06805_),
    .ZN(_06810_)
  );
  INV_X1 _16873_ (
    .A(_06810_),
    .ZN(_06811_)
  );
  AND2_X1 _16874_ (
    .A1(_06809_),
    .A2(_06811_),
    .ZN(_06813_)
  );
  INV_X1 _16875_ (
    .A(_06813_),
    .ZN(_06814_)
  );
  AND2_X1 _16876_ (
    .A1(_06802_),
    .A2(_06813_),
    .ZN(_06815_)
  );
  INV_X1 _16877_ (
    .A(_06815_),
    .ZN(_06816_)
  );
  AND2_X1 _16878_ (
    .A1(_06803_),
    .A2(_06814_),
    .ZN(_06817_)
  );
  INV_X1 _16879_ (
    .A(_06817_),
    .ZN(_06818_)
  );
  AND2_X1 _16880_ (
    .A1(_06816_),
    .A2(_06818_),
    .ZN(_06819_)
  );
  INV_X1 _16881_ (
    .A(_06819_),
    .ZN(_06820_)
  );
  AND2_X1 _16882_ (
    .A1(_06520_),
    .A2(_06819_),
    .ZN(_06821_)
  );
  INV_X1 _16883_ (
    .A(_06821_),
    .ZN(_06822_)
  );
  AND2_X1 _16884_ (
    .A1(_06521_),
    .A2(_06820_),
    .ZN(_06823_)
  );
  INV_X1 _16885_ (
    .A(_06823_),
    .ZN(_06824_)
  );
  AND2_X1 _16886_ (
    .A1(_06822_),
    .A2(_06824_),
    .ZN(_06825_)
  );
  INV_X1 _16887_ (
    .A(_06825_),
    .ZN(_06826_)
  );
  AND2_X1 _16888_ (
    .A1(divisor[19]),
    .A2(remainder[5]),
    .ZN(_06827_)
  );
  INV_X1 _16889_ (
    .A(_06827_),
    .ZN(_06828_)
  );
  AND2_X1 _16890_ (
    .A1(divisor[20]),
    .A2(remainder[4]),
    .ZN(_06829_)
  );
  INV_X1 _16891_ (
    .A(_06829_),
    .ZN(_06830_)
  );
  AND2_X1 _16892_ (
    .A1(divisor[21]),
    .A2(remainder[4]),
    .ZN(_06831_)
  );
  INV_X1 _16893_ (
    .A(_06831_),
    .ZN(_06832_)
  );
  AND2_X1 _16894_ (
    .A1(_06531_),
    .A2(_06829_),
    .ZN(_06834_)
  );
  INV_X1 _16895_ (
    .A(_06834_),
    .ZN(_06835_)
  );
  AND2_X1 _16896_ (
    .A1(_06532_),
    .A2(_06830_),
    .ZN(_06836_)
  );
  INV_X1 _16897_ (
    .A(_06836_),
    .ZN(_06837_)
  );
  AND2_X1 _16898_ (
    .A1(_06835_),
    .A2(_06837_),
    .ZN(_06838_)
  );
  INV_X1 _16899_ (
    .A(_06838_),
    .ZN(_06839_)
  );
  AND2_X1 _16900_ (
    .A1(_06827_),
    .A2(_06838_),
    .ZN(_06840_)
  );
  INV_X1 _16901_ (
    .A(_06840_),
    .ZN(_06841_)
  );
  AND2_X1 _16902_ (
    .A1(_06828_),
    .A2(_06839_),
    .ZN(_06842_)
  );
  INV_X1 _16903_ (
    .A(_06842_),
    .ZN(_06843_)
  );
  AND2_X1 _16904_ (
    .A1(_06841_),
    .A2(_06843_),
    .ZN(_06845_)
  );
  INV_X1 _16905_ (
    .A(_06845_),
    .ZN(_06846_)
  );
  AND2_X1 _16906_ (
    .A1(_06825_),
    .A2(_06845_),
    .ZN(_06847_)
  );
  INV_X1 _16907_ (
    .A(_06847_),
    .ZN(_06848_)
  );
  AND2_X1 _16908_ (
    .A1(_06826_),
    .A2(_06846_),
    .ZN(_06849_)
  );
  INV_X1 _16909_ (
    .A(_06849_),
    .ZN(_06850_)
  );
  AND2_X1 _16910_ (
    .A1(_06848_),
    .A2(_06850_),
    .ZN(_06851_)
  );
  INV_X1 _16911_ (
    .A(_06851_),
    .ZN(_06852_)
  );
  AND2_X1 _16912_ (
    .A1(_06698_),
    .A2(_06852_),
    .ZN(_06853_)
  );
  INV_X1 _16913_ (
    .A(_06853_),
    .ZN(_06854_)
  );
  AND2_X1 _16914_ (
    .A1(_06699_),
    .A2(_06851_),
    .ZN(_06856_)
  );
  INV_X1 _16915_ (
    .A(_06856_),
    .ZN(_06857_)
  );
  AND2_X1 _16916_ (
    .A1(_06699_),
    .A2(_06852_),
    .ZN(_06858_)
  );
  INV_X1 _16917_ (
    .A(_06858_),
    .ZN(_06859_)
  );
  AND2_X1 _16918_ (
    .A1(_06698_),
    .A2(_06851_),
    .ZN(_06860_)
  );
  INV_X1 _16919_ (
    .A(_06860_),
    .ZN(_06861_)
  );
  AND2_X1 _16920_ (
    .A1(_06854_),
    .A2(_06857_),
    .ZN(_06862_)
  );
  AND2_X1 _16921_ (
    .A1(_06859_),
    .A2(_06861_),
    .ZN(_06863_)
  );
  AND2_X1 _16922_ (
    .A1(_06799_),
    .A2(_06863_),
    .ZN(_06864_)
  );
  INV_X1 _16923_ (
    .A(_06864_),
    .ZN(_06865_)
  );
  AND2_X1 _16924_ (
    .A1(_06800_),
    .A2(_06862_),
    .ZN(_06867_)
  );
  INV_X1 _16925_ (
    .A(_06867_),
    .ZN(_06868_)
  );
  AND2_X1 _16926_ (
    .A1(_06865_),
    .A2(_06868_),
    .ZN(_06869_)
  );
  INV_X1 _16927_ (
    .A(_06869_),
    .ZN(_06870_)
  );
  AND2_X1 _16928_ (
    .A1(_06704_),
    .A2(_06869_),
    .ZN(_06871_)
  );
  INV_X1 _16929_ (
    .A(_06871_),
    .ZN(_06872_)
  );
  AND2_X1 _16930_ (
    .A1(_06703_),
    .A2(_06870_),
    .ZN(_06873_)
  );
  INV_X1 _16931_ (
    .A(_06873_),
    .ZN(_06874_)
  );
  AND2_X1 _16932_ (
    .A1(_06872_),
    .A2(_06874_),
    .ZN(_06875_)
  );
  INV_X1 _16933_ (
    .A(_06875_),
    .ZN(_06876_)
  );
  AND2_X1 _16934_ (
    .A1(_06599_),
    .A2(_06606_),
    .ZN(_06878_)
  );
  INV_X1 _16935_ (
    .A(_06878_),
    .ZN(_06879_)
  );
  AND2_X1 _16936_ (
    .A1(_06586_),
    .A2(_06592_),
    .ZN(_06880_)
  );
  INV_X1 _16937_ (
    .A(_06880_),
    .ZN(_06881_)
  );
  AND2_X1 _16938_ (
    .A1(_06428_),
    .A2(_06435_),
    .ZN(_06882_)
  );
  INV_X1 _16939_ (
    .A(_06882_),
    .ZN(_06883_)
  );
  AND2_X1 _16940_ (
    .A1(_06266_),
    .A2(_06883_),
    .ZN(_06884_)
  );
  INV_X1 _16941_ (
    .A(_06884_),
    .ZN(_06885_)
  );
  AND2_X1 _16942_ (
    .A1(_06268_),
    .A2(_06882_),
    .ZN(_06886_)
  );
  INV_X1 _16943_ (
    .A(_06886_),
    .ZN(_06887_)
  );
  AND2_X1 _16944_ (
    .A1(_06885_),
    .A2(_06887_),
    .ZN(_06889_)
  );
  INV_X1 _16945_ (
    .A(_06889_),
    .ZN(_06890_)
  );
  AND2_X1 _16946_ (
    .A1(_06581_),
    .A2(_06889_),
    .ZN(_06891_)
  );
  INV_X1 _16947_ (
    .A(_06891_),
    .ZN(_06892_)
  );
  AND2_X1 _16948_ (
    .A1(_06580_),
    .A2(_06890_),
    .ZN(_06893_)
  );
  INV_X1 _16949_ (
    .A(_06893_),
    .ZN(_06894_)
  );
  AND2_X1 _16950_ (
    .A1(_06892_),
    .A2(_06894_),
    .ZN(_06895_)
  );
  INV_X1 _16951_ (
    .A(_06895_),
    .ZN(_06896_)
  );
  AND2_X1 _16952_ (
    .A1(_06881_),
    .A2(_06895_),
    .ZN(_06897_)
  );
  INV_X1 _16953_ (
    .A(_06897_),
    .ZN(_06898_)
  );
  AND2_X1 _16954_ (
    .A1(_06880_),
    .A2(_06896_),
    .ZN(_06900_)
  );
  INV_X1 _16955_ (
    .A(_06900_),
    .ZN(_06901_)
  );
  AND2_X1 _16956_ (
    .A1(_06898_),
    .A2(_06901_),
    .ZN(_06902_)
  );
  INV_X1 _16957_ (
    .A(_06902_),
    .ZN(_06903_)
  );
  AND2_X1 _16958_ (
    .A1(_03170_),
    .A2(_06902_),
    .ZN(_06904_)
  );
  INV_X1 _16959_ (
    .A(_06904_),
    .ZN(_06905_)
  );
  AND2_X1 _16960_ (
    .A1(_03169_),
    .A2(_06903_),
    .ZN(_06906_)
  );
  INV_X1 _16961_ (
    .A(_06906_),
    .ZN(_06907_)
  );
  AND2_X1 _16962_ (
    .A1(_06905_),
    .A2(_06907_),
    .ZN(_06908_)
  );
  INV_X1 _16963_ (
    .A(_06908_),
    .ZN(_06909_)
  );
  AND2_X1 _16964_ (
    .A1(_06507_),
    .A2(_06908_),
    .ZN(_06911_)
  );
  INV_X1 _16965_ (
    .A(_06911_),
    .ZN(_06912_)
  );
  AND2_X1 _16966_ (
    .A1(_06508_),
    .A2(_06909_),
    .ZN(_06913_)
  );
  INV_X1 _16967_ (
    .A(_06913_),
    .ZN(_06914_)
  );
  AND2_X1 _16968_ (
    .A1(_06912_),
    .A2(_06914_),
    .ZN(_06915_)
  );
  INV_X1 _16969_ (
    .A(_06915_),
    .ZN(_06916_)
  );
  AND2_X1 _16970_ (
    .A1(_06879_),
    .A2(_06915_),
    .ZN(_06917_)
  );
  INV_X1 _16971_ (
    .A(_06917_),
    .ZN(_06918_)
  );
  AND2_X1 _16972_ (
    .A1(_06878_),
    .A2(_06916_),
    .ZN(_06919_)
  );
  INV_X1 _16973_ (
    .A(_06919_),
    .ZN(_06920_)
  );
  AND2_X1 _16974_ (
    .A1(_06918_),
    .A2(_06920_),
    .ZN(_06922_)
  );
  INV_X1 _16975_ (
    .A(_06922_),
    .ZN(_06923_)
  );
  AND2_X1 _16976_ (
    .A1(_06875_),
    .A2(_06922_),
    .ZN(_06924_)
  );
  INV_X1 _16977_ (
    .A(_06924_),
    .ZN(_06925_)
  );
  AND2_X1 _16978_ (
    .A1(_06876_),
    .A2(_06923_),
    .ZN(_06926_)
  );
  INV_X1 _16979_ (
    .A(_06926_),
    .ZN(_06927_)
  );
  AND2_X1 _16980_ (
    .A1(_06925_),
    .A2(_06927_),
    .ZN(_06928_)
  );
  INV_X1 _16981_ (
    .A(_06928_),
    .ZN(_06929_)
  );
  AND2_X1 _16982_ (
    .A1(_06697_),
    .A2(_06928_),
    .ZN(_06930_)
  );
  INV_X1 _16983_ (
    .A(_06930_),
    .ZN(_06931_)
  );
  AND2_X1 _16984_ (
    .A1(_06696_),
    .A2(_06929_),
    .ZN(_06933_)
  );
  INV_X1 _16985_ (
    .A(_06933_),
    .ZN(_06934_)
  );
  AND2_X1 _16986_ (
    .A1(_06931_),
    .A2(_06934_),
    .ZN(_06935_)
  );
  INV_X1 _16987_ (
    .A(_06935_),
    .ZN(_06936_)
  );
  AND2_X1 _16988_ (
    .A1(_06695_),
    .A2(_06935_),
    .ZN(_06937_)
  );
  INV_X1 _16989_ (
    .A(_06937_),
    .ZN(_06938_)
  );
  AND2_X1 _16990_ (
    .A1(_06694_),
    .A2(_06936_),
    .ZN(_06939_)
  );
  INV_X1 _16991_ (
    .A(_06939_),
    .ZN(_06940_)
  );
  AND2_X1 _16992_ (
    .A1(_06938_),
    .A2(_06940_),
    .ZN(_06941_)
  );
  INV_X1 _16993_ (
    .A(_06941_),
    .ZN(_06942_)
  );
  AND2_X1 _16994_ (
    .A1(_06693_),
    .A2(_06941_),
    .ZN(_06944_)
  );
  INV_X1 _16995_ (
    .A(_06944_),
    .ZN(_06945_)
  );
  AND2_X1 _16996_ (
    .A1(_06692_),
    .A2(_06942_),
    .ZN(_06946_)
  );
  INV_X1 _16997_ (
    .A(_06946_),
    .ZN(_06947_)
  );
  AND2_X1 _16998_ (
    .A1(_06945_),
    .A2(_06947_),
    .ZN(_06948_)
  );
  INV_X1 _16999_ (
    .A(_06948_),
    .ZN(_06949_)
  );
  AND2_X1 _17000_ (
    .A1(_06644_),
    .A2(_06948_),
    .ZN(_06950_)
  );
  INV_X1 _17001_ (
    .A(_06950_),
    .ZN(_06951_)
  );
  AND2_X1 _17002_ (
    .A1(_06645_),
    .A2(_06949_),
    .ZN(_06952_)
  );
  INV_X1 _17003_ (
    .A(_06952_),
    .ZN(_06953_)
  );
  AND2_X1 _17004_ (
    .A1(_06951_),
    .A2(_06953_),
    .ZN(_06955_)
  );
  INV_X1 _17005_ (
    .A(_06955_),
    .ZN(_06956_)
  );
  AND2_X1 _17006_ (
    .A1(_06388_),
    .A2(_06652_),
    .ZN(_06957_)
  );
  INV_X1 _17007_ (
    .A(_06957_),
    .ZN(_06958_)
  );
  AND2_X1 _17008_ (
    .A1(_06652_),
    .A2(_06661_),
    .ZN(_06959_)
  );
  AND2_X1 _17009_ (
    .A1(_06654_),
    .A2(_06958_),
    .ZN(_06960_)
  );
  AND2_X1 _17010_ (
    .A1(_06955_),
    .A2(_06960_),
    .ZN(_06961_)
  );
  INV_X1 _17011_ (
    .A(_06961_),
    .ZN(_06962_)
  );
  AND2_X1 _17012_ (
    .A1(_06956_),
    .A2(_06959_),
    .ZN(_06963_)
  );
  INV_X1 _17013_ (
    .A(_06963_),
    .ZN(_06964_)
  );
  AND2_X1 _17014_ (
    .A1(_06962_),
    .A2(_06964_),
    .ZN(_06966_)
  );
  INV_X1 _17015_ (
    .A(_06966_),
    .ZN(_06967_)
  );
  AND2_X1 _17016_ (
    .A1(remainder[57]),
    .A2(_06966_),
    .ZN(_06968_)
  );
  INV_X1 _17017_ (
    .A(_06968_),
    .ZN(_06969_)
  );
  AND2_X1 _17018_ (
    .A1(_04492_),
    .A2(_06967_),
    .ZN(_06970_)
  );
  INV_X1 _17019_ (
    .A(_06970_),
    .ZN(_06971_)
  );
  AND2_X1 _17020_ (
    .A1(_06969_),
    .A2(_06971_),
    .ZN(_06972_)
  );
  INV_X1 _17021_ (
    .A(_06972_),
    .ZN(_06973_)
  );
  AND2_X1 _17022_ (
    .A1(_06690_),
    .A2(_06972_),
    .ZN(_06974_)
  );
  INV_X1 _17023_ (
    .A(_06974_),
    .ZN(_06975_)
  );
  AND2_X1 _17024_ (
    .A1(_06689_),
    .A2(_06973_),
    .ZN(_06977_)
  );
  INV_X1 _17025_ (
    .A(_06977_),
    .ZN(_06978_)
  );
  AND2_X1 _17026_ (
    .A1(_02082_),
    .A2(_06978_),
    .ZN(_06979_)
  );
  AND2_X1 _17027_ (
    .A1(_06975_),
    .A2(_06979_),
    .ZN(_06980_)
  );
  INV_X1 _17028_ (
    .A(_06980_),
    .ZN(_06981_)
  );
  AND2_X1 _17029_ (
    .A1(remainder[49]),
    .A2(_02077_),
    .ZN(_06982_)
  );
  INV_X1 _17030_ (
    .A(_06982_),
    .ZN(_06983_)
  );
  AND2_X1 _17031_ (
    .A1(_06688_),
    .A2(_06983_),
    .ZN(_06984_)
  );
  AND2_X1 _17032_ (
    .A1(_06981_),
    .A2(_06984_),
    .ZN(_06985_)
  );
  INV_X1 _17033_ (
    .A(_06985_),
    .ZN(_06986_)
  );
  AND2_X1 _17034_ (
    .A1(_06201_),
    .A2(_06986_),
    .ZN(_00070_)
  );
  MUX2_X1 _17035_ (
    .A(remainder[49]),
    .B(_01862_),
    .S(_10462_),
    .Z(_06988_)
  );
  AND2_X1 _17036_ (
    .A1(_05983_),
    .A2(_06988_),
    .ZN(_06989_)
  );
  INV_X1 _17037_ (
    .A(_06989_),
    .ZN(_06990_)
  );
  AND2_X1 _17038_ (
    .A1(remainder[50]),
    .A2(_02077_),
    .ZN(_06991_)
  );
  INV_X1 _17039_ (
    .A(_06991_),
    .ZN(_06992_)
  );
  AND2_X1 _17040_ (
    .A1(_06969_),
    .A2(_06975_),
    .ZN(_06993_)
  );
  INV_X1 _17041_ (
    .A(_06993_),
    .ZN(_06994_)
  );
  AND2_X1 _17042_ (
    .A1(_06951_),
    .A2(_06962_),
    .ZN(_06995_)
  );
  INV_X1 _17043_ (
    .A(_06995_),
    .ZN(_06996_)
  );
  AND2_X1 _17044_ (
    .A1(_06931_),
    .A2(_06938_),
    .ZN(_06998_)
  );
  INV_X1 _17045_ (
    .A(_06998_),
    .ZN(_06999_)
  );
  AND2_X1 _17046_ (
    .A1(_06912_),
    .A2(_06918_),
    .ZN(_07000_)
  );
  INV_X1 _17047_ (
    .A(_07000_),
    .ZN(_07001_)
  );
  AND2_X1 _17048_ (
    .A1(_06872_),
    .A2(_06925_),
    .ZN(_07002_)
  );
  INV_X1 _17049_ (
    .A(_07002_),
    .ZN(_07003_)
  );
  AND2_X1 _17050_ (
    .A1(_03249_),
    .A2(_06852_),
    .ZN(_07004_)
  );
  INV_X1 _17051_ (
    .A(_07004_),
    .ZN(_07005_)
  );
  AND2_X1 _17052_ (
    .A1(_06550_),
    .A2(_07004_),
    .ZN(_07006_)
  );
  INV_X1 _17053_ (
    .A(_07006_),
    .ZN(_07007_)
  );
  AND2_X1 _17054_ (
    .A1(_06865_),
    .A2(_07007_),
    .ZN(_07009_)
  );
  INV_X1 _17055_ (
    .A(_07009_),
    .ZN(_07010_)
  );
  AND2_X1 _17056_ (
    .A1(_06763_),
    .A2(_06789_),
    .ZN(_07011_)
  );
  INV_X1 _17057_ (
    .A(_07011_),
    .ZN(_07012_)
  );
  AND2_X1 _17058_ (
    .A1(_06750_),
    .A2(_06756_),
    .ZN(_07013_)
  );
  INV_X1 _17059_ (
    .A(_07013_),
    .ZN(_07014_)
  );
  AND2_X1 _17060_ (
    .A1(_06737_),
    .A2(_06743_),
    .ZN(_07015_)
  );
  INV_X1 _17061_ (
    .A(_07015_),
    .ZN(_07016_)
  );
  AND2_X1 _17062_ (
    .A1(_06822_),
    .A2(_06848_),
    .ZN(_07017_)
  );
  INV_X1 _17063_ (
    .A(_07017_),
    .ZN(_07018_)
  );
  AND2_X1 _17064_ (
    .A1(_06723_),
    .A2(_06730_),
    .ZN(_07020_)
  );
  INV_X1 _17065_ (
    .A(_07020_),
    .ZN(_07021_)
  );
  AND2_X1 _17066_ (
    .A1(_06835_),
    .A2(_06841_),
    .ZN(_07022_)
  );
  INV_X1 _17067_ (
    .A(_07022_),
    .ZN(_07023_)
  );
  AND2_X1 _17068_ (
    .A1(remainder[32]),
    .A2(divisor[18]),
    .ZN(_07024_)
  );
  AND2_X1 _17069_ (
    .A1(remainder[32]),
    .A2(divisor[17]),
    .ZN(_07025_)
  );
  INV_X1 _17070_ (
    .A(_07025_),
    .ZN(_07026_)
  );
  AND2_X1 _17071_ (
    .A1(divisor[18]),
    .A2(_07025_),
    .ZN(_07027_)
  );
  INV_X1 _17072_ (
    .A(_07027_),
    .ZN(_07028_)
  );
  AND2_X1 _17073_ (
    .A1(_06720_),
    .A2(_07025_),
    .ZN(_07029_)
  );
  INV_X1 _17074_ (
    .A(_07029_),
    .ZN(_07031_)
  );
  AND2_X1 _17075_ (
    .A1(_06721_),
    .A2(_07026_),
    .ZN(_07032_)
  );
  INV_X1 _17076_ (
    .A(_07032_),
    .ZN(_07033_)
  );
  AND2_X1 _17077_ (
    .A1(_07031_),
    .A2(_07033_),
    .ZN(_07034_)
  );
  INV_X1 _17078_ (
    .A(_07034_),
    .ZN(_07035_)
  );
  AND2_X1 _17079_ (
    .A1(_06716_),
    .A2(_07034_),
    .ZN(_07036_)
  );
  INV_X1 _17080_ (
    .A(_07036_),
    .ZN(_07037_)
  );
  AND2_X1 _17081_ (
    .A1(_06717_),
    .A2(_07035_),
    .ZN(_07038_)
  );
  INV_X1 _17082_ (
    .A(_07038_),
    .ZN(_07039_)
  );
  AND2_X1 _17083_ (
    .A1(_07037_),
    .A2(_07039_),
    .ZN(_07040_)
  );
  INV_X1 _17084_ (
    .A(_07040_),
    .ZN(_07042_)
  );
  AND2_X1 _17085_ (
    .A1(_07023_),
    .A2(_07040_),
    .ZN(_07043_)
  );
  INV_X1 _17086_ (
    .A(_07043_),
    .ZN(_07044_)
  );
  AND2_X1 _17087_ (
    .A1(_07022_),
    .A2(_07042_),
    .ZN(_07045_)
  );
  INV_X1 _17088_ (
    .A(_07045_),
    .ZN(_07046_)
  );
  AND2_X1 _17089_ (
    .A1(_07044_),
    .A2(_07046_),
    .ZN(_07047_)
  );
  INV_X1 _17090_ (
    .A(_07047_),
    .ZN(_07048_)
  );
  AND2_X1 _17091_ (
    .A1(_07021_),
    .A2(_07047_),
    .ZN(_07049_)
  );
  INV_X1 _17092_ (
    .A(_07049_),
    .ZN(_07050_)
  );
  AND2_X1 _17093_ (
    .A1(_07020_),
    .A2(_07048_),
    .ZN(_07051_)
  );
  INV_X1 _17094_ (
    .A(_07051_),
    .ZN(_07053_)
  );
  AND2_X1 _17095_ (
    .A1(_07050_),
    .A2(_07053_),
    .ZN(_07054_)
  );
  INV_X1 _17096_ (
    .A(_07054_),
    .ZN(_07055_)
  );
  AND2_X1 _17097_ (
    .A1(_07018_),
    .A2(_07054_),
    .ZN(_07056_)
  );
  INV_X1 _17098_ (
    .A(_07056_),
    .ZN(_07057_)
  );
  AND2_X1 _17099_ (
    .A1(_07017_),
    .A2(_07055_),
    .ZN(_07058_)
  );
  INV_X1 _17100_ (
    .A(_07058_),
    .ZN(_07059_)
  );
  AND2_X1 _17101_ (
    .A1(_07057_),
    .A2(_07059_),
    .ZN(_07060_)
  );
  INV_X1 _17102_ (
    .A(_07060_),
    .ZN(_07061_)
  );
  AND2_X1 _17103_ (
    .A1(_07016_),
    .A2(_07060_),
    .ZN(_07062_)
  );
  INV_X1 _17104_ (
    .A(_07062_),
    .ZN(_07064_)
  );
  AND2_X1 _17105_ (
    .A1(_07015_),
    .A2(_07061_),
    .ZN(_07065_)
  );
  INV_X1 _17106_ (
    .A(_07065_),
    .ZN(_07066_)
  );
  AND2_X1 _17107_ (
    .A1(_07064_),
    .A2(_07066_),
    .ZN(_07067_)
  );
  INV_X1 _17108_ (
    .A(_07067_),
    .ZN(_07068_)
  );
  AND2_X1 _17109_ (
    .A1(_07014_),
    .A2(_07067_),
    .ZN(_07069_)
  );
  INV_X1 _17110_ (
    .A(_07069_),
    .ZN(_07070_)
  );
  AND2_X1 _17111_ (
    .A1(_07013_),
    .A2(_07068_),
    .ZN(_07071_)
  );
  INV_X1 _17112_ (
    .A(_07071_),
    .ZN(_07072_)
  );
  AND2_X1 _17113_ (
    .A1(_07070_),
    .A2(_07072_),
    .ZN(_07073_)
  );
  INV_X1 _17114_ (
    .A(_07073_),
    .ZN(_07075_)
  );
  AND2_X1 _17115_ (
    .A1(_06772_),
    .A2(_06778_),
    .ZN(_07076_)
  );
  INV_X1 _17116_ (
    .A(_07076_),
    .ZN(_07077_)
  );
  AND2_X1 _17117_ (
    .A1(_05813_),
    .A2(_07076_),
    .ZN(_07078_)
  );
  INV_X1 _17118_ (
    .A(_07078_),
    .ZN(_07079_)
  );
  AND2_X1 _17119_ (
    .A1(_05814_),
    .A2(_07077_),
    .ZN(_07080_)
  );
  INV_X1 _17120_ (
    .A(_07080_),
    .ZN(_07081_)
  );
  AND2_X1 _17121_ (
    .A1(_07079_),
    .A2(_07081_),
    .ZN(_07082_)
  );
  INV_X1 _17122_ (
    .A(_07082_),
    .ZN(_07083_)
  );
  AND2_X1 _17123_ (
    .A1(_07073_),
    .A2(_07082_),
    .ZN(_07084_)
  );
  INV_X1 _17124_ (
    .A(_07084_),
    .ZN(_07086_)
  );
  AND2_X1 _17125_ (
    .A1(_07075_),
    .A2(_07083_),
    .ZN(_07087_)
  );
  INV_X1 _17126_ (
    .A(_07087_),
    .ZN(_07088_)
  );
  AND2_X1 _17127_ (
    .A1(_07086_),
    .A2(_07088_),
    .ZN(_07089_)
  );
  INV_X1 _17128_ (
    .A(_07089_),
    .ZN(_07090_)
  );
  AND2_X1 _17129_ (
    .A1(_07012_),
    .A2(_07089_),
    .ZN(_07091_)
  );
  INV_X1 _17130_ (
    .A(_07091_),
    .ZN(_07092_)
  );
  AND2_X1 _17131_ (
    .A1(_07011_),
    .A2(_07090_),
    .ZN(_07093_)
  );
  INV_X1 _17132_ (
    .A(_07093_),
    .ZN(_07094_)
  );
  AND2_X1 _17133_ (
    .A1(_07092_),
    .A2(_07094_),
    .ZN(_07095_)
  );
  INV_X1 _17134_ (
    .A(_07095_),
    .ZN(_07097_)
  );
  AND2_X1 _17135_ (
    .A1(divisor[25]),
    .A2(remainder[0]),
    .ZN(_07098_)
  );
  INV_X1 _17136_ (
    .A(_07098_),
    .ZN(_07099_)
  );
  AND2_X1 _17137_ (
    .A1(_06809_),
    .A2(_06816_),
    .ZN(_07100_)
  );
  INV_X1 _17138_ (
    .A(_07100_),
    .ZN(_07101_)
  );
  AND2_X1 _17139_ (
    .A1(divisor[22]),
    .A2(remainder[3]),
    .ZN(_07102_)
  );
  INV_X1 _17140_ (
    .A(_07102_),
    .ZN(_07103_)
  );
  AND2_X1 _17141_ (
    .A1(divisor[23]),
    .A2(remainder[2]),
    .ZN(_07104_)
  );
  INV_X1 _17142_ (
    .A(_07104_),
    .ZN(_07105_)
  );
  AND2_X1 _17143_ (
    .A1(divisor[24]),
    .A2(remainder[2]),
    .ZN(_07106_)
  );
  INV_X1 _17144_ (
    .A(_07106_),
    .ZN(_07108_)
  );
  AND2_X1 _17145_ (
    .A1(_06518_),
    .A2(_07106_),
    .ZN(_07109_)
  );
  INV_X1 _17146_ (
    .A(_07109_),
    .ZN(_07110_)
  );
  AND2_X1 _17147_ (
    .A1(_06807_),
    .A2(_07105_),
    .ZN(_07111_)
  );
  INV_X1 _17148_ (
    .A(_07111_),
    .ZN(_07112_)
  );
  AND2_X1 _17149_ (
    .A1(_07110_),
    .A2(_07112_),
    .ZN(_07113_)
  );
  INV_X1 _17150_ (
    .A(_07113_),
    .ZN(_07114_)
  );
  AND2_X1 _17151_ (
    .A1(_07102_),
    .A2(_07113_),
    .ZN(_07115_)
  );
  INV_X1 _17152_ (
    .A(_07115_),
    .ZN(_07116_)
  );
  AND2_X1 _17153_ (
    .A1(_07103_),
    .A2(_07114_),
    .ZN(_07117_)
  );
  INV_X1 _17154_ (
    .A(_07117_),
    .ZN(_07119_)
  );
  AND2_X1 _17155_ (
    .A1(_07116_),
    .A2(_07119_),
    .ZN(_07120_)
  );
  INV_X1 _17156_ (
    .A(_07120_),
    .ZN(_07121_)
  );
  AND2_X1 _17157_ (
    .A1(_07101_),
    .A2(_07120_),
    .ZN(_07122_)
  );
  INV_X1 _17158_ (
    .A(_07122_),
    .ZN(_07123_)
  );
  AND2_X1 _17159_ (
    .A1(_07100_),
    .A2(_07121_),
    .ZN(_07124_)
  );
  INV_X1 _17160_ (
    .A(_07124_),
    .ZN(_07125_)
  );
  AND2_X1 _17161_ (
    .A1(_07123_),
    .A2(_07125_),
    .ZN(_07126_)
  );
  INV_X1 _17162_ (
    .A(_07126_),
    .ZN(_07127_)
  );
  AND2_X1 _17163_ (
    .A1(divisor[19]),
    .A2(remainder[6]),
    .ZN(_07128_)
  );
  INV_X1 _17164_ (
    .A(_07128_),
    .ZN(_07130_)
  );
  AND2_X1 _17165_ (
    .A1(divisor[20]),
    .A2(remainder[5]),
    .ZN(_07131_)
  );
  INV_X1 _17166_ (
    .A(_07131_),
    .ZN(_07132_)
  );
  AND2_X1 _17167_ (
    .A1(divisor[21]),
    .A2(remainder[5]),
    .ZN(_07133_)
  );
  INV_X1 _17168_ (
    .A(_07133_),
    .ZN(_07134_)
  );
  AND2_X1 _17169_ (
    .A1(_06831_),
    .A2(_07131_),
    .ZN(_07135_)
  );
  INV_X1 _17170_ (
    .A(_07135_),
    .ZN(_07136_)
  );
  AND2_X1 _17171_ (
    .A1(_06832_),
    .A2(_07132_),
    .ZN(_07137_)
  );
  INV_X1 _17172_ (
    .A(_07137_),
    .ZN(_07138_)
  );
  AND2_X1 _17173_ (
    .A1(_07136_),
    .A2(_07138_),
    .ZN(_07139_)
  );
  INV_X1 _17174_ (
    .A(_07139_),
    .ZN(_07141_)
  );
  AND2_X1 _17175_ (
    .A1(_07128_),
    .A2(_07139_),
    .ZN(_07142_)
  );
  INV_X1 _17176_ (
    .A(_07142_),
    .ZN(_07143_)
  );
  AND2_X1 _17177_ (
    .A1(_07130_),
    .A2(_07141_),
    .ZN(_07144_)
  );
  INV_X1 _17178_ (
    .A(_07144_),
    .ZN(_07145_)
  );
  AND2_X1 _17179_ (
    .A1(_07143_),
    .A2(_07145_),
    .ZN(_07146_)
  );
  INV_X1 _17180_ (
    .A(_07146_),
    .ZN(_07147_)
  );
  AND2_X1 _17181_ (
    .A1(_07126_),
    .A2(_07146_),
    .ZN(_07148_)
  );
  INV_X1 _17182_ (
    .A(_07148_),
    .ZN(_07149_)
  );
  AND2_X1 _17183_ (
    .A1(_07127_),
    .A2(_07147_),
    .ZN(_07150_)
  );
  INV_X1 _17184_ (
    .A(_07150_),
    .ZN(_07152_)
  );
  AND2_X1 _17185_ (
    .A1(_07149_),
    .A2(_07152_),
    .ZN(_07153_)
  );
  INV_X1 _17186_ (
    .A(_07153_),
    .ZN(_07154_)
  );
  AND2_X1 _17187_ (
    .A1(_07098_),
    .A2(_07153_),
    .ZN(_07155_)
  );
  INV_X1 _17188_ (
    .A(_07155_),
    .ZN(_07156_)
  );
  AND2_X1 _17189_ (
    .A1(_07099_),
    .A2(_07154_),
    .ZN(_07157_)
  );
  INV_X1 _17190_ (
    .A(_07157_),
    .ZN(_07158_)
  );
  AND2_X1 _17191_ (
    .A1(_07156_),
    .A2(_07158_),
    .ZN(_07159_)
  );
  INV_X1 _17192_ (
    .A(_07159_),
    .ZN(_07160_)
  );
  AND2_X1 _17193_ (
    .A1(_07005_),
    .A2(_07160_),
    .ZN(_07161_)
  );
  INV_X1 _17194_ (
    .A(_07161_),
    .ZN(_07163_)
  );
  AND2_X1 _17195_ (
    .A1(_07004_),
    .A2(_07159_),
    .ZN(_07164_)
  );
  INV_X1 _17196_ (
    .A(_07164_),
    .ZN(_07165_)
  );
  AND2_X1 _17197_ (
    .A1(_07005_),
    .A2(_07159_),
    .ZN(_07166_)
  );
  INV_X1 _17198_ (
    .A(_07166_),
    .ZN(_07167_)
  );
  AND2_X1 _17199_ (
    .A1(_07004_),
    .A2(_07160_),
    .ZN(_07168_)
  );
  INV_X1 _17200_ (
    .A(_07168_),
    .ZN(_07169_)
  );
  AND2_X1 _17201_ (
    .A1(_07163_),
    .A2(_07165_),
    .ZN(_07170_)
  );
  AND2_X1 _17202_ (
    .A1(_07167_),
    .A2(_07169_),
    .ZN(_07171_)
  );
  AND2_X1 _17203_ (
    .A1(_07095_),
    .A2(_07170_),
    .ZN(_07172_)
  );
  INV_X1 _17204_ (
    .A(_07172_),
    .ZN(_07174_)
  );
  AND2_X1 _17205_ (
    .A1(_07097_),
    .A2(_07171_),
    .ZN(_07175_)
  );
  INV_X1 _17206_ (
    .A(_07175_),
    .ZN(_07176_)
  );
  AND2_X1 _17207_ (
    .A1(_07174_),
    .A2(_07176_),
    .ZN(_07177_)
  );
  INV_X1 _17208_ (
    .A(_07177_),
    .ZN(_07178_)
  );
  AND2_X1 _17209_ (
    .A1(_07010_),
    .A2(_07177_),
    .ZN(_07179_)
  );
  INV_X1 _17210_ (
    .A(_07179_),
    .ZN(_07180_)
  );
  AND2_X1 _17211_ (
    .A1(_07009_),
    .A2(_07178_),
    .ZN(_07181_)
  );
  INV_X1 _17212_ (
    .A(_07181_),
    .ZN(_07182_)
  );
  AND2_X1 _17213_ (
    .A1(_07180_),
    .A2(_07182_),
    .ZN(_07183_)
  );
  INV_X1 _17214_ (
    .A(_07183_),
    .ZN(_07185_)
  );
  AND2_X1 _17215_ (
    .A1(_06898_),
    .A2(_06905_),
    .ZN(_07186_)
  );
  INV_X1 _17216_ (
    .A(_07186_),
    .ZN(_07187_)
  );
  AND2_X1 _17217_ (
    .A1(_06885_),
    .A2(_06892_),
    .ZN(_07188_)
  );
  INV_X1 _17218_ (
    .A(_07188_),
    .ZN(_07189_)
  );
  AND2_X1 _17219_ (
    .A1(_06778_),
    .A2(_06783_),
    .ZN(_07190_)
  );
  INV_X1 _17220_ (
    .A(_07190_),
    .ZN(_07191_)
  );
  AND2_X1 _17221_ (
    .A1(_06266_),
    .A2(_07191_),
    .ZN(_07192_)
  );
  INV_X1 _17222_ (
    .A(_07192_),
    .ZN(_07193_)
  );
  AND2_X1 _17223_ (
    .A1(_06268_),
    .A2(_07190_),
    .ZN(_07194_)
  );
  INV_X1 _17224_ (
    .A(_07194_),
    .ZN(_07196_)
  );
  AND2_X1 _17225_ (
    .A1(_07193_),
    .A2(_07196_),
    .ZN(_07197_)
  );
  INV_X1 _17226_ (
    .A(_07197_),
    .ZN(_07198_)
  );
  AND2_X1 _17227_ (
    .A1(_06581_),
    .A2(_07197_),
    .ZN(_07199_)
  );
  INV_X1 _17228_ (
    .A(_07199_),
    .ZN(_07200_)
  );
  AND2_X1 _17229_ (
    .A1(_06580_),
    .A2(_07198_),
    .ZN(_07201_)
  );
  INV_X1 _17230_ (
    .A(_07201_),
    .ZN(_07202_)
  );
  AND2_X1 _17231_ (
    .A1(_07200_),
    .A2(_07202_),
    .ZN(_07203_)
  );
  INV_X1 _17232_ (
    .A(_07203_),
    .ZN(_07204_)
  );
  AND2_X1 _17233_ (
    .A1(_07189_),
    .A2(_07203_),
    .ZN(_07205_)
  );
  INV_X1 _17234_ (
    .A(_07205_),
    .ZN(_07207_)
  );
  AND2_X1 _17235_ (
    .A1(_07188_),
    .A2(_07204_),
    .ZN(_07208_)
  );
  INV_X1 _17236_ (
    .A(_07208_),
    .ZN(_07209_)
  );
  AND2_X1 _17237_ (
    .A1(_07207_),
    .A2(_07209_),
    .ZN(_07210_)
  );
  INV_X1 _17238_ (
    .A(_07210_),
    .ZN(_07211_)
  );
  AND2_X1 _17239_ (
    .A1(_03170_),
    .A2(_07210_),
    .ZN(_07212_)
  );
  INV_X1 _17240_ (
    .A(_07212_),
    .ZN(_07213_)
  );
  AND2_X1 _17241_ (
    .A1(_03169_),
    .A2(_07211_),
    .ZN(_07214_)
  );
  INV_X1 _17242_ (
    .A(_07214_),
    .ZN(_07215_)
  );
  AND2_X1 _17243_ (
    .A1(_07213_),
    .A2(_07215_),
    .ZN(_07216_)
  );
  INV_X1 _17244_ (
    .A(_07216_),
    .ZN(_07218_)
  );
  AND2_X1 _17245_ (
    .A1(_06795_),
    .A2(_07216_),
    .ZN(_07219_)
  );
  INV_X1 _17246_ (
    .A(_07219_),
    .ZN(_07220_)
  );
  AND2_X1 _17247_ (
    .A1(_06796_),
    .A2(_07218_),
    .ZN(_07221_)
  );
  INV_X1 _17248_ (
    .A(_07221_),
    .ZN(_07222_)
  );
  AND2_X1 _17249_ (
    .A1(_07220_),
    .A2(_07222_),
    .ZN(_07223_)
  );
  INV_X1 _17250_ (
    .A(_07223_),
    .ZN(_07224_)
  );
  AND2_X1 _17251_ (
    .A1(_07187_),
    .A2(_07223_),
    .ZN(_07225_)
  );
  INV_X1 _17252_ (
    .A(_07225_),
    .ZN(_07226_)
  );
  AND2_X1 _17253_ (
    .A1(_07186_),
    .A2(_07224_),
    .ZN(_07227_)
  );
  INV_X1 _17254_ (
    .A(_07227_),
    .ZN(_07229_)
  );
  AND2_X1 _17255_ (
    .A1(_07226_),
    .A2(_07229_),
    .ZN(_07230_)
  );
  INV_X1 _17256_ (
    .A(_07230_),
    .ZN(_07231_)
  );
  AND2_X1 _17257_ (
    .A1(_07183_),
    .A2(_07230_),
    .ZN(_07232_)
  );
  INV_X1 _17258_ (
    .A(_07232_),
    .ZN(_07233_)
  );
  AND2_X1 _17259_ (
    .A1(_07185_),
    .A2(_07231_),
    .ZN(_07234_)
  );
  INV_X1 _17260_ (
    .A(_07234_),
    .ZN(_07235_)
  );
  AND2_X1 _17261_ (
    .A1(_07233_),
    .A2(_07235_),
    .ZN(_07236_)
  );
  INV_X1 _17262_ (
    .A(_07236_),
    .ZN(_07237_)
  );
  AND2_X1 _17263_ (
    .A1(_07003_),
    .A2(_07236_),
    .ZN(_07238_)
  );
  INV_X1 _17264_ (
    .A(_07238_),
    .ZN(_07240_)
  );
  AND2_X1 _17265_ (
    .A1(_07002_),
    .A2(_07237_),
    .ZN(_07241_)
  );
  INV_X1 _17266_ (
    .A(_07241_),
    .ZN(_07242_)
  );
  AND2_X1 _17267_ (
    .A1(_07240_),
    .A2(_07242_),
    .ZN(_07243_)
  );
  INV_X1 _17268_ (
    .A(_07243_),
    .ZN(_07244_)
  );
  AND2_X1 _17269_ (
    .A1(_07001_),
    .A2(_07243_),
    .ZN(_07245_)
  );
  INV_X1 _17270_ (
    .A(_07245_),
    .ZN(_07246_)
  );
  AND2_X1 _17271_ (
    .A1(_07000_),
    .A2(_07244_),
    .ZN(_07247_)
  );
  INV_X1 _17272_ (
    .A(_07247_),
    .ZN(_07248_)
  );
  AND2_X1 _17273_ (
    .A1(_07246_),
    .A2(_07248_),
    .ZN(_07249_)
  );
  INV_X1 _17274_ (
    .A(_07249_),
    .ZN(_07251_)
  );
  AND2_X1 _17275_ (
    .A1(_06999_),
    .A2(_07249_),
    .ZN(_07252_)
  );
  INV_X1 _17276_ (
    .A(_07252_),
    .ZN(_07253_)
  );
  AND2_X1 _17277_ (
    .A1(_06998_),
    .A2(_07251_),
    .ZN(_07254_)
  );
  INV_X1 _17278_ (
    .A(_07254_),
    .ZN(_07255_)
  );
  AND2_X1 _17279_ (
    .A1(_07253_),
    .A2(_07255_),
    .ZN(_07256_)
  );
  INV_X1 _17280_ (
    .A(_07256_),
    .ZN(_07257_)
  );
  AND2_X1 _17281_ (
    .A1(_06944_),
    .A2(_07256_),
    .ZN(_07258_)
  );
  INV_X1 _17282_ (
    .A(_07258_),
    .ZN(_07259_)
  );
  AND2_X1 _17283_ (
    .A1(_06945_),
    .A2(_07257_),
    .ZN(_07260_)
  );
  INV_X1 _17284_ (
    .A(_07260_),
    .ZN(_07262_)
  );
  AND2_X1 _17285_ (
    .A1(_07259_),
    .A2(_07262_),
    .ZN(_07263_)
  );
  INV_X1 _17286_ (
    .A(_07263_),
    .ZN(_07264_)
  );
  AND2_X1 _17287_ (
    .A1(_06995_),
    .A2(_07264_),
    .ZN(_07265_)
  );
  INV_X1 _17288_ (
    .A(_07265_),
    .ZN(_07266_)
  );
  AND2_X1 _17289_ (
    .A1(_06996_),
    .A2(_07263_),
    .ZN(_07267_)
  );
  INV_X1 _17290_ (
    .A(_07267_),
    .ZN(_07268_)
  );
  AND2_X1 _17291_ (
    .A1(_07266_),
    .A2(_07268_),
    .ZN(_07269_)
  );
  INV_X1 _17292_ (
    .A(_07269_),
    .ZN(_07270_)
  );
  AND2_X1 _17293_ (
    .A1(remainder[58]),
    .A2(_07269_),
    .ZN(_07271_)
  );
  INV_X1 _17294_ (
    .A(_07271_),
    .ZN(_07273_)
  );
  AND2_X1 _17295_ (
    .A1(_04481_),
    .A2(_07270_),
    .ZN(_07274_)
  );
  INV_X1 _17296_ (
    .A(_07274_),
    .ZN(_07275_)
  );
  AND2_X1 _17297_ (
    .A1(_07273_),
    .A2(_07275_),
    .ZN(_07276_)
  );
  INV_X1 _17298_ (
    .A(_07276_),
    .ZN(_07277_)
  );
  AND2_X1 _17299_ (
    .A1(_06993_),
    .A2(_07277_),
    .ZN(_07278_)
  );
  INV_X1 _17300_ (
    .A(_07278_),
    .ZN(_07279_)
  );
  AND2_X1 _17301_ (
    .A1(_06994_),
    .A2(_07276_),
    .ZN(_07280_)
  );
  INV_X1 _17302_ (
    .A(_07280_),
    .ZN(_07281_)
  );
  AND2_X1 _17303_ (
    .A1(_02082_),
    .A2(_07281_),
    .ZN(_07282_)
  );
  AND2_X1 _17304_ (
    .A1(_07279_),
    .A2(_07282_),
    .ZN(_07284_)
  );
  INV_X1 _17305_ (
    .A(_07284_),
    .ZN(_07285_)
  );
  AND2_X1 _17306_ (
    .A1(_06990_),
    .A2(_07285_),
    .ZN(_07286_)
  );
  AND2_X1 _17307_ (
    .A1(_06992_),
    .A2(_07286_),
    .ZN(_07287_)
  );
  INV_X1 _17308_ (
    .A(_07287_),
    .ZN(_07288_)
  );
  AND2_X1 _17309_ (
    .A1(_06201_),
    .A2(_07288_),
    .ZN(_00071_)
  );
  AND2_X1 _17310_ (
    .A1(_07240_),
    .A2(_07246_),
    .ZN(_07289_)
  );
  INV_X1 _17311_ (
    .A(_07289_),
    .ZN(_07290_)
  );
  AND2_X1 _17312_ (
    .A1(_07220_),
    .A2(_07226_),
    .ZN(_07291_)
  );
  INV_X1 _17313_ (
    .A(_07291_),
    .ZN(_07292_)
  );
  AND2_X1 _17314_ (
    .A1(_07180_),
    .A2(_07233_),
    .ZN(_07294_)
  );
  INV_X1 _17315_ (
    .A(_07294_),
    .ZN(_07295_)
  );
  AND2_X1 _17316_ (
    .A1(_03249_),
    .A2(_07160_),
    .ZN(_07296_)
  );
  INV_X1 _17317_ (
    .A(_07296_),
    .ZN(_07297_)
  );
  AND2_X1 _17318_ (
    .A1(_06851_),
    .A2(_07296_),
    .ZN(_07298_)
  );
  INV_X1 _17319_ (
    .A(_07298_),
    .ZN(_07299_)
  );
  AND2_X1 _17320_ (
    .A1(_07174_),
    .A2(_07299_),
    .ZN(_07300_)
  );
  INV_X1 _17321_ (
    .A(_07300_),
    .ZN(_07301_)
  );
  AND2_X1 _17322_ (
    .A1(_07070_),
    .A2(_07086_),
    .ZN(_07302_)
  );
  INV_X1 _17323_ (
    .A(_07302_),
    .ZN(_07303_)
  );
  AND2_X1 _17324_ (
    .A1(_07057_),
    .A2(_07064_),
    .ZN(_07305_)
  );
  INV_X1 _17325_ (
    .A(_07305_),
    .ZN(_07306_)
  );
  AND2_X1 _17326_ (
    .A1(_07044_),
    .A2(_07050_),
    .ZN(_07307_)
  );
  INV_X1 _17327_ (
    .A(_07307_),
    .ZN(_07308_)
  );
  AND2_X1 _17328_ (
    .A1(_07123_),
    .A2(_07149_),
    .ZN(_07309_)
  );
  INV_X1 _17329_ (
    .A(_07309_),
    .ZN(_07310_)
  );
  AND2_X1 _17330_ (
    .A1(_07031_),
    .A2(_07037_),
    .ZN(_07311_)
  );
  INV_X1 _17331_ (
    .A(_07311_),
    .ZN(_07312_)
  );
  AND2_X1 _17332_ (
    .A1(_07136_),
    .A2(_07143_),
    .ZN(_07313_)
  );
  INV_X1 _17333_ (
    .A(_07313_),
    .ZN(_07314_)
  );
  MUX2_X1 _17334_ (
    .A(_07025_),
    .B(_04974_),
    .S(_07024_),
    .Z(_07316_)
  );
  AND2_X1 _17335_ (
    .A1(divisor[16]),
    .A2(_07316_),
    .ZN(_07317_)
  );
  INV_X1 _17336_ (
    .A(_07317_),
    .ZN(_07318_)
  );
  MUX2_X1 _17337_ (
    .A(_06716_),
    .B(_04963_),
    .S(_07316_),
    .Z(_07319_)
  );
  MUX2_X1 _17338_ (
    .A(_06717_),
    .B(divisor[16]),
    .S(_07316_),
    .Z(_07320_)
  );
  AND2_X1 _17339_ (
    .A1(_07314_),
    .A2(_07319_),
    .ZN(_07321_)
  );
  INV_X1 _17340_ (
    .A(_07321_),
    .ZN(_07322_)
  );
  AND2_X1 _17341_ (
    .A1(_07313_),
    .A2(_07320_),
    .ZN(_07323_)
  );
  INV_X1 _17342_ (
    .A(_07323_),
    .ZN(_07324_)
  );
  AND2_X1 _17343_ (
    .A1(_07322_),
    .A2(_07324_),
    .ZN(_07325_)
  );
  INV_X1 _17344_ (
    .A(_07325_),
    .ZN(_07327_)
  );
  AND2_X1 _17345_ (
    .A1(_07312_),
    .A2(_07325_),
    .ZN(_07328_)
  );
  INV_X1 _17346_ (
    .A(_07328_),
    .ZN(_07329_)
  );
  AND2_X1 _17347_ (
    .A1(_07311_),
    .A2(_07327_),
    .ZN(_07330_)
  );
  INV_X1 _17348_ (
    .A(_07330_),
    .ZN(_07331_)
  );
  AND2_X1 _17349_ (
    .A1(_07329_),
    .A2(_07331_),
    .ZN(_07332_)
  );
  INV_X1 _17350_ (
    .A(_07332_),
    .ZN(_07333_)
  );
  AND2_X1 _17351_ (
    .A1(_07310_),
    .A2(_07332_),
    .ZN(_07334_)
  );
  INV_X1 _17352_ (
    .A(_07334_),
    .ZN(_07335_)
  );
  AND2_X1 _17353_ (
    .A1(_07309_),
    .A2(_07333_),
    .ZN(_07336_)
  );
  INV_X1 _17354_ (
    .A(_07336_),
    .ZN(_07338_)
  );
  AND2_X1 _17355_ (
    .A1(_07335_),
    .A2(_07338_),
    .ZN(_07339_)
  );
  INV_X1 _17356_ (
    .A(_07339_),
    .ZN(_07340_)
  );
  AND2_X1 _17357_ (
    .A1(_07308_),
    .A2(_07339_),
    .ZN(_07341_)
  );
  INV_X1 _17358_ (
    .A(_07341_),
    .ZN(_07342_)
  );
  AND2_X1 _17359_ (
    .A1(_07307_),
    .A2(_07340_),
    .ZN(_07343_)
  );
  INV_X1 _17360_ (
    .A(_07343_),
    .ZN(_07344_)
  );
  AND2_X1 _17361_ (
    .A1(_07342_),
    .A2(_07344_),
    .ZN(_07345_)
  );
  INV_X1 _17362_ (
    .A(_07345_),
    .ZN(_07346_)
  );
  AND2_X1 _17363_ (
    .A1(_07306_),
    .A2(_07345_),
    .ZN(_07347_)
  );
  INV_X1 _17364_ (
    .A(_07347_),
    .ZN(_07349_)
  );
  AND2_X1 _17365_ (
    .A1(_07305_),
    .A2(_07346_),
    .ZN(_07350_)
  );
  INV_X1 _17366_ (
    .A(_07350_),
    .ZN(_07351_)
  );
  AND2_X1 _17367_ (
    .A1(_07349_),
    .A2(_07351_),
    .ZN(_07352_)
  );
  INV_X1 _17368_ (
    .A(_07352_),
    .ZN(_07353_)
  );
  AND2_X1 _17369_ (
    .A1(_07082_),
    .A2(_07352_),
    .ZN(_07354_)
  );
  INV_X1 _17370_ (
    .A(_07354_),
    .ZN(_07355_)
  );
  AND2_X1 _17371_ (
    .A1(_07083_),
    .A2(_07353_),
    .ZN(_07356_)
  );
  INV_X1 _17372_ (
    .A(_07356_),
    .ZN(_07357_)
  );
  AND2_X1 _17373_ (
    .A1(_07355_),
    .A2(_07357_),
    .ZN(_07358_)
  );
  INV_X1 _17374_ (
    .A(_07358_),
    .ZN(_07360_)
  );
  AND2_X1 _17375_ (
    .A1(_07303_),
    .A2(_07358_),
    .ZN(_07361_)
  );
  INV_X1 _17376_ (
    .A(_07361_),
    .ZN(_07362_)
  );
  AND2_X1 _17377_ (
    .A1(_07302_),
    .A2(_07360_),
    .ZN(_07363_)
  );
  INV_X1 _17378_ (
    .A(_07363_),
    .ZN(_07364_)
  );
  AND2_X1 _17379_ (
    .A1(_07362_),
    .A2(_07364_),
    .ZN(_07365_)
  );
  INV_X1 _17380_ (
    .A(_07365_),
    .ZN(_07366_)
  );
  AND2_X1 _17381_ (
    .A1(divisor[26]),
    .A2(remainder[0]),
    .ZN(_07367_)
  );
  INV_X1 _17382_ (
    .A(_07367_),
    .ZN(_07368_)
  );
  AND2_X1 _17383_ (
    .A1(divisor[25]),
    .A2(remainder[1]),
    .ZN(_07369_)
  );
  INV_X1 _17384_ (
    .A(_07369_),
    .ZN(_07371_)
  );
  AND2_X1 _17385_ (
    .A1(divisor[26]),
    .A2(remainder[1]),
    .ZN(_07372_)
  );
  INV_X1 _17386_ (
    .A(_07372_),
    .ZN(_07373_)
  );
  AND2_X1 _17387_ (
    .A1(_07098_),
    .A2(_07372_),
    .ZN(_07374_)
  );
  INV_X1 _17388_ (
    .A(_07374_),
    .ZN(_07375_)
  );
  AND2_X1 _17389_ (
    .A1(_07368_),
    .A2(_07371_),
    .ZN(_07376_)
  );
  INV_X1 _17390_ (
    .A(_07376_),
    .ZN(_07377_)
  );
  AND2_X1 _17391_ (
    .A1(_07375_),
    .A2(_07377_),
    .ZN(_07378_)
  );
  INV_X1 _17392_ (
    .A(_07378_),
    .ZN(_07379_)
  );
  AND2_X1 _17393_ (
    .A1(_07110_),
    .A2(_07116_),
    .ZN(_07380_)
  );
  INV_X1 _17394_ (
    .A(_07380_),
    .ZN(_07382_)
  );
  AND2_X1 _17395_ (
    .A1(divisor[22]),
    .A2(remainder[4]),
    .ZN(_07383_)
  );
  INV_X1 _17396_ (
    .A(_07383_),
    .ZN(_07384_)
  );
  AND2_X1 _17397_ (
    .A1(divisor[23]),
    .A2(remainder[3]),
    .ZN(_07385_)
  );
  INV_X1 _17398_ (
    .A(_07385_),
    .ZN(_07386_)
  );
  AND2_X1 _17399_ (
    .A1(divisor[24]),
    .A2(remainder[3]),
    .ZN(_07387_)
  );
  INV_X1 _17400_ (
    .A(_07387_),
    .ZN(_07388_)
  );
  AND2_X1 _17401_ (
    .A1(_07106_),
    .A2(_07385_),
    .ZN(_07389_)
  );
  INV_X1 _17402_ (
    .A(_07389_),
    .ZN(_07390_)
  );
  AND2_X1 _17403_ (
    .A1(_07108_),
    .A2(_07386_),
    .ZN(_07391_)
  );
  INV_X1 _17404_ (
    .A(_07391_),
    .ZN(_07393_)
  );
  AND2_X1 _17405_ (
    .A1(_07390_),
    .A2(_07393_),
    .ZN(_07394_)
  );
  INV_X1 _17406_ (
    .A(_07394_),
    .ZN(_07395_)
  );
  AND2_X1 _17407_ (
    .A1(_07383_),
    .A2(_07394_),
    .ZN(_07396_)
  );
  INV_X1 _17408_ (
    .A(_07396_),
    .ZN(_07397_)
  );
  AND2_X1 _17409_ (
    .A1(_07384_),
    .A2(_07395_),
    .ZN(_07398_)
  );
  INV_X1 _17410_ (
    .A(_07398_),
    .ZN(_07399_)
  );
  AND2_X1 _17411_ (
    .A1(_07397_),
    .A2(_07399_),
    .ZN(_07400_)
  );
  INV_X1 _17412_ (
    .A(_07400_),
    .ZN(_07401_)
  );
  AND2_X1 _17413_ (
    .A1(_07382_),
    .A2(_07400_),
    .ZN(_07402_)
  );
  INV_X1 _17414_ (
    .A(_07402_),
    .ZN(_07404_)
  );
  AND2_X1 _17415_ (
    .A1(_07380_),
    .A2(_07401_),
    .ZN(_07405_)
  );
  INV_X1 _17416_ (
    .A(_07405_),
    .ZN(_07406_)
  );
  AND2_X1 _17417_ (
    .A1(_07404_),
    .A2(_07406_),
    .ZN(_07407_)
  );
  INV_X1 _17418_ (
    .A(_07407_),
    .ZN(_07408_)
  );
  AND2_X1 _17419_ (
    .A1(divisor[19]),
    .A2(remainder[7]),
    .ZN(_07409_)
  );
  INV_X1 _17420_ (
    .A(_07409_),
    .ZN(_07410_)
  );
  AND2_X1 _17421_ (
    .A1(divisor[20]),
    .A2(remainder[6]),
    .ZN(_07411_)
  );
  INV_X1 _17422_ (
    .A(_07411_),
    .ZN(_07412_)
  );
  AND2_X1 _17423_ (
    .A1(divisor[21]),
    .A2(remainder[6]),
    .ZN(_07413_)
  );
  INV_X1 _17424_ (
    .A(_07413_),
    .ZN(_07415_)
  );
  AND2_X1 _17425_ (
    .A1(_07133_),
    .A2(_07411_),
    .ZN(_07416_)
  );
  INV_X1 _17426_ (
    .A(_07416_),
    .ZN(_07417_)
  );
  AND2_X1 _17427_ (
    .A1(_07134_),
    .A2(_07412_),
    .ZN(_07418_)
  );
  INV_X1 _17428_ (
    .A(_07418_),
    .ZN(_07419_)
  );
  AND2_X1 _17429_ (
    .A1(_07417_),
    .A2(_07419_),
    .ZN(_07420_)
  );
  INV_X1 _17430_ (
    .A(_07420_),
    .ZN(_07421_)
  );
  AND2_X1 _17431_ (
    .A1(_07409_),
    .A2(_07420_),
    .ZN(_07422_)
  );
  INV_X1 _17432_ (
    .A(_07422_),
    .ZN(_07423_)
  );
  AND2_X1 _17433_ (
    .A1(_07410_),
    .A2(_07421_),
    .ZN(_07424_)
  );
  INV_X1 _17434_ (
    .A(_07424_),
    .ZN(_07426_)
  );
  AND2_X1 _17435_ (
    .A1(_07423_),
    .A2(_07426_),
    .ZN(_07427_)
  );
  INV_X1 _17436_ (
    .A(_07427_),
    .ZN(_07428_)
  );
  AND2_X1 _17437_ (
    .A1(_07407_),
    .A2(_07427_),
    .ZN(_07429_)
  );
  INV_X1 _17438_ (
    .A(_07429_),
    .ZN(_07430_)
  );
  AND2_X1 _17439_ (
    .A1(_07408_),
    .A2(_07428_),
    .ZN(_07431_)
  );
  INV_X1 _17440_ (
    .A(_07431_),
    .ZN(_07432_)
  );
  AND2_X1 _17441_ (
    .A1(_07430_),
    .A2(_07432_),
    .ZN(_07433_)
  );
  INV_X1 _17442_ (
    .A(_07433_),
    .ZN(_07434_)
  );
  AND2_X1 _17443_ (
    .A1(_07378_),
    .A2(_07433_),
    .ZN(_07435_)
  );
  INV_X1 _17444_ (
    .A(_07435_),
    .ZN(_07437_)
  );
  AND2_X1 _17445_ (
    .A1(_07379_),
    .A2(_07434_),
    .ZN(_07438_)
  );
  INV_X1 _17446_ (
    .A(_07438_),
    .ZN(_07439_)
  );
  AND2_X1 _17447_ (
    .A1(_07437_),
    .A2(_07439_),
    .ZN(_07440_)
  );
  INV_X1 _17448_ (
    .A(_07440_),
    .ZN(_07441_)
  );
  AND2_X1 _17449_ (
    .A1(_07155_),
    .A2(_07440_),
    .ZN(_07442_)
  );
  INV_X1 _17450_ (
    .A(_07442_),
    .ZN(_07443_)
  );
  AND2_X1 _17451_ (
    .A1(_07156_),
    .A2(_07441_),
    .ZN(_07444_)
  );
  INV_X1 _17452_ (
    .A(_07444_),
    .ZN(_07445_)
  );
  AND2_X1 _17453_ (
    .A1(_07443_),
    .A2(_07445_),
    .ZN(_07446_)
  );
  INV_X1 _17454_ (
    .A(_07446_),
    .ZN(_07448_)
  );
  AND2_X1 _17455_ (
    .A1(_07296_),
    .A2(_07448_),
    .ZN(_07449_)
  );
  INV_X1 _17456_ (
    .A(_07449_),
    .ZN(_07450_)
  );
  AND2_X1 _17457_ (
    .A1(_07297_),
    .A2(_07446_),
    .ZN(_07451_)
  );
  INV_X1 _17458_ (
    .A(_07451_),
    .ZN(_07452_)
  );
  AND2_X1 _17459_ (
    .A1(_07450_),
    .A2(_07452_),
    .ZN(_07453_)
  );
  INV_X1 _17460_ (
    .A(_07453_),
    .ZN(_07454_)
  );
  AND2_X1 _17461_ (
    .A1(_07365_),
    .A2(_07454_),
    .ZN(_07455_)
  );
  INV_X1 _17462_ (
    .A(_07455_),
    .ZN(_07456_)
  );
  AND2_X1 _17463_ (
    .A1(_07366_),
    .A2(_07453_),
    .ZN(_07457_)
  );
  INV_X1 _17464_ (
    .A(_07457_),
    .ZN(_07459_)
  );
  AND2_X1 _17465_ (
    .A1(_07456_),
    .A2(_07459_),
    .ZN(_07460_)
  );
  INV_X1 _17466_ (
    .A(_07460_),
    .ZN(_07461_)
  );
  AND2_X1 _17467_ (
    .A1(_07301_),
    .A2(_07460_),
    .ZN(_07462_)
  );
  INV_X1 _17468_ (
    .A(_07462_),
    .ZN(_07463_)
  );
  AND2_X1 _17469_ (
    .A1(_07300_),
    .A2(_07461_),
    .ZN(_07464_)
  );
  INV_X1 _17470_ (
    .A(_07464_),
    .ZN(_07465_)
  );
  AND2_X1 _17471_ (
    .A1(_07463_),
    .A2(_07465_),
    .ZN(_07466_)
  );
  INV_X1 _17472_ (
    .A(_07466_),
    .ZN(_07467_)
  );
  AND2_X1 _17473_ (
    .A1(_07207_),
    .A2(_07213_),
    .ZN(_07468_)
  );
  INV_X1 _17474_ (
    .A(_07468_),
    .ZN(_07470_)
  );
  AND2_X1 _17475_ (
    .A1(_07193_),
    .A2(_07200_),
    .ZN(_07471_)
  );
  INV_X1 _17476_ (
    .A(_07471_),
    .ZN(_07472_)
  );
  AND2_X1 _17477_ (
    .A1(_06778_),
    .A2(_07079_),
    .ZN(_07473_)
  );
  INV_X1 _17478_ (
    .A(_07473_),
    .ZN(_07474_)
  );
  AND2_X1 _17479_ (
    .A1(_06266_),
    .A2(_07474_),
    .ZN(_07475_)
  );
  INV_X1 _17480_ (
    .A(_07475_),
    .ZN(_07476_)
  );
  AND2_X1 _17481_ (
    .A1(_06268_),
    .A2(_07473_),
    .ZN(_07477_)
  );
  INV_X1 _17482_ (
    .A(_07477_),
    .ZN(_07478_)
  );
  AND2_X1 _17483_ (
    .A1(_07476_),
    .A2(_07478_),
    .ZN(_07479_)
  );
  INV_X1 _17484_ (
    .A(_07479_),
    .ZN(_07481_)
  );
  AND2_X1 _17485_ (
    .A1(_06580_),
    .A2(_07481_),
    .ZN(_07482_)
  );
  INV_X1 _17486_ (
    .A(_07482_),
    .ZN(_07483_)
  );
  AND2_X1 _17487_ (
    .A1(_06581_),
    .A2(_07479_),
    .ZN(_07484_)
  );
  INV_X1 _17488_ (
    .A(_07484_),
    .ZN(_07485_)
  );
  AND2_X1 _17489_ (
    .A1(_06580_),
    .A2(_07479_),
    .ZN(_07486_)
  );
  INV_X1 _17490_ (
    .A(_07486_),
    .ZN(_07487_)
  );
  AND2_X1 _17491_ (
    .A1(_06581_),
    .A2(_07481_),
    .ZN(_07488_)
  );
  INV_X1 _17492_ (
    .A(_07488_),
    .ZN(_07489_)
  );
  AND2_X1 _17493_ (
    .A1(_07483_),
    .A2(_07485_),
    .ZN(_07490_)
  );
  AND2_X1 _17494_ (
    .A1(_07487_),
    .A2(_07489_),
    .ZN(_07492_)
  );
  AND2_X1 _17495_ (
    .A1(_07472_),
    .A2(_07490_),
    .ZN(_07493_)
  );
  INV_X1 _17496_ (
    .A(_07493_),
    .ZN(_07494_)
  );
  AND2_X1 _17497_ (
    .A1(_07471_),
    .A2(_07492_),
    .ZN(_07495_)
  );
  INV_X1 _17498_ (
    .A(_07495_),
    .ZN(_07496_)
  );
  AND2_X1 _17499_ (
    .A1(_07494_),
    .A2(_07496_),
    .ZN(_07497_)
  );
  INV_X1 _17500_ (
    .A(_07497_),
    .ZN(_07498_)
  );
  AND2_X1 _17501_ (
    .A1(_03170_),
    .A2(_07497_),
    .ZN(_07499_)
  );
  INV_X1 _17502_ (
    .A(_07499_),
    .ZN(_07500_)
  );
  AND2_X1 _17503_ (
    .A1(_03169_),
    .A2(_07498_),
    .ZN(_07501_)
  );
  INV_X1 _17504_ (
    .A(_07501_),
    .ZN(_07503_)
  );
  AND2_X1 _17505_ (
    .A1(_07500_),
    .A2(_07503_),
    .ZN(_07504_)
  );
  INV_X1 _17506_ (
    .A(_07504_),
    .ZN(_07505_)
  );
  AND2_X1 _17507_ (
    .A1(_07091_),
    .A2(_07504_),
    .ZN(_07506_)
  );
  INV_X1 _17508_ (
    .A(_07506_),
    .ZN(_07507_)
  );
  AND2_X1 _17509_ (
    .A1(_07092_),
    .A2(_07505_),
    .ZN(_07508_)
  );
  INV_X1 _17510_ (
    .A(_07508_),
    .ZN(_07509_)
  );
  AND2_X1 _17511_ (
    .A1(_07507_),
    .A2(_07509_),
    .ZN(_07510_)
  );
  INV_X1 _17512_ (
    .A(_07510_),
    .ZN(_07511_)
  );
  AND2_X1 _17513_ (
    .A1(_07470_),
    .A2(_07510_),
    .ZN(_07512_)
  );
  INV_X1 _17514_ (
    .A(_07512_),
    .ZN(_07514_)
  );
  AND2_X1 _17515_ (
    .A1(_07468_),
    .A2(_07511_),
    .ZN(_07515_)
  );
  INV_X1 _17516_ (
    .A(_07515_),
    .ZN(_07516_)
  );
  AND2_X1 _17517_ (
    .A1(_07514_),
    .A2(_07516_),
    .ZN(_07517_)
  );
  INV_X1 _17518_ (
    .A(_07517_),
    .ZN(_07518_)
  );
  AND2_X1 _17519_ (
    .A1(_07466_),
    .A2(_07517_),
    .ZN(_07519_)
  );
  INV_X1 _17520_ (
    .A(_07519_),
    .ZN(_07520_)
  );
  AND2_X1 _17521_ (
    .A1(_07467_),
    .A2(_07518_),
    .ZN(_07521_)
  );
  INV_X1 _17522_ (
    .A(_07521_),
    .ZN(_07522_)
  );
  AND2_X1 _17523_ (
    .A1(_07520_),
    .A2(_07522_),
    .ZN(_07523_)
  );
  INV_X1 _17524_ (
    .A(_07523_),
    .ZN(_07525_)
  );
  AND2_X1 _17525_ (
    .A1(_07295_),
    .A2(_07523_),
    .ZN(_07526_)
  );
  INV_X1 _17526_ (
    .A(_07526_),
    .ZN(_07527_)
  );
  AND2_X1 _17527_ (
    .A1(_07294_),
    .A2(_07525_),
    .ZN(_07528_)
  );
  INV_X1 _17528_ (
    .A(_07528_),
    .ZN(_07529_)
  );
  AND2_X1 _17529_ (
    .A1(_07527_),
    .A2(_07529_),
    .ZN(_07530_)
  );
  INV_X1 _17530_ (
    .A(_07530_),
    .ZN(_07531_)
  );
  AND2_X1 _17531_ (
    .A1(_07292_),
    .A2(_07530_),
    .ZN(_07532_)
  );
  INV_X1 _17532_ (
    .A(_07532_),
    .ZN(_07533_)
  );
  AND2_X1 _17533_ (
    .A1(_07291_),
    .A2(_07531_),
    .ZN(_07534_)
  );
  INV_X1 _17534_ (
    .A(_07534_),
    .ZN(_07536_)
  );
  AND2_X1 _17535_ (
    .A1(_07533_),
    .A2(_07536_),
    .ZN(_07537_)
  );
  INV_X1 _17536_ (
    .A(_07537_),
    .ZN(_07538_)
  );
  AND2_X1 _17537_ (
    .A1(_07290_),
    .A2(_07537_),
    .ZN(_07539_)
  );
  INV_X1 _17538_ (
    .A(_07539_),
    .ZN(_07540_)
  );
  AND2_X1 _17539_ (
    .A1(_07289_),
    .A2(_07538_),
    .ZN(_07541_)
  );
  INV_X1 _17540_ (
    .A(_07541_),
    .ZN(_07542_)
  );
  AND2_X1 _17541_ (
    .A1(_07540_),
    .A2(_07542_),
    .ZN(_07543_)
  );
  INV_X1 _17542_ (
    .A(_07543_),
    .ZN(_07544_)
  );
  AND2_X1 _17543_ (
    .A1(_07252_),
    .A2(_07543_),
    .ZN(_07545_)
  );
  INV_X1 _17544_ (
    .A(_07545_),
    .ZN(_07547_)
  );
  AND2_X1 _17545_ (
    .A1(_07253_),
    .A2(_07544_),
    .ZN(_07548_)
  );
  INV_X1 _17546_ (
    .A(_07548_),
    .ZN(_07549_)
  );
  AND2_X1 _17547_ (
    .A1(_07547_),
    .A2(_07549_),
    .ZN(_07550_)
  );
  INV_X1 _17548_ (
    .A(_07550_),
    .ZN(_07551_)
  );
  AND2_X1 _17549_ (
    .A1(_06995_),
    .A2(_07259_),
    .ZN(_07552_)
  );
  INV_X1 _17550_ (
    .A(_07552_),
    .ZN(_07553_)
  );
  AND2_X1 _17551_ (
    .A1(_07259_),
    .A2(_07268_),
    .ZN(_07554_)
  );
  AND2_X1 _17552_ (
    .A1(_07262_),
    .A2(_07553_),
    .ZN(_07555_)
  );
  AND2_X1 _17553_ (
    .A1(_07550_),
    .A2(_07555_),
    .ZN(_07556_)
  );
  INV_X1 _17554_ (
    .A(_07556_),
    .ZN(_07558_)
  );
  AND2_X1 _17555_ (
    .A1(_07551_),
    .A2(_07554_),
    .ZN(_07559_)
  );
  INV_X1 _17556_ (
    .A(_07559_),
    .ZN(_07560_)
  );
  AND2_X1 _17557_ (
    .A1(_07558_),
    .A2(_07560_),
    .ZN(_07561_)
  );
  INV_X1 _17558_ (
    .A(_07561_),
    .ZN(_07562_)
  );
  AND2_X1 _17559_ (
    .A1(remainder[59]),
    .A2(_07561_),
    .ZN(_07563_)
  );
  INV_X1 _17560_ (
    .A(_07563_),
    .ZN(_07564_)
  );
  AND2_X1 _17561_ (
    .A1(_04470_),
    .A2(_07562_),
    .ZN(_07565_)
  );
  INV_X1 _17562_ (
    .A(_07565_),
    .ZN(_07566_)
  );
  AND2_X1 _17563_ (
    .A1(_07564_),
    .A2(_07566_),
    .ZN(_07567_)
  );
  INV_X1 _17564_ (
    .A(_07567_),
    .ZN(_07569_)
  );
  AND2_X1 _17565_ (
    .A1(_06993_),
    .A2(_07273_),
    .ZN(_07570_)
  );
  INV_X1 _17566_ (
    .A(_07570_),
    .ZN(_07571_)
  );
  AND2_X1 _17567_ (
    .A1(_06994_),
    .A2(_07275_),
    .ZN(_07572_)
  );
  INV_X1 _17568_ (
    .A(_07572_),
    .ZN(_07573_)
  );
  AND2_X1 _17569_ (
    .A1(_07275_),
    .A2(_07571_),
    .ZN(_07574_)
  );
  AND2_X1 _17570_ (
    .A1(_07273_),
    .A2(_07573_),
    .ZN(_07575_)
  );
  AND2_X1 _17571_ (
    .A1(_07567_),
    .A2(_07574_),
    .ZN(_07576_)
  );
  INV_X1 _17572_ (
    .A(_07576_),
    .ZN(_07577_)
  );
  AND2_X1 _17573_ (
    .A1(_07569_),
    .A2(_07575_),
    .ZN(_07578_)
  );
  INV_X1 _17574_ (
    .A(_07578_),
    .ZN(_07580_)
  );
  AND2_X1 _17575_ (
    .A1(_02082_),
    .A2(_07577_),
    .ZN(_07581_)
  );
  AND2_X1 _17576_ (
    .A1(_07580_),
    .A2(_07581_),
    .ZN(_07582_)
  );
  INV_X1 _17577_ (
    .A(_07582_),
    .ZN(_07583_)
  );
  AND2_X1 _17578_ (
    .A1(remainder[51]),
    .A2(_02077_),
    .ZN(_07584_)
  );
  INV_X1 _17579_ (
    .A(_07584_),
    .ZN(_07585_)
  );
  MUX2_X1 _17580_ (
    .A(remainder[50]),
    .B(_01873_),
    .S(_10462_),
    .Z(_07586_)
  );
  AND2_X1 _17581_ (
    .A1(_05983_),
    .A2(_07586_),
    .ZN(_07587_)
  );
  INV_X1 _17582_ (
    .A(_07587_),
    .ZN(_07588_)
  );
  AND2_X1 _17583_ (
    .A1(_07585_),
    .A2(_07588_),
    .ZN(_07589_)
  );
  AND2_X1 _17584_ (
    .A1(_07583_),
    .A2(_07589_),
    .ZN(_07591_)
  );
  INV_X1 _17585_ (
    .A(_07591_),
    .ZN(_07592_)
  );
  AND2_X1 _17586_ (
    .A1(_06201_),
    .A2(_07592_),
    .ZN(_00072_)
  );
  AND2_X1 _17587_ (
    .A1(_07564_),
    .A2(_07577_),
    .ZN(_07593_)
  );
  INV_X1 _17588_ (
    .A(_07593_),
    .ZN(_07594_)
  );
  AND2_X1 _17589_ (
    .A1(_07547_),
    .A2(_07558_),
    .ZN(_07595_)
  );
  INV_X1 _17590_ (
    .A(_07595_),
    .ZN(_07596_)
  );
  AND2_X1 _17591_ (
    .A1(_07527_),
    .A2(_07533_),
    .ZN(_07597_)
  );
  INV_X1 _17592_ (
    .A(_07597_),
    .ZN(_07598_)
  );
  AND2_X1 _17593_ (
    .A1(_07507_),
    .A2(_07514_),
    .ZN(_07599_)
  );
  INV_X1 _17594_ (
    .A(_07599_),
    .ZN(_07601_)
  );
  AND2_X1 _17595_ (
    .A1(_07463_),
    .A2(_07520_),
    .ZN(_07602_)
  );
  INV_X1 _17596_ (
    .A(_07602_),
    .ZN(_07603_)
  );
  AND2_X1 _17597_ (
    .A1(_03249_),
    .A2(_07448_),
    .ZN(_07604_)
  );
  INV_X1 _17598_ (
    .A(_07604_),
    .ZN(_07605_)
  );
  AND2_X1 _17599_ (
    .A1(_07159_),
    .A2(_07604_),
    .ZN(_07606_)
  );
  INV_X1 _17600_ (
    .A(_07606_),
    .ZN(_07607_)
  );
  AND2_X1 _17601_ (
    .A1(_07456_),
    .A2(_07607_),
    .ZN(_07608_)
  );
  INV_X1 _17602_ (
    .A(_07608_),
    .ZN(_07609_)
  );
  AND2_X1 _17603_ (
    .A1(_07349_),
    .A2(_07355_),
    .ZN(_07610_)
  );
  INV_X1 _17604_ (
    .A(_07610_),
    .ZN(_07612_)
  );
  AND2_X1 _17605_ (
    .A1(_07335_),
    .A2(_07342_),
    .ZN(_07613_)
  );
  INV_X1 _17606_ (
    .A(_07613_),
    .ZN(_07614_)
  );
  AND2_X1 _17607_ (
    .A1(_07322_),
    .A2(_07329_),
    .ZN(_07615_)
  );
  INV_X1 _17608_ (
    .A(_07615_),
    .ZN(_07616_)
  );
  AND2_X1 _17609_ (
    .A1(_07404_),
    .A2(_07430_),
    .ZN(_07617_)
  );
  INV_X1 _17610_ (
    .A(_07617_),
    .ZN(_07618_)
  );
  AND2_X1 _17611_ (
    .A1(_07028_),
    .A2(_07318_),
    .ZN(_07619_)
  );
  INV_X1 _17612_ (
    .A(_07619_),
    .ZN(_07620_)
  );
  AND2_X1 _17613_ (
    .A1(_07417_),
    .A2(_07423_),
    .ZN(_07621_)
  );
  INV_X1 _17614_ (
    .A(_07621_),
    .ZN(_07623_)
  );
  AND2_X1 _17615_ (
    .A1(_07319_),
    .A2(_07623_),
    .ZN(_07624_)
  );
  INV_X1 _17616_ (
    .A(_07624_),
    .ZN(_07625_)
  );
  AND2_X1 _17617_ (
    .A1(_07320_),
    .A2(_07621_),
    .ZN(_07626_)
  );
  INV_X1 _17618_ (
    .A(_07626_),
    .ZN(_07627_)
  );
  AND2_X1 _17619_ (
    .A1(_07625_),
    .A2(_07627_),
    .ZN(_07628_)
  );
  INV_X1 _17620_ (
    .A(_07628_),
    .ZN(_07629_)
  );
  AND2_X1 _17621_ (
    .A1(_07620_),
    .A2(_07628_),
    .ZN(_07630_)
  );
  INV_X1 _17622_ (
    .A(_07630_),
    .ZN(_07631_)
  );
  AND2_X1 _17623_ (
    .A1(_07619_),
    .A2(_07629_),
    .ZN(_07632_)
  );
  INV_X1 _17624_ (
    .A(_07632_),
    .ZN(_07634_)
  );
  AND2_X1 _17625_ (
    .A1(_07631_),
    .A2(_07634_),
    .ZN(_07635_)
  );
  INV_X1 _17626_ (
    .A(_07635_),
    .ZN(_07636_)
  );
  AND2_X1 _17627_ (
    .A1(_07618_),
    .A2(_07635_),
    .ZN(_07637_)
  );
  INV_X1 _17628_ (
    .A(_07637_),
    .ZN(_07638_)
  );
  AND2_X1 _17629_ (
    .A1(_07617_),
    .A2(_07636_),
    .ZN(_07639_)
  );
  INV_X1 _17630_ (
    .A(_07639_),
    .ZN(_07640_)
  );
  AND2_X1 _17631_ (
    .A1(_07638_),
    .A2(_07640_),
    .ZN(_07641_)
  );
  INV_X1 _17632_ (
    .A(_07641_),
    .ZN(_07642_)
  );
  AND2_X1 _17633_ (
    .A1(_07616_),
    .A2(_07641_),
    .ZN(_07643_)
  );
  INV_X1 _17634_ (
    .A(_07643_),
    .ZN(_07645_)
  );
  AND2_X1 _17635_ (
    .A1(_07615_),
    .A2(_07642_),
    .ZN(_07646_)
  );
  INV_X1 _17636_ (
    .A(_07646_),
    .ZN(_07647_)
  );
  AND2_X1 _17637_ (
    .A1(_07645_),
    .A2(_07647_),
    .ZN(_07648_)
  );
  INV_X1 _17638_ (
    .A(_07648_),
    .ZN(_07649_)
  );
  AND2_X1 _17639_ (
    .A1(_07614_),
    .A2(_07648_),
    .ZN(_07650_)
  );
  INV_X1 _17640_ (
    .A(_07650_),
    .ZN(_07651_)
  );
  AND2_X1 _17641_ (
    .A1(_07613_),
    .A2(_07649_),
    .ZN(_07652_)
  );
  INV_X1 _17642_ (
    .A(_07652_),
    .ZN(_07653_)
  );
  AND2_X1 _17643_ (
    .A1(_07651_),
    .A2(_07653_),
    .ZN(_07654_)
  );
  INV_X1 _17644_ (
    .A(_07654_),
    .ZN(_07656_)
  );
  AND2_X1 _17645_ (
    .A1(_07082_),
    .A2(_07654_),
    .ZN(_07657_)
  );
  INV_X1 _17646_ (
    .A(_07657_),
    .ZN(_07658_)
  );
  AND2_X1 _17647_ (
    .A1(_07083_),
    .A2(_07656_),
    .ZN(_07659_)
  );
  INV_X1 _17648_ (
    .A(_07659_),
    .ZN(_07660_)
  );
  AND2_X1 _17649_ (
    .A1(_07658_),
    .A2(_07660_),
    .ZN(_07661_)
  );
  INV_X1 _17650_ (
    .A(_07661_),
    .ZN(_07662_)
  );
  AND2_X1 _17651_ (
    .A1(_07442_),
    .A2(_07661_),
    .ZN(_07663_)
  );
  INV_X1 _17652_ (
    .A(_07663_),
    .ZN(_07664_)
  );
  AND2_X1 _17653_ (
    .A1(_07443_),
    .A2(_07662_),
    .ZN(_07665_)
  );
  INV_X1 _17654_ (
    .A(_07665_),
    .ZN(_07667_)
  );
  AND2_X1 _17655_ (
    .A1(_07664_),
    .A2(_07667_),
    .ZN(_07668_)
  );
  INV_X1 _17656_ (
    .A(_07668_),
    .ZN(_07669_)
  );
  AND2_X1 _17657_ (
    .A1(_07612_),
    .A2(_07668_),
    .ZN(_07670_)
  );
  INV_X1 _17658_ (
    .A(_07670_),
    .ZN(_07671_)
  );
  AND2_X1 _17659_ (
    .A1(_07610_),
    .A2(_07669_),
    .ZN(_07672_)
  );
  INV_X1 _17660_ (
    .A(_07672_),
    .ZN(_07673_)
  );
  AND2_X1 _17661_ (
    .A1(_07671_),
    .A2(_07673_),
    .ZN(_07674_)
  );
  INV_X1 _17662_ (
    .A(_07674_),
    .ZN(_07675_)
  );
  AND2_X1 _17663_ (
    .A1(divisor[25]),
    .A2(remainder[2]),
    .ZN(_07676_)
  );
  INV_X1 _17664_ (
    .A(_07676_),
    .ZN(_07678_)
  );
  AND2_X1 _17665_ (
    .A1(divisor[27]),
    .A2(remainder[0]),
    .ZN(_07679_)
  );
  INV_X1 _17666_ (
    .A(_07679_),
    .ZN(_07680_)
  );
  AND2_X1 _17667_ (
    .A1(divisor[27]),
    .A2(remainder[1]),
    .ZN(_07681_)
  );
  INV_X1 _17668_ (
    .A(_07681_),
    .ZN(_07682_)
  );
  AND2_X1 _17669_ (
    .A1(_07367_),
    .A2(_07681_),
    .ZN(_07683_)
  );
  INV_X1 _17670_ (
    .A(_07683_),
    .ZN(_07684_)
  );
  AND2_X1 _17671_ (
    .A1(_07373_),
    .A2(_07680_),
    .ZN(_07685_)
  );
  INV_X1 _17672_ (
    .A(_07685_),
    .ZN(_07686_)
  );
  AND2_X1 _17673_ (
    .A1(_07684_),
    .A2(_07686_),
    .ZN(_07687_)
  );
  INV_X1 _17674_ (
    .A(_07687_),
    .ZN(_07689_)
  );
  AND2_X1 _17675_ (
    .A1(_07676_),
    .A2(_07687_),
    .ZN(_07690_)
  );
  INV_X1 _17676_ (
    .A(_07690_),
    .ZN(_07691_)
  );
  AND2_X1 _17677_ (
    .A1(_07678_),
    .A2(_07689_),
    .ZN(_07692_)
  );
  INV_X1 _17678_ (
    .A(_07692_),
    .ZN(_07693_)
  );
  AND2_X1 _17679_ (
    .A1(_07691_),
    .A2(_07693_),
    .ZN(_07694_)
  );
  INV_X1 _17680_ (
    .A(_07694_),
    .ZN(_07695_)
  );
  AND2_X1 _17681_ (
    .A1(_07374_),
    .A2(_07694_),
    .ZN(_07696_)
  );
  INV_X1 _17682_ (
    .A(_07696_),
    .ZN(_07697_)
  );
  AND2_X1 _17683_ (
    .A1(_07375_),
    .A2(_07695_),
    .ZN(_07698_)
  );
  INV_X1 _17684_ (
    .A(_07698_),
    .ZN(_07700_)
  );
  AND2_X1 _17685_ (
    .A1(_07697_),
    .A2(_07700_),
    .ZN(_07701_)
  );
  INV_X1 _17686_ (
    .A(_07701_),
    .ZN(_07702_)
  );
  AND2_X1 _17687_ (
    .A1(_07390_),
    .A2(_07397_),
    .ZN(_07703_)
  );
  INV_X1 _17688_ (
    .A(_07703_),
    .ZN(_07704_)
  );
  AND2_X1 _17689_ (
    .A1(divisor[22]),
    .A2(remainder[5]),
    .ZN(_07705_)
  );
  INV_X1 _17690_ (
    .A(_07705_),
    .ZN(_07706_)
  );
  AND2_X1 _17691_ (
    .A1(divisor[23]),
    .A2(remainder[4]),
    .ZN(_07707_)
  );
  INV_X1 _17692_ (
    .A(_07707_),
    .ZN(_07708_)
  );
  AND2_X1 _17693_ (
    .A1(divisor[24]),
    .A2(remainder[4]),
    .ZN(_07709_)
  );
  INV_X1 _17694_ (
    .A(_07709_),
    .ZN(_07711_)
  );
  AND2_X1 _17695_ (
    .A1(_07387_),
    .A2(_07707_),
    .ZN(_07712_)
  );
  INV_X1 _17696_ (
    .A(_07712_),
    .ZN(_07713_)
  );
  AND2_X1 _17697_ (
    .A1(_07388_),
    .A2(_07708_),
    .ZN(_07714_)
  );
  INV_X1 _17698_ (
    .A(_07714_),
    .ZN(_07715_)
  );
  AND2_X1 _17699_ (
    .A1(_07713_),
    .A2(_07715_),
    .ZN(_07716_)
  );
  INV_X1 _17700_ (
    .A(_07716_),
    .ZN(_07717_)
  );
  AND2_X1 _17701_ (
    .A1(_07705_),
    .A2(_07716_),
    .ZN(_07718_)
  );
  INV_X1 _17702_ (
    .A(_07718_),
    .ZN(_07719_)
  );
  AND2_X1 _17703_ (
    .A1(_07706_),
    .A2(_07717_),
    .ZN(_07720_)
  );
  INV_X1 _17704_ (
    .A(_07720_),
    .ZN(_07722_)
  );
  AND2_X1 _17705_ (
    .A1(_07719_),
    .A2(_07722_),
    .ZN(_07723_)
  );
  INV_X1 _17706_ (
    .A(_07723_),
    .ZN(_07724_)
  );
  AND2_X1 _17707_ (
    .A1(_07704_),
    .A2(_07723_),
    .ZN(_07725_)
  );
  INV_X1 _17708_ (
    .A(_07725_),
    .ZN(_07726_)
  );
  AND2_X1 _17709_ (
    .A1(_07703_),
    .A2(_07724_),
    .ZN(_07727_)
  );
  INV_X1 _17710_ (
    .A(_07727_),
    .ZN(_07728_)
  );
  AND2_X1 _17711_ (
    .A1(_07726_),
    .A2(_07728_),
    .ZN(_07729_)
  );
  INV_X1 _17712_ (
    .A(_07729_),
    .ZN(_07730_)
  );
  AND2_X1 _17713_ (
    .A1(divisor[20]),
    .A2(remainder[7]),
    .ZN(_07731_)
  );
  INV_X1 _17714_ (
    .A(_07731_),
    .ZN(_07733_)
  );
  AND2_X1 _17715_ (
    .A1(divisor[21]),
    .A2(remainder[7]),
    .ZN(_07734_)
  );
  INV_X1 _17716_ (
    .A(_07734_),
    .ZN(_07735_)
  );
  AND2_X1 _17717_ (
    .A1(_07411_),
    .A2(_07734_),
    .ZN(_07736_)
  );
  INV_X1 _17718_ (
    .A(_07736_),
    .ZN(_07737_)
  );
  AND2_X1 _17719_ (
    .A1(_07415_),
    .A2(_07733_),
    .ZN(_07738_)
  );
  INV_X1 _17720_ (
    .A(_07738_),
    .ZN(_07739_)
  );
  AND2_X1 _17721_ (
    .A1(_07737_),
    .A2(_07739_),
    .ZN(_07740_)
  );
  INV_X1 _17722_ (
    .A(_07740_),
    .ZN(_07741_)
  );
  AND2_X1 _17723_ (
    .A1(_05269_),
    .A2(_07740_),
    .ZN(_07742_)
  );
  INV_X1 _17724_ (
    .A(_07742_),
    .ZN(_07744_)
  );
  AND2_X1 _17725_ (
    .A1(_05271_),
    .A2(_07741_),
    .ZN(_07745_)
  );
  INV_X1 _17726_ (
    .A(_07745_),
    .ZN(_07746_)
  );
  AND2_X1 _17727_ (
    .A1(_07744_),
    .A2(_07746_),
    .ZN(_07747_)
  );
  INV_X1 _17728_ (
    .A(_07747_),
    .ZN(_07748_)
  );
  AND2_X1 _17729_ (
    .A1(_07729_),
    .A2(_07747_),
    .ZN(_07749_)
  );
  INV_X1 _17730_ (
    .A(_07749_),
    .ZN(_07750_)
  );
  AND2_X1 _17731_ (
    .A1(_07730_),
    .A2(_07748_),
    .ZN(_07751_)
  );
  INV_X1 _17732_ (
    .A(_07751_),
    .ZN(_07752_)
  );
  AND2_X1 _17733_ (
    .A1(_07750_),
    .A2(_07752_),
    .ZN(_07753_)
  );
  INV_X1 _17734_ (
    .A(_07753_),
    .ZN(_07755_)
  );
  AND2_X1 _17735_ (
    .A1(_07701_),
    .A2(_07753_),
    .ZN(_07756_)
  );
  INV_X1 _17736_ (
    .A(_07756_),
    .ZN(_07757_)
  );
  AND2_X1 _17737_ (
    .A1(_07702_),
    .A2(_07755_),
    .ZN(_07758_)
  );
  INV_X1 _17738_ (
    .A(_07758_),
    .ZN(_07759_)
  );
  AND2_X1 _17739_ (
    .A1(_07757_),
    .A2(_07759_),
    .ZN(_07760_)
  );
  INV_X1 _17740_ (
    .A(_07760_),
    .ZN(_07761_)
  );
  AND2_X1 _17741_ (
    .A1(_07435_),
    .A2(_07760_),
    .ZN(_07762_)
  );
  INV_X1 _17742_ (
    .A(_07762_),
    .ZN(_07763_)
  );
  AND2_X1 _17743_ (
    .A1(_07437_),
    .A2(_07761_),
    .ZN(_07764_)
  );
  INV_X1 _17744_ (
    .A(_07764_),
    .ZN(_07766_)
  );
  AND2_X1 _17745_ (
    .A1(_07763_),
    .A2(_07766_),
    .ZN(_07767_)
  );
  INV_X1 _17746_ (
    .A(_07767_),
    .ZN(_07768_)
  );
  AND2_X1 _17747_ (
    .A1(_07605_),
    .A2(_07768_),
    .ZN(_07769_)
  );
  INV_X1 _17748_ (
    .A(_07769_),
    .ZN(_07770_)
  );
  AND2_X1 _17749_ (
    .A1(_07604_),
    .A2(_07767_),
    .ZN(_07771_)
  );
  INV_X1 _17750_ (
    .A(_07771_),
    .ZN(_07772_)
  );
  AND2_X1 _17751_ (
    .A1(_07605_),
    .A2(_07767_),
    .ZN(_07773_)
  );
  INV_X1 _17752_ (
    .A(_07773_),
    .ZN(_07774_)
  );
  AND2_X1 _17753_ (
    .A1(_07604_),
    .A2(_07768_),
    .ZN(_07775_)
  );
  INV_X1 _17754_ (
    .A(_07775_),
    .ZN(_07777_)
  );
  AND2_X1 _17755_ (
    .A1(_07770_),
    .A2(_07772_),
    .ZN(_07778_)
  );
  AND2_X1 _17756_ (
    .A1(_07774_),
    .A2(_07777_),
    .ZN(_07779_)
  );
  AND2_X1 _17757_ (
    .A1(_07674_),
    .A2(_07778_),
    .ZN(_07780_)
  );
  INV_X1 _17758_ (
    .A(_07780_),
    .ZN(_07781_)
  );
  AND2_X1 _17759_ (
    .A1(_07675_),
    .A2(_07779_),
    .ZN(_07782_)
  );
  INV_X1 _17760_ (
    .A(_07782_),
    .ZN(_07783_)
  );
  AND2_X1 _17761_ (
    .A1(_07781_),
    .A2(_07783_),
    .ZN(_07784_)
  );
  INV_X1 _17762_ (
    .A(_07784_),
    .ZN(_07785_)
  );
  AND2_X1 _17763_ (
    .A1(_07609_),
    .A2(_07784_),
    .ZN(_07786_)
  );
  INV_X1 _17764_ (
    .A(_07786_),
    .ZN(_07788_)
  );
  AND2_X1 _17765_ (
    .A1(_07608_),
    .A2(_07785_),
    .ZN(_07789_)
  );
  INV_X1 _17766_ (
    .A(_07789_),
    .ZN(_07790_)
  );
  AND2_X1 _17767_ (
    .A1(_07788_),
    .A2(_07790_),
    .ZN(_07791_)
  );
  INV_X1 _17768_ (
    .A(_07791_),
    .ZN(_07792_)
  );
  AND2_X1 _17769_ (
    .A1(_07494_),
    .A2(_07500_),
    .ZN(_07793_)
  );
  INV_X1 _17770_ (
    .A(_07793_),
    .ZN(_07794_)
  );
  AND2_X1 _17771_ (
    .A1(_06580_),
    .A2(_07477_),
    .ZN(_07795_)
  );
  INV_X1 _17772_ (
    .A(_07795_),
    .ZN(_07796_)
  );
  AND2_X1 _17773_ (
    .A1(_07494_),
    .A2(_07796_),
    .ZN(_07797_)
  );
  INV_X1 _17774_ (
    .A(_07797_),
    .ZN(_07799_)
  );
  AND2_X1 _17775_ (
    .A1(_03170_),
    .A2(_07797_),
    .ZN(_07800_)
  );
  INV_X1 _17776_ (
    .A(_07800_),
    .ZN(_07801_)
  );
  AND2_X1 _17777_ (
    .A1(_03169_),
    .A2(_07799_),
    .ZN(_07802_)
  );
  INV_X1 _17778_ (
    .A(_07802_),
    .ZN(_07803_)
  );
  AND2_X1 _17779_ (
    .A1(_07801_),
    .A2(_07803_),
    .ZN(_07804_)
  );
  INV_X1 _17780_ (
    .A(_07804_),
    .ZN(_07805_)
  );
  AND2_X1 _17781_ (
    .A1(_07361_),
    .A2(_07804_),
    .ZN(_07806_)
  );
  INV_X1 _17782_ (
    .A(_07806_),
    .ZN(_07807_)
  );
  AND2_X1 _17783_ (
    .A1(_07362_),
    .A2(_07805_),
    .ZN(_07808_)
  );
  INV_X1 _17784_ (
    .A(_07808_),
    .ZN(_07810_)
  );
  AND2_X1 _17785_ (
    .A1(_07807_),
    .A2(_07810_),
    .ZN(_07811_)
  );
  INV_X1 _17786_ (
    .A(_07811_),
    .ZN(_07812_)
  );
  AND2_X1 _17787_ (
    .A1(_07794_),
    .A2(_07811_),
    .ZN(_07813_)
  );
  INV_X1 _17788_ (
    .A(_07813_),
    .ZN(_07814_)
  );
  AND2_X1 _17789_ (
    .A1(_07793_),
    .A2(_07812_),
    .ZN(_07815_)
  );
  INV_X1 _17790_ (
    .A(_07815_),
    .ZN(_07816_)
  );
  AND2_X1 _17791_ (
    .A1(_07814_),
    .A2(_07816_),
    .ZN(_07817_)
  );
  INV_X1 _17792_ (
    .A(_07817_),
    .ZN(_07818_)
  );
  AND2_X1 _17793_ (
    .A1(_07791_),
    .A2(_07817_),
    .ZN(_07819_)
  );
  INV_X1 _17794_ (
    .A(_07819_),
    .ZN(_07821_)
  );
  AND2_X1 _17795_ (
    .A1(_07792_),
    .A2(_07818_),
    .ZN(_07822_)
  );
  INV_X1 _17796_ (
    .A(_07822_),
    .ZN(_07823_)
  );
  AND2_X1 _17797_ (
    .A1(_07821_),
    .A2(_07823_),
    .ZN(_07824_)
  );
  INV_X1 _17798_ (
    .A(_07824_),
    .ZN(_07825_)
  );
  AND2_X1 _17799_ (
    .A1(_07603_),
    .A2(_07824_),
    .ZN(_07826_)
  );
  INV_X1 _17800_ (
    .A(_07826_),
    .ZN(_07827_)
  );
  AND2_X1 _17801_ (
    .A1(_07602_),
    .A2(_07825_),
    .ZN(_07828_)
  );
  INV_X1 _17802_ (
    .A(_07828_),
    .ZN(_07829_)
  );
  AND2_X1 _17803_ (
    .A1(_07827_),
    .A2(_07829_),
    .ZN(_07830_)
  );
  INV_X1 _17804_ (
    .A(_07830_),
    .ZN(_07832_)
  );
  AND2_X1 _17805_ (
    .A1(_07601_),
    .A2(_07830_),
    .ZN(_07833_)
  );
  INV_X1 _17806_ (
    .A(_07833_),
    .ZN(_07834_)
  );
  AND2_X1 _17807_ (
    .A1(_07599_),
    .A2(_07832_),
    .ZN(_07835_)
  );
  INV_X1 _17808_ (
    .A(_07835_),
    .ZN(_07836_)
  );
  AND2_X1 _17809_ (
    .A1(_07834_),
    .A2(_07836_),
    .ZN(_07837_)
  );
  INV_X1 _17810_ (
    .A(_07837_),
    .ZN(_07838_)
  );
  AND2_X1 _17811_ (
    .A1(_07598_),
    .A2(_07837_),
    .ZN(_07839_)
  );
  INV_X1 _17812_ (
    .A(_07839_),
    .ZN(_07840_)
  );
  AND2_X1 _17813_ (
    .A1(_07597_),
    .A2(_07838_),
    .ZN(_07841_)
  );
  INV_X1 _17814_ (
    .A(_07841_),
    .ZN(_07843_)
  );
  AND2_X1 _17815_ (
    .A1(_07840_),
    .A2(_07843_),
    .ZN(_07844_)
  );
  INV_X1 _17816_ (
    .A(_07844_),
    .ZN(_07845_)
  );
  AND2_X1 _17817_ (
    .A1(_07539_),
    .A2(_07844_),
    .ZN(_07846_)
  );
  INV_X1 _17818_ (
    .A(_07846_),
    .ZN(_07847_)
  );
  AND2_X1 _17819_ (
    .A1(_07540_),
    .A2(_07845_),
    .ZN(_07848_)
  );
  INV_X1 _17820_ (
    .A(_07848_),
    .ZN(_07849_)
  );
  AND2_X1 _17821_ (
    .A1(_07847_),
    .A2(_07849_),
    .ZN(_07850_)
  );
  INV_X1 _17822_ (
    .A(_07850_),
    .ZN(_07851_)
  );
  AND2_X1 _17823_ (
    .A1(_07595_),
    .A2(_07851_),
    .ZN(_07852_)
  );
  INV_X1 _17824_ (
    .A(_07852_),
    .ZN(_07854_)
  );
  AND2_X1 _17825_ (
    .A1(_07596_),
    .A2(_07850_),
    .ZN(_07855_)
  );
  INV_X1 _17826_ (
    .A(_07855_),
    .ZN(_07856_)
  );
  AND2_X1 _17827_ (
    .A1(_07854_),
    .A2(_07856_),
    .ZN(_07857_)
  );
  INV_X1 _17828_ (
    .A(_07857_),
    .ZN(_07858_)
  );
  AND2_X1 _17829_ (
    .A1(remainder[60]),
    .A2(_07857_),
    .ZN(_07859_)
  );
  INV_X1 _17830_ (
    .A(_07859_),
    .ZN(_07860_)
  );
  AND2_X1 _17831_ (
    .A1(_04459_),
    .A2(_07858_),
    .ZN(_07861_)
  );
  INV_X1 _17832_ (
    .A(_07861_),
    .ZN(_07862_)
  );
  AND2_X1 _17833_ (
    .A1(_07860_),
    .A2(_07862_),
    .ZN(_07863_)
  );
  INV_X1 _17834_ (
    .A(_07863_),
    .ZN(_07865_)
  );
  AND2_X1 _17835_ (
    .A1(_07593_),
    .A2(_07865_),
    .ZN(_07866_)
  );
  INV_X1 _17836_ (
    .A(_07866_),
    .ZN(_07867_)
  );
  AND2_X1 _17837_ (
    .A1(_07594_),
    .A2(_07863_),
    .ZN(_07868_)
  );
  INV_X1 _17838_ (
    .A(_07868_),
    .ZN(_07869_)
  );
  AND2_X1 _17839_ (
    .A1(_07867_),
    .A2(_07869_),
    .ZN(_07870_)
  );
  AND2_X1 _17840_ (
    .A1(_02082_),
    .A2(_07870_),
    .ZN(_07871_)
  );
  INV_X1 _17841_ (
    .A(_07871_),
    .ZN(_07872_)
  );
  AND2_X1 _17842_ (
    .A1(remainder[52]),
    .A2(_02077_),
    .ZN(_07873_)
  );
  INV_X1 _17843_ (
    .A(_07873_),
    .ZN(_07874_)
  );
  AND2_X1 _17844_ (
    .A1(_04557_),
    .A2(_10451_),
    .ZN(_07876_)
  );
  INV_X1 _17845_ (
    .A(_07876_),
    .ZN(_07877_)
  );
  AND2_X1 _17846_ (
    .A1(_10462_),
    .A2(_01892_),
    .ZN(_07878_)
  );
  INV_X1 _17847_ (
    .A(_07878_),
    .ZN(_07879_)
  );
  AND2_X1 _17848_ (
    .A1(_05983_),
    .A2(_07879_),
    .ZN(_07880_)
  );
  AND2_X1 _17849_ (
    .A1(_07877_),
    .A2(_07880_),
    .ZN(_07881_)
  );
  INV_X1 _17850_ (
    .A(_07881_),
    .ZN(_07882_)
  );
  AND2_X1 _17851_ (
    .A1(_07874_),
    .A2(_07882_),
    .ZN(_07883_)
  );
  AND2_X1 _17852_ (
    .A1(_07872_),
    .A2(_07883_),
    .ZN(_07884_)
  );
  INV_X1 _17853_ (
    .A(_07884_),
    .ZN(_07885_)
  );
  AND2_X1 _17854_ (
    .A1(_06201_),
    .A2(_07885_),
    .ZN(_00073_)
  );
  AND2_X1 _17855_ (
    .A1(_07827_),
    .A2(_07834_),
    .ZN(_07887_)
  );
  INV_X1 _17856_ (
    .A(_07887_),
    .ZN(_07888_)
  );
  AND2_X1 _17857_ (
    .A1(_07807_),
    .A2(_07814_),
    .ZN(_07889_)
  );
  INV_X1 _17858_ (
    .A(_07889_),
    .ZN(_07890_)
  );
  AND2_X1 _17859_ (
    .A1(_07788_),
    .A2(_07821_),
    .ZN(_07891_)
  );
  INV_X1 _17860_ (
    .A(_07891_),
    .ZN(_07892_)
  );
  AND2_X1 _17861_ (
    .A1(_03249_),
    .A2(_07446_),
    .ZN(_07893_)
  );
  AND2_X1 _17862_ (
    .A1(_07768_),
    .A2(_07893_),
    .ZN(_07894_)
  );
  INV_X1 _17863_ (
    .A(_07894_),
    .ZN(_07895_)
  );
  AND2_X1 _17864_ (
    .A1(_07781_),
    .A2(_07895_),
    .ZN(_07897_)
  );
  INV_X1 _17865_ (
    .A(_07897_),
    .ZN(_07898_)
  );
  AND2_X1 _17866_ (
    .A1(_03249_),
    .A2(_07767_),
    .ZN(_07899_)
  );
  INV_X1 _17867_ (
    .A(_07899_),
    .ZN(_07900_)
  );
  AND2_X1 _17868_ (
    .A1(_07684_),
    .A2(_07691_),
    .ZN(_07901_)
  );
  INV_X1 _17869_ (
    .A(_07901_),
    .ZN(_07902_)
  );
  AND2_X1 _17870_ (
    .A1(divisor[25]),
    .A2(remainder[3]),
    .ZN(_07903_)
  );
  INV_X1 _17871_ (
    .A(_07903_),
    .ZN(_07904_)
  );
  AND2_X1 _17872_ (
    .A1(divisor[26]),
    .A2(remainder[2]),
    .ZN(_07905_)
  );
  INV_X1 _17873_ (
    .A(_07905_),
    .ZN(_07906_)
  );
  AND2_X1 _17874_ (
    .A1(divisor[27]),
    .A2(remainder[2]),
    .ZN(_07908_)
  );
  INV_X1 _17875_ (
    .A(_07908_),
    .ZN(_07909_)
  );
  AND2_X1 _17876_ (
    .A1(_07372_),
    .A2(_07908_),
    .ZN(_07910_)
  );
  INV_X1 _17877_ (
    .A(_07910_),
    .ZN(_07911_)
  );
  AND2_X1 _17878_ (
    .A1(_07682_),
    .A2(_07906_),
    .ZN(_07912_)
  );
  INV_X1 _17879_ (
    .A(_07912_),
    .ZN(_07913_)
  );
  AND2_X1 _17880_ (
    .A1(_07911_),
    .A2(_07913_),
    .ZN(_07914_)
  );
  INV_X1 _17881_ (
    .A(_07914_),
    .ZN(_07915_)
  );
  AND2_X1 _17882_ (
    .A1(_07903_),
    .A2(_07914_),
    .ZN(_07916_)
  );
  INV_X1 _17883_ (
    .A(_07916_),
    .ZN(_07917_)
  );
  AND2_X1 _17884_ (
    .A1(_07904_),
    .A2(_07915_),
    .ZN(_07919_)
  );
  INV_X1 _17885_ (
    .A(_07919_),
    .ZN(_07920_)
  );
  AND2_X1 _17886_ (
    .A1(_07917_),
    .A2(_07920_),
    .ZN(_07921_)
  );
  INV_X1 _17887_ (
    .A(_07921_),
    .ZN(_07922_)
  );
  AND2_X1 _17888_ (
    .A1(_07902_),
    .A2(_07921_),
    .ZN(_07923_)
  );
  INV_X1 _17889_ (
    .A(_07923_),
    .ZN(_07924_)
  );
  AND2_X1 _17890_ (
    .A1(_07901_),
    .A2(_07922_),
    .ZN(_07925_)
  );
  INV_X1 _17891_ (
    .A(_07925_),
    .ZN(_07926_)
  );
  AND2_X1 _17892_ (
    .A1(_07924_),
    .A2(_07926_),
    .ZN(_07927_)
  );
  INV_X1 _17893_ (
    .A(_07927_),
    .ZN(_07928_)
  );
  AND2_X1 _17894_ (
    .A1(_07696_),
    .A2(_07927_),
    .ZN(_07930_)
  );
  INV_X1 _17895_ (
    .A(_07930_),
    .ZN(_07931_)
  );
  AND2_X1 _17896_ (
    .A1(_07697_),
    .A2(_07928_),
    .ZN(_07932_)
  );
  INV_X1 _17897_ (
    .A(_07932_),
    .ZN(_07933_)
  );
  AND2_X1 _17898_ (
    .A1(_07931_),
    .A2(_07933_),
    .ZN(_07934_)
  );
  INV_X1 _17899_ (
    .A(_07934_),
    .ZN(_07935_)
  );
  AND2_X1 _17900_ (
    .A1(_07713_),
    .A2(_07719_),
    .ZN(_07936_)
  );
  INV_X1 _17901_ (
    .A(_07936_),
    .ZN(_07937_)
  );
  AND2_X1 _17902_ (
    .A1(divisor[22]),
    .A2(remainder[6]),
    .ZN(_07938_)
  );
  INV_X1 _17903_ (
    .A(_07938_),
    .ZN(_07939_)
  );
  AND2_X1 _17904_ (
    .A1(divisor[23]),
    .A2(remainder[5]),
    .ZN(_07941_)
  );
  INV_X1 _17905_ (
    .A(_07941_),
    .ZN(_07942_)
  );
  AND2_X1 _17906_ (
    .A1(divisor[24]),
    .A2(remainder[5]),
    .ZN(_07943_)
  );
  INV_X1 _17907_ (
    .A(_07943_),
    .ZN(_07944_)
  );
  AND2_X1 _17908_ (
    .A1(_07709_),
    .A2(_07941_),
    .ZN(_07945_)
  );
  INV_X1 _17909_ (
    .A(_07945_),
    .ZN(_07946_)
  );
  AND2_X1 _17910_ (
    .A1(_07711_),
    .A2(_07942_),
    .ZN(_07947_)
  );
  INV_X1 _17911_ (
    .A(_07947_),
    .ZN(_07948_)
  );
  AND2_X1 _17912_ (
    .A1(_07946_),
    .A2(_07948_),
    .ZN(_07949_)
  );
  INV_X1 _17913_ (
    .A(_07949_),
    .ZN(_07950_)
  );
  AND2_X1 _17914_ (
    .A1(_07938_),
    .A2(_07949_),
    .ZN(_07952_)
  );
  INV_X1 _17915_ (
    .A(_07952_),
    .ZN(_07953_)
  );
  AND2_X1 _17916_ (
    .A1(_07939_),
    .A2(_07950_),
    .ZN(_07954_)
  );
  INV_X1 _17917_ (
    .A(_07954_),
    .ZN(_07955_)
  );
  AND2_X1 _17918_ (
    .A1(_07953_),
    .A2(_07955_),
    .ZN(_07956_)
  );
  INV_X1 _17919_ (
    .A(_07956_),
    .ZN(_07957_)
  );
  AND2_X1 _17920_ (
    .A1(_07937_),
    .A2(_07956_),
    .ZN(_07958_)
  );
  INV_X1 _17921_ (
    .A(_07958_),
    .ZN(_07959_)
  );
  AND2_X1 _17922_ (
    .A1(_07936_),
    .A2(_07957_),
    .ZN(_07960_)
  );
  INV_X1 _17923_ (
    .A(_07960_),
    .ZN(_07961_)
  );
  AND2_X1 _17924_ (
    .A1(_07959_),
    .A2(_07961_),
    .ZN(_07963_)
  );
  INV_X1 _17925_ (
    .A(_07963_),
    .ZN(_07964_)
  );
  AND2_X1 _17926_ (
    .A1(remainder[32]),
    .A2(divisor[21]),
    .ZN(_07965_)
  );
  AND2_X1 _17927_ (
    .A1(remainder[32]),
    .A2(divisor[20]),
    .ZN(_07966_)
  );
  INV_X1 _17928_ (
    .A(_07966_),
    .ZN(_07967_)
  );
  AND2_X1 _17929_ (
    .A1(divisor[21]),
    .A2(_07966_),
    .ZN(_07968_)
  );
  INV_X1 _17930_ (
    .A(_07968_),
    .ZN(_07969_)
  );
  AND2_X1 _17931_ (
    .A1(_07734_),
    .A2(_07966_),
    .ZN(_07970_)
  );
  INV_X1 _17932_ (
    .A(_07970_),
    .ZN(_07971_)
  );
  AND2_X1 _17933_ (
    .A1(_07735_),
    .A2(_07967_),
    .ZN(_07972_)
  );
  INV_X1 _17934_ (
    .A(_07972_),
    .ZN(_07974_)
  );
  AND2_X1 _17935_ (
    .A1(_07971_),
    .A2(_07974_),
    .ZN(_07975_)
  );
  INV_X1 _17936_ (
    .A(_07975_),
    .ZN(_07976_)
  );
  AND2_X1 _17937_ (
    .A1(_05269_),
    .A2(_07975_),
    .ZN(_07977_)
  );
  INV_X1 _17938_ (
    .A(_07977_),
    .ZN(_07978_)
  );
  AND2_X1 _17939_ (
    .A1(_05271_),
    .A2(_07976_),
    .ZN(_07979_)
  );
  INV_X1 _17940_ (
    .A(_07979_),
    .ZN(_07980_)
  );
  AND2_X1 _17941_ (
    .A1(_07978_),
    .A2(_07980_),
    .ZN(_07981_)
  );
  INV_X1 _17942_ (
    .A(_07981_),
    .ZN(_07982_)
  );
  AND2_X1 _17943_ (
    .A1(_07963_),
    .A2(_07981_),
    .ZN(_07983_)
  );
  INV_X1 _17944_ (
    .A(_07983_),
    .ZN(_07985_)
  );
  AND2_X1 _17945_ (
    .A1(_07964_),
    .A2(_07982_),
    .ZN(_07986_)
  );
  INV_X1 _17946_ (
    .A(_07986_),
    .ZN(_07987_)
  );
  AND2_X1 _17947_ (
    .A1(_07985_),
    .A2(_07987_),
    .ZN(_07988_)
  );
  INV_X1 _17948_ (
    .A(_07988_),
    .ZN(_07989_)
  );
  AND2_X1 _17949_ (
    .A1(_07934_),
    .A2(_07988_),
    .ZN(_07990_)
  );
  INV_X1 _17950_ (
    .A(_07990_),
    .ZN(_07991_)
  );
  AND2_X1 _17951_ (
    .A1(_07935_),
    .A2(_07989_),
    .ZN(_07992_)
  );
  INV_X1 _17952_ (
    .A(_07992_),
    .ZN(_07993_)
  );
  AND2_X1 _17953_ (
    .A1(_07991_),
    .A2(_07993_),
    .ZN(_07994_)
  );
  INV_X1 _17954_ (
    .A(_07994_),
    .ZN(_07996_)
  );
  AND2_X1 _17955_ (
    .A1(_07756_),
    .A2(_07994_),
    .ZN(_07997_)
  );
  INV_X1 _17956_ (
    .A(_07997_),
    .ZN(_07998_)
  );
  AND2_X1 _17957_ (
    .A1(_07757_),
    .A2(_07996_),
    .ZN(_07999_)
  );
  INV_X1 _17958_ (
    .A(_07999_),
    .ZN(_08000_)
  );
  AND2_X1 _17959_ (
    .A1(_07998_),
    .A2(_08000_),
    .ZN(_08001_)
  );
  INV_X1 _17960_ (
    .A(_08001_),
    .ZN(_08002_)
  );
  AND2_X1 _17961_ (
    .A1(divisor[28]),
    .A2(remainder[0]),
    .ZN(_08003_)
  );
  INV_X1 _17962_ (
    .A(_08003_),
    .ZN(_08004_)
  );
  AND2_X1 _17963_ (
    .A1(remainder[32]),
    .A2(divisor[28]),
    .ZN(_08005_)
  );
  INV_X1 _17964_ (
    .A(_08005_),
    .ZN(_08007_)
  );
  AND2_X1 _17965_ (
    .A1(_03249_),
    .A2(_08003_),
    .ZN(_08008_)
  );
  AND2_X1 _17966_ (
    .A1(_03249_),
    .A2(_08004_),
    .ZN(_08009_)
  );
  INV_X1 _17967_ (
    .A(_08009_),
    .ZN(_08010_)
  );
  AND2_X1 _17968_ (
    .A1(_03250_),
    .A2(_08003_),
    .ZN(_08011_)
  );
  INV_X1 _17969_ (
    .A(_08011_),
    .ZN(_08012_)
  );
  AND2_X1 _17970_ (
    .A1(_08010_),
    .A2(_08012_),
    .ZN(_08013_)
  );
  INV_X1 _17971_ (
    .A(_08013_),
    .ZN(_08014_)
  );
  AND2_X1 _17972_ (
    .A1(_08001_),
    .A2(_08014_),
    .ZN(_08015_)
  );
  INV_X1 _17973_ (
    .A(_08015_),
    .ZN(_08016_)
  );
  AND2_X1 _17974_ (
    .A1(_08002_),
    .A2(_08013_),
    .ZN(_08018_)
  );
  INV_X1 _17975_ (
    .A(_08018_),
    .ZN(_08019_)
  );
  AND2_X1 _17976_ (
    .A1(_08016_),
    .A2(_08019_),
    .ZN(_08020_)
  );
  INV_X1 _17977_ (
    .A(_08020_),
    .ZN(_08021_)
  );
  AND2_X1 _17978_ (
    .A1(_07899_),
    .A2(_08020_),
    .ZN(_08022_)
  );
  INV_X1 _17979_ (
    .A(_08022_),
    .ZN(_08023_)
  );
  AND2_X1 _17980_ (
    .A1(_07900_),
    .A2(_08021_),
    .ZN(_08024_)
  );
  INV_X1 _17981_ (
    .A(_08024_),
    .ZN(_08025_)
  );
  AND2_X1 _17982_ (
    .A1(_08023_),
    .A2(_08025_),
    .ZN(_08026_)
  );
  INV_X1 _17983_ (
    .A(_08026_),
    .ZN(_08027_)
  );
  AND2_X1 _17984_ (
    .A1(_07651_),
    .A2(_07658_),
    .ZN(_08029_)
  );
  INV_X1 _17985_ (
    .A(_08029_),
    .ZN(_08030_)
  );
  AND2_X1 _17986_ (
    .A1(_07638_),
    .A2(_07645_),
    .ZN(_08031_)
  );
  INV_X1 _17987_ (
    .A(_08031_),
    .ZN(_08032_)
  );
  AND2_X1 _17988_ (
    .A1(_07625_),
    .A2(_07631_),
    .ZN(_08033_)
  );
  INV_X1 _17989_ (
    .A(_08033_),
    .ZN(_08034_)
  );
  AND2_X1 _17990_ (
    .A1(_07726_),
    .A2(_07750_),
    .ZN(_08035_)
  );
  INV_X1 _17991_ (
    .A(_08035_),
    .ZN(_08036_)
  );
  AND2_X1 _17992_ (
    .A1(_07737_),
    .A2(_07744_),
    .ZN(_08037_)
  );
  INV_X1 _17993_ (
    .A(_08037_),
    .ZN(_08038_)
  );
  AND2_X1 _17994_ (
    .A1(_07319_),
    .A2(_08038_),
    .ZN(_08040_)
  );
  INV_X1 _17995_ (
    .A(_08040_),
    .ZN(_08041_)
  );
  AND2_X1 _17996_ (
    .A1(_07320_),
    .A2(_08037_),
    .ZN(_08042_)
  );
  INV_X1 _17997_ (
    .A(_08042_),
    .ZN(_08043_)
  );
  AND2_X1 _17998_ (
    .A1(_08041_),
    .A2(_08043_),
    .ZN(_08044_)
  );
  INV_X1 _17999_ (
    .A(_08044_),
    .ZN(_08045_)
  );
  AND2_X1 _18000_ (
    .A1(_07620_),
    .A2(_08044_),
    .ZN(_08046_)
  );
  INV_X1 _18001_ (
    .A(_08046_),
    .ZN(_08047_)
  );
  AND2_X1 _18002_ (
    .A1(_07619_),
    .A2(_08045_),
    .ZN(_08048_)
  );
  INV_X1 _18003_ (
    .A(_08048_),
    .ZN(_08049_)
  );
  AND2_X1 _18004_ (
    .A1(_08047_),
    .A2(_08049_),
    .ZN(_08051_)
  );
  INV_X1 _18005_ (
    .A(_08051_),
    .ZN(_08052_)
  );
  AND2_X1 _18006_ (
    .A1(_08036_),
    .A2(_08051_),
    .ZN(_08053_)
  );
  INV_X1 _18007_ (
    .A(_08053_),
    .ZN(_08054_)
  );
  AND2_X1 _18008_ (
    .A1(_08035_),
    .A2(_08052_),
    .ZN(_08055_)
  );
  INV_X1 _18009_ (
    .A(_08055_),
    .ZN(_08056_)
  );
  AND2_X1 _18010_ (
    .A1(_08054_),
    .A2(_08056_),
    .ZN(_08057_)
  );
  INV_X1 _18011_ (
    .A(_08057_),
    .ZN(_08058_)
  );
  AND2_X1 _18012_ (
    .A1(_08034_),
    .A2(_08057_),
    .ZN(_08059_)
  );
  INV_X1 _18013_ (
    .A(_08059_),
    .ZN(_08060_)
  );
  AND2_X1 _18014_ (
    .A1(_08033_),
    .A2(_08058_),
    .ZN(_08062_)
  );
  INV_X1 _18015_ (
    .A(_08062_),
    .ZN(_08063_)
  );
  AND2_X1 _18016_ (
    .A1(_08060_),
    .A2(_08063_),
    .ZN(_08064_)
  );
  INV_X1 _18017_ (
    .A(_08064_),
    .ZN(_08065_)
  );
  AND2_X1 _18018_ (
    .A1(_08032_),
    .A2(_08064_),
    .ZN(_08066_)
  );
  INV_X1 _18019_ (
    .A(_08066_),
    .ZN(_08067_)
  );
  AND2_X1 _18020_ (
    .A1(_08031_),
    .A2(_08065_),
    .ZN(_08068_)
  );
  INV_X1 _18021_ (
    .A(_08068_),
    .ZN(_08069_)
  );
  AND2_X1 _18022_ (
    .A1(_08067_),
    .A2(_08069_),
    .ZN(_08070_)
  );
  INV_X1 _18023_ (
    .A(_08070_),
    .ZN(_08071_)
  );
  AND2_X1 _18024_ (
    .A1(_07082_),
    .A2(_08070_),
    .ZN(_08073_)
  );
  INV_X1 _18025_ (
    .A(_08073_),
    .ZN(_08074_)
  );
  AND2_X1 _18026_ (
    .A1(_07083_),
    .A2(_08071_),
    .ZN(_08075_)
  );
  INV_X1 _18027_ (
    .A(_08075_),
    .ZN(_08076_)
  );
  AND2_X1 _18028_ (
    .A1(_08074_),
    .A2(_08076_),
    .ZN(_08077_)
  );
  INV_X1 _18029_ (
    .A(_08077_),
    .ZN(_08078_)
  );
  AND2_X1 _18030_ (
    .A1(_07762_),
    .A2(_08077_),
    .ZN(_08079_)
  );
  INV_X1 _18031_ (
    .A(_08079_),
    .ZN(_08080_)
  );
  AND2_X1 _18032_ (
    .A1(_07763_),
    .A2(_08078_),
    .ZN(_08081_)
  );
  INV_X1 _18033_ (
    .A(_08081_),
    .ZN(_08082_)
  );
  AND2_X1 _18034_ (
    .A1(_08080_),
    .A2(_08082_),
    .ZN(_08084_)
  );
  INV_X1 _18035_ (
    .A(_08084_),
    .ZN(_08085_)
  );
  AND2_X1 _18036_ (
    .A1(_08030_),
    .A2(_08084_),
    .ZN(_08086_)
  );
  INV_X1 _18037_ (
    .A(_08086_),
    .ZN(_08087_)
  );
  AND2_X1 _18038_ (
    .A1(_08029_),
    .A2(_08085_),
    .ZN(_08088_)
  );
  INV_X1 _18039_ (
    .A(_08088_),
    .ZN(_08089_)
  );
  AND2_X1 _18040_ (
    .A1(_08087_),
    .A2(_08089_),
    .ZN(_08090_)
  );
  INV_X1 _18041_ (
    .A(_08090_),
    .ZN(_08091_)
  );
  AND2_X1 _18042_ (
    .A1(_08026_),
    .A2(_08090_),
    .ZN(_08092_)
  );
  INV_X1 _18043_ (
    .A(_08092_),
    .ZN(_08093_)
  );
  AND2_X1 _18044_ (
    .A1(_08027_),
    .A2(_08091_),
    .ZN(_08095_)
  );
  INV_X1 _18045_ (
    .A(_08095_),
    .ZN(_08096_)
  );
  AND2_X1 _18046_ (
    .A1(_08093_),
    .A2(_08096_),
    .ZN(_08097_)
  );
  INV_X1 _18047_ (
    .A(_08097_),
    .ZN(_08098_)
  );
  AND2_X1 _18048_ (
    .A1(_07898_),
    .A2(_08097_),
    .ZN(_08099_)
  );
  INV_X1 _18049_ (
    .A(_08099_),
    .ZN(_08100_)
  );
  AND2_X1 _18050_ (
    .A1(_07897_),
    .A2(_08098_),
    .ZN(_08101_)
  );
  INV_X1 _18051_ (
    .A(_08101_),
    .ZN(_08102_)
  );
  AND2_X1 _18052_ (
    .A1(_08100_),
    .A2(_08102_),
    .ZN(_08103_)
  );
  INV_X1 _18053_ (
    .A(_08103_),
    .ZN(_08104_)
  );
  AND2_X1 _18054_ (
    .A1(_07494_),
    .A2(_07801_),
    .ZN(_08106_)
  );
  INV_X1 _18055_ (
    .A(_08106_),
    .ZN(_08107_)
  );
  AND2_X1 _18056_ (
    .A1(_07664_),
    .A2(_07671_),
    .ZN(_08108_)
  );
  INV_X1 _18057_ (
    .A(_08108_),
    .ZN(_08109_)
  );
  AND2_X1 _18058_ (
    .A1(_07804_),
    .A2(_08109_),
    .ZN(_08110_)
  );
  INV_X1 _18059_ (
    .A(_08110_),
    .ZN(_08111_)
  );
  AND2_X1 _18060_ (
    .A1(_07805_),
    .A2(_08108_),
    .ZN(_08112_)
  );
  INV_X1 _18061_ (
    .A(_08112_),
    .ZN(_08113_)
  );
  AND2_X1 _18062_ (
    .A1(_08111_),
    .A2(_08113_),
    .ZN(_08114_)
  );
  INV_X1 _18063_ (
    .A(_08114_),
    .ZN(_08115_)
  );
  AND2_X1 _18064_ (
    .A1(_08107_),
    .A2(_08114_),
    .ZN(_08117_)
  );
  INV_X1 _18065_ (
    .A(_08117_),
    .ZN(_08118_)
  );
  AND2_X1 _18066_ (
    .A1(_08106_),
    .A2(_08115_),
    .ZN(_08119_)
  );
  INV_X1 _18067_ (
    .A(_08119_),
    .ZN(_08120_)
  );
  AND2_X1 _18068_ (
    .A1(_08118_),
    .A2(_08120_),
    .ZN(_08121_)
  );
  INV_X1 _18069_ (
    .A(_08121_),
    .ZN(_08122_)
  );
  AND2_X1 _18070_ (
    .A1(_08103_),
    .A2(_08121_),
    .ZN(_08123_)
  );
  INV_X1 _18071_ (
    .A(_08123_),
    .ZN(_08124_)
  );
  AND2_X1 _18072_ (
    .A1(_08104_),
    .A2(_08122_),
    .ZN(_08125_)
  );
  INV_X1 _18073_ (
    .A(_08125_),
    .ZN(_08126_)
  );
  AND2_X1 _18074_ (
    .A1(_08124_),
    .A2(_08126_),
    .ZN(_08128_)
  );
  INV_X1 _18075_ (
    .A(_08128_),
    .ZN(_08129_)
  );
  AND2_X1 _18076_ (
    .A1(_07892_),
    .A2(_08128_),
    .ZN(_08130_)
  );
  INV_X1 _18077_ (
    .A(_08130_),
    .ZN(_08131_)
  );
  AND2_X1 _18078_ (
    .A1(_07891_),
    .A2(_08129_),
    .ZN(_08132_)
  );
  INV_X1 _18079_ (
    .A(_08132_),
    .ZN(_08133_)
  );
  AND2_X1 _18080_ (
    .A1(_08131_),
    .A2(_08133_),
    .ZN(_08134_)
  );
  INV_X1 _18081_ (
    .A(_08134_),
    .ZN(_08135_)
  );
  AND2_X1 _18082_ (
    .A1(_07890_),
    .A2(_08134_),
    .ZN(_08136_)
  );
  INV_X1 _18083_ (
    .A(_08136_),
    .ZN(_08137_)
  );
  AND2_X1 _18084_ (
    .A1(_07889_),
    .A2(_08135_),
    .ZN(_08139_)
  );
  INV_X1 _18085_ (
    .A(_08139_),
    .ZN(_08140_)
  );
  AND2_X1 _18086_ (
    .A1(_08137_),
    .A2(_08140_),
    .ZN(_08141_)
  );
  INV_X1 _18087_ (
    .A(_08141_),
    .ZN(_08142_)
  );
  AND2_X1 _18088_ (
    .A1(_07888_),
    .A2(_08141_),
    .ZN(_08143_)
  );
  INV_X1 _18089_ (
    .A(_08143_),
    .ZN(_08144_)
  );
  AND2_X1 _18090_ (
    .A1(_07887_),
    .A2(_08142_),
    .ZN(_08145_)
  );
  INV_X1 _18091_ (
    .A(_08145_),
    .ZN(_08146_)
  );
  AND2_X1 _18092_ (
    .A1(_08144_),
    .A2(_08146_),
    .ZN(_08147_)
  );
  INV_X1 _18093_ (
    .A(_08147_),
    .ZN(_08148_)
  );
  AND2_X1 _18094_ (
    .A1(_07839_),
    .A2(_08147_),
    .ZN(_08150_)
  );
  INV_X1 _18095_ (
    .A(_08150_),
    .ZN(_08151_)
  );
  AND2_X1 _18096_ (
    .A1(_07840_),
    .A2(_08148_),
    .ZN(_08152_)
  );
  INV_X1 _18097_ (
    .A(_08152_),
    .ZN(_08153_)
  );
  AND2_X1 _18098_ (
    .A1(_08151_),
    .A2(_08153_),
    .ZN(_08154_)
  );
  INV_X1 _18099_ (
    .A(_08154_),
    .ZN(_08155_)
  );
  AND2_X1 _18100_ (
    .A1(_07595_),
    .A2(_07847_),
    .ZN(_08156_)
  );
  INV_X1 _18101_ (
    .A(_08156_),
    .ZN(_08157_)
  );
  AND2_X1 _18102_ (
    .A1(_07847_),
    .A2(_07856_),
    .ZN(_08158_)
  );
  AND2_X1 _18103_ (
    .A1(_07849_),
    .A2(_08157_),
    .ZN(_08159_)
  );
  AND2_X1 _18104_ (
    .A1(_08154_),
    .A2(_08159_),
    .ZN(_08161_)
  );
  INV_X1 _18105_ (
    .A(_08161_),
    .ZN(_08162_)
  );
  AND2_X1 _18106_ (
    .A1(_08155_),
    .A2(_08158_),
    .ZN(_08163_)
  );
  INV_X1 _18107_ (
    .A(_08163_),
    .ZN(_08164_)
  );
  AND2_X1 _18108_ (
    .A1(_08162_),
    .A2(_08164_),
    .ZN(_08165_)
  );
  INV_X1 _18109_ (
    .A(_08165_),
    .ZN(_08166_)
  );
  AND2_X1 _18110_ (
    .A1(remainder[61]),
    .A2(_08165_),
    .ZN(_08167_)
  );
  INV_X1 _18111_ (
    .A(_08167_),
    .ZN(_08168_)
  );
  AND2_X1 _18112_ (
    .A1(_04448_),
    .A2(_08166_),
    .ZN(_08169_)
  );
  INV_X1 _18113_ (
    .A(_08169_),
    .ZN(_08170_)
  );
  AND2_X1 _18114_ (
    .A1(_08168_),
    .A2(_08170_),
    .ZN(_08172_)
  );
  INV_X1 _18115_ (
    .A(_08172_),
    .ZN(_08173_)
  );
  AND2_X1 _18116_ (
    .A1(_07593_),
    .A2(_07860_),
    .ZN(_08174_)
  );
  INV_X1 _18117_ (
    .A(_08174_),
    .ZN(_08175_)
  );
  AND2_X1 _18118_ (
    .A1(_07862_),
    .A2(_08175_),
    .ZN(_08176_)
  );
  INV_X1 _18119_ (
    .A(_08176_),
    .ZN(_08177_)
  );
  AND2_X1 _18120_ (
    .A1(_08173_),
    .A2(_08177_),
    .ZN(_08178_)
  );
  INV_X1 _18121_ (
    .A(_08178_),
    .ZN(_08179_)
  );
  AND2_X1 _18122_ (
    .A1(_08172_),
    .A2(_08176_),
    .ZN(_08180_)
  );
  INV_X1 _18123_ (
    .A(_08180_),
    .ZN(_08181_)
  );
  AND2_X1 _18124_ (
    .A1(_02082_),
    .A2(_08181_),
    .ZN(_08183_)
  );
  AND2_X1 _18125_ (
    .A1(_08179_),
    .A2(_08183_),
    .ZN(_08184_)
  );
  INV_X1 _18126_ (
    .A(_08184_),
    .ZN(_08185_)
  );
  AND2_X1 _18127_ (
    .A1(remainder[53]),
    .A2(_02077_),
    .ZN(_08186_)
  );
  INV_X1 _18128_ (
    .A(_08186_),
    .ZN(_08187_)
  );
  AND2_X1 _18129_ (
    .A1(_10462_),
    .A2(_01905_),
    .ZN(_08188_)
  );
  INV_X1 _18130_ (
    .A(_08188_),
    .ZN(_08189_)
  );
  AND2_X1 _18131_ (
    .A1(_04546_),
    .A2(_10451_),
    .ZN(_08190_)
  );
  INV_X1 _18132_ (
    .A(_08190_),
    .ZN(_08191_)
  );
  AND2_X1 _18133_ (
    .A1(_05983_),
    .A2(_08189_),
    .ZN(_08192_)
  );
  AND2_X1 _18134_ (
    .A1(_08191_),
    .A2(_08192_),
    .ZN(_08194_)
  );
  INV_X1 _18135_ (
    .A(_08194_),
    .ZN(_08195_)
  );
  AND2_X1 _18136_ (
    .A1(_08187_),
    .A2(_08195_),
    .ZN(_08196_)
  );
  AND2_X1 _18137_ (
    .A1(_08185_),
    .A2(_08196_),
    .ZN(_08197_)
  );
  INV_X1 _18138_ (
    .A(_08197_),
    .ZN(_08198_)
  );
  AND2_X1 _18139_ (
    .A1(_06201_),
    .A2(_08198_),
    .ZN(_00074_)
  );
  AND2_X1 _18140_ (
    .A1(_08168_),
    .A2(_08181_),
    .ZN(_08199_)
  );
  INV_X1 _18141_ (
    .A(_08199_),
    .ZN(_08200_)
  );
  AND2_X1 _18142_ (
    .A1(_08151_),
    .A2(_08162_),
    .ZN(_08201_)
  );
  INV_X1 _18143_ (
    .A(_08201_),
    .ZN(_08202_)
  );
  AND2_X1 _18144_ (
    .A1(_08131_),
    .A2(_08137_),
    .ZN(_08204_)
  );
  INV_X1 _18145_ (
    .A(_08204_),
    .ZN(_08205_)
  );
  AND2_X1 _18146_ (
    .A1(_08111_),
    .A2(_08118_),
    .ZN(_08206_)
  );
  INV_X1 _18147_ (
    .A(_08206_),
    .ZN(_08207_)
  );
  AND2_X1 _18148_ (
    .A1(_08100_),
    .A2(_08124_),
    .ZN(_08208_)
  );
  INV_X1 _18149_ (
    .A(_08208_),
    .ZN(_08209_)
  );
  AND2_X1 _18150_ (
    .A1(_08023_),
    .A2(_08093_),
    .ZN(_08210_)
  );
  INV_X1 _18151_ (
    .A(_08210_),
    .ZN(_08211_)
  );
  AND2_X1 _18152_ (
    .A1(_07931_),
    .A2(_07991_),
    .ZN(_08212_)
  );
  INV_X1 _18153_ (
    .A(_08212_),
    .ZN(_08213_)
  );
  AND2_X1 _18154_ (
    .A1(_07911_),
    .A2(_07917_),
    .ZN(_08215_)
  );
  INV_X1 _18155_ (
    .A(_08215_),
    .ZN(_08216_)
  );
  AND2_X1 _18156_ (
    .A1(divisor[25]),
    .A2(remainder[4]),
    .ZN(_08217_)
  );
  INV_X1 _18157_ (
    .A(_08217_),
    .ZN(_08218_)
  );
  AND2_X1 _18158_ (
    .A1(divisor[26]),
    .A2(remainder[3]),
    .ZN(_08219_)
  );
  INV_X1 _18159_ (
    .A(_08219_),
    .ZN(_08220_)
  );
  AND2_X1 _18160_ (
    .A1(divisor[27]),
    .A2(remainder[3]),
    .ZN(_08221_)
  );
  INV_X1 _18161_ (
    .A(_08221_),
    .ZN(_08222_)
  );
  AND2_X1 _18162_ (
    .A1(_07908_),
    .A2(_08219_),
    .ZN(_08223_)
  );
  INV_X1 _18163_ (
    .A(_08223_),
    .ZN(_08224_)
  );
  AND2_X1 _18164_ (
    .A1(_07909_),
    .A2(_08220_),
    .ZN(_08226_)
  );
  INV_X1 _18165_ (
    .A(_08226_),
    .ZN(_08227_)
  );
  AND2_X1 _18166_ (
    .A1(_08224_),
    .A2(_08227_),
    .ZN(_08228_)
  );
  INV_X1 _18167_ (
    .A(_08228_),
    .ZN(_08229_)
  );
  AND2_X1 _18168_ (
    .A1(_08217_),
    .A2(_08228_),
    .ZN(_08230_)
  );
  INV_X1 _18169_ (
    .A(_08230_),
    .ZN(_08231_)
  );
  AND2_X1 _18170_ (
    .A1(_08218_),
    .A2(_08229_),
    .ZN(_08232_)
  );
  INV_X1 _18171_ (
    .A(_08232_),
    .ZN(_08233_)
  );
  AND2_X1 _18172_ (
    .A1(_08231_),
    .A2(_08233_),
    .ZN(_08234_)
  );
  INV_X1 _18173_ (
    .A(_08234_),
    .ZN(_08235_)
  );
  AND2_X1 _18174_ (
    .A1(_08216_),
    .A2(_08234_),
    .ZN(_08237_)
  );
  INV_X1 _18175_ (
    .A(_08237_),
    .ZN(_08238_)
  );
  AND2_X1 _18176_ (
    .A1(_08215_),
    .A2(_08235_),
    .ZN(_08239_)
  );
  INV_X1 _18177_ (
    .A(_08239_),
    .ZN(_08240_)
  );
  AND2_X1 _18178_ (
    .A1(_08238_),
    .A2(_08240_),
    .ZN(_08241_)
  );
  INV_X1 _18179_ (
    .A(_08241_),
    .ZN(_08242_)
  );
  AND2_X1 _18180_ (
    .A1(_07923_),
    .A2(_08241_),
    .ZN(_08243_)
  );
  INV_X1 _18181_ (
    .A(_08243_),
    .ZN(_08244_)
  );
  AND2_X1 _18182_ (
    .A1(_07924_),
    .A2(_08242_),
    .ZN(_08245_)
  );
  INV_X1 _18183_ (
    .A(_08245_),
    .ZN(_08246_)
  );
  AND2_X1 _18184_ (
    .A1(_08244_),
    .A2(_08246_),
    .ZN(_08248_)
  );
  INV_X1 _18185_ (
    .A(_08248_),
    .ZN(_08249_)
  );
  AND2_X1 _18186_ (
    .A1(_07946_),
    .A2(_07953_),
    .ZN(_08250_)
  );
  INV_X1 _18187_ (
    .A(_08250_),
    .ZN(_08251_)
  );
  AND2_X1 _18188_ (
    .A1(divisor[22]),
    .A2(remainder[7]),
    .ZN(_08252_)
  );
  INV_X1 _18189_ (
    .A(_08252_),
    .ZN(_08253_)
  );
  AND2_X1 _18190_ (
    .A1(divisor[23]),
    .A2(remainder[6]),
    .ZN(_08254_)
  );
  INV_X1 _18191_ (
    .A(_08254_),
    .ZN(_08255_)
  );
  AND2_X1 _18192_ (
    .A1(divisor[24]),
    .A2(remainder[6]),
    .ZN(_08256_)
  );
  INV_X1 _18193_ (
    .A(_08256_),
    .ZN(_08257_)
  );
  AND2_X1 _18194_ (
    .A1(_07943_),
    .A2(_08254_),
    .ZN(_08259_)
  );
  INV_X1 _18195_ (
    .A(_08259_),
    .ZN(_08260_)
  );
  AND2_X1 _18196_ (
    .A1(_07944_),
    .A2(_08255_),
    .ZN(_08261_)
  );
  INV_X1 _18197_ (
    .A(_08261_),
    .ZN(_08262_)
  );
  AND2_X1 _18198_ (
    .A1(_08260_),
    .A2(_08262_),
    .ZN(_08263_)
  );
  INV_X1 _18199_ (
    .A(_08263_),
    .ZN(_08264_)
  );
  AND2_X1 _18200_ (
    .A1(_08252_),
    .A2(_08263_),
    .ZN(_08265_)
  );
  INV_X1 _18201_ (
    .A(_08265_),
    .ZN(_08266_)
  );
  AND2_X1 _18202_ (
    .A1(_08253_),
    .A2(_08264_),
    .ZN(_08267_)
  );
  INV_X1 _18203_ (
    .A(_08267_),
    .ZN(_08268_)
  );
  AND2_X1 _18204_ (
    .A1(_08266_),
    .A2(_08268_),
    .ZN(_08270_)
  );
  INV_X1 _18205_ (
    .A(_08270_),
    .ZN(_08271_)
  );
  AND2_X1 _18206_ (
    .A1(_08251_),
    .A2(_08270_),
    .ZN(_08272_)
  );
  INV_X1 _18207_ (
    .A(_08272_),
    .ZN(_08273_)
  );
  AND2_X1 _18208_ (
    .A1(_08250_),
    .A2(_08271_),
    .ZN(_08274_)
  );
  INV_X1 _18209_ (
    .A(_08274_),
    .ZN(_08275_)
  );
  AND2_X1 _18210_ (
    .A1(_08273_),
    .A2(_08275_),
    .ZN(_08276_)
  );
  INV_X1 _18211_ (
    .A(_08276_),
    .ZN(_08277_)
  );
  MUX2_X1 _18212_ (
    .A(_07966_),
    .B(_04996_),
    .S(_07965_),
    .Z(_08278_)
  );
  AND2_X1 _18213_ (
    .A1(divisor[19]),
    .A2(_08278_),
    .ZN(_08279_)
  );
  INV_X1 _18214_ (
    .A(_08279_),
    .ZN(_08281_)
  );
  MUX2_X1 _18215_ (
    .A(_05269_),
    .B(_04985_),
    .S(_08278_),
    .Z(_08282_)
  );
  MUX2_X1 _18216_ (
    .A(_05271_),
    .B(divisor[19]),
    .S(_08278_),
    .Z(_08283_)
  );
  AND2_X1 _18217_ (
    .A1(_08276_),
    .A2(_08282_),
    .ZN(_08284_)
  );
  INV_X1 _18218_ (
    .A(_08284_),
    .ZN(_08285_)
  );
  AND2_X1 _18219_ (
    .A1(_08277_),
    .A2(_08283_),
    .ZN(_08286_)
  );
  INV_X1 _18220_ (
    .A(_08286_),
    .ZN(_08287_)
  );
  AND2_X1 _18221_ (
    .A1(_08285_),
    .A2(_08287_),
    .ZN(_08288_)
  );
  INV_X1 _18222_ (
    .A(_08288_),
    .ZN(_08289_)
  );
  AND2_X1 _18223_ (
    .A1(_08248_),
    .A2(_08288_),
    .ZN(_08290_)
  );
  INV_X1 _18224_ (
    .A(_08290_),
    .ZN(_08292_)
  );
  AND2_X1 _18225_ (
    .A1(_08249_),
    .A2(_08289_),
    .ZN(_08293_)
  );
  INV_X1 _18226_ (
    .A(_08293_),
    .ZN(_08294_)
  );
  AND2_X1 _18227_ (
    .A1(_08292_),
    .A2(_08294_),
    .ZN(_08295_)
  );
  INV_X1 _18228_ (
    .A(_08295_),
    .ZN(_08296_)
  );
  AND2_X1 _18229_ (
    .A1(_08213_),
    .A2(_08295_),
    .ZN(_08297_)
  );
  INV_X1 _18230_ (
    .A(_08297_),
    .ZN(_08298_)
  );
  AND2_X1 _18231_ (
    .A1(_08212_),
    .A2(_08296_),
    .ZN(_08299_)
  );
  INV_X1 _18232_ (
    .A(_08299_),
    .ZN(_08300_)
  );
  AND2_X1 _18233_ (
    .A1(_08298_),
    .A2(_08300_),
    .ZN(_08301_)
  );
  INV_X1 _18234_ (
    .A(_08301_),
    .ZN(_08303_)
  );
  AND2_X1 _18235_ (
    .A1(divisor[29]),
    .A2(remainder[0]),
    .ZN(_08304_)
  );
  INV_X1 _18236_ (
    .A(_08304_),
    .ZN(_08305_)
  );
  AND2_X1 _18237_ (
    .A1(divisor[28]),
    .A2(remainder[1]),
    .ZN(_08306_)
  );
  INV_X1 _18238_ (
    .A(_08306_),
    .ZN(_08307_)
  );
  AND2_X1 _18239_ (
    .A1(divisor[29]),
    .A2(remainder[1]),
    .ZN(_08308_)
  );
  INV_X1 _18240_ (
    .A(_08308_),
    .ZN(_08309_)
  );
  AND2_X1 _18241_ (
    .A1(_08003_),
    .A2(_08308_),
    .ZN(_08310_)
  );
  INV_X1 _18242_ (
    .A(_08310_),
    .ZN(_08311_)
  );
  AND2_X1 _18243_ (
    .A1(_08305_),
    .A2(_08307_),
    .ZN(_08312_)
  );
  INV_X1 _18244_ (
    .A(_08312_),
    .ZN(_08314_)
  );
  AND2_X1 _18245_ (
    .A1(_08311_),
    .A2(_08314_),
    .ZN(_08315_)
  );
  INV_X1 _18246_ (
    .A(_08315_),
    .ZN(_08316_)
  );
  AND2_X1 _18247_ (
    .A1(_08009_),
    .A2(_08316_),
    .ZN(_08317_)
  );
  INV_X1 _18248_ (
    .A(_08317_),
    .ZN(_08318_)
  );
  AND2_X1 _18249_ (
    .A1(_08010_),
    .A2(_08315_),
    .ZN(_08319_)
  );
  INV_X1 _18250_ (
    .A(_08319_),
    .ZN(_08320_)
  );
  AND2_X1 _18251_ (
    .A1(_08009_),
    .A2(_08315_),
    .ZN(_08321_)
  );
  INV_X1 _18252_ (
    .A(_08321_),
    .ZN(_08322_)
  );
  AND2_X1 _18253_ (
    .A1(_08010_),
    .A2(_08316_),
    .ZN(_08323_)
  );
  INV_X1 _18254_ (
    .A(_08323_),
    .ZN(_08325_)
  );
  AND2_X1 _18255_ (
    .A1(_08318_),
    .A2(_08320_),
    .ZN(_08326_)
  );
  AND2_X1 _18256_ (
    .A1(_08322_),
    .A2(_08325_),
    .ZN(_08327_)
  );
  AND2_X1 _18257_ (
    .A1(_08301_),
    .A2(_08327_),
    .ZN(_08328_)
  );
  INV_X1 _18258_ (
    .A(_08328_),
    .ZN(_08329_)
  );
  AND2_X1 _18259_ (
    .A1(_08303_),
    .A2(_08326_),
    .ZN(_08330_)
  );
  INV_X1 _18260_ (
    .A(_08330_),
    .ZN(_08331_)
  );
  AND2_X1 _18261_ (
    .A1(_08329_),
    .A2(_08331_),
    .ZN(_08332_)
  );
  INV_X1 _18262_ (
    .A(_08332_),
    .ZN(_08333_)
  );
  AND2_X1 _18263_ (
    .A1(_08015_),
    .A2(_08332_),
    .ZN(_08334_)
  );
  INV_X1 _18264_ (
    .A(_08334_),
    .ZN(_08336_)
  );
  AND2_X1 _18265_ (
    .A1(_08016_),
    .A2(_08333_),
    .ZN(_08337_)
  );
  INV_X1 _18266_ (
    .A(_08337_),
    .ZN(_08338_)
  );
  AND2_X1 _18267_ (
    .A1(_08336_),
    .A2(_08338_),
    .ZN(_08339_)
  );
  INV_X1 _18268_ (
    .A(_08339_),
    .ZN(_08340_)
  );
  AND2_X1 _18269_ (
    .A1(_08067_),
    .A2(_08074_),
    .ZN(_08341_)
  );
  INV_X1 _18270_ (
    .A(_08341_),
    .ZN(_08342_)
  );
  AND2_X1 _18271_ (
    .A1(_08054_),
    .A2(_08060_),
    .ZN(_08343_)
  );
  INV_X1 _18272_ (
    .A(_08343_),
    .ZN(_08344_)
  );
  AND2_X1 _18273_ (
    .A1(_08041_),
    .A2(_08047_),
    .ZN(_08345_)
  );
  INV_X1 _18274_ (
    .A(_08345_),
    .ZN(_08347_)
  );
  AND2_X1 _18275_ (
    .A1(_07959_),
    .A2(_07985_),
    .ZN(_08348_)
  );
  INV_X1 _18276_ (
    .A(_08348_),
    .ZN(_08349_)
  );
  AND2_X1 _18277_ (
    .A1(_07971_),
    .A2(_07978_),
    .ZN(_08350_)
  );
  INV_X1 _18278_ (
    .A(_08350_),
    .ZN(_08351_)
  );
  AND2_X1 _18279_ (
    .A1(_07319_),
    .A2(_08351_),
    .ZN(_08352_)
  );
  INV_X1 _18280_ (
    .A(_08352_),
    .ZN(_08353_)
  );
  AND2_X1 _18281_ (
    .A1(_07320_),
    .A2(_08350_),
    .ZN(_08354_)
  );
  INV_X1 _18282_ (
    .A(_08354_),
    .ZN(_08355_)
  );
  AND2_X1 _18283_ (
    .A1(_08353_),
    .A2(_08355_),
    .ZN(_08356_)
  );
  INV_X1 _18284_ (
    .A(_08356_),
    .ZN(_08358_)
  );
  AND2_X1 _18285_ (
    .A1(_07620_),
    .A2(_08356_),
    .ZN(_08359_)
  );
  INV_X1 _18286_ (
    .A(_08359_),
    .ZN(_08360_)
  );
  AND2_X1 _18287_ (
    .A1(_07619_),
    .A2(_08358_),
    .ZN(_08361_)
  );
  INV_X1 _18288_ (
    .A(_08361_),
    .ZN(_08362_)
  );
  AND2_X1 _18289_ (
    .A1(_08360_),
    .A2(_08362_),
    .ZN(_08363_)
  );
  INV_X1 _18290_ (
    .A(_08363_),
    .ZN(_08364_)
  );
  AND2_X1 _18291_ (
    .A1(_08349_),
    .A2(_08363_),
    .ZN(_08365_)
  );
  INV_X1 _18292_ (
    .A(_08365_),
    .ZN(_08366_)
  );
  AND2_X1 _18293_ (
    .A1(_08348_),
    .A2(_08364_),
    .ZN(_08367_)
  );
  INV_X1 _18294_ (
    .A(_08367_),
    .ZN(_08369_)
  );
  AND2_X1 _18295_ (
    .A1(_08366_),
    .A2(_08369_),
    .ZN(_08370_)
  );
  INV_X1 _18296_ (
    .A(_08370_),
    .ZN(_08371_)
  );
  AND2_X1 _18297_ (
    .A1(_08347_),
    .A2(_08370_),
    .ZN(_08372_)
  );
  INV_X1 _18298_ (
    .A(_08372_),
    .ZN(_08373_)
  );
  AND2_X1 _18299_ (
    .A1(_08345_),
    .A2(_08371_),
    .ZN(_08374_)
  );
  INV_X1 _18300_ (
    .A(_08374_),
    .ZN(_08375_)
  );
  AND2_X1 _18301_ (
    .A1(_08373_),
    .A2(_08375_),
    .ZN(_08376_)
  );
  INV_X1 _18302_ (
    .A(_08376_),
    .ZN(_08377_)
  );
  AND2_X1 _18303_ (
    .A1(_08344_),
    .A2(_08376_),
    .ZN(_08378_)
  );
  INV_X1 _18304_ (
    .A(_08378_),
    .ZN(_08380_)
  );
  AND2_X1 _18305_ (
    .A1(_08343_),
    .A2(_08377_),
    .ZN(_08381_)
  );
  INV_X1 _18306_ (
    .A(_08381_),
    .ZN(_08382_)
  );
  AND2_X1 _18307_ (
    .A1(_08380_),
    .A2(_08382_),
    .ZN(_08383_)
  );
  INV_X1 _18308_ (
    .A(_08383_),
    .ZN(_08384_)
  );
  AND2_X1 _18309_ (
    .A1(_07082_),
    .A2(_08383_),
    .ZN(_08385_)
  );
  INV_X1 _18310_ (
    .A(_08385_),
    .ZN(_08386_)
  );
  AND2_X1 _18311_ (
    .A1(_07083_),
    .A2(_08384_),
    .ZN(_08387_)
  );
  INV_X1 _18312_ (
    .A(_08387_),
    .ZN(_08388_)
  );
  AND2_X1 _18313_ (
    .A1(_08386_),
    .A2(_08388_),
    .ZN(_08389_)
  );
  INV_X1 _18314_ (
    .A(_08389_),
    .ZN(_08391_)
  );
  AND2_X1 _18315_ (
    .A1(_07997_),
    .A2(_08389_),
    .ZN(_08392_)
  );
  INV_X1 _18316_ (
    .A(_08392_),
    .ZN(_08393_)
  );
  AND2_X1 _18317_ (
    .A1(_07998_),
    .A2(_08391_),
    .ZN(_08394_)
  );
  INV_X1 _18318_ (
    .A(_08394_),
    .ZN(_08395_)
  );
  AND2_X1 _18319_ (
    .A1(_08393_),
    .A2(_08395_),
    .ZN(_08396_)
  );
  INV_X1 _18320_ (
    .A(_08396_),
    .ZN(_08397_)
  );
  AND2_X1 _18321_ (
    .A1(_08342_),
    .A2(_08396_),
    .ZN(_08398_)
  );
  INV_X1 _18322_ (
    .A(_08398_),
    .ZN(_08399_)
  );
  AND2_X1 _18323_ (
    .A1(_08341_),
    .A2(_08397_),
    .ZN(_08400_)
  );
  INV_X1 _18324_ (
    .A(_08400_),
    .ZN(_08402_)
  );
  AND2_X1 _18325_ (
    .A1(_08399_),
    .A2(_08402_),
    .ZN(_08403_)
  );
  INV_X1 _18326_ (
    .A(_08403_),
    .ZN(_08404_)
  );
  AND2_X1 _18327_ (
    .A1(_08339_),
    .A2(_08403_),
    .ZN(_08405_)
  );
  INV_X1 _18328_ (
    .A(_08405_),
    .ZN(_08406_)
  );
  AND2_X1 _18329_ (
    .A1(_08340_),
    .A2(_08404_),
    .ZN(_08407_)
  );
  INV_X1 _18330_ (
    .A(_08407_),
    .ZN(_08408_)
  );
  AND2_X1 _18331_ (
    .A1(_08406_),
    .A2(_08408_),
    .ZN(_08409_)
  );
  INV_X1 _18332_ (
    .A(_08409_),
    .ZN(_08410_)
  );
  AND2_X1 _18333_ (
    .A1(_08211_),
    .A2(_08409_),
    .ZN(_08411_)
  );
  INV_X1 _18334_ (
    .A(_08411_),
    .ZN(_08413_)
  );
  AND2_X1 _18335_ (
    .A1(_08210_),
    .A2(_08410_),
    .ZN(_08414_)
  );
  INV_X1 _18336_ (
    .A(_08414_),
    .ZN(_08415_)
  );
  AND2_X1 _18337_ (
    .A1(_08413_),
    .A2(_08415_),
    .ZN(_08416_)
  );
  INV_X1 _18338_ (
    .A(_08416_),
    .ZN(_08417_)
  );
  AND2_X1 _18339_ (
    .A1(_08080_),
    .A2(_08087_),
    .ZN(_08418_)
  );
  INV_X1 _18340_ (
    .A(_08418_),
    .ZN(_08419_)
  );
  AND2_X1 _18341_ (
    .A1(_07804_),
    .A2(_08419_),
    .ZN(_08420_)
  );
  INV_X1 _18342_ (
    .A(_08420_),
    .ZN(_08421_)
  );
  AND2_X1 _18343_ (
    .A1(_07805_),
    .A2(_08418_),
    .ZN(_08422_)
  );
  INV_X1 _18344_ (
    .A(_08422_),
    .ZN(_08424_)
  );
  AND2_X1 _18345_ (
    .A1(_08421_),
    .A2(_08424_),
    .ZN(_08425_)
  );
  INV_X1 _18346_ (
    .A(_08425_),
    .ZN(_08426_)
  );
  AND2_X1 _18347_ (
    .A1(_08107_),
    .A2(_08425_),
    .ZN(_08427_)
  );
  INV_X1 _18348_ (
    .A(_08427_),
    .ZN(_08428_)
  );
  AND2_X1 _18349_ (
    .A1(_08106_),
    .A2(_08426_),
    .ZN(_08429_)
  );
  INV_X1 _18350_ (
    .A(_08429_),
    .ZN(_08430_)
  );
  AND2_X1 _18351_ (
    .A1(_08428_),
    .A2(_08430_),
    .ZN(_08431_)
  );
  INV_X1 _18352_ (
    .A(_08431_),
    .ZN(_08432_)
  );
  AND2_X1 _18353_ (
    .A1(_08416_),
    .A2(_08431_),
    .ZN(_08433_)
  );
  INV_X1 _18354_ (
    .A(_08433_),
    .ZN(_08435_)
  );
  AND2_X1 _18355_ (
    .A1(_08417_),
    .A2(_08432_),
    .ZN(_08436_)
  );
  INV_X1 _18356_ (
    .A(_08436_),
    .ZN(_08437_)
  );
  AND2_X1 _18357_ (
    .A1(_08435_),
    .A2(_08437_),
    .ZN(_08438_)
  );
  INV_X1 _18358_ (
    .A(_08438_),
    .ZN(_08439_)
  );
  AND2_X1 _18359_ (
    .A1(_08209_),
    .A2(_08438_),
    .ZN(_08440_)
  );
  INV_X1 _18360_ (
    .A(_08440_),
    .ZN(_08441_)
  );
  AND2_X1 _18361_ (
    .A1(_08208_),
    .A2(_08439_),
    .ZN(_08442_)
  );
  INV_X1 _18362_ (
    .A(_08442_),
    .ZN(_08443_)
  );
  AND2_X1 _18363_ (
    .A1(_08441_),
    .A2(_08443_),
    .ZN(_08444_)
  );
  INV_X1 _18364_ (
    .A(_08444_),
    .ZN(_08446_)
  );
  AND2_X1 _18365_ (
    .A1(_08207_),
    .A2(_08444_),
    .ZN(_08447_)
  );
  INV_X1 _18366_ (
    .A(_08447_),
    .ZN(_08448_)
  );
  AND2_X1 _18367_ (
    .A1(_08206_),
    .A2(_08446_),
    .ZN(_08449_)
  );
  INV_X1 _18368_ (
    .A(_08449_),
    .ZN(_08450_)
  );
  AND2_X1 _18369_ (
    .A1(_08448_),
    .A2(_08450_),
    .ZN(_08451_)
  );
  INV_X1 _18370_ (
    .A(_08451_),
    .ZN(_08452_)
  );
  AND2_X1 _18371_ (
    .A1(_08205_),
    .A2(_08451_),
    .ZN(_08453_)
  );
  INV_X1 _18372_ (
    .A(_08453_),
    .ZN(_08454_)
  );
  AND2_X1 _18373_ (
    .A1(_08204_),
    .A2(_08452_),
    .ZN(_08455_)
  );
  INV_X1 _18374_ (
    .A(_08455_),
    .ZN(_08457_)
  );
  AND2_X1 _18375_ (
    .A1(_08454_),
    .A2(_08457_),
    .ZN(_08458_)
  );
  INV_X1 _18376_ (
    .A(_08458_),
    .ZN(_08459_)
  );
  AND2_X1 _18377_ (
    .A1(_08143_),
    .A2(_08458_),
    .ZN(_08460_)
  );
  INV_X1 _18378_ (
    .A(_08460_),
    .ZN(_08461_)
  );
  AND2_X1 _18379_ (
    .A1(_08144_),
    .A2(_08459_),
    .ZN(_08462_)
  );
  INV_X1 _18380_ (
    .A(_08462_),
    .ZN(_08463_)
  );
  AND2_X1 _18381_ (
    .A1(_08461_),
    .A2(_08463_),
    .ZN(_08464_)
  );
  INV_X1 _18382_ (
    .A(_08464_),
    .ZN(_08465_)
  );
  AND2_X1 _18383_ (
    .A1(_08202_),
    .A2(_08465_),
    .ZN(_08466_)
  );
  INV_X1 _18384_ (
    .A(_08466_),
    .ZN(_08468_)
  );
  AND2_X1 _18385_ (
    .A1(_08201_),
    .A2(_08464_),
    .ZN(_08469_)
  );
  INV_X1 _18386_ (
    .A(_08469_),
    .ZN(_08470_)
  );
  AND2_X1 _18387_ (
    .A1(_08468_),
    .A2(_08470_),
    .ZN(_08471_)
  );
  INV_X1 _18388_ (
    .A(_08471_),
    .ZN(_08472_)
  );
  AND2_X1 _18389_ (
    .A1(remainder[62]),
    .A2(_08472_),
    .ZN(_08473_)
  );
  INV_X1 _18390_ (
    .A(_08473_),
    .ZN(_08474_)
  );
  AND2_X1 _18391_ (
    .A1(_04437_),
    .A2(_08471_),
    .ZN(_08475_)
  );
  INV_X1 _18392_ (
    .A(_08475_),
    .ZN(_08476_)
  );
  AND2_X1 _18393_ (
    .A1(_08474_),
    .A2(_08476_),
    .ZN(_08477_)
  );
  INV_X1 _18394_ (
    .A(_08477_),
    .ZN(_08479_)
  );
  AND2_X1 _18395_ (
    .A1(_08199_),
    .A2(_08479_),
    .ZN(_08480_)
  );
  INV_X1 _18396_ (
    .A(_08480_),
    .ZN(_08481_)
  );
  AND2_X1 _18397_ (
    .A1(_08200_),
    .A2(_08477_),
    .ZN(_08482_)
  );
  INV_X1 _18398_ (
    .A(_08482_),
    .ZN(_08483_)
  );
  AND2_X1 _18399_ (
    .A1(_08481_),
    .A2(_08483_),
    .ZN(_08484_)
  );
  AND2_X1 _18400_ (
    .A1(_02082_),
    .A2(_08484_),
    .ZN(_08485_)
  );
  INV_X1 _18401_ (
    .A(_08485_),
    .ZN(_08486_)
  );
  AND2_X1 _18402_ (
    .A1(remainder[54]),
    .A2(_02077_),
    .ZN(_08487_)
  );
  INV_X1 _18403_ (
    .A(_08487_),
    .ZN(_08488_)
  );
  AND2_X1 _18404_ (
    .A1(_10462_),
    .A2(_01924_),
    .ZN(_08490_)
  );
  INV_X1 _18405_ (
    .A(_08490_),
    .ZN(_08491_)
  );
  AND2_X1 _18406_ (
    .A1(_04536_),
    .A2(_10451_),
    .ZN(_08492_)
  );
  INV_X1 _18407_ (
    .A(_08492_),
    .ZN(_08493_)
  );
  AND2_X1 _18408_ (
    .A1(_05983_),
    .A2(_08491_),
    .ZN(_08494_)
  );
  AND2_X1 _18409_ (
    .A1(_08493_),
    .A2(_08494_),
    .ZN(_08495_)
  );
  INV_X1 _18410_ (
    .A(_08495_),
    .ZN(_08496_)
  );
  AND2_X1 _18411_ (
    .A1(_08488_),
    .A2(_08496_),
    .ZN(_08497_)
  );
  AND2_X1 _18412_ (
    .A1(_08486_),
    .A2(_08497_),
    .ZN(_08498_)
  );
  INV_X1 _18413_ (
    .A(_08498_),
    .ZN(_08499_)
  );
  AND2_X1 _18414_ (
    .A1(_06201_),
    .A2(_08499_),
    .ZN(_00075_)
  );
  AND2_X1 _18415_ (
    .A1(_08441_),
    .A2(_08448_),
    .ZN(_08501_)
  );
  INV_X1 _18416_ (
    .A(_08501_),
    .ZN(_08502_)
  );
  AND2_X1 _18417_ (
    .A1(_08421_),
    .A2(_08428_),
    .ZN(_08503_)
  );
  INV_X1 _18418_ (
    .A(_08503_),
    .ZN(_08504_)
  );
  AND2_X1 _18419_ (
    .A1(_08413_),
    .A2(_08435_),
    .ZN(_08505_)
  );
  INV_X1 _18420_ (
    .A(_08505_),
    .ZN(_08506_)
  );
  AND2_X1 _18421_ (
    .A1(_08336_),
    .A2(_08406_),
    .ZN(_08507_)
  );
  INV_X1 _18422_ (
    .A(_08507_),
    .ZN(_08508_)
  );
  AND2_X1 _18423_ (
    .A1(_08008_),
    .A2(_08316_),
    .ZN(_08509_)
  );
  INV_X1 _18424_ (
    .A(_08509_),
    .ZN(_08511_)
  );
  AND2_X1 _18425_ (
    .A1(_08329_),
    .A2(_08511_),
    .ZN(_08512_)
  );
  INV_X1 _18426_ (
    .A(_08512_),
    .ZN(_08513_)
  );
  AND2_X1 _18427_ (
    .A1(_08244_),
    .A2(_08292_),
    .ZN(_08514_)
  );
  INV_X1 _18428_ (
    .A(_08514_),
    .ZN(_08515_)
  );
  AND2_X1 _18429_ (
    .A1(_08224_),
    .A2(_08231_),
    .ZN(_08516_)
  );
  INV_X1 _18430_ (
    .A(_08516_),
    .ZN(_08517_)
  );
  AND2_X1 _18431_ (
    .A1(divisor[25]),
    .A2(remainder[5]),
    .ZN(_08518_)
  );
  INV_X1 _18432_ (
    .A(_08518_),
    .ZN(_08519_)
  );
  AND2_X1 _18433_ (
    .A1(divisor[26]),
    .A2(remainder[4]),
    .ZN(_08520_)
  );
  INV_X1 _18434_ (
    .A(_08520_),
    .ZN(_08522_)
  );
  AND2_X1 _18435_ (
    .A1(divisor[27]),
    .A2(remainder[4]),
    .ZN(_08523_)
  );
  INV_X1 _18436_ (
    .A(_08523_),
    .ZN(_08524_)
  );
  AND2_X1 _18437_ (
    .A1(_08221_),
    .A2(_08520_),
    .ZN(_08525_)
  );
  INV_X1 _18438_ (
    .A(_08525_),
    .ZN(_08526_)
  );
  AND2_X1 _18439_ (
    .A1(_08222_),
    .A2(_08522_),
    .ZN(_08527_)
  );
  INV_X1 _18440_ (
    .A(_08527_),
    .ZN(_08528_)
  );
  AND2_X1 _18441_ (
    .A1(_08526_),
    .A2(_08528_),
    .ZN(_08529_)
  );
  INV_X1 _18442_ (
    .A(_08529_),
    .ZN(_08530_)
  );
  AND2_X1 _18443_ (
    .A1(_08518_),
    .A2(_08529_),
    .ZN(_08531_)
  );
  INV_X1 _18444_ (
    .A(_08531_),
    .ZN(_08533_)
  );
  AND2_X1 _18445_ (
    .A1(_08519_),
    .A2(_08530_),
    .ZN(_08534_)
  );
  INV_X1 _18446_ (
    .A(_08534_),
    .ZN(_08535_)
  );
  AND2_X1 _18447_ (
    .A1(_08533_),
    .A2(_08535_),
    .ZN(_08536_)
  );
  INV_X1 _18448_ (
    .A(_08536_),
    .ZN(_08537_)
  );
  AND2_X1 _18449_ (
    .A1(_08310_),
    .A2(_08536_),
    .ZN(_08538_)
  );
  INV_X1 _18450_ (
    .A(_08538_),
    .ZN(_08539_)
  );
  AND2_X1 _18451_ (
    .A1(_08311_),
    .A2(_08537_),
    .ZN(_08540_)
  );
  INV_X1 _18452_ (
    .A(_08540_),
    .ZN(_08541_)
  );
  AND2_X1 _18453_ (
    .A1(_08539_),
    .A2(_08541_),
    .ZN(_08542_)
  );
  INV_X1 _18454_ (
    .A(_08542_),
    .ZN(_08544_)
  );
  AND2_X1 _18455_ (
    .A1(_08517_),
    .A2(_08542_),
    .ZN(_08545_)
  );
  INV_X1 _18456_ (
    .A(_08545_),
    .ZN(_08546_)
  );
  AND2_X1 _18457_ (
    .A1(_08516_),
    .A2(_08544_),
    .ZN(_08547_)
  );
  INV_X1 _18458_ (
    .A(_08547_),
    .ZN(_08548_)
  );
  AND2_X1 _18459_ (
    .A1(_08546_),
    .A2(_08548_),
    .ZN(_08549_)
  );
  INV_X1 _18460_ (
    .A(_08549_),
    .ZN(_08550_)
  );
  AND2_X1 _18461_ (
    .A1(_08237_),
    .A2(_08549_),
    .ZN(_08551_)
  );
  INV_X1 _18462_ (
    .A(_08551_),
    .ZN(_08552_)
  );
  AND2_X1 _18463_ (
    .A1(_08238_),
    .A2(_08550_),
    .ZN(_08553_)
  );
  INV_X1 _18464_ (
    .A(_08553_),
    .ZN(_08555_)
  );
  AND2_X1 _18465_ (
    .A1(_08552_),
    .A2(_08555_),
    .ZN(_08556_)
  );
  INV_X1 _18466_ (
    .A(_08556_),
    .ZN(_08557_)
  );
  AND2_X1 _18467_ (
    .A1(_08260_),
    .A2(_08266_),
    .ZN(_08558_)
  );
  INV_X1 _18468_ (
    .A(_08558_),
    .ZN(_08559_)
  );
  AND2_X1 _18469_ (
    .A1(remainder[32]),
    .A2(divisor[22]),
    .ZN(_08560_)
  );
  INV_X1 _18470_ (
    .A(_08560_),
    .ZN(_08561_)
  );
  AND2_X1 _18471_ (
    .A1(divisor[23]),
    .A2(remainder[7]),
    .ZN(_08562_)
  );
  INV_X1 _18472_ (
    .A(_08562_),
    .ZN(_08563_)
  );
  AND2_X1 _18473_ (
    .A1(divisor[24]),
    .A2(remainder[7]),
    .ZN(_08564_)
  );
  INV_X1 _18474_ (
    .A(_08564_),
    .ZN(_08566_)
  );
  AND2_X1 _18475_ (
    .A1(_08254_),
    .A2(_08564_),
    .ZN(_08567_)
  );
  INV_X1 _18476_ (
    .A(_08567_),
    .ZN(_08568_)
  );
  AND2_X1 _18477_ (
    .A1(_08257_),
    .A2(_08563_),
    .ZN(_08569_)
  );
  INV_X1 _18478_ (
    .A(_08569_),
    .ZN(_08570_)
  );
  AND2_X1 _18479_ (
    .A1(_08568_),
    .A2(_08570_),
    .ZN(_08571_)
  );
  INV_X1 _18480_ (
    .A(_08571_),
    .ZN(_08572_)
  );
  AND2_X1 _18481_ (
    .A1(_08560_),
    .A2(_08571_),
    .ZN(_08573_)
  );
  INV_X1 _18482_ (
    .A(_08573_),
    .ZN(_08574_)
  );
  AND2_X1 _18483_ (
    .A1(_08561_),
    .A2(_08572_),
    .ZN(_08575_)
  );
  INV_X1 _18484_ (
    .A(_08575_),
    .ZN(_08577_)
  );
  AND2_X1 _18485_ (
    .A1(_08574_),
    .A2(_08577_),
    .ZN(_08578_)
  );
  INV_X1 _18486_ (
    .A(_08578_),
    .ZN(_08579_)
  );
  AND2_X1 _18487_ (
    .A1(_08559_),
    .A2(_08578_),
    .ZN(_08580_)
  );
  INV_X1 _18488_ (
    .A(_08580_),
    .ZN(_08581_)
  );
  AND2_X1 _18489_ (
    .A1(_08558_),
    .A2(_08579_),
    .ZN(_08582_)
  );
  INV_X1 _18490_ (
    .A(_08582_),
    .ZN(_08583_)
  );
  AND2_X1 _18491_ (
    .A1(_08581_),
    .A2(_08583_),
    .ZN(_08584_)
  );
  INV_X1 _18492_ (
    .A(_08584_),
    .ZN(_08585_)
  );
  AND2_X1 _18493_ (
    .A1(_08282_),
    .A2(_08584_),
    .ZN(_08586_)
  );
  INV_X1 _18494_ (
    .A(_08586_),
    .ZN(_08588_)
  );
  AND2_X1 _18495_ (
    .A1(_08283_),
    .A2(_08585_),
    .ZN(_08589_)
  );
  INV_X1 _18496_ (
    .A(_08589_),
    .ZN(_08590_)
  );
  AND2_X1 _18497_ (
    .A1(_08588_),
    .A2(_08590_),
    .ZN(_08591_)
  );
  INV_X1 _18498_ (
    .A(_08591_),
    .ZN(_08592_)
  );
  AND2_X1 _18499_ (
    .A1(_08556_),
    .A2(_08591_),
    .ZN(_08593_)
  );
  INV_X1 _18500_ (
    .A(_08593_),
    .ZN(_08594_)
  );
  AND2_X1 _18501_ (
    .A1(_08557_),
    .A2(_08592_),
    .ZN(_08595_)
  );
  INV_X1 _18502_ (
    .A(_08595_),
    .ZN(_08596_)
  );
  AND2_X1 _18503_ (
    .A1(_08594_),
    .A2(_08596_),
    .ZN(_08597_)
  );
  INV_X1 _18504_ (
    .A(_08597_),
    .ZN(_08599_)
  );
  AND2_X1 _18505_ (
    .A1(_08515_),
    .A2(_08597_),
    .ZN(_08600_)
  );
  INV_X1 _18506_ (
    .A(_08600_),
    .ZN(_08601_)
  );
  AND2_X1 _18507_ (
    .A1(_08514_),
    .A2(_08599_),
    .ZN(_08602_)
  );
  INV_X1 _18508_ (
    .A(_08602_),
    .ZN(_08603_)
  );
  AND2_X1 _18509_ (
    .A1(_08601_),
    .A2(_08603_),
    .ZN(_08604_)
  );
  INV_X1 _18510_ (
    .A(_08604_),
    .ZN(_08605_)
  );
  AND2_X1 _18511_ (
    .A1(divisor[28]),
    .A2(remainder[2]),
    .ZN(_08606_)
  );
  INV_X1 _18512_ (
    .A(_08606_),
    .ZN(_08607_)
  );
  AND2_X1 _18513_ (
    .A1(divisor[30]),
    .A2(remainder[0]),
    .ZN(_08608_)
  );
  INV_X1 _18514_ (
    .A(_08608_),
    .ZN(_08610_)
  );
  AND2_X1 _18515_ (
    .A1(divisor[30]),
    .A2(remainder[1]),
    .ZN(_08611_)
  );
  INV_X1 _18516_ (
    .A(_08611_),
    .ZN(_08612_)
  );
  AND2_X1 _18517_ (
    .A1(_08304_),
    .A2(_08611_),
    .ZN(_08613_)
  );
  INV_X1 _18518_ (
    .A(_08613_),
    .ZN(_08614_)
  );
  AND2_X1 _18519_ (
    .A1(_08309_),
    .A2(_08610_),
    .ZN(_08615_)
  );
  INV_X1 _18520_ (
    .A(_08615_),
    .ZN(_08616_)
  );
  AND2_X1 _18521_ (
    .A1(_08614_),
    .A2(_08616_),
    .ZN(_08617_)
  );
  INV_X1 _18522_ (
    .A(_08617_),
    .ZN(_08618_)
  );
  AND2_X1 _18523_ (
    .A1(_08606_),
    .A2(_08617_),
    .ZN(_08619_)
  );
  INV_X1 _18524_ (
    .A(_08619_),
    .ZN(_08621_)
  );
  AND2_X1 _18525_ (
    .A1(_08607_),
    .A2(_08618_),
    .ZN(_08622_)
  );
  INV_X1 _18526_ (
    .A(_08622_),
    .ZN(_08623_)
  );
  AND2_X1 _18527_ (
    .A1(_08621_),
    .A2(_08623_),
    .ZN(_08624_)
  );
  INV_X1 _18528_ (
    .A(_08624_),
    .ZN(_08625_)
  );
  AND2_X1 _18529_ (
    .A1(_03249_),
    .A2(_08316_),
    .ZN(_08626_)
  );
  INV_X1 _18530_ (
    .A(_08626_),
    .ZN(_08627_)
  );
  AND2_X1 _18531_ (
    .A1(_08625_),
    .A2(_08627_),
    .ZN(_08628_)
  );
  INV_X1 _18532_ (
    .A(_08628_),
    .ZN(_08629_)
  );
  AND2_X1 _18533_ (
    .A1(_08624_),
    .A2(_08626_),
    .ZN(_08630_)
  );
  INV_X1 _18534_ (
    .A(_08630_),
    .ZN(_08632_)
  );
  AND2_X1 _18535_ (
    .A1(_08624_),
    .A2(_08627_),
    .ZN(_08633_)
  );
  INV_X1 _18536_ (
    .A(_08633_),
    .ZN(_08634_)
  );
  AND2_X1 _18537_ (
    .A1(_08625_),
    .A2(_08626_),
    .ZN(_08635_)
  );
  INV_X1 _18538_ (
    .A(_08635_),
    .ZN(_08636_)
  );
  AND2_X1 _18539_ (
    .A1(_08629_),
    .A2(_08632_),
    .ZN(_08637_)
  );
  AND2_X1 _18540_ (
    .A1(_08634_),
    .A2(_08636_),
    .ZN(_08638_)
  );
  AND2_X1 _18541_ (
    .A1(_08604_),
    .A2(_08637_),
    .ZN(_08639_)
  );
  INV_X1 _18542_ (
    .A(_08639_),
    .ZN(_08640_)
  );
  AND2_X1 _18543_ (
    .A1(_08605_),
    .A2(_08638_),
    .ZN(_08641_)
  );
  INV_X1 _18544_ (
    .A(_08641_),
    .ZN(_08643_)
  );
  AND2_X1 _18545_ (
    .A1(_08640_),
    .A2(_08643_),
    .ZN(_08644_)
  );
  INV_X1 _18546_ (
    .A(_08644_),
    .ZN(_08645_)
  );
  AND2_X1 _18547_ (
    .A1(_08513_),
    .A2(_08644_),
    .ZN(_08646_)
  );
  INV_X1 _18548_ (
    .A(_08646_),
    .ZN(_08647_)
  );
  AND2_X1 _18549_ (
    .A1(_08512_),
    .A2(_08645_),
    .ZN(_08648_)
  );
  INV_X1 _18550_ (
    .A(_08648_),
    .ZN(_08649_)
  );
  AND2_X1 _18551_ (
    .A1(_08647_),
    .A2(_08649_),
    .ZN(_08650_)
  );
  INV_X1 _18552_ (
    .A(_08650_),
    .ZN(_08651_)
  );
  AND2_X1 _18553_ (
    .A1(_08380_),
    .A2(_08386_),
    .ZN(_08652_)
  );
  INV_X1 _18554_ (
    .A(_08652_),
    .ZN(_08654_)
  );
  AND2_X1 _18555_ (
    .A1(_08366_),
    .A2(_08373_),
    .ZN(_08655_)
  );
  INV_X1 _18556_ (
    .A(_08655_),
    .ZN(_08656_)
  );
  AND2_X1 _18557_ (
    .A1(_08353_),
    .A2(_08360_),
    .ZN(_08657_)
  );
  INV_X1 _18558_ (
    .A(_08657_),
    .ZN(_08658_)
  );
  AND2_X1 _18559_ (
    .A1(_08273_),
    .A2(_08285_),
    .ZN(_08659_)
  );
  INV_X1 _18560_ (
    .A(_08659_),
    .ZN(_08660_)
  );
  AND2_X1 _18561_ (
    .A1(_07969_),
    .A2(_08281_),
    .ZN(_08661_)
  );
  INV_X1 _18562_ (
    .A(_08661_),
    .ZN(_08662_)
  );
  AND2_X1 _18563_ (
    .A1(_07319_),
    .A2(_08662_),
    .ZN(_08663_)
  );
  INV_X1 _18564_ (
    .A(_08663_),
    .ZN(_08665_)
  );
  AND2_X1 _18565_ (
    .A1(_07320_),
    .A2(_08661_),
    .ZN(_08666_)
  );
  INV_X1 _18566_ (
    .A(_08666_),
    .ZN(_08667_)
  );
  AND2_X1 _18567_ (
    .A1(_08665_),
    .A2(_08667_),
    .ZN(_08668_)
  );
  INV_X1 _18568_ (
    .A(_08668_),
    .ZN(_08669_)
  );
  AND2_X1 _18569_ (
    .A1(_07620_),
    .A2(_08668_),
    .ZN(_08670_)
  );
  INV_X1 _18570_ (
    .A(_08670_),
    .ZN(_08671_)
  );
  AND2_X1 _18571_ (
    .A1(_07619_),
    .A2(_08669_),
    .ZN(_08672_)
  );
  INV_X1 _18572_ (
    .A(_08672_),
    .ZN(_08673_)
  );
  AND2_X1 _18573_ (
    .A1(_08671_),
    .A2(_08673_),
    .ZN(_08674_)
  );
  INV_X1 _18574_ (
    .A(_08674_),
    .ZN(_08676_)
  );
  AND2_X1 _18575_ (
    .A1(_08660_),
    .A2(_08674_),
    .ZN(_08677_)
  );
  INV_X1 _18576_ (
    .A(_08677_),
    .ZN(_08678_)
  );
  AND2_X1 _18577_ (
    .A1(_08659_),
    .A2(_08676_),
    .ZN(_08679_)
  );
  INV_X1 _18578_ (
    .A(_08679_),
    .ZN(_08680_)
  );
  AND2_X1 _18579_ (
    .A1(_08678_),
    .A2(_08680_),
    .ZN(_08681_)
  );
  INV_X1 _18580_ (
    .A(_08681_),
    .ZN(_08682_)
  );
  AND2_X1 _18581_ (
    .A1(_08658_),
    .A2(_08681_),
    .ZN(_08683_)
  );
  INV_X1 _18582_ (
    .A(_08683_),
    .ZN(_08684_)
  );
  AND2_X1 _18583_ (
    .A1(_08657_),
    .A2(_08682_),
    .ZN(_08685_)
  );
  INV_X1 _18584_ (
    .A(_08685_),
    .ZN(_08687_)
  );
  AND2_X1 _18585_ (
    .A1(_08684_),
    .A2(_08687_),
    .ZN(_08688_)
  );
  INV_X1 _18586_ (
    .A(_08688_),
    .ZN(_08689_)
  );
  AND2_X1 _18587_ (
    .A1(_08656_),
    .A2(_08688_),
    .ZN(_08690_)
  );
  INV_X1 _18588_ (
    .A(_08690_),
    .ZN(_08691_)
  );
  AND2_X1 _18589_ (
    .A1(_08655_),
    .A2(_08689_),
    .ZN(_08692_)
  );
  INV_X1 _18590_ (
    .A(_08692_),
    .ZN(_08693_)
  );
  AND2_X1 _18591_ (
    .A1(_08691_),
    .A2(_08693_),
    .ZN(_08694_)
  );
  INV_X1 _18592_ (
    .A(_08694_),
    .ZN(_08695_)
  );
  AND2_X1 _18593_ (
    .A1(_07082_),
    .A2(_08694_),
    .ZN(_08696_)
  );
  INV_X1 _18594_ (
    .A(_08696_),
    .ZN(_08698_)
  );
  AND2_X1 _18595_ (
    .A1(_07083_),
    .A2(_08695_),
    .ZN(_08699_)
  );
  INV_X1 _18596_ (
    .A(_08699_),
    .ZN(_08700_)
  );
  AND2_X1 _18597_ (
    .A1(_08698_),
    .A2(_08700_),
    .ZN(_08701_)
  );
  INV_X1 _18598_ (
    .A(_08701_),
    .ZN(_08702_)
  );
  AND2_X1 _18599_ (
    .A1(_08297_),
    .A2(_08701_),
    .ZN(_08703_)
  );
  INV_X1 _18600_ (
    .A(_08703_),
    .ZN(_08704_)
  );
  AND2_X1 _18601_ (
    .A1(_08298_),
    .A2(_08702_),
    .ZN(_08705_)
  );
  INV_X1 _18602_ (
    .A(_08705_),
    .ZN(_08706_)
  );
  AND2_X1 _18603_ (
    .A1(_08704_),
    .A2(_08706_),
    .ZN(_08707_)
  );
  INV_X1 _18604_ (
    .A(_08707_),
    .ZN(_08709_)
  );
  AND2_X1 _18605_ (
    .A1(_08654_),
    .A2(_08707_),
    .ZN(_08710_)
  );
  INV_X1 _18606_ (
    .A(_08710_),
    .ZN(_08711_)
  );
  AND2_X1 _18607_ (
    .A1(_08652_),
    .A2(_08709_),
    .ZN(_08712_)
  );
  INV_X1 _18608_ (
    .A(_08712_),
    .ZN(_08713_)
  );
  AND2_X1 _18609_ (
    .A1(_08711_),
    .A2(_08713_),
    .ZN(_08714_)
  );
  INV_X1 _18610_ (
    .A(_08714_),
    .ZN(_08715_)
  );
  AND2_X1 _18611_ (
    .A1(_08650_),
    .A2(_08714_),
    .ZN(_08716_)
  );
  INV_X1 _18612_ (
    .A(_08716_),
    .ZN(_08717_)
  );
  AND2_X1 _18613_ (
    .A1(_08651_),
    .A2(_08715_),
    .ZN(_08718_)
  );
  INV_X1 _18614_ (
    .A(_08718_),
    .ZN(_08720_)
  );
  AND2_X1 _18615_ (
    .A1(_08717_),
    .A2(_08720_),
    .ZN(_08721_)
  );
  INV_X1 _18616_ (
    .A(_08721_),
    .ZN(_08722_)
  );
  AND2_X1 _18617_ (
    .A1(_08508_),
    .A2(_08721_),
    .ZN(_08723_)
  );
  INV_X1 _18618_ (
    .A(_08723_),
    .ZN(_08724_)
  );
  AND2_X1 _18619_ (
    .A1(_08507_),
    .A2(_08722_),
    .ZN(_08725_)
  );
  INV_X1 _18620_ (
    .A(_08725_),
    .ZN(_08726_)
  );
  AND2_X1 _18621_ (
    .A1(_08724_),
    .A2(_08726_),
    .ZN(_08727_)
  );
  INV_X1 _18622_ (
    .A(_08727_),
    .ZN(_08728_)
  );
  AND2_X1 _18623_ (
    .A1(_08393_),
    .A2(_08399_),
    .ZN(_08729_)
  );
  INV_X1 _18624_ (
    .A(_08729_),
    .ZN(_08731_)
  );
  AND2_X1 _18625_ (
    .A1(_07804_),
    .A2(_08731_),
    .ZN(_08732_)
  );
  INV_X1 _18626_ (
    .A(_08732_),
    .ZN(_08733_)
  );
  AND2_X1 _18627_ (
    .A1(_07805_),
    .A2(_08729_),
    .ZN(_08734_)
  );
  INV_X1 _18628_ (
    .A(_08734_),
    .ZN(_08735_)
  );
  AND2_X1 _18629_ (
    .A1(_08733_),
    .A2(_08735_),
    .ZN(_08736_)
  );
  INV_X1 _18630_ (
    .A(_08736_),
    .ZN(_08737_)
  );
  AND2_X1 _18631_ (
    .A1(_08107_),
    .A2(_08736_),
    .ZN(_08738_)
  );
  INV_X1 _18632_ (
    .A(_08738_),
    .ZN(_08739_)
  );
  AND2_X1 _18633_ (
    .A1(_08106_),
    .A2(_08737_),
    .ZN(_08740_)
  );
  INV_X1 _18634_ (
    .A(_08740_),
    .ZN(_08742_)
  );
  AND2_X1 _18635_ (
    .A1(_08739_),
    .A2(_08742_),
    .ZN(_08743_)
  );
  INV_X1 _18636_ (
    .A(_08743_),
    .ZN(_08744_)
  );
  AND2_X1 _18637_ (
    .A1(_08727_),
    .A2(_08743_),
    .ZN(_08745_)
  );
  INV_X1 _18638_ (
    .A(_08745_),
    .ZN(_08746_)
  );
  AND2_X1 _18639_ (
    .A1(_08728_),
    .A2(_08744_),
    .ZN(_08747_)
  );
  INV_X1 _18640_ (
    .A(_08747_),
    .ZN(_08748_)
  );
  AND2_X1 _18641_ (
    .A1(_08746_),
    .A2(_08748_),
    .ZN(_08749_)
  );
  INV_X1 _18642_ (
    .A(_08749_),
    .ZN(_08750_)
  );
  AND2_X1 _18643_ (
    .A1(_08506_),
    .A2(_08749_),
    .ZN(_08751_)
  );
  INV_X1 _18644_ (
    .A(_08751_),
    .ZN(_08753_)
  );
  AND2_X1 _18645_ (
    .A1(_08505_),
    .A2(_08750_),
    .ZN(_08754_)
  );
  INV_X1 _18646_ (
    .A(_08754_),
    .ZN(_08755_)
  );
  AND2_X1 _18647_ (
    .A1(_08753_),
    .A2(_08755_),
    .ZN(_08756_)
  );
  INV_X1 _18648_ (
    .A(_08756_),
    .ZN(_08757_)
  );
  AND2_X1 _18649_ (
    .A1(_08504_),
    .A2(_08756_),
    .ZN(_08758_)
  );
  INV_X1 _18650_ (
    .A(_08758_),
    .ZN(_08759_)
  );
  AND2_X1 _18651_ (
    .A1(_08503_),
    .A2(_08757_),
    .ZN(_08760_)
  );
  INV_X1 _18652_ (
    .A(_08760_),
    .ZN(_08761_)
  );
  AND2_X1 _18653_ (
    .A1(_08759_),
    .A2(_08761_),
    .ZN(_08762_)
  );
  INV_X1 _18654_ (
    .A(_08762_),
    .ZN(_08764_)
  );
  AND2_X1 _18655_ (
    .A1(_08502_),
    .A2(_08762_),
    .ZN(_08765_)
  );
  INV_X1 _18656_ (
    .A(_08765_),
    .ZN(_08766_)
  );
  AND2_X1 _18657_ (
    .A1(_08501_),
    .A2(_08764_),
    .ZN(_08767_)
  );
  INV_X1 _18658_ (
    .A(_08767_),
    .ZN(_08768_)
  );
  AND2_X1 _18659_ (
    .A1(_08766_),
    .A2(_08768_),
    .ZN(_08769_)
  );
  INV_X1 _18660_ (
    .A(_08769_),
    .ZN(_08770_)
  );
  AND2_X1 _18661_ (
    .A1(_08453_),
    .A2(_08769_),
    .ZN(_08771_)
  );
  INV_X1 _18662_ (
    .A(_08771_),
    .ZN(_08772_)
  );
  AND2_X1 _18663_ (
    .A1(_08454_),
    .A2(_08770_),
    .ZN(_08773_)
  );
  INV_X1 _18664_ (
    .A(_08773_),
    .ZN(_08775_)
  );
  AND2_X1 _18665_ (
    .A1(_08772_),
    .A2(_08775_),
    .ZN(_08776_)
  );
  INV_X1 _18666_ (
    .A(_08776_),
    .ZN(_08777_)
  );
  AND2_X1 _18667_ (
    .A1(_08161_),
    .A2(_08464_),
    .ZN(_08778_)
  );
  INV_X1 _18668_ (
    .A(_08778_),
    .ZN(_08779_)
  );
  AND2_X1 _18669_ (
    .A1(_08150_),
    .A2(_08463_),
    .ZN(_08780_)
  );
  INV_X1 _18670_ (
    .A(_08780_),
    .ZN(_08781_)
  );
  AND2_X1 _18671_ (
    .A1(_08461_),
    .A2(_08781_),
    .ZN(_08782_)
  );
  AND2_X1 _18672_ (
    .A1(_08779_),
    .A2(_08782_),
    .ZN(_08783_)
  );
  INV_X1 _18673_ (
    .A(_08783_),
    .ZN(_08784_)
  );
  AND2_X1 _18674_ (
    .A1(_08776_),
    .A2(_08784_),
    .ZN(_08786_)
  );
  INV_X1 _18675_ (
    .A(_08786_),
    .ZN(_08787_)
  );
  AND2_X1 _18676_ (
    .A1(_08777_),
    .A2(_08783_),
    .ZN(_08788_)
  );
  INV_X1 _18677_ (
    .A(_08788_),
    .ZN(_08789_)
  );
  AND2_X1 _18678_ (
    .A1(_08787_),
    .A2(_08789_),
    .ZN(_08790_)
  );
  INV_X1 _18679_ (
    .A(_08790_),
    .ZN(_08791_)
  );
  AND2_X1 _18680_ (
    .A1(remainder[63]),
    .A2(_08790_),
    .ZN(_08792_)
  );
  INV_X1 _18681_ (
    .A(_08792_),
    .ZN(_08793_)
  );
  AND2_X1 _18682_ (
    .A1(_04426_),
    .A2(_08791_),
    .ZN(_08794_)
  );
  INV_X1 _18683_ (
    .A(_08794_),
    .ZN(_08795_)
  );
  AND2_X1 _18684_ (
    .A1(_08793_),
    .A2(_08795_),
    .ZN(_08797_)
  );
  INV_X1 _18685_ (
    .A(_08797_),
    .ZN(_08798_)
  );
  AND2_X1 _18686_ (
    .A1(_08199_),
    .A2(_08474_),
    .ZN(_08799_)
  );
  INV_X1 _18687_ (
    .A(_08799_),
    .ZN(_08800_)
  );
  AND2_X1 _18688_ (
    .A1(_08200_),
    .A2(_08476_),
    .ZN(_08801_)
  );
  INV_X1 _18689_ (
    .A(_08801_),
    .ZN(_08802_)
  );
  AND2_X1 _18690_ (
    .A1(_08476_),
    .A2(_08800_),
    .ZN(_08803_)
  );
  AND2_X1 _18691_ (
    .A1(_08474_),
    .A2(_08802_),
    .ZN(_08804_)
  );
  AND2_X1 _18692_ (
    .A1(_08797_),
    .A2(_08803_),
    .ZN(_08805_)
  );
  INV_X1 _18693_ (
    .A(_08805_),
    .ZN(_08806_)
  );
  AND2_X1 _18694_ (
    .A1(_08798_),
    .A2(_08804_),
    .ZN(_08808_)
  );
  INV_X1 _18695_ (
    .A(_08808_),
    .ZN(_08809_)
  );
  AND2_X1 _18696_ (
    .A1(_02082_),
    .A2(_08806_),
    .ZN(_08810_)
  );
  AND2_X1 _18697_ (
    .A1(_08809_),
    .A2(_08810_),
    .ZN(_08811_)
  );
  INV_X1 _18698_ (
    .A(_08811_),
    .ZN(_08812_)
  );
  AND2_X1 _18699_ (
    .A1(remainder[55]),
    .A2(_02077_),
    .ZN(_08813_)
  );
  INV_X1 _18700_ (
    .A(_08813_),
    .ZN(_08814_)
  );
  AND2_X1 _18701_ (
    .A1(_04525_),
    .A2(_10451_),
    .ZN(_08815_)
  );
  INV_X1 _18702_ (
    .A(_08815_),
    .ZN(_08816_)
  );
  AND2_X1 _18703_ (
    .A1(_10462_),
    .A2(_01937_),
    .ZN(_08817_)
  );
  INV_X1 _18704_ (
    .A(_08817_),
    .ZN(_08819_)
  );
  AND2_X1 _18705_ (
    .A1(_05983_),
    .A2(_08819_),
    .ZN(_08820_)
  );
  AND2_X1 _18706_ (
    .A1(_08816_),
    .A2(_08820_),
    .ZN(_08821_)
  );
  INV_X1 _18707_ (
    .A(_08821_),
    .ZN(_08822_)
  );
  AND2_X1 _18708_ (
    .A1(_08814_),
    .A2(_08822_),
    .ZN(_08823_)
  );
  AND2_X1 _18709_ (
    .A1(_08812_),
    .A2(_08823_),
    .ZN(_08824_)
  );
  INV_X1 _18710_ (
    .A(_08824_),
    .ZN(_08825_)
  );
  AND2_X1 _18711_ (
    .A1(_06201_),
    .A2(_08825_),
    .ZN(_00076_)
  );
  AND2_X1 _18712_ (
    .A1(_08793_),
    .A2(_08806_),
    .ZN(_08826_)
  );
  INV_X1 _18713_ (
    .A(_08826_),
    .ZN(_08827_)
  );
  AND2_X1 _18714_ (
    .A1(_08772_),
    .A2(_08787_),
    .ZN(_08829_)
  );
  INV_X1 _18715_ (
    .A(_08829_),
    .ZN(_08830_)
  );
  AND2_X1 _18716_ (
    .A1(_08753_),
    .A2(_08759_),
    .ZN(_08831_)
  );
  INV_X1 _18717_ (
    .A(_08831_),
    .ZN(_08832_)
  );
  AND2_X1 _18718_ (
    .A1(_08733_),
    .A2(_08739_),
    .ZN(_08833_)
  );
  INV_X1 _18719_ (
    .A(_08833_),
    .ZN(_08834_)
  );
  AND2_X1 _18720_ (
    .A1(_08724_),
    .A2(_08746_),
    .ZN(_08835_)
  );
  INV_X1 _18721_ (
    .A(_08835_),
    .ZN(_08836_)
  );
  AND2_X1 _18722_ (
    .A1(_08647_),
    .A2(_08717_),
    .ZN(_08837_)
  );
  INV_X1 _18723_ (
    .A(_08837_),
    .ZN(_08838_)
  );
  AND2_X1 _18724_ (
    .A1(_03249_),
    .A2(_08625_),
    .ZN(_08840_)
  );
  INV_X1 _18725_ (
    .A(_08840_),
    .ZN(_08841_)
  );
  AND2_X1 _18726_ (
    .A1(_08315_),
    .A2(_08840_),
    .ZN(_08842_)
  );
  INV_X1 _18727_ (
    .A(_08842_),
    .ZN(_08843_)
  );
  AND2_X1 _18728_ (
    .A1(_08640_),
    .A2(_08843_),
    .ZN(_08844_)
  );
  INV_X1 _18729_ (
    .A(_08844_),
    .ZN(_08845_)
  );
  AND2_X1 _18730_ (
    .A1(_08552_),
    .A2(_08594_),
    .ZN(_08846_)
  );
  INV_X1 _18731_ (
    .A(_08846_),
    .ZN(_08847_)
  );
  AND2_X1 _18732_ (
    .A1(_08539_),
    .A2(_08546_),
    .ZN(_08848_)
  );
  INV_X1 _18733_ (
    .A(_08848_),
    .ZN(_08849_)
  );
  AND2_X1 _18734_ (
    .A1(_08526_),
    .A2(_08533_),
    .ZN(_08851_)
  );
  INV_X1 _18735_ (
    .A(_08851_),
    .ZN(_08852_)
  );
  AND2_X1 _18736_ (
    .A1(_08614_),
    .A2(_08621_),
    .ZN(_08853_)
  );
  INV_X1 _18737_ (
    .A(_08853_),
    .ZN(_08854_)
  );
  AND2_X1 _18738_ (
    .A1(divisor[25]),
    .A2(remainder[6]),
    .ZN(_08855_)
  );
  INV_X1 _18739_ (
    .A(_08855_),
    .ZN(_08856_)
  );
  AND2_X1 _18740_ (
    .A1(divisor[26]),
    .A2(remainder[5]),
    .ZN(_08857_)
  );
  INV_X1 _18741_ (
    .A(_08857_),
    .ZN(_08858_)
  );
  AND2_X1 _18742_ (
    .A1(divisor[27]),
    .A2(remainder[5]),
    .ZN(_08859_)
  );
  INV_X1 _18743_ (
    .A(_08859_),
    .ZN(_08860_)
  );
  AND2_X1 _18744_ (
    .A1(_08523_),
    .A2(_08857_),
    .ZN(_08862_)
  );
  INV_X1 _18745_ (
    .A(_08862_),
    .ZN(_08863_)
  );
  AND2_X1 _18746_ (
    .A1(_08524_),
    .A2(_08858_),
    .ZN(_08864_)
  );
  INV_X1 _18747_ (
    .A(_08864_),
    .ZN(_08865_)
  );
  AND2_X1 _18748_ (
    .A1(_08863_),
    .A2(_08865_),
    .ZN(_08866_)
  );
  INV_X1 _18749_ (
    .A(_08866_),
    .ZN(_08867_)
  );
  AND2_X1 _18750_ (
    .A1(_08855_),
    .A2(_08866_),
    .ZN(_08868_)
  );
  INV_X1 _18751_ (
    .A(_08868_),
    .ZN(_08869_)
  );
  AND2_X1 _18752_ (
    .A1(_08856_),
    .A2(_08867_),
    .ZN(_08870_)
  );
  INV_X1 _18753_ (
    .A(_08870_),
    .ZN(_08871_)
  );
  AND2_X1 _18754_ (
    .A1(_08869_),
    .A2(_08871_),
    .ZN(_08873_)
  );
  INV_X1 _18755_ (
    .A(_08873_),
    .ZN(_08874_)
  );
  AND2_X1 _18756_ (
    .A1(_08854_),
    .A2(_08873_),
    .ZN(_08875_)
  );
  INV_X1 _18757_ (
    .A(_08875_),
    .ZN(_08876_)
  );
  AND2_X1 _18758_ (
    .A1(_08853_),
    .A2(_08874_),
    .ZN(_08877_)
  );
  INV_X1 _18759_ (
    .A(_08877_),
    .ZN(_08878_)
  );
  AND2_X1 _18760_ (
    .A1(_08876_),
    .A2(_08878_),
    .ZN(_08879_)
  );
  INV_X1 _18761_ (
    .A(_08879_),
    .ZN(_08880_)
  );
  AND2_X1 _18762_ (
    .A1(_08852_),
    .A2(_08879_),
    .ZN(_08881_)
  );
  INV_X1 _18763_ (
    .A(_08881_),
    .ZN(_08882_)
  );
  AND2_X1 _18764_ (
    .A1(_08851_),
    .A2(_08880_),
    .ZN(_08884_)
  );
  INV_X1 _18765_ (
    .A(_08884_),
    .ZN(_08885_)
  );
  AND2_X1 _18766_ (
    .A1(_08882_),
    .A2(_08885_),
    .ZN(_08886_)
  );
  INV_X1 _18767_ (
    .A(_08886_),
    .ZN(_08887_)
  );
  AND2_X1 _18768_ (
    .A1(_08849_),
    .A2(_08886_),
    .ZN(_08888_)
  );
  INV_X1 _18769_ (
    .A(_08888_),
    .ZN(_08889_)
  );
  AND2_X1 _18770_ (
    .A1(_08848_),
    .A2(_08887_),
    .ZN(_08890_)
  );
  INV_X1 _18771_ (
    .A(_08890_),
    .ZN(_08891_)
  );
  AND2_X1 _18772_ (
    .A1(_08889_),
    .A2(_08891_),
    .ZN(_08892_)
  );
  INV_X1 _18773_ (
    .A(_08892_),
    .ZN(_08893_)
  );
  AND2_X1 _18774_ (
    .A1(_08568_),
    .A2(_08574_),
    .ZN(_08895_)
  );
  INV_X1 _18775_ (
    .A(_08895_),
    .ZN(_08896_)
  );
  AND2_X1 _18776_ (
    .A1(remainder[32]),
    .A2(divisor[24]),
    .ZN(_08897_)
  );
  INV_X1 _18777_ (
    .A(_08897_),
    .ZN(_08898_)
  );
  AND2_X1 _18778_ (
    .A1(remainder[32]),
    .A2(divisor[23]),
    .ZN(_08899_)
  );
  INV_X1 _18779_ (
    .A(_08899_),
    .ZN(_08900_)
  );
  AND2_X1 _18780_ (
    .A1(_08564_),
    .A2(_08899_),
    .ZN(_08901_)
  );
  INV_X1 _18781_ (
    .A(_08901_),
    .ZN(_08902_)
  );
  AND2_X1 _18782_ (
    .A1(_08566_),
    .A2(_08900_),
    .ZN(_08903_)
  );
  INV_X1 _18783_ (
    .A(_08903_),
    .ZN(_08904_)
  );
  AND2_X1 _18784_ (
    .A1(_08902_),
    .A2(_08904_),
    .ZN(_08906_)
  );
  INV_X1 _18785_ (
    .A(_08906_),
    .ZN(_08907_)
  );
  AND2_X1 _18786_ (
    .A1(_08560_),
    .A2(_08906_),
    .ZN(_08908_)
  );
  INV_X1 _18787_ (
    .A(_08908_),
    .ZN(_08909_)
  );
  AND2_X1 _18788_ (
    .A1(_08561_),
    .A2(_08907_),
    .ZN(_08910_)
  );
  INV_X1 _18789_ (
    .A(_08910_),
    .ZN(_08911_)
  );
  AND2_X1 _18790_ (
    .A1(_08909_),
    .A2(_08911_),
    .ZN(_08912_)
  );
  INV_X1 _18791_ (
    .A(_08912_),
    .ZN(_08913_)
  );
  AND2_X1 _18792_ (
    .A1(_08896_),
    .A2(_08912_),
    .ZN(_08914_)
  );
  INV_X1 _18793_ (
    .A(_08914_),
    .ZN(_08915_)
  );
  AND2_X1 _18794_ (
    .A1(_08895_),
    .A2(_08913_),
    .ZN(_08917_)
  );
  INV_X1 _18795_ (
    .A(_08917_),
    .ZN(_08918_)
  );
  AND2_X1 _18796_ (
    .A1(_08915_),
    .A2(_08918_),
    .ZN(_08919_)
  );
  INV_X1 _18797_ (
    .A(_08919_),
    .ZN(_08920_)
  );
  AND2_X1 _18798_ (
    .A1(_08282_),
    .A2(_08919_),
    .ZN(_08921_)
  );
  INV_X1 _18799_ (
    .A(_08921_),
    .ZN(_08922_)
  );
  AND2_X1 _18800_ (
    .A1(_08283_),
    .A2(_08920_),
    .ZN(_08923_)
  );
  INV_X1 _18801_ (
    .A(_08923_),
    .ZN(_08924_)
  );
  AND2_X1 _18802_ (
    .A1(_08922_),
    .A2(_08924_),
    .ZN(_08925_)
  );
  INV_X1 _18803_ (
    .A(_08925_),
    .ZN(_08926_)
  );
  AND2_X1 _18804_ (
    .A1(_08892_),
    .A2(_08925_),
    .ZN(_08928_)
  );
  INV_X1 _18805_ (
    .A(_08928_),
    .ZN(_08929_)
  );
  AND2_X1 _18806_ (
    .A1(_08893_),
    .A2(_08926_),
    .ZN(_08930_)
  );
  INV_X1 _18807_ (
    .A(_08930_),
    .ZN(_08931_)
  );
  AND2_X1 _18808_ (
    .A1(_08929_),
    .A2(_08931_),
    .ZN(_08932_)
  );
  INV_X1 _18809_ (
    .A(_08932_),
    .ZN(_08933_)
  );
  AND2_X1 _18810_ (
    .A1(_08847_),
    .A2(_08932_),
    .ZN(_08934_)
  );
  INV_X1 _18811_ (
    .A(_08934_),
    .ZN(_08935_)
  );
  AND2_X1 _18812_ (
    .A1(_08846_),
    .A2(_08933_),
    .ZN(_08936_)
  );
  INV_X1 _18813_ (
    .A(_08936_),
    .ZN(_08937_)
  );
  AND2_X1 _18814_ (
    .A1(_08935_),
    .A2(_08937_),
    .ZN(_08939_)
  );
  INV_X1 _18815_ (
    .A(_08939_),
    .ZN(_08940_)
  );
  AND2_X1 _18816_ (
    .A1(divisor[31]),
    .A2(remainder[0]),
    .ZN(_08941_)
  );
  INV_X1 _18817_ (
    .A(_08941_),
    .ZN(_08942_)
  );
  AND2_X1 _18818_ (
    .A1(divisor[28]),
    .A2(remainder[3]),
    .ZN(_08943_)
  );
  INV_X1 _18819_ (
    .A(_08943_),
    .ZN(_08944_)
  );
  AND2_X1 _18820_ (
    .A1(divisor[29]),
    .A2(remainder[2]),
    .ZN(_08945_)
  );
  INV_X1 _18821_ (
    .A(_08945_),
    .ZN(_08946_)
  );
  AND2_X1 _18822_ (
    .A1(divisor[30]),
    .A2(remainder[2]),
    .ZN(_08947_)
  );
  INV_X1 _18823_ (
    .A(_08947_),
    .ZN(_08948_)
  );
  AND2_X1 _18824_ (
    .A1(_08308_),
    .A2(_08947_),
    .ZN(_08950_)
  );
  INV_X1 _18825_ (
    .A(_08950_),
    .ZN(_08951_)
  );
  AND2_X1 _18826_ (
    .A1(_08612_),
    .A2(_08946_),
    .ZN(_08952_)
  );
  INV_X1 _18827_ (
    .A(_08952_),
    .ZN(_08953_)
  );
  AND2_X1 _18828_ (
    .A1(_08951_),
    .A2(_08953_),
    .ZN(_08954_)
  );
  INV_X1 _18829_ (
    .A(_08954_),
    .ZN(_08955_)
  );
  AND2_X1 _18830_ (
    .A1(_08943_),
    .A2(_08954_),
    .ZN(_08956_)
  );
  INV_X1 _18831_ (
    .A(_08956_),
    .ZN(_08957_)
  );
  AND2_X1 _18832_ (
    .A1(_08944_),
    .A2(_08955_),
    .ZN(_08958_)
  );
  INV_X1 _18833_ (
    .A(_08958_),
    .ZN(_08959_)
  );
  AND2_X1 _18834_ (
    .A1(_08957_),
    .A2(_08959_),
    .ZN(_08961_)
  );
  INV_X1 _18835_ (
    .A(_08961_),
    .ZN(_08962_)
  );
  AND2_X1 _18836_ (
    .A1(_08941_),
    .A2(_08961_),
    .ZN(_08963_)
  );
  INV_X1 _18837_ (
    .A(_08963_),
    .ZN(_08964_)
  );
  AND2_X1 _18838_ (
    .A1(_08942_),
    .A2(_08962_),
    .ZN(_08965_)
  );
  INV_X1 _18839_ (
    .A(_08965_),
    .ZN(_08966_)
  );
  AND2_X1 _18840_ (
    .A1(_08964_),
    .A2(_08966_),
    .ZN(_08967_)
  );
  INV_X1 _18841_ (
    .A(_08967_),
    .ZN(_08968_)
  );
  AND2_X1 _18842_ (
    .A1(_08841_),
    .A2(_08968_),
    .ZN(_08969_)
  );
  INV_X1 _18843_ (
    .A(_08969_),
    .ZN(_08970_)
  );
  AND2_X1 _18844_ (
    .A1(_08840_),
    .A2(_08967_),
    .ZN(_08972_)
  );
  INV_X1 _18845_ (
    .A(_08972_),
    .ZN(_08973_)
  );
  AND2_X1 _18846_ (
    .A1(_08840_),
    .A2(_08968_),
    .ZN(_08974_)
  );
  INV_X1 _18847_ (
    .A(_08974_),
    .ZN(_08975_)
  );
  AND2_X1 _18848_ (
    .A1(_08841_),
    .A2(_08967_),
    .ZN(_08976_)
  );
  INV_X1 _18849_ (
    .A(_08976_),
    .ZN(_08977_)
  );
  AND2_X1 _18850_ (
    .A1(_08970_),
    .A2(_08973_),
    .ZN(_08978_)
  );
  AND2_X1 _18851_ (
    .A1(_08975_),
    .A2(_08977_),
    .ZN(_08979_)
  );
  AND2_X1 _18852_ (
    .A1(_08939_),
    .A2(_08978_),
    .ZN(_08980_)
  );
  INV_X1 _18853_ (
    .A(_08980_),
    .ZN(_08981_)
  );
  AND2_X1 _18854_ (
    .A1(_08940_),
    .A2(_08979_),
    .ZN(_08983_)
  );
  INV_X1 _18855_ (
    .A(_08983_),
    .ZN(_08984_)
  );
  AND2_X1 _18856_ (
    .A1(_08981_),
    .A2(_08984_),
    .ZN(_08985_)
  );
  INV_X1 _18857_ (
    .A(_08985_),
    .ZN(_08986_)
  );
  AND2_X1 _18858_ (
    .A1(_08845_),
    .A2(_08985_),
    .ZN(_08987_)
  );
  INV_X1 _18859_ (
    .A(_08987_),
    .ZN(_08988_)
  );
  AND2_X1 _18860_ (
    .A1(_08844_),
    .A2(_08986_),
    .ZN(_08989_)
  );
  INV_X1 _18861_ (
    .A(_08989_),
    .ZN(_08990_)
  );
  AND2_X1 _18862_ (
    .A1(_08988_),
    .A2(_08990_),
    .ZN(_08991_)
  );
  INV_X1 _18863_ (
    .A(_08991_),
    .ZN(_08992_)
  );
  AND2_X1 _18864_ (
    .A1(_08691_),
    .A2(_08698_),
    .ZN(_08994_)
  );
  INV_X1 _18865_ (
    .A(_08994_),
    .ZN(_08995_)
  );
  AND2_X1 _18866_ (
    .A1(_08678_),
    .A2(_08684_),
    .ZN(_08996_)
  );
  INV_X1 _18867_ (
    .A(_08996_),
    .ZN(_08997_)
  );
  AND2_X1 _18868_ (
    .A1(_08665_),
    .A2(_08671_),
    .ZN(_08998_)
  );
  INV_X1 _18869_ (
    .A(_08998_),
    .ZN(_08999_)
  );
  AND2_X1 _18870_ (
    .A1(_08581_),
    .A2(_08588_),
    .ZN(_09000_)
  );
  INV_X1 _18871_ (
    .A(_09000_),
    .ZN(_09001_)
  );
  AND2_X1 _18872_ (
    .A1(_08674_),
    .A2(_09001_),
    .ZN(_09002_)
  );
  INV_X1 _18873_ (
    .A(_09002_),
    .ZN(_09003_)
  );
  AND2_X1 _18874_ (
    .A1(_08676_),
    .A2(_09000_),
    .ZN(_09005_)
  );
  INV_X1 _18875_ (
    .A(_09005_),
    .ZN(_09006_)
  );
  AND2_X1 _18876_ (
    .A1(_09003_),
    .A2(_09006_),
    .ZN(_09007_)
  );
  INV_X1 _18877_ (
    .A(_09007_),
    .ZN(_09008_)
  );
  AND2_X1 _18878_ (
    .A1(_08999_),
    .A2(_09007_),
    .ZN(_09009_)
  );
  INV_X1 _18879_ (
    .A(_09009_),
    .ZN(_09010_)
  );
  AND2_X1 _18880_ (
    .A1(_08998_),
    .A2(_09008_),
    .ZN(_09011_)
  );
  INV_X1 _18881_ (
    .A(_09011_),
    .ZN(_09012_)
  );
  AND2_X1 _18882_ (
    .A1(_09010_),
    .A2(_09012_),
    .ZN(_09013_)
  );
  INV_X1 _18883_ (
    .A(_09013_),
    .ZN(_09014_)
  );
  AND2_X1 _18884_ (
    .A1(_08997_),
    .A2(_09013_),
    .ZN(_09016_)
  );
  INV_X1 _18885_ (
    .A(_09016_),
    .ZN(_09017_)
  );
  AND2_X1 _18886_ (
    .A1(_08996_),
    .A2(_09014_),
    .ZN(_09018_)
  );
  INV_X1 _18887_ (
    .A(_09018_),
    .ZN(_09019_)
  );
  AND2_X1 _18888_ (
    .A1(_09017_),
    .A2(_09019_),
    .ZN(_09020_)
  );
  INV_X1 _18889_ (
    .A(_09020_),
    .ZN(_09021_)
  );
  AND2_X1 _18890_ (
    .A1(_07082_),
    .A2(_09020_),
    .ZN(_09022_)
  );
  INV_X1 _18891_ (
    .A(_09022_),
    .ZN(_09023_)
  );
  AND2_X1 _18892_ (
    .A1(_07083_),
    .A2(_09021_),
    .ZN(_09024_)
  );
  INV_X1 _18893_ (
    .A(_09024_),
    .ZN(_09025_)
  );
  AND2_X1 _18894_ (
    .A1(_09023_),
    .A2(_09025_),
    .ZN(_09027_)
  );
  INV_X1 _18895_ (
    .A(_09027_),
    .ZN(_09028_)
  );
  AND2_X1 _18896_ (
    .A1(_08600_),
    .A2(_09027_),
    .ZN(_09029_)
  );
  INV_X1 _18897_ (
    .A(_09029_),
    .ZN(_09030_)
  );
  AND2_X1 _18898_ (
    .A1(_08601_),
    .A2(_09028_),
    .ZN(_09031_)
  );
  INV_X1 _18899_ (
    .A(_09031_),
    .ZN(_09032_)
  );
  AND2_X1 _18900_ (
    .A1(_09030_),
    .A2(_09032_),
    .ZN(_09033_)
  );
  INV_X1 _18901_ (
    .A(_09033_),
    .ZN(_09034_)
  );
  AND2_X1 _18902_ (
    .A1(_08995_),
    .A2(_09033_),
    .ZN(_09035_)
  );
  INV_X1 _18903_ (
    .A(_09035_),
    .ZN(_09036_)
  );
  AND2_X1 _18904_ (
    .A1(_08994_),
    .A2(_09034_),
    .ZN(_09038_)
  );
  INV_X1 _18905_ (
    .A(_09038_),
    .ZN(_09039_)
  );
  AND2_X1 _18906_ (
    .A1(_09036_),
    .A2(_09039_),
    .ZN(_09040_)
  );
  INV_X1 _18907_ (
    .A(_09040_),
    .ZN(_09041_)
  );
  AND2_X1 _18908_ (
    .A1(_08991_),
    .A2(_09040_),
    .ZN(_09042_)
  );
  INV_X1 _18909_ (
    .A(_09042_),
    .ZN(_09043_)
  );
  AND2_X1 _18910_ (
    .A1(_08992_),
    .A2(_09041_),
    .ZN(_09044_)
  );
  INV_X1 _18911_ (
    .A(_09044_),
    .ZN(_09045_)
  );
  AND2_X1 _18912_ (
    .A1(_09043_),
    .A2(_09045_),
    .ZN(_09046_)
  );
  INV_X1 _18913_ (
    .A(_09046_),
    .ZN(_09047_)
  );
  AND2_X1 _18914_ (
    .A1(_08838_),
    .A2(_09046_),
    .ZN(_09049_)
  );
  INV_X1 _18915_ (
    .A(_09049_),
    .ZN(_09050_)
  );
  AND2_X1 _18916_ (
    .A1(_08837_),
    .A2(_09047_),
    .ZN(_09051_)
  );
  INV_X1 _18917_ (
    .A(_09051_),
    .ZN(_09052_)
  );
  AND2_X1 _18918_ (
    .A1(_09050_),
    .A2(_09052_),
    .ZN(_09053_)
  );
  INV_X1 _18919_ (
    .A(_09053_),
    .ZN(_09054_)
  );
  AND2_X1 _18920_ (
    .A1(_08704_),
    .A2(_08711_),
    .ZN(_09055_)
  );
  INV_X1 _18921_ (
    .A(_09055_),
    .ZN(_09056_)
  );
  AND2_X1 _18922_ (
    .A1(_07804_),
    .A2(_09056_),
    .ZN(_09057_)
  );
  INV_X1 _18923_ (
    .A(_09057_),
    .ZN(_09058_)
  );
  AND2_X1 _18924_ (
    .A1(_07805_),
    .A2(_09055_),
    .ZN(_09060_)
  );
  INV_X1 _18925_ (
    .A(_09060_),
    .ZN(_09061_)
  );
  AND2_X1 _18926_ (
    .A1(_09058_),
    .A2(_09061_),
    .ZN(_09062_)
  );
  INV_X1 _18927_ (
    .A(_09062_),
    .ZN(_09063_)
  );
  AND2_X1 _18928_ (
    .A1(_08107_),
    .A2(_09062_),
    .ZN(_09064_)
  );
  INV_X1 _18929_ (
    .A(_09064_),
    .ZN(_09065_)
  );
  AND2_X1 _18930_ (
    .A1(_08106_),
    .A2(_09063_),
    .ZN(_09066_)
  );
  INV_X1 _18931_ (
    .A(_09066_),
    .ZN(_09067_)
  );
  AND2_X1 _18932_ (
    .A1(_09065_),
    .A2(_09067_),
    .ZN(_09068_)
  );
  INV_X1 _18933_ (
    .A(_09068_),
    .ZN(_09069_)
  );
  AND2_X1 _18934_ (
    .A1(_09053_),
    .A2(_09068_),
    .ZN(_09071_)
  );
  INV_X1 _18935_ (
    .A(_09071_),
    .ZN(_09072_)
  );
  AND2_X1 _18936_ (
    .A1(_09054_),
    .A2(_09069_),
    .ZN(_09073_)
  );
  INV_X1 _18937_ (
    .A(_09073_),
    .ZN(_09074_)
  );
  AND2_X1 _18938_ (
    .A1(_09072_),
    .A2(_09074_),
    .ZN(_09075_)
  );
  INV_X1 _18939_ (
    .A(_09075_),
    .ZN(_09076_)
  );
  AND2_X1 _18940_ (
    .A1(_08836_),
    .A2(_09075_),
    .ZN(_09077_)
  );
  INV_X1 _18941_ (
    .A(_09077_),
    .ZN(_09078_)
  );
  AND2_X1 _18942_ (
    .A1(_08835_),
    .A2(_09076_),
    .ZN(_09079_)
  );
  INV_X1 _18943_ (
    .A(_09079_),
    .ZN(_09080_)
  );
  AND2_X1 _18944_ (
    .A1(_09078_),
    .A2(_09080_),
    .ZN(_09082_)
  );
  INV_X1 _18945_ (
    .A(_09082_),
    .ZN(_09083_)
  );
  AND2_X1 _18946_ (
    .A1(_08834_),
    .A2(_09082_),
    .ZN(_09084_)
  );
  INV_X1 _18947_ (
    .A(_09084_),
    .ZN(_09085_)
  );
  AND2_X1 _18948_ (
    .A1(_08833_),
    .A2(_09083_),
    .ZN(_09086_)
  );
  INV_X1 _18949_ (
    .A(_09086_),
    .ZN(_09087_)
  );
  AND2_X1 _18950_ (
    .A1(_09085_),
    .A2(_09087_),
    .ZN(_09088_)
  );
  INV_X1 _18951_ (
    .A(_09088_),
    .ZN(_09089_)
  );
  AND2_X1 _18952_ (
    .A1(_08832_),
    .A2(_09088_),
    .ZN(_09090_)
  );
  INV_X1 _18953_ (
    .A(_09090_),
    .ZN(_09091_)
  );
  AND2_X1 _18954_ (
    .A1(_08831_),
    .A2(_09089_),
    .ZN(_09093_)
  );
  INV_X1 _18955_ (
    .A(_09093_),
    .ZN(_09094_)
  );
  AND2_X1 _18956_ (
    .A1(_09091_),
    .A2(_09094_),
    .ZN(_09095_)
  );
  INV_X1 _18957_ (
    .A(_09095_),
    .ZN(_09096_)
  );
  AND2_X1 _18958_ (
    .A1(_08765_),
    .A2(_09095_),
    .ZN(_09097_)
  );
  INV_X1 _18959_ (
    .A(_09097_),
    .ZN(_09098_)
  );
  AND2_X1 _18960_ (
    .A1(_08766_),
    .A2(_09096_),
    .ZN(_09099_)
  );
  INV_X1 _18961_ (
    .A(_09099_),
    .ZN(_09100_)
  );
  AND2_X1 _18962_ (
    .A1(_09098_),
    .A2(_09100_),
    .ZN(_09101_)
  );
  INV_X1 _18963_ (
    .A(_09101_),
    .ZN(_09102_)
  );
  AND2_X1 _18964_ (
    .A1(_08829_),
    .A2(_09102_),
    .ZN(_09104_)
  );
  INV_X1 _18965_ (
    .A(_09104_),
    .ZN(_09105_)
  );
  AND2_X1 _18966_ (
    .A1(_08830_),
    .A2(_09101_),
    .ZN(_09106_)
  );
  INV_X1 _18967_ (
    .A(_09106_),
    .ZN(_09107_)
  );
  AND2_X1 _18968_ (
    .A1(_09105_),
    .A2(_09107_),
    .ZN(_09108_)
  );
  INV_X1 _18969_ (
    .A(_09108_),
    .ZN(_09109_)
  );
  AND2_X1 _18970_ (
    .A1(remainder[64]),
    .A2(_09108_),
    .ZN(_09110_)
  );
  INV_X1 _18971_ (
    .A(_09110_),
    .ZN(_09111_)
  );
  AND2_X1 _18972_ (
    .A1(_04415_),
    .A2(_09109_),
    .ZN(_09112_)
  );
  INV_X1 _18973_ (
    .A(_09112_),
    .ZN(_09113_)
  );
  AND2_X1 _18974_ (
    .A1(_09111_),
    .A2(_09113_),
    .ZN(_09115_)
  );
  INV_X1 _18975_ (
    .A(_09115_),
    .ZN(_09116_)
  );
  AND2_X1 _18976_ (
    .A1(_08827_),
    .A2(_09115_),
    .ZN(_09117_)
  );
  INV_X1 _18977_ (
    .A(_09117_),
    .ZN(_09118_)
  );
  AND2_X1 _18978_ (
    .A1(_08826_),
    .A2(_09116_),
    .ZN(_09119_)
  );
  INV_X1 _18979_ (
    .A(_09119_),
    .ZN(_09120_)
  );
  AND2_X1 _18980_ (
    .A1(_02082_),
    .A2(_09120_),
    .ZN(_09121_)
  );
  AND2_X1 _18981_ (
    .A1(_09118_),
    .A2(_09121_),
    .ZN(_09122_)
  );
  INV_X1 _18982_ (
    .A(_09122_),
    .ZN(_09123_)
  );
  AND2_X1 _18983_ (
    .A1(remainder[56]),
    .A2(_02077_),
    .ZN(_09124_)
  );
  INV_X1 _18984_ (
    .A(_09124_),
    .ZN(_09126_)
  );
  MUX2_X1 _18985_ (
    .A(remainder[55]),
    .B(_01952_),
    .S(_10462_),
    .Z(_09127_)
  );
  AND2_X1 _18986_ (
    .A1(_05983_),
    .A2(_09127_),
    .ZN(_09128_)
  );
  INV_X1 _18987_ (
    .A(_09128_),
    .ZN(_09129_)
  );
  AND2_X1 _18988_ (
    .A1(_09126_),
    .A2(_09129_),
    .ZN(_09130_)
  );
  AND2_X1 _18989_ (
    .A1(_09123_),
    .A2(_09130_),
    .ZN(_09131_)
  );
  INV_X1 _18990_ (
    .A(_09131_),
    .ZN(_09132_)
  );
  AND2_X1 _18991_ (
    .A1(_06201_),
    .A2(_09132_),
    .ZN(_00077_)
  );
  AND2_X1 _18992_ (
    .A1(_09111_),
    .A2(_09118_),
    .ZN(_09133_)
  );
  INV_X1 _18993_ (
    .A(_09133_),
    .ZN(_09134_)
  );
  AND2_X1 _18994_ (
    .A1(_09078_),
    .A2(_09085_),
    .ZN(_09136_)
  );
  INV_X1 _18995_ (
    .A(_09136_),
    .ZN(_09137_)
  );
  AND2_X1 _18996_ (
    .A1(_09058_),
    .A2(_09065_),
    .ZN(_09138_)
  );
  INV_X1 _18997_ (
    .A(_09138_),
    .ZN(_09139_)
  );
  AND2_X1 _18998_ (
    .A1(_09050_),
    .A2(_09072_),
    .ZN(_09140_)
  );
  INV_X1 _18999_ (
    .A(_09140_),
    .ZN(_09141_)
  );
  AND2_X1 _19000_ (
    .A1(_08988_),
    .A2(_09043_),
    .ZN(_09142_)
  );
  INV_X1 _19001_ (
    .A(_09142_),
    .ZN(_09143_)
  );
  AND2_X1 _19002_ (
    .A1(_03249_),
    .A2(_08968_),
    .ZN(_09144_)
  );
  INV_X1 _19003_ (
    .A(_09144_),
    .ZN(_09145_)
  );
  AND2_X1 _19004_ (
    .A1(_08624_),
    .A2(_09144_),
    .ZN(_09147_)
  );
  INV_X1 _19005_ (
    .A(_09147_),
    .ZN(_09148_)
  );
  AND2_X1 _19006_ (
    .A1(_08981_),
    .A2(_09148_),
    .ZN(_09149_)
  );
  INV_X1 _19007_ (
    .A(_09149_),
    .ZN(_09150_)
  );
  AND2_X1 _19008_ (
    .A1(_08889_),
    .A2(_08929_),
    .ZN(_09151_)
  );
  INV_X1 _19009_ (
    .A(_09151_),
    .ZN(_09152_)
  );
  AND2_X1 _19010_ (
    .A1(_08876_),
    .A2(_08882_),
    .ZN(_09153_)
  );
  INV_X1 _19011_ (
    .A(_09153_),
    .ZN(_09154_)
  );
  AND2_X1 _19012_ (
    .A1(_08863_),
    .A2(_08869_),
    .ZN(_09155_)
  );
  INV_X1 _19013_ (
    .A(_09155_),
    .ZN(_09156_)
  );
  AND2_X1 _19014_ (
    .A1(_08951_),
    .A2(_08957_),
    .ZN(_09158_)
  );
  INV_X1 _19015_ (
    .A(_09158_),
    .ZN(_09159_)
  );
  AND2_X1 _19016_ (
    .A1(divisor[25]),
    .A2(remainder[7]),
    .ZN(_09160_)
  );
  INV_X1 _19017_ (
    .A(_09160_),
    .ZN(_09161_)
  );
  AND2_X1 _19018_ (
    .A1(divisor[26]),
    .A2(remainder[6]),
    .ZN(_09162_)
  );
  INV_X1 _19019_ (
    .A(_09162_),
    .ZN(_09163_)
  );
  AND2_X1 _19020_ (
    .A1(divisor[27]),
    .A2(remainder[6]),
    .ZN(_09164_)
  );
  INV_X1 _19021_ (
    .A(_09164_),
    .ZN(_09165_)
  );
  AND2_X1 _19022_ (
    .A1(_08859_),
    .A2(_09162_),
    .ZN(_09166_)
  );
  INV_X1 _19023_ (
    .A(_09166_),
    .ZN(_09167_)
  );
  AND2_X1 _19024_ (
    .A1(_08860_),
    .A2(_09163_),
    .ZN(_09169_)
  );
  INV_X1 _19025_ (
    .A(_09169_),
    .ZN(_09170_)
  );
  AND2_X1 _19026_ (
    .A1(_09167_),
    .A2(_09170_),
    .ZN(_09171_)
  );
  INV_X1 _19027_ (
    .A(_09171_),
    .ZN(_09172_)
  );
  AND2_X1 _19028_ (
    .A1(_09160_),
    .A2(_09171_),
    .ZN(_09173_)
  );
  INV_X1 _19029_ (
    .A(_09173_),
    .ZN(_09174_)
  );
  AND2_X1 _19030_ (
    .A1(_09161_),
    .A2(_09172_),
    .ZN(_09175_)
  );
  INV_X1 _19031_ (
    .A(_09175_),
    .ZN(_09176_)
  );
  AND2_X1 _19032_ (
    .A1(_09174_),
    .A2(_09176_),
    .ZN(_09177_)
  );
  INV_X1 _19033_ (
    .A(_09177_),
    .ZN(_09178_)
  );
  AND2_X1 _19034_ (
    .A1(_09159_),
    .A2(_09177_),
    .ZN(_09180_)
  );
  INV_X1 _19035_ (
    .A(_09180_),
    .ZN(_09181_)
  );
  AND2_X1 _19036_ (
    .A1(_09158_),
    .A2(_09178_),
    .ZN(_09182_)
  );
  INV_X1 _19037_ (
    .A(_09182_),
    .ZN(_09183_)
  );
  AND2_X1 _19038_ (
    .A1(_09181_),
    .A2(_09183_),
    .ZN(_09184_)
  );
  INV_X1 _19039_ (
    .A(_09184_),
    .ZN(_09185_)
  );
  AND2_X1 _19040_ (
    .A1(_09156_),
    .A2(_09184_),
    .ZN(_09186_)
  );
  INV_X1 _19041_ (
    .A(_09186_),
    .ZN(_09187_)
  );
  AND2_X1 _19042_ (
    .A1(_09155_),
    .A2(_09185_),
    .ZN(_09188_)
  );
  INV_X1 _19043_ (
    .A(_09188_),
    .ZN(_09189_)
  );
  AND2_X1 _19044_ (
    .A1(_09187_),
    .A2(_09189_),
    .ZN(_09191_)
  );
  INV_X1 _19045_ (
    .A(_09191_),
    .ZN(_09192_)
  );
  AND2_X1 _19046_ (
    .A1(_09154_),
    .A2(_09191_),
    .ZN(_09193_)
  );
  INV_X1 _19047_ (
    .A(_09193_),
    .ZN(_09194_)
  );
  AND2_X1 _19048_ (
    .A1(_09153_),
    .A2(_09192_),
    .ZN(_09195_)
  );
  INV_X1 _19049_ (
    .A(_09195_),
    .ZN(_09196_)
  );
  AND2_X1 _19050_ (
    .A1(_09194_),
    .A2(_09196_),
    .ZN(_09197_)
  );
  INV_X1 _19051_ (
    .A(_09197_),
    .ZN(_09198_)
  );
  AND2_X1 _19052_ (
    .A1(_08902_),
    .A2(_08909_),
    .ZN(_09199_)
  );
  INV_X1 _19053_ (
    .A(_09199_),
    .ZN(_09200_)
  );
  AND2_X1 _19054_ (
    .A1(_08898_),
    .A2(_08900_),
    .ZN(_09202_)
  );
  MUX2_X1 _19055_ (
    .A(_08899_),
    .B(_05018_),
    .S(_08897_),
    .Z(_09203_)
  );
  MUX2_X1 _19056_ (
    .A(_08560_),
    .B(_05007_),
    .S(_09203_),
    .Z(_09204_)
  );
  MUX2_X1 _19057_ (
    .A(_08561_),
    .B(divisor[22]),
    .S(_09203_),
    .Z(_09205_)
  );
  AND2_X1 _19058_ (
    .A1(_09200_),
    .A2(_09204_),
    .ZN(_09206_)
  );
  INV_X1 _19059_ (
    .A(_09206_),
    .ZN(_09207_)
  );
  AND2_X1 _19060_ (
    .A1(_09199_),
    .A2(_09205_),
    .ZN(_09208_)
  );
  INV_X1 _19061_ (
    .A(_09208_),
    .ZN(_09209_)
  );
  AND2_X1 _19062_ (
    .A1(_09207_),
    .A2(_09209_),
    .ZN(_09210_)
  );
  INV_X1 _19063_ (
    .A(_09210_),
    .ZN(_09211_)
  );
  AND2_X1 _19064_ (
    .A1(_08282_),
    .A2(_09210_),
    .ZN(_09213_)
  );
  INV_X1 _19065_ (
    .A(_09213_),
    .ZN(_09214_)
  );
  AND2_X1 _19066_ (
    .A1(_08283_),
    .A2(_09211_),
    .ZN(_09215_)
  );
  INV_X1 _19067_ (
    .A(_09215_),
    .ZN(_09216_)
  );
  AND2_X1 _19068_ (
    .A1(_09214_),
    .A2(_09216_),
    .ZN(_09217_)
  );
  INV_X1 _19069_ (
    .A(_09217_),
    .ZN(_09218_)
  );
  AND2_X1 _19070_ (
    .A1(_09197_),
    .A2(_09217_),
    .ZN(_09219_)
  );
  INV_X1 _19071_ (
    .A(_09219_),
    .ZN(_09220_)
  );
  AND2_X1 _19072_ (
    .A1(_09198_),
    .A2(_09218_),
    .ZN(_09221_)
  );
  INV_X1 _19073_ (
    .A(_09221_),
    .ZN(_09222_)
  );
  AND2_X1 _19074_ (
    .A1(_09220_),
    .A2(_09222_),
    .ZN(_09224_)
  );
  INV_X1 _19075_ (
    .A(_09224_),
    .ZN(_09225_)
  );
  AND2_X1 _19076_ (
    .A1(_09152_),
    .A2(_09224_),
    .ZN(_09226_)
  );
  INV_X1 _19077_ (
    .A(_09226_),
    .ZN(_09227_)
  );
  AND2_X1 _19078_ (
    .A1(_09151_),
    .A2(_09225_),
    .ZN(_09228_)
  );
  INV_X1 _19079_ (
    .A(_09228_),
    .ZN(_09229_)
  );
  AND2_X1 _19080_ (
    .A1(_09227_),
    .A2(_09229_),
    .ZN(_09230_)
  );
  INV_X1 _19081_ (
    .A(_09230_),
    .ZN(_09231_)
  );
  AND2_X1 _19082_ (
    .A1(divisor[32]),
    .A2(remainder[0]),
    .ZN(_09232_)
  );
  INV_X1 _19083_ (
    .A(_09232_),
    .ZN(_09233_)
  );
  AND2_X1 _19084_ (
    .A1(divisor[31]),
    .A2(remainder[1]),
    .ZN(_09235_)
  );
  INV_X1 _19085_ (
    .A(_09235_),
    .ZN(_09236_)
  );
  AND2_X1 _19086_ (
    .A1(divisor[32]),
    .A2(remainder[1]),
    .ZN(_09237_)
  );
  AND2_X1 _19087_ (
    .A1(_08941_),
    .A2(_09237_),
    .ZN(_09238_)
  );
  INV_X1 _19088_ (
    .A(_09238_),
    .ZN(_09239_)
  );
  AND2_X1 _19089_ (
    .A1(_09233_),
    .A2(_09236_),
    .ZN(_09240_)
  );
  INV_X1 _19090_ (
    .A(_09240_),
    .ZN(_09241_)
  );
  AND2_X1 _19091_ (
    .A1(_09239_),
    .A2(_09241_),
    .ZN(_09242_)
  );
  INV_X1 _19092_ (
    .A(_09242_),
    .ZN(_09243_)
  );
  AND2_X1 _19093_ (
    .A1(divisor[28]),
    .A2(remainder[4]),
    .ZN(_09244_)
  );
  INV_X1 _19094_ (
    .A(_09244_),
    .ZN(_09246_)
  );
  AND2_X1 _19095_ (
    .A1(divisor[29]),
    .A2(remainder[3]),
    .ZN(_09247_)
  );
  INV_X1 _19096_ (
    .A(_09247_),
    .ZN(_09248_)
  );
  AND2_X1 _19097_ (
    .A1(divisor[30]),
    .A2(remainder[3]),
    .ZN(_09249_)
  );
  INV_X1 _19098_ (
    .A(_09249_),
    .ZN(_09250_)
  );
  AND2_X1 _19099_ (
    .A1(_08947_),
    .A2(_09247_),
    .ZN(_09251_)
  );
  INV_X1 _19100_ (
    .A(_09251_),
    .ZN(_09252_)
  );
  AND2_X1 _19101_ (
    .A1(_08948_),
    .A2(_09248_),
    .ZN(_09253_)
  );
  INV_X1 _19102_ (
    .A(_09253_),
    .ZN(_09254_)
  );
  AND2_X1 _19103_ (
    .A1(_09252_),
    .A2(_09254_),
    .ZN(_09255_)
  );
  INV_X1 _19104_ (
    .A(_09255_),
    .ZN(_09257_)
  );
  AND2_X1 _19105_ (
    .A1(_09244_),
    .A2(_09255_),
    .ZN(_09258_)
  );
  INV_X1 _19106_ (
    .A(_09258_),
    .ZN(_09259_)
  );
  AND2_X1 _19107_ (
    .A1(_09246_),
    .A2(_09257_),
    .ZN(_09260_)
  );
  INV_X1 _19108_ (
    .A(_09260_),
    .ZN(_09261_)
  );
  AND2_X1 _19109_ (
    .A1(_09259_),
    .A2(_09261_),
    .ZN(_09262_)
  );
  INV_X1 _19110_ (
    .A(_09262_),
    .ZN(_09263_)
  );
  AND2_X1 _19111_ (
    .A1(_09242_),
    .A2(_09262_),
    .ZN(_09264_)
  );
  INV_X1 _19112_ (
    .A(_09264_),
    .ZN(_09265_)
  );
  AND2_X1 _19113_ (
    .A1(_09243_),
    .A2(_09263_),
    .ZN(_09266_)
  );
  INV_X1 _19114_ (
    .A(_09266_),
    .ZN(_09268_)
  );
  AND2_X1 _19115_ (
    .A1(_09265_),
    .A2(_09268_),
    .ZN(_09269_)
  );
  INV_X1 _19116_ (
    .A(_09269_),
    .ZN(_09270_)
  );
  AND2_X1 _19117_ (
    .A1(_08963_),
    .A2(_09269_),
    .ZN(_09271_)
  );
  INV_X1 _19118_ (
    .A(_09271_),
    .ZN(_09272_)
  );
  AND2_X1 _19119_ (
    .A1(_08964_),
    .A2(_09270_),
    .ZN(_09273_)
  );
  INV_X1 _19120_ (
    .A(_09273_),
    .ZN(_09274_)
  );
  AND2_X1 _19121_ (
    .A1(_09272_),
    .A2(_09274_),
    .ZN(_09275_)
  );
  INV_X1 _19122_ (
    .A(_09275_),
    .ZN(_09276_)
  );
  AND2_X1 _19123_ (
    .A1(_09144_),
    .A2(_09276_),
    .ZN(_09277_)
  );
  INV_X1 _19124_ (
    .A(_09277_),
    .ZN(_09279_)
  );
  AND2_X1 _19125_ (
    .A1(_09145_),
    .A2(_09275_),
    .ZN(_09280_)
  );
  INV_X1 _19126_ (
    .A(_09280_),
    .ZN(_09281_)
  );
  AND2_X1 _19127_ (
    .A1(_09279_),
    .A2(_09281_),
    .ZN(_09282_)
  );
  INV_X1 _19128_ (
    .A(_09282_),
    .ZN(_09283_)
  );
  AND2_X1 _19129_ (
    .A1(_09230_),
    .A2(_09283_),
    .ZN(_09284_)
  );
  INV_X1 _19130_ (
    .A(_09284_),
    .ZN(_09285_)
  );
  AND2_X1 _19131_ (
    .A1(_09231_),
    .A2(_09282_),
    .ZN(_09286_)
  );
  INV_X1 _19132_ (
    .A(_09286_),
    .ZN(_09287_)
  );
  AND2_X1 _19133_ (
    .A1(_09285_),
    .A2(_09287_),
    .ZN(_09288_)
  );
  INV_X1 _19134_ (
    .A(_09288_),
    .ZN(_09290_)
  );
  AND2_X1 _19135_ (
    .A1(_09150_),
    .A2(_09288_),
    .ZN(_09291_)
  );
  INV_X1 _19136_ (
    .A(_09291_),
    .ZN(_09292_)
  );
  AND2_X1 _19137_ (
    .A1(_09149_),
    .A2(_09290_),
    .ZN(_09293_)
  );
  INV_X1 _19138_ (
    .A(_09293_),
    .ZN(_09294_)
  );
  AND2_X1 _19139_ (
    .A1(_09292_),
    .A2(_09294_),
    .ZN(_09295_)
  );
  INV_X1 _19140_ (
    .A(_09295_),
    .ZN(_09296_)
  );
  AND2_X1 _19141_ (
    .A1(_09017_),
    .A2(_09023_),
    .ZN(_09297_)
  );
  INV_X1 _19142_ (
    .A(_09297_),
    .ZN(_09298_)
  );
  AND2_X1 _19143_ (
    .A1(_09003_),
    .A2(_09010_),
    .ZN(_09299_)
  );
  INV_X1 _19144_ (
    .A(_09299_),
    .ZN(_09301_)
  );
  AND2_X1 _19145_ (
    .A1(_08915_),
    .A2(_08922_),
    .ZN(_09302_)
  );
  INV_X1 _19146_ (
    .A(_09302_),
    .ZN(_09303_)
  );
  AND2_X1 _19147_ (
    .A1(_08674_),
    .A2(_09303_),
    .ZN(_09304_)
  );
  INV_X1 _19148_ (
    .A(_09304_),
    .ZN(_09305_)
  );
  AND2_X1 _19149_ (
    .A1(_08676_),
    .A2(_09302_),
    .ZN(_09306_)
  );
  INV_X1 _19150_ (
    .A(_09306_),
    .ZN(_09307_)
  );
  AND2_X1 _19151_ (
    .A1(_09305_),
    .A2(_09307_),
    .ZN(_09308_)
  );
  INV_X1 _19152_ (
    .A(_09308_),
    .ZN(_09309_)
  );
  AND2_X1 _19153_ (
    .A1(_08999_),
    .A2(_09308_),
    .ZN(_09310_)
  );
  INV_X1 _19154_ (
    .A(_09310_),
    .ZN(_09312_)
  );
  AND2_X1 _19155_ (
    .A1(_08998_),
    .A2(_09309_),
    .ZN(_09313_)
  );
  INV_X1 _19156_ (
    .A(_09313_),
    .ZN(_09314_)
  );
  AND2_X1 _19157_ (
    .A1(_09312_),
    .A2(_09314_),
    .ZN(_09315_)
  );
  INV_X1 _19158_ (
    .A(_09315_),
    .ZN(_09316_)
  );
  AND2_X1 _19159_ (
    .A1(_09301_),
    .A2(_09315_),
    .ZN(_09317_)
  );
  INV_X1 _19160_ (
    .A(_09317_),
    .ZN(_09318_)
  );
  AND2_X1 _19161_ (
    .A1(_09299_),
    .A2(_09316_),
    .ZN(_09319_)
  );
  INV_X1 _19162_ (
    .A(_09319_),
    .ZN(_09320_)
  );
  AND2_X1 _19163_ (
    .A1(_09318_),
    .A2(_09320_),
    .ZN(_09321_)
  );
  INV_X1 _19164_ (
    .A(_09321_),
    .ZN(_09323_)
  );
  AND2_X1 _19165_ (
    .A1(_07082_),
    .A2(_09321_),
    .ZN(_09324_)
  );
  INV_X1 _19166_ (
    .A(_09324_),
    .ZN(_09325_)
  );
  AND2_X1 _19167_ (
    .A1(_07083_),
    .A2(_09323_),
    .ZN(_09326_)
  );
  INV_X1 _19168_ (
    .A(_09326_),
    .ZN(_09327_)
  );
  AND2_X1 _19169_ (
    .A1(_09325_),
    .A2(_09327_),
    .ZN(_09328_)
  );
  INV_X1 _19170_ (
    .A(_09328_),
    .ZN(_09329_)
  );
  AND2_X1 _19171_ (
    .A1(_08934_),
    .A2(_09328_),
    .ZN(_09330_)
  );
  INV_X1 _19172_ (
    .A(_09330_),
    .ZN(_09331_)
  );
  AND2_X1 _19173_ (
    .A1(_08935_),
    .A2(_09329_),
    .ZN(_09332_)
  );
  INV_X1 _19174_ (
    .A(_09332_),
    .ZN(_09334_)
  );
  AND2_X1 _19175_ (
    .A1(_09331_),
    .A2(_09334_),
    .ZN(_09335_)
  );
  INV_X1 _19176_ (
    .A(_09335_),
    .ZN(_09336_)
  );
  AND2_X1 _19177_ (
    .A1(_09298_),
    .A2(_09335_),
    .ZN(_09337_)
  );
  INV_X1 _19178_ (
    .A(_09337_),
    .ZN(_09338_)
  );
  AND2_X1 _19179_ (
    .A1(_09297_),
    .A2(_09336_),
    .ZN(_09339_)
  );
  INV_X1 _19180_ (
    .A(_09339_),
    .ZN(_09340_)
  );
  AND2_X1 _19181_ (
    .A1(_09338_),
    .A2(_09340_),
    .ZN(_09341_)
  );
  INV_X1 _19182_ (
    .A(_09341_),
    .ZN(_09342_)
  );
  AND2_X1 _19183_ (
    .A1(_09295_),
    .A2(_09341_),
    .ZN(_09343_)
  );
  INV_X1 _19184_ (
    .A(_09343_),
    .ZN(_09345_)
  );
  AND2_X1 _19185_ (
    .A1(_09296_),
    .A2(_09342_),
    .ZN(_09346_)
  );
  INV_X1 _19186_ (
    .A(_09346_),
    .ZN(_09347_)
  );
  AND2_X1 _19187_ (
    .A1(_09345_),
    .A2(_09347_),
    .ZN(_09348_)
  );
  INV_X1 _19188_ (
    .A(_09348_),
    .ZN(_09349_)
  );
  AND2_X1 _19189_ (
    .A1(_09143_),
    .A2(_09348_),
    .ZN(_09350_)
  );
  INV_X1 _19190_ (
    .A(_09350_),
    .ZN(_09351_)
  );
  AND2_X1 _19191_ (
    .A1(_09142_),
    .A2(_09349_),
    .ZN(_09352_)
  );
  INV_X1 _19192_ (
    .A(_09352_),
    .ZN(_09353_)
  );
  AND2_X1 _19193_ (
    .A1(_09351_),
    .A2(_09353_),
    .ZN(_09354_)
  );
  INV_X1 _19194_ (
    .A(_09354_),
    .ZN(_09356_)
  );
  AND2_X1 _19195_ (
    .A1(_09030_),
    .A2(_09036_),
    .ZN(_09357_)
  );
  INV_X1 _19196_ (
    .A(_09357_),
    .ZN(_09358_)
  );
  AND2_X1 _19197_ (
    .A1(_07804_),
    .A2(_09358_),
    .ZN(_09359_)
  );
  INV_X1 _19198_ (
    .A(_09359_),
    .ZN(_09360_)
  );
  AND2_X1 _19199_ (
    .A1(_07805_),
    .A2(_09357_),
    .ZN(_09361_)
  );
  INV_X1 _19200_ (
    .A(_09361_),
    .ZN(_09362_)
  );
  AND2_X1 _19201_ (
    .A1(_09360_),
    .A2(_09362_),
    .ZN(_09363_)
  );
  INV_X1 _19202_ (
    .A(_09363_),
    .ZN(_09364_)
  );
  AND2_X1 _19203_ (
    .A1(_08107_),
    .A2(_09363_),
    .ZN(_09365_)
  );
  INV_X1 _19204_ (
    .A(_09365_),
    .ZN(_09367_)
  );
  AND2_X1 _19205_ (
    .A1(_08106_),
    .A2(_09364_),
    .ZN(_09368_)
  );
  INV_X1 _19206_ (
    .A(_09368_),
    .ZN(_09369_)
  );
  AND2_X1 _19207_ (
    .A1(_09367_),
    .A2(_09369_),
    .ZN(_09370_)
  );
  INV_X1 _19208_ (
    .A(_09370_),
    .ZN(_09371_)
  );
  AND2_X1 _19209_ (
    .A1(_09354_),
    .A2(_09370_),
    .ZN(_09372_)
  );
  INV_X1 _19210_ (
    .A(_09372_),
    .ZN(_09373_)
  );
  AND2_X1 _19211_ (
    .A1(_09356_),
    .A2(_09371_),
    .ZN(_09374_)
  );
  INV_X1 _19212_ (
    .A(_09374_),
    .ZN(_09375_)
  );
  AND2_X1 _19213_ (
    .A1(_09373_),
    .A2(_09375_),
    .ZN(_09376_)
  );
  INV_X1 _19214_ (
    .A(_09376_),
    .ZN(_09378_)
  );
  AND2_X1 _19215_ (
    .A1(_09141_),
    .A2(_09376_),
    .ZN(_09379_)
  );
  INV_X1 _19216_ (
    .A(_09379_),
    .ZN(_09380_)
  );
  AND2_X1 _19217_ (
    .A1(_09140_),
    .A2(_09378_),
    .ZN(_09381_)
  );
  INV_X1 _19218_ (
    .A(_09381_),
    .ZN(_09382_)
  );
  AND2_X1 _19219_ (
    .A1(_09380_),
    .A2(_09382_),
    .ZN(_09383_)
  );
  INV_X1 _19220_ (
    .A(_09383_),
    .ZN(_09384_)
  );
  AND2_X1 _19221_ (
    .A1(_09139_),
    .A2(_09383_),
    .ZN(_09385_)
  );
  INV_X1 _19222_ (
    .A(_09385_),
    .ZN(_09386_)
  );
  AND2_X1 _19223_ (
    .A1(_09138_),
    .A2(_09384_),
    .ZN(_09387_)
  );
  INV_X1 _19224_ (
    .A(_09387_),
    .ZN(_09389_)
  );
  AND2_X1 _19225_ (
    .A1(_09386_),
    .A2(_09389_),
    .ZN(_09390_)
  );
  INV_X1 _19226_ (
    .A(_09390_),
    .ZN(_09391_)
  );
  AND2_X1 _19227_ (
    .A1(_09137_),
    .A2(_09390_),
    .ZN(_09392_)
  );
  INV_X1 _19228_ (
    .A(_09392_),
    .ZN(_09393_)
  );
  AND2_X1 _19229_ (
    .A1(_09136_),
    .A2(_09391_),
    .ZN(_09394_)
  );
  INV_X1 _19230_ (
    .A(_09394_),
    .ZN(_09395_)
  );
  AND2_X1 _19231_ (
    .A1(_09393_),
    .A2(_09395_),
    .ZN(_09396_)
  );
  INV_X1 _19232_ (
    .A(_09396_),
    .ZN(_09397_)
  );
  AND2_X1 _19233_ (
    .A1(_09090_),
    .A2(_09396_),
    .ZN(_09398_)
  );
  INV_X1 _19234_ (
    .A(_09398_),
    .ZN(_09400_)
  );
  AND2_X1 _19235_ (
    .A1(_09091_),
    .A2(_09397_),
    .ZN(_09401_)
  );
  INV_X1 _19236_ (
    .A(_09401_),
    .ZN(_09402_)
  );
  AND2_X1 _19237_ (
    .A1(_09400_),
    .A2(_09402_),
    .ZN(_09403_)
  );
  INV_X1 _19238_ (
    .A(_09403_),
    .ZN(_09404_)
  );
  AND2_X1 _19239_ (
    .A1(_08829_),
    .A2(_09098_),
    .ZN(_09405_)
  );
  INV_X1 _19240_ (
    .A(_09405_),
    .ZN(_09406_)
  );
  AND2_X1 _19241_ (
    .A1(_09100_),
    .A2(_09406_),
    .ZN(_09407_)
  );
  AND2_X1 _19242_ (
    .A1(_09098_),
    .A2(_09107_),
    .ZN(_09408_)
  );
  AND2_X1 _19243_ (
    .A1(_09403_),
    .A2(_09407_),
    .ZN(_09409_)
  );
  INV_X1 _19244_ (
    .A(_09409_),
    .ZN(_09411_)
  );
  AND2_X1 _19245_ (
    .A1(_09404_),
    .A2(_09408_),
    .ZN(_09412_)
  );
  INV_X1 _19246_ (
    .A(_09412_),
    .ZN(_09413_)
  );
  AND2_X1 _19247_ (
    .A1(_09411_),
    .A2(_09413_),
    .ZN(_09414_)
  );
  INV_X1 _19248_ (
    .A(_09414_),
    .ZN(_09415_)
  );
  AND2_X1 _19249_ (
    .A1(remainder[65]),
    .A2(_09414_),
    .ZN(_09416_)
  );
  INV_X1 _19250_ (
    .A(_09416_),
    .ZN(_09417_)
  );
  AND2_X1 _19251_ (
    .A1(_04404_),
    .A2(_09415_),
    .ZN(_09418_)
  );
  INV_X1 _19252_ (
    .A(_09418_),
    .ZN(_09419_)
  );
  AND2_X1 _19253_ (
    .A1(_09417_),
    .A2(_09419_),
    .ZN(_09420_)
  );
  INV_X1 _19254_ (
    .A(_09420_),
    .ZN(_09422_)
  );
  AND2_X1 _19255_ (
    .A1(_09134_),
    .A2(_09420_),
    .ZN(_09423_)
  );
  INV_X1 _19256_ (
    .A(_09423_),
    .ZN(_09424_)
  );
  AND2_X1 _19257_ (
    .A1(_09133_),
    .A2(_09422_),
    .ZN(_09425_)
  );
  INV_X1 _19258_ (
    .A(_09425_),
    .ZN(_09426_)
  );
  AND2_X1 _19259_ (
    .A1(_02082_),
    .A2(_09426_),
    .ZN(_09427_)
  );
  AND2_X1 _19260_ (
    .A1(_09424_),
    .A2(_09427_),
    .ZN(_09428_)
  );
  INV_X1 _19261_ (
    .A(_09428_),
    .ZN(_09429_)
  );
  AND2_X1 _19262_ (
    .A1(remainder[57]),
    .A2(_02077_),
    .ZN(_09430_)
  );
  INV_X1 _19263_ (
    .A(_09430_),
    .ZN(_09431_)
  );
  AND2_X1 _19264_ (
    .A1(_04503_),
    .A2(_10451_),
    .ZN(_09433_)
  );
  INV_X1 _19265_ (
    .A(_09433_),
    .ZN(_09434_)
  );
  AND2_X1 _19266_ (
    .A1(_10462_),
    .A2(_01964_),
    .ZN(_09435_)
  );
  INV_X1 _19267_ (
    .A(_09435_),
    .ZN(_09436_)
  );
  AND2_X1 _19268_ (
    .A1(_05983_),
    .A2(_09436_),
    .ZN(_09437_)
  );
  AND2_X1 _19269_ (
    .A1(_09434_),
    .A2(_09437_),
    .ZN(_09438_)
  );
  INV_X1 _19270_ (
    .A(_09438_),
    .ZN(_09439_)
  );
  AND2_X1 _19271_ (
    .A1(_09431_),
    .A2(_09439_),
    .ZN(_09440_)
  );
  AND2_X1 _19272_ (
    .A1(_09429_),
    .A2(_09440_),
    .ZN(_09441_)
  );
  INV_X1 _19273_ (
    .A(_09441_),
    .ZN(_09442_)
  );
  AND2_X1 _19274_ (
    .A1(_06201_),
    .A2(_09442_),
    .ZN(_00078_)
  );
  AND2_X1 _19275_ (
    .A1(_09417_),
    .A2(_09424_),
    .ZN(_09444_)
  );
  INV_X1 _19276_ (
    .A(_09444_),
    .ZN(_09445_)
  );
  AND2_X1 _19277_ (
    .A1(_09400_),
    .A2(_09411_),
    .ZN(_09446_)
  );
  INV_X1 _19278_ (
    .A(_09446_),
    .ZN(_09447_)
  );
  AND2_X1 _19279_ (
    .A1(_09380_),
    .A2(_09386_),
    .ZN(_09448_)
  );
  INV_X1 _19280_ (
    .A(_09448_),
    .ZN(_09449_)
  );
  AND2_X1 _19281_ (
    .A1(_09360_),
    .A2(_09367_),
    .ZN(_09450_)
  );
  INV_X1 _19282_ (
    .A(_09450_),
    .ZN(_09451_)
  );
  AND2_X1 _19283_ (
    .A1(_09351_),
    .A2(_09373_),
    .ZN(_09452_)
  );
  INV_X1 _19284_ (
    .A(_09452_),
    .ZN(_09454_)
  );
  AND2_X1 _19285_ (
    .A1(_09292_),
    .A2(_09345_),
    .ZN(_09455_)
  );
  INV_X1 _19286_ (
    .A(_09455_),
    .ZN(_09456_)
  );
  AND2_X1 _19287_ (
    .A1(_03249_),
    .A2(_09276_),
    .ZN(_09457_)
  );
  INV_X1 _19288_ (
    .A(_09457_),
    .ZN(_09458_)
  );
  AND2_X1 _19289_ (
    .A1(_08967_),
    .A2(_09457_),
    .ZN(_09459_)
  );
  INV_X1 _19290_ (
    .A(_09459_),
    .ZN(_09460_)
  );
  AND2_X1 _19291_ (
    .A1(_09285_),
    .A2(_09460_),
    .ZN(_09461_)
  );
  INV_X1 _19292_ (
    .A(_09461_),
    .ZN(_09462_)
  );
  AND2_X1 _19293_ (
    .A1(_09194_),
    .A2(_09220_),
    .ZN(_09463_)
  );
  INV_X1 _19294_ (
    .A(_09463_),
    .ZN(_09465_)
  );
  AND2_X1 _19295_ (
    .A1(_09181_),
    .A2(_09187_),
    .ZN(_09466_)
  );
  INV_X1 _19296_ (
    .A(_09466_),
    .ZN(_09467_)
  );
  AND2_X1 _19297_ (
    .A1(_09167_),
    .A2(_09174_),
    .ZN(_09468_)
  );
  INV_X1 _19298_ (
    .A(_09468_),
    .ZN(_09469_)
  );
  AND2_X1 _19299_ (
    .A1(_09252_),
    .A2(_09259_),
    .ZN(_09470_)
  );
  INV_X1 _19300_ (
    .A(_09470_),
    .ZN(_09471_)
  );
  AND2_X1 _19301_ (
    .A1(remainder[32]),
    .A2(divisor[25]),
    .ZN(_09472_)
  );
  INV_X1 _19302_ (
    .A(_09472_),
    .ZN(_09473_)
  );
  AND2_X1 _19303_ (
    .A1(divisor[26]),
    .A2(remainder[7]),
    .ZN(_09474_)
  );
  INV_X1 _19304_ (
    .A(_09474_),
    .ZN(_09476_)
  );
  AND2_X1 _19305_ (
    .A1(divisor[27]),
    .A2(remainder[7]),
    .ZN(_09477_)
  );
  INV_X1 _19306_ (
    .A(_09477_),
    .ZN(_09478_)
  );
  AND2_X1 _19307_ (
    .A1(_09162_),
    .A2(_09477_),
    .ZN(_09479_)
  );
  INV_X1 _19308_ (
    .A(_09479_),
    .ZN(_09480_)
  );
  AND2_X1 _19309_ (
    .A1(_09165_),
    .A2(_09476_),
    .ZN(_09481_)
  );
  INV_X1 _19310_ (
    .A(_09481_),
    .ZN(_09482_)
  );
  AND2_X1 _19311_ (
    .A1(_09480_),
    .A2(_09482_),
    .ZN(_09483_)
  );
  INV_X1 _19312_ (
    .A(_09483_),
    .ZN(_09484_)
  );
  AND2_X1 _19313_ (
    .A1(_09472_),
    .A2(_09483_),
    .ZN(_09485_)
  );
  INV_X1 _19314_ (
    .A(_09485_),
    .ZN(_09487_)
  );
  AND2_X1 _19315_ (
    .A1(_09473_),
    .A2(_09484_),
    .ZN(_09488_)
  );
  INV_X1 _19316_ (
    .A(_09488_),
    .ZN(_09489_)
  );
  AND2_X1 _19317_ (
    .A1(_09487_),
    .A2(_09489_),
    .ZN(_09490_)
  );
  INV_X1 _19318_ (
    .A(_09490_),
    .ZN(_09491_)
  );
  AND2_X1 _19319_ (
    .A1(_09471_),
    .A2(_09490_),
    .ZN(_09492_)
  );
  INV_X1 _19320_ (
    .A(_09492_),
    .ZN(_09493_)
  );
  AND2_X1 _19321_ (
    .A1(_09470_),
    .A2(_09491_),
    .ZN(_09494_)
  );
  INV_X1 _19322_ (
    .A(_09494_),
    .ZN(_09495_)
  );
  AND2_X1 _19323_ (
    .A1(_09493_),
    .A2(_09495_),
    .ZN(_09496_)
  );
  INV_X1 _19324_ (
    .A(_09496_),
    .ZN(_09498_)
  );
  AND2_X1 _19325_ (
    .A1(_09469_),
    .A2(_09496_),
    .ZN(_09499_)
  );
  INV_X1 _19326_ (
    .A(_09499_),
    .ZN(_09500_)
  );
  AND2_X1 _19327_ (
    .A1(_09468_),
    .A2(_09498_),
    .ZN(_09501_)
  );
  INV_X1 _19328_ (
    .A(_09501_),
    .ZN(_09502_)
  );
  AND2_X1 _19329_ (
    .A1(_09500_),
    .A2(_09502_),
    .ZN(_09503_)
  );
  INV_X1 _19330_ (
    .A(_09503_),
    .ZN(_09504_)
  );
  AND2_X1 _19331_ (
    .A1(_09467_),
    .A2(_09503_),
    .ZN(_09505_)
  );
  INV_X1 _19332_ (
    .A(_09505_),
    .ZN(_09506_)
  );
  AND2_X1 _19333_ (
    .A1(_09466_),
    .A2(_09504_),
    .ZN(_09507_)
  );
  INV_X1 _19334_ (
    .A(_09507_),
    .ZN(_09509_)
  );
  AND2_X1 _19335_ (
    .A1(_09506_),
    .A2(_09509_),
    .ZN(_09510_)
  );
  INV_X1 _19336_ (
    .A(_09510_),
    .ZN(_09511_)
  );
  AND2_X1 _19337_ (
    .A1(_08561_),
    .A2(_09202_),
    .ZN(_09512_)
  );
  INV_X1 _19338_ (
    .A(_09512_),
    .ZN(_09513_)
  );
  AND2_X1 _19339_ (
    .A1(_09207_),
    .A2(_09513_),
    .ZN(_09514_)
  );
  INV_X1 _19340_ (
    .A(_09514_),
    .ZN(_09515_)
  );
  AND2_X1 _19341_ (
    .A1(_08282_),
    .A2(_09514_),
    .ZN(_09516_)
  );
  INV_X1 _19342_ (
    .A(_09516_),
    .ZN(_09517_)
  );
  AND2_X1 _19343_ (
    .A1(_08283_),
    .A2(_09515_),
    .ZN(_09518_)
  );
  INV_X1 _19344_ (
    .A(_09518_),
    .ZN(_09520_)
  );
  AND2_X1 _19345_ (
    .A1(_09517_),
    .A2(_09520_),
    .ZN(_09521_)
  );
  INV_X1 _19346_ (
    .A(_09521_),
    .ZN(_09522_)
  );
  AND2_X1 _19347_ (
    .A1(_09510_),
    .A2(_09521_),
    .ZN(_09523_)
  );
  INV_X1 _19348_ (
    .A(_09523_),
    .ZN(_09524_)
  );
  AND2_X1 _19349_ (
    .A1(_09511_),
    .A2(_09522_),
    .ZN(_09525_)
  );
  INV_X1 _19350_ (
    .A(_09525_),
    .ZN(_09526_)
  );
  AND2_X1 _19351_ (
    .A1(_09524_),
    .A2(_09526_),
    .ZN(_09527_)
  );
  INV_X1 _19352_ (
    .A(_09527_),
    .ZN(_09528_)
  );
  AND2_X1 _19353_ (
    .A1(_09271_),
    .A2(_09527_),
    .ZN(_09529_)
  );
  INV_X1 _19354_ (
    .A(_09529_),
    .ZN(_09531_)
  );
  AND2_X1 _19355_ (
    .A1(_09272_),
    .A2(_09528_),
    .ZN(_09532_)
  );
  INV_X1 _19356_ (
    .A(_09532_),
    .ZN(_09533_)
  );
  AND2_X1 _19357_ (
    .A1(_09531_),
    .A2(_09533_),
    .ZN(_09534_)
  );
  INV_X1 _19358_ (
    .A(_09534_),
    .ZN(_09535_)
  );
  AND2_X1 _19359_ (
    .A1(_09465_),
    .A2(_09534_),
    .ZN(_09536_)
  );
  INV_X1 _19360_ (
    .A(_09536_),
    .ZN(_09537_)
  );
  AND2_X1 _19361_ (
    .A1(_09463_),
    .A2(_09535_),
    .ZN(_09538_)
  );
  INV_X1 _19362_ (
    .A(_09538_),
    .ZN(_09539_)
  );
  AND2_X1 _19363_ (
    .A1(_09537_),
    .A2(_09539_),
    .ZN(_09540_)
  );
  INV_X1 _19364_ (
    .A(_09540_),
    .ZN(_09542_)
  );
  AND2_X1 _19365_ (
    .A1(divisor[31]),
    .A2(remainder[2]),
    .ZN(_09543_)
  );
  INV_X1 _19366_ (
    .A(_09543_),
    .ZN(_09544_)
  );
  AND2_X1 _19367_ (
    .A1(remainder[1]),
    .A2(_09232_),
    .ZN(_09545_)
  );
  INV_X1 _19368_ (
    .A(_09545_),
    .ZN(_09546_)
  );
  MUX2_X1 _19369_ (
    .A(_09232_),
    .B(_05073_),
    .S(_09237_),
    .Z(_09547_)
  );
  MUX2_X1 _19370_ (
    .A(_09233_),
    .B(remainder[0]),
    .S(_09237_),
    .Z(_09548_)
  );
  AND2_X1 _19371_ (
    .A1(_09543_),
    .A2(_09547_),
    .ZN(_09549_)
  );
  INV_X1 _19372_ (
    .A(_09549_),
    .ZN(_09550_)
  );
  AND2_X1 _19373_ (
    .A1(_09544_),
    .A2(_09548_),
    .ZN(_09551_)
  );
  INV_X1 _19374_ (
    .A(_09551_),
    .ZN(_09553_)
  );
  AND2_X1 _19375_ (
    .A1(_09550_),
    .A2(_09553_),
    .ZN(_09554_)
  );
  INV_X1 _19376_ (
    .A(_09554_),
    .ZN(_09555_)
  );
  AND2_X1 _19377_ (
    .A1(_09238_),
    .A2(_09554_),
    .ZN(_09556_)
  );
  INV_X1 _19378_ (
    .A(_09556_),
    .ZN(_09557_)
  );
  AND2_X1 _19379_ (
    .A1(_09239_),
    .A2(_09555_),
    .ZN(_09558_)
  );
  INV_X1 _19380_ (
    .A(_09558_),
    .ZN(_09559_)
  );
  AND2_X1 _19381_ (
    .A1(_09557_),
    .A2(_09559_),
    .ZN(_09560_)
  );
  INV_X1 _19382_ (
    .A(_09560_),
    .ZN(_09561_)
  );
  AND2_X1 _19383_ (
    .A1(divisor[28]),
    .A2(remainder[5]),
    .ZN(_09562_)
  );
  INV_X1 _19384_ (
    .A(_09562_),
    .ZN(_09564_)
  );
  AND2_X1 _19385_ (
    .A1(divisor[29]),
    .A2(remainder[4]),
    .ZN(_09565_)
  );
  INV_X1 _19386_ (
    .A(_09565_),
    .ZN(_09566_)
  );
  AND2_X1 _19387_ (
    .A1(divisor[30]),
    .A2(remainder[4]),
    .ZN(_09567_)
  );
  INV_X1 _19388_ (
    .A(_09567_),
    .ZN(_09568_)
  );
  AND2_X1 _19389_ (
    .A1(_09249_),
    .A2(_09565_),
    .ZN(_09569_)
  );
  INV_X1 _19390_ (
    .A(_09569_),
    .ZN(_09570_)
  );
  AND2_X1 _19391_ (
    .A1(_09250_),
    .A2(_09566_),
    .ZN(_09571_)
  );
  INV_X1 _19392_ (
    .A(_09571_),
    .ZN(_09572_)
  );
  AND2_X1 _19393_ (
    .A1(_09570_),
    .A2(_09572_),
    .ZN(_09573_)
  );
  INV_X1 _19394_ (
    .A(_09573_),
    .ZN(_09575_)
  );
  AND2_X1 _19395_ (
    .A1(_09562_),
    .A2(_09573_),
    .ZN(_09576_)
  );
  INV_X1 _19396_ (
    .A(_09576_),
    .ZN(_09577_)
  );
  AND2_X1 _19397_ (
    .A1(_09564_),
    .A2(_09575_),
    .ZN(_09578_)
  );
  INV_X1 _19398_ (
    .A(_09578_),
    .ZN(_09579_)
  );
  AND2_X1 _19399_ (
    .A1(_09577_),
    .A2(_09579_),
    .ZN(_09580_)
  );
  INV_X1 _19400_ (
    .A(_09580_),
    .ZN(_09581_)
  );
  AND2_X1 _19401_ (
    .A1(_09560_),
    .A2(_09580_),
    .ZN(_09582_)
  );
  INV_X1 _19402_ (
    .A(_09582_),
    .ZN(_09583_)
  );
  AND2_X1 _19403_ (
    .A1(_09561_),
    .A2(_09581_),
    .ZN(_09584_)
  );
  INV_X1 _19404_ (
    .A(_09584_),
    .ZN(_09586_)
  );
  AND2_X1 _19405_ (
    .A1(_09583_),
    .A2(_09586_),
    .ZN(_09587_)
  );
  INV_X1 _19406_ (
    .A(_09587_),
    .ZN(_09588_)
  );
  AND2_X1 _19407_ (
    .A1(_09264_),
    .A2(_09587_),
    .ZN(_09589_)
  );
  INV_X1 _19408_ (
    .A(_09589_),
    .ZN(_09590_)
  );
  AND2_X1 _19409_ (
    .A1(_09265_),
    .A2(_09588_),
    .ZN(_09591_)
  );
  INV_X1 _19410_ (
    .A(_09591_),
    .ZN(_09592_)
  );
  AND2_X1 _19411_ (
    .A1(_09590_),
    .A2(_09592_),
    .ZN(_09593_)
  );
  INV_X1 _19412_ (
    .A(_09593_),
    .ZN(_09594_)
  );
  AND2_X1 _19413_ (
    .A1(_09458_),
    .A2(_09594_),
    .ZN(_09595_)
  );
  INV_X1 _19414_ (
    .A(_09595_),
    .ZN(_09597_)
  );
  AND2_X1 _19415_ (
    .A1(_09457_),
    .A2(_09593_),
    .ZN(_09598_)
  );
  INV_X1 _19416_ (
    .A(_09598_),
    .ZN(_09599_)
  );
  AND2_X1 _19417_ (
    .A1(_09458_),
    .A2(_09593_),
    .ZN(_09600_)
  );
  INV_X1 _19418_ (
    .A(_09600_),
    .ZN(_09601_)
  );
  AND2_X1 _19419_ (
    .A1(_09457_),
    .A2(_09594_),
    .ZN(_09602_)
  );
  INV_X1 _19420_ (
    .A(_09602_),
    .ZN(_09603_)
  );
  AND2_X1 _19421_ (
    .A1(_09597_),
    .A2(_09599_),
    .ZN(_09604_)
  );
  AND2_X1 _19422_ (
    .A1(_09601_),
    .A2(_09603_),
    .ZN(_09605_)
  );
  AND2_X1 _19423_ (
    .A1(_09540_),
    .A2(_09604_),
    .ZN(_09606_)
  );
  INV_X1 _19424_ (
    .A(_09606_),
    .ZN(_09608_)
  );
  AND2_X1 _19425_ (
    .A1(_09542_),
    .A2(_09605_),
    .ZN(_09609_)
  );
  INV_X1 _19426_ (
    .A(_09609_),
    .ZN(_09610_)
  );
  AND2_X1 _19427_ (
    .A1(_09608_),
    .A2(_09610_),
    .ZN(_09611_)
  );
  INV_X1 _19428_ (
    .A(_09611_),
    .ZN(_09612_)
  );
  AND2_X1 _19429_ (
    .A1(_09462_),
    .A2(_09611_),
    .ZN(_09613_)
  );
  INV_X1 _19430_ (
    .A(_09613_),
    .ZN(_09614_)
  );
  AND2_X1 _19431_ (
    .A1(_09461_),
    .A2(_09612_),
    .ZN(_09615_)
  );
  INV_X1 _19432_ (
    .A(_09615_),
    .ZN(_09616_)
  );
  AND2_X1 _19433_ (
    .A1(_09614_),
    .A2(_09616_),
    .ZN(_09617_)
  );
  INV_X1 _19434_ (
    .A(_09617_),
    .ZN(_09619_)
  );
  AND2_X1 _19435_ (
    .A1(_09318_),
    .A2(_09325_),
    .ZN(_09620_)
  );
  INV_X1 _19436_ (
    .A(_09620_),
    .ZN(_09621_)
  );
  AND2_X1 _19437_ (
    .A1(_09305_),
    .A2(_09312_),
    .ZN(_09622_)
  );
  INV_X1 _19438_ (
    .A(_09622_),
    .ZN(_09623_)
  );
  AND2_X1 _19439_ (
    .A1(_09207_),
    .A2(_09214_),
    .ZN(_09624_)
  );
  INV_X1 _19440_ (
    .A(_09624_),
    .ZN(_09625_)
  );
  AND2_X1 _19441_ (
    .A1(_08674_),
    .A2(_09625_),
    .ZN(_09626_)
  );
  INV_X1 _19442_ (
    .A(_09626_),
    .ZN(_09627_)
  );
  AND2_X1 _19443_ (
    .A1(_08676_),
    .A2(_09624_),
    .ZN(_09628_)
  );
  INV_X1 _19444_ (
    .A(_09628_),
    .ZN(_09630_)
  );
  AND2_X1 _19445_ (
    .A1(_09627_),
    .A2(_09630_),
    .ZN(_09631_)
  );
  INV_X1 _19446_ (
    .A(_09631_),
    .ZN(_09632_)
  );
  AND2_X1 _19447_ (
    .A1(_08999_),
    .A2(_09631_),
    .ZN(_09633_)
  );
  INV_X1 _19448_ (
    .A(_09633_),
    .ZN(_09634_)
  );
  AND2_X1 _19449_ (
    .A1(_08998_),
    .A2(_09632_),
    .ZN(_09635_)
  );
  INV_X1 _19450_ (
    .A(_09635_),
    .ZN(_09636_)
  );
  AND2_X1 _19451_ (
    .A1(_09634_),
    .A2(_09636_),
    .ZN(_09637_)
  );
  INV_X1 _19452_ (
    .A(_09637_),
    .ZN(_09638_)
  );
  AND2_X1 _19453_ (
    .A1(_09623_),
    .A2(_09637_),
    .ZN(_09639_)
  );
  INV_X1 _19454_ (
    .A(_09639_),
    .ZN(_09641_)
  );
  AND2_X1 _19455_ (
    .A1(_09622_),
    .A2(_09638_),
    .ZN(_09642_)
  );
  INV_X1 _19456_ (
    .A(_09642_),
    .ZN(_09643_)
  );
  AND2_X1 _19457_ (
    .A1(_09641_),
    .A2(_09643_),
    .ZN(_09644_)
  );
  INV_X1 _19458_ (
    .A(_09644_),
    .ZN(_09645_)
  );
  AND2_X1 _19459_ (
    .A1(_07082_),
    .A2(_09644_),
    .ZN(_09646_)
  );
  INV_X1 _19460_ (
    .A(_09646_),
    .ZN(_09647_)
  );
  AND2_X1 _19461_ (
    .A1(_07083_),
    .A2(_09645_),
    .ZN(_09648_)
  );
  INV_X1 _19462_ (
    .A(_09648_),
    .ZN(_09649_)
  );
  AND2_X1 _19463_ (
    .A1(_09647_),
    .A2(_09649_),
    .ZN(_09650_)
  );
  INV_X1 _19464_ (
    .A(_09650_),
    .ZN(_09652_)
  );
  AND2_X1 _19465_ (
    .A1(_09226_),
    .A2(_09650_),
    .ZN(_09653_)
  );
  INV_X1 _19466_ (
    .A(_09653_),
    .ZN(_09654_)
  );
  AND2_X1 _19467_ (
    .A1(_09227_),
    .A2(_09652_),
    .ZN(_09655_)
  );
  INV_X1 _19468_ (
    .A(_09655_),
    .ZN(_09656_)
  );
  AND2_X1 _19469_ (
    .A1(_09654_),
    .A2(_09656_),
    .ZN(_09657_)
  );
  INV_X1 _19470_ (
    .A(_09657_),
    .ZN(_09658_)
  );
  AND2_X1 _19471_ (
    .A1(_09621_),
    .A2(_09657_),
    .ZN(_09659_)
  );
  INV_X1 _19472_ (
    .A(_09659_),
    .ZN(_09660_)
  );
  AND2_X1 _19473_ (
    .A1(_09620_),
    .A2(_09658_),
    .ZN(_09661_)
  );
  INV_X1 _19474_ (
    .A(_09661_),
    .ZN(_09663_)
  );
  AND2_X1 _19475_ (
    .A1(_09660_),
    .A2(_09663_),
    .ZN(_09664_)
  );
  INV_X1 _19476_ (
    .A(_09664_),
    .ZN(_09665_)
  );
  AND2_X1 _19477_ (
    .A1(_09617_),
    .A2(_09664_),
    .ZN(_09666_)
  );
  INV_X1 _19478_ (
    .A(_09666_),
    .ZN(_09667_)
  );
  AND2_X1 _19479_ (
    .A1(_09619_),
    .A2(_09665_),
    .ZN(_09668_)
  );
  INV_X1 _19480_ (
    .A(_09668_),
    .ZN(_09669_)
  );
  AND2_X1 _19481_ (
    .A1(_09667_),
    .A2(_09669_),
    .ZN(_09670_)
  );
  INV_X1 _19482_ (
    .A(_09670_),
    .ZN(_09671_)
  );
  AND2_X1 _19483_ (
    .A1(_09456_),
    .A2(_09670_),
    .ZN(_09672_)
  );
  INV_X1 _19484_ (
    .A(_09672_),
    .ZN(_09674_)
  );
  AND2_X1 _19485_ (
    .A1(_09455_),
    .A2(_09671_),
    .ZN(_09675_)
  );
  INV_X1 _19486_ (
    .A(_09675_),
    .ZN(_09676_)
  );
  AND2_X1 _19487_ (
    .A1(_09674_),
    .A2(_09676_),
    .ZN(_09677_)
  );
  INV_X1 _19488_ (
    .A(_09677_),
    .ZN(_09678_)
  );
  AND2_X1 _19489_ (
    .A1(_09331_),
    .A2(_09338_),
    .ZN(_09679_)
  );
  INV_X1 _19490_ (
    .A(_09679_),
    .ZN(_09680_)
  );
  AND2_X1 _19491_ (
    .A1(_07804_),
    .A2(_09680_),
    .ZN(_09681_)
  );
  INV_X1 _19492_ (
    .A(_09681_),
    .ZN(_09682_)
  );
  AND2_X1 _19493_ (
    .A1(_07805_),
    .A2(_09679_),
    .ZN(_09683_)
  );
  INV_X1 _19494_ (
    .A(_09683_),
    .ZN(_09685_)
  );
  AND2_X1 _19495_ (
    .A1(_09682_),
    .A2(_09685_),
    .ZN(_09686_)
  );
  INV_X1 _19496_ (
    .A(_09686_),
    .ZN(_09687_)
  );
  AND2_X1 _19497_ (
    .A1(_08107_),
    .A2(_09686_),
    .ZN(_09688_)
  );
  INV_X1 _19498_ (
    .A(_09688_),
    .ZN(_09689_)
  );
  AND2_X1 _19499_ (
    .A1(_08106_),
    .A2(_09687_),
    .ZN(_09690_)
  );
  INV_X1 _19500_ (
    .A(_09690_),
    .ZN(_09691_)
  );
  AND2_X1 _19501_ (
    .A1(_09689_),
    .A2(_09691_),
    .ZN(_09692_)
  );
  INV_X1 _19502_ (
    .A(_09692_),
    .ZN(_09693_)
  );
  AND2_X1 _19503_ (
    .A1(_09677_),
    .A2(_09692_),
    .ZN(_09694_)
  );
  INV_X1 _19504_ (
    .A(_09694_),
    .ZN(_09696_)
  );
  AND2_X1 _19505_ (
    .A1(_09678_),
    .A2(_09693_),
    .ZN(_09697_)
  );
  INV_X1 _19506_ (
    .A(_09697_),
    .ZN(_09698_)
  );
  AND2_X1 _19507_ (
    .A1(_09696_),
    .A2(_09698_),
    .ZN(_09699_)
  );
  INV_X1 _19508_ (
    .A(_09699_),
    .ZN(_09700_)
  );
  AND2_X1 _19509_ (
    .A1(_09454_),
    .A2(_09699_),
    .ZN(_09701_)
  );
  INV_X1 _19510_ (
    .A(_09701_),
    .ZN(_09702_)
  );
  AND2_X1 _19511_ (
    .A1(_09452_),
    .A2(_09700_),
    .ZN(_09703_)
  );
  INV_X1 _19512_ (
    .A(_09703_),
    .ZN(_09704_)
  );
  AND2_X1 _19513_ (
    .A1(_09702_),
    .A2(_09704_),
    .ZN(_09705_)
  );
  INV_X1 _19514_ (
    .A(_09705_),
    .ZN(_09707_)
  );
  AND2_X1 _19515_ (
    .A1(_09451_),
    .A2(_09705_),
    .ZN(_09708_)
  );
  INV_X1 _19516_ (
    .A(_09708_),
    .ZN(_09709_)
  );
  AND2_X1 _19517_ (
    .A1(_09450_),
    .A2(_09707_),
    .ZN(_09710_)
  );
  INV_X1 _19518_ (
    .A(_09710_),
    .ZN(_09711_)
  );
  AND2_X1 _19519_ (
    .A1(_09709_),
    .A2(_09711_),
    .ZN(_09712_)
  );
  INV_X1 _19520_ (
    .A(_09712_),
    .ZN(_09713_)
  );
  AND2_X1 _19521_ (
    .A1(_09449_),
    .A2(_09712_),
    .ZN(_09714_)
  );
  INV_X1 _19522_ (
    .A(_09714_),
    .ZN(_09715_)
  );
  AND2_X1 _19523_ (
    .A1(_09448_),
    .A2(_09713_),
    .ZN(_09716_)
  );
  INV_X1 _19524_ (
    .A(_09716_),
    .ZN(_09718_)
  );
  AND2_X1 _19525_ (
    .A1(_09715_),
    .A2(_09718_),
    .ZN(_09719_)
  );
  INV_X1 _19526_ (
    .A(_09719_),
    .ZN(_09720_)
  );
  AND2_X1 _19527_ (
    .A1(_09392_),
    .A2(_09719_),
    .ZN(_09721_)
  );
  INV_X1 _19528_ (
    .A(_09721_),
    .ZN(_09722_)
  );
  AND2_X1 _19529_ (
    .A1(_09393_),
    .A2(_09720_),
    .ZN(_09723_)
  );
  INV_X1 _19530_ (
    .A(_09723_),
    .ZN(_09724_)
  );
  AND2_X1 _19531_ (
    .A1(_09722_),
    .A2(_09724_),
    .ZN(_09725_)
  );
  INV_X1 _19532_ (
    .A(_09725_),
    .ZN(_09726_)
  );
  AND2_X1 _19533_ (
    .A1(_09446_),
    .A2(_09726_),
    .ZN(_09727_)
  );
  INV_X1 _19534_ (
    .A(_09727_),
    .ZN(_09729_)
  );
  AND2_X1 _19535_ (
    .A1(_09447_),
    .A2(_09725_),
    .ZN(_09730_)
  );
  INV_X1 _19536_ (
    .A(_09730_),
    .ZN(_09731_)
  );
  AND2_X1 _19537_ (
    .A1(_09729_),
    .A2(_09731_),
    .ZN(_09732_)
  );
  INV_X1 _19538_ (
    .A(_09732_),
    .ZN(_09733_)
  );
  AND2_X1 _19539_ (
    .A1(_04404_),
    .A2(_09733_),
    .ZN(_09734_)
  );
  INV_X1 _19540_ (
    .A(_09734_),
    .ZN(_09735_)
  );
  AND2_X1 _19541_ (
    .A1(remainder[65]),
    .A2(_09732_),
    .ZN(_09736_)
  );
  INV_X1 _19542_ (
    .A(_09736_),
    .ZN(_09737_)
  );
  AND2_X1 _19543_ (
    .A1(_09735_),
    .A2(_09737_),
    .ZN(_09738_)
  );
  INV_X1 _19544_ (
    .A(_09738_),
    .ZN(_09740_)
  );
  AND2_X1 _19545_ (
    .A1(_09444_),
    .A2(_09740_),
    .ZN(_09741_)
  );
  INV_X1 _19546_ (
    .A(_09741_),
    .ZN(_09742_)
  );
  AND2_X1 _19547_ (
    .A1(_09445_),
    .A2(_09738_),
    .ZN(_09743_)
  );
  INV_X1 _19548_ (
    .A(_09743_),
    .ZN(_09744_)
  );
  AND2_X1 _19549_ (
    .A1(_09742_),
    .A2(_09744_),
    .ZN(_09745_)
  );
  AND2_X1 _19550_ (
    .A1(_02082_),
    .A2(_09745_),
    .ZN(_09746_)
  );
  INV_X1 _19551_ (
    .A(_09746_),
    .ZN(_09747_)
  );
  AND2_X1 _19552_ (
    .A1(remainder[58]),
    .A2(_02077_),
    .ZN(_09748_)
  );
  INV_X1 _19553_ (
    .A(_09748_),
    .ZN(_09749_)
  );
  MUX2_X1 _19554_ (
    .A(remainder[57]),
    .B(_01979_),
    .S(_10462_),
    .Z(_09751_)
  );
  AND2_X1 _19555_ (
    .A1(_05983_),
    .A2(_09751_),
    .ZN(_09752_)
  );
  INV_X1 _19556_ (
    .A(_09752_),
    .ZN(_09753_)
  );
  AND2_X1 _19557_ (
    .A1(_09749_),
    .A2(_09753_),
    .ZN(_09754_)
  );
  AND2_X1 _19558_ (
    .A1(_09747_),
    .A2(_09754_),
    .ZN(_09755_)
  );
  INV_X1 _19559_ (
    .A(_09755_),
    .ZN(_09756_)
  );
  AND2_X1 _19560_ (
    .A1(_06201_),
    .A2(_09756_),
    .ZN(_00079_)
  );
  AND2_X1 _19561_ (
    .A1(_09423_),
    .A2(_09738_),
    .ZN(_09757_)
  );
  INV_X1 _19562_ (
    .A(_09757_),
    .ZN(_09758_)
  );
  AND2_X1 _19563_ (
    .A1(_09417_),
    .A2(_09737_),
    .ZN(_09759_)
  );
  AND2_X1 _19564_ (
    .A1(_09758_),
    .A2(_09759_),
    .ZN(_09761_)
  );
  INV_X1 _19565_ (
    .A(_09761_),
    .ZN(_09762_)
  );
  AND2_X1 _19566_ (
    .A1(_09702_),
    .A2(_09709_),
    .ZN(_09763_)
  );
  INV_X1 _19567_ (
    .A(_09763_),
    .ZN(_09764_)
  );
  AND2_X1 _19568_ (
    .A1(_09682_),
    .A2(_09689_),
    .ZN(_09765_)
  );
  INV_X1 _19569_ (
    .A(_09765_),
    .ZN(_09766_)
  );
  AND2_X1 _19570_ (
    .A1(_09674_),
    .A2(_09696_),
    .ZN(_09767_)
  );
  INV_X1 _19571_ (
    .A(_09767_),
    .ZN(_09768_)
  );
  AND2_X1 _19572_ (
    .A1(_09614_),
    .A2(_09667_),
    .ZN(_09769_)
  );
  INV_X1 _19573_ (
    .A(_09769_),
    .ZN(_09770_)
  );
  AND2_X1 _19574_ (
    .A1(_03249_),
    .A2(_09275_),
    .ZN(_09772_)
  );
  AND2_X1 _19575_ (
    .A1(_09594_),
    .A2(_09772_),
    .ZN(_09773_)
  );
  INV_X1 _19576_ (
    .A(_09773_),
    .ZN(_09774_)
  );
  AND2_X1 _19577_ (
    .A1(_09608_),
    .A2(_09774_),
    .ZN(_09775_)
  );
  INV_X1 _19578_ (
    .A(_09775_),
    .ZN(_09776_)
  );
  AND2_X1 _19579_ (
    .A1(_03249_),
    .A2(_09593_),
    .ZN(_09777_)
  );
  INV_X1 _19580_ (
    .A(_09777_),
    .ZN(_09778_)
  );
  AND2_X1 _19581_ (
    .A1(_03249_),
    .A2(_09232_),
    .ZN(_09779_)
  );
  INV_X1 _19582_ (
    .A(_09779_),
    .ZN(_09780_)
  );
  AND2_X1 _19583_ (
    .A1(_03250_),
    .A2(_09233_),
    .ZN(_09781_)
  );
  INV_X1 _19584_ (
    .A(_09781_),
    .ZN(_09783_)
  );
  AND2_X1 _19585_ (
    .A1(_09780_),
    .A2(_09783_),
    .ZN(_09784_)
  );
  INV_X1 _19586_ (
    .A(_09784_),
    .ZN(_09785_)
  );
  AND2_X1 _19587_ (
    .A1(_09557_),
    .A2(_09583_),
    .ZN(_09786_)
  );
  INV_X1 _19588_ (
    .A(_09786_),
    .ZN(_09787_)
  );
  AND2_X1 _19589_ (
    .A1(_09546_),
    .A2(_09550_),
    .ZN(_09788_)
  );
  INV_X1 _19590_ (
    .A(_09788_),
    .ZN(_09789_)
  );
  AND2_X1 _19591_ (
    .A1(divisor[31]),
    .A2(remainder[3]),
    .ZN(_09790_)
  );
  INV_X1 _19592_ (
    .A(_09790_),
    .ZN(_09791_)
  );
  AND2_X1 _19593_ (
    .A1(divisor[32]),
    .A2(remainder[2]),
    .ZN(_09792_)
  );
  INV_X1 _19594_ (
    .A(_09792_),
    .ZN(_09794_)
  );
  AND2_X1 _19595_ (
    .A1(remainder[1]),
    .A2(_09792_),
    .ZN(_09795_)
  );
  INV_X1 _19596_ (
    .A(_09795_),
    .ZN(_09796_)
  );
  MUX2_X1 _19597_ (
    .A(_09792_),
    .B(_05095_),
    .S(_09237_),
    .Z(_09797_)
  );
  MUX2_X1 _19598_ (
    .A(_09794_),
    .B(remainder[2]),
    .S(_09237_),
    .Z(_09798_)
  );
  AND2_X1 _19599_ (
    .A1(_09790_),
    .A2(_09797_),
    .ZN(_09799_)
  );
  INV_X1 _19600_ (
    .A(_09799_),
    .ZN(_09800_)
  );
  AND2_X1 _19601_ (
    .A1(_09791_),
    .A2(_09798_),
    .ZN(_09801_)
  );
  INV_X1 _19602_ (
    .A(_09801_),
    .ZN(_09802_)
  );
  AND2_X1 _19603_ (
    .A1(_09800_),
    .A2(_09802_),
    .ZN(_09803_)
  );
  INV_X1 _19604_ (
    .A(_09803_),
    .ZN(_09805_)
  );
  AND2_X1 _19605_ (
    .A1(_09789_),
    .A2(_09803_),
    .ZN(_09806_)
  );
  INV_X1 _19606_ (
    .A(_09806_),
    .ZN(_09807_)
  );
  AND2_X1 _19607_ (
    .A1(_09788_),
    .A2(_09805_),
    .ZN(_09808_)
  );
  INV_X1 _19608_ (
    .A(_09808_),
    .ZN(_09809_)
  );
  AND2_X1 _19609_ (
    .A1(_09807_),
    .A2(_09809_),
    .ZN(_09810_)
  );
  INV_X1 _19610_ (
    .A(_09810_),
    .ZN(_09811_)
  );
  AND2_X1 _19611_ (
    .A1(divisor[28]),
    .A2(remainder[6]),
    .ZN(_09812_)
  );
  INV_X1 _19612_ (
    .A(_09812_),
    .ZN(_09813_)
  );
  AND2_X1 _19613_ (
    .A1(divisor[29]),
    .A2(remainder[5]),
    .ZN(_09814_)
  );
  INV_X1 _19614_ (
    .A(_09814_),
    .ZN(_09816_)
  );
  AND2_X1 _19615_ (
    .A1(divisor[30]),
    .A2(remainder[5]),
    .ZN(_09817_)
  );
  INV_X1 _19616_ (
    .A(_09817_),
    .ZN(_09818_)
  );
  AND2_X1 _19617_ (
    .A1(_09567_),
    .A2(_09814_),
    .ZN(_09819_)
  );
  INV_X1 _19618_ (
    .A(_09819_),
    .ZN(_09820_)
  );
  AND2_X1 _19619_ (
    .A1(_09568_),
    .A2(_09816_),
    .ZN(_09821_)
  );
  INV_X1 _19620_ (
    .A(_09821_),
    .ZN(_09822_)
  );
  AND2_X1 _19621_ (
    .A1(_09820_),
    .A2(_09822_),
    .ZN(_09823_)
  );
  INV_X1 _19622_ (
    .A(_09823_),
    .ZN(_09824_)
  );
  AND2_X1 _19623_ (
    .A1(_09812_),
    .A2(_09823_),
    .ZN(_09825_)
  );
  INV_X1 _19624_ (
    .A(_09825_),
    .ZN(_09827_)
  );
  AND2_X1 _19625_ (
    .A1(_09813_),
    .A2(_09824_),
    .ZN(_09828_)
  );
  INV_X1 _19626_ (
    .A(_09828_),
    .ZN(_09829_)
  );
  AND2_X1 _19627_ (
    .A1(_09827_),
    .A2(_09829_),
    .ZN(_09830_)
  );
  INV_X1 _19628_ (
    .A(_09830_),
    .ZN(_09831_)
  );
  AND2_X1 _19629_ (
    .A1(_09810_),
    .A2(_09830_),
    .ZN(_09832_)
  );
  INV_X1 _19630_ (
    .A(_09832_),
    .ZN(_09833_)
  );
  AND2_X1 _19631_ (
    .A1(_09811_),
    .A2(_09831_),
    .ZN(_09834_)
  );
  INV_X1 _19632_ (
    .A(_09834_),
    .ZN(_09835_)
  );
  AND2_X1 _19633_ (
    .A1(_09833_),
    .A2(_09835_),
    .ZN(_09836_)
  );
  INV_X1 _19634_ (
    .A(_09836_),
    .ZN(_09838_)
  );
  AND2_X1 _19635_ (
    .A1(_09787_),
    .A2(_09836_),
    .ZN(_09839_)
  );
  INV_X1 _19636_ (
    .A(_09839_),
    .ZN(_09840_)
  );
  AND2_X1 _19637_ (
    .A1(_09786_),
    .A2(_09838_),
    .ZN(_09841_)
  );
  INV_X1 _19638_ (
    .A(_09841_),
    .ZN(_09842_)
  );
  AND2_X1 _19639_ (
    .A1(_09840_),
    .A2(_09842_),
    .ZN(_09843_)
  );
  INV_X1 _19640_ (
    .A(_09843_),
    .ZN(_09844_)
  );
  AND2_X1 _19641_ (
    .A1(_09784_),
    .A2(_09843_),
    .ZN(_09845_)
  );
  INV_X1 _19642_ (
    .A(_09845_),
    .ZN(_09846_)
  );
  AND2_X1 _19643_ (
    .A1(_09785_),
    .A2(_09844_),
    .ZN(_09847_)
  );
  INV_X1 _19644_ (
    .A(_09847_),
    .ZN(_09849_)
  );
  AND2_X1 _19645_ (
    .A1(_09846_),
    .A2(_09849_),
    .ZN(_09850_)
  );
  INV_X1 _19646_ (
    .A(_09850_),
    .ZN(_09851_)
  );
  AND2_X1 _19647_ (
    .A1(_09777_),
    .A2(_09850_),
    .ZN(_09852_)
  );
  INV_X1 _19648_ (
    .A(_09852_),
    .ZN(_09853_)
  );
  AND2_X1 _19649_ (
    .A1(_09778_),
    .A2(_09851_),
    .ZN(_09854_)
  );
  INV_X1 _19650_ (
    .A(_09854_),
    .ZN(_09855_)
  );
  AND2_X1 _19651_ (
    .A1(_09853_),
    .A2(_09855_),
    .ZN(_09856_)
  );
  INV_X1 _19652_ (
    .A(_09856_),
    .ZN(_09857_)
  );
  AND2_X1 _19653_ (
    .A1(_09506_),
    .A2(_09524_),
    .ZN(_09858_)
  );
  INV_X1 _19654_ (
    .A(_09858_),
    .ZN(_09860_)
  );
  AND2_X1 _19655_ (
    .A1(_09493_),
    .A2(_09500_),
    .ZN(_09861_)
  );
  INV_X1 _19656_ (
    .A(_09861_),
    .ZN(_09862_)
  );
  AND2_X1 _19657_ (
    .A1(_09480_),
    .A2(_09487_),
    .ZN(_09863_)
  );
  INV_X1 _19658_ (
    .A(_09863_),
    .ZN(_09864_)
  );
  AND2_X1 _19659_ (
    .A1(_09570_),
    .A2(_09577_),
    .ZN(_09865_)
  );
  INV_X1 _19660_ (
    .A(_09865_),
    .ZN(_09866_)
  );
  AND2_X1 _19661_ (
    .A1(remainder[32]),
    .A2(divisor[27]),
    .ZN(_09867_)
  );
  AND2_X1 _19662_ (
    .A1(remainder[32]),
    .A2(divisor[26]),
    .ZN(_09868_)
  );
  INV_X1 _19663_ (
    .A(_09868_),
    .ZN(_09869_)
  );
  AND2_X1 _19664_ (
    .A1(divisor[27]),
    .A2(_09868_),
    .ZN(_09871_)
  );
  INV_X1 _19665_ (
    .A(_09871_),
    .ZN(_09872_)
  );
  AND2_X1 _19666_ (
    .A1(_09477_),
    .A2(_09868_),
    .ZN(_09873_)
  );
  INV_X1 _19667_ (
    .A(_09873_),
    .ZN(_09874_)
  );
  AND2_X1 _19668_ (
    .A1(_09478_),
    .A2(_09869_),
    .ZN(_09875_)
  );
  INV_X1 _19669_ (
    .A(_09875_),
    .ZN(_09876_)
  );
  AND2_X1 _19670_ (
    .A1(_09874_),
    .A2(_09876_),
    .ZN(_09877_)
  );
  INV_X1 _19671_ (
    .A(_09877_),
    .ZN(_09878_)
  );
  AND2_X1 _19672_ (
    .A1(_09472_),
    .A2(_09877_),
    .ZN(_09879_)
  );
  INV_X1 _19673_ (
    .A(_09879_),
    .ZN(_09880_)
  );
  AND2_X1 _19674_ (
    .A1(_09473_),
    .A2(_09878_),
    .ZN(_09882_)
  );
  INV_X1 _19675_ (
    .A(_09882_),
    .ZN(_09883_)
  );
  AND2_X1 _19676_ (
    .A1(_09880_),
    .A2(_09883_),
    .ZN(_09884_)
  );
  INV_X1 _19677_ (
    .A(_09884_),
    .ZN(_09885_)
  );
  AND2_X1 _19678_ (
    .A1(_09866_),
    .A2(_09884_),
    .ZN(_09886_)
  );
  INV_X1 _19679_ (
    .A(_09886_),
    .ZN(_09887_)
  );
  AND2_X1 _19680_ (
    .A1(_09865_),
    .A2(_09885_),
    .ZN(_09888_)
  );
  INV_X1 _19681_ (
    .A(_09888_),
    .ZN(_09889_)
  );
  AND2_X1 _19682_ (
    .A1(_09887_),
    .A2(_09889_),
    .ZN(_09890_)
  );
  INV_X1 _19683_ (
    .A(_09890_),
    .ZN(_09891_)
  );
  AND2_X1 _19684_ (
    .A1(_09864_),
    .A2(_09890_),
    .ZN(_09893_)
  );
  INV_X1 _19685_ (
    .A(_09893_),
    .ZN(_09894_)
  );
  AND2_X1 _19686_ (
    .A1(_09863_),
    .A2(_09891_),
    .ZN(_09895_)
  );
  INV_X1 _19687_ (
    .A(_09895_),
    .ZN(_09896_)
  );
  AND2_X1 _19688_ (
    .A1(_09894_),
    .A2(_09896_),
    .ZN(_09897_)
  );
  INV_X1 _19689_ (
    .A(_09897_),
    .ZN(_09898_)
  );
  AND2_X1 _19690_ (
    .A1(_09862_),
    .A2(_09897_),
    .ZN(_09899_)
  );
  INV_X1 _19691_ (
    .A(_09899_),
    .ZN(_09900_)
  );
  AND2_X1 _19692_ (
    .A1(_09861_),
    .A2(_09898_),
    .ZN(_09901_)
  );
  INV_X1 _19693_ (
    .A(_09901_),
    .ZN(_09902_)
  );
  AND2_X1 _19694_ (
    .A1(_09900_),
    .A2(_09902_),
    .ZN(_09904_)
  );
  INV_X1 _19695_ (
    .A(_09904_),
    .ZN(_09905_)
  );
  AND2_X1 _19696_ (
    .A1(_09521_),
    .A2(_09904_),
    .ZN(_09906_)
  );
  INV_X1 _19697_ (
    .A(_09906_),
    .ZN(_09907_)
  );
  AND2_X1 _19698_ (
    .A1(_09522_),
    .A2(_09905_),
    .ZN(_09908_)
  );
  INV_X1 _19699_ (
    .A(_09908_),
    .ZN(_09909_)
  );
  AND2_X1 _19700_ (
    .A1(_09907_),
    .A2(_09909_),
    .ZN(_09910_)
  );
  INV_X1 _19701_ (
    .A(_09910_),
    .ZN(_09911_)
  );
  AND2_X1 _19702_ (
    .A1(_09589_),
    .A2(_09910_),
    .ZN(_09912_)
  );
  INV_X1 _19703_ (
    .A(_09912_),
    .ZN(_09913_)
  );
  AND2_X1 _19704_ (
    .A1(_09590_),
    .A2(_09911_),
    .ZN(_09915_)
  );
  INV_X1 _19705_ (
    .A(_09915_),
    .ZN(_09916_)
  );
  AND2_X1 _19706_ (
    .A1(_09913_),
    .A2(_09916_),
    .ZN(_09917_)
  );
  INV_X1 _19707_ (
    .A(_09917_),
    .ZN(_09918_)
  );
  AND2_X1 _19708_ (
    .A1(_09860_),
    .A2(_09917_),
    .ZN(_09919_)
  );
  INV_X1 _19709_ (
    .A(_09919_),
    .ZN(_09920_)
  );
  AND2_X1 _19710_ (
    .A1(_09858_),
    .A2(_09918_),
    .ZN(_09921_)
  );
  INV_X1 _19711_ (
    .A(_09921_),
    .ZN(_09922_)
  );
  AND2_X1 _19712_ (
    .A1(_09920_),
    .A2(_09922_),
    .ZN(_09923_)
  );
  INV_X1 _19713_ (
    .A(_09923_),
    .ZN(_09924_)
  );
  AND2_X1 _19714_ (
    .A1(_09856_),
    .A2(_09923_),
    .ZN(_09926_)
  );
  INV_X1 _19715_ (
    .A(_09926_),
    .ZN(_09927_)
  );
  AND2_X1 _19716_ (
    .A1(_09857_),
    .A2(_09924_),
    .ZN(_09928_)
  );
  INV_X1 _19717_ (
    .A(_09928_),
    .ZN(_09929_)
  );
  AND2_X1 _19718_ (
    .A1(_09927_),
    .A2(_09929_),
    .ZN(_09930_)
  );
  INV_X1 _19719_ (
    .A(_09930_),
    .ZN(_09931_)
  );
  AND2_X1 _19720_ (
    .A1(_09776_),
    .A2(_09930_),
    .ZN(_09932_)
  );
  INV_X1 _19721_ (
    .A(_09932_),
    .ZN(_09933_)
  );
  AND2_X1 _19722_ (
    .A1(_09775_),
    .A2(_09931_),
    .ZN(_09934_)
  );
  INV_X1 _19723_ (
    .A(_09934_),
    .ZN(_09935_)
  );
  AND2_X1 _19724_ (
    .A1(_09933_),
    .A2(_09935_),
    .ZN(_09937_)
  );
  INV_X1 _19725_ (
    .A(_09937_),
    .ZN(_09938_)
  );
  AND2_X1 _19726_ (
    .A1(_09641_),
    .A2(_09647_),
    .ZN(_09939_)
  );
  INV_X1 _19727_ (
    .A(_09939_),
    .ZN(_09940_)
  );
  AND2_X1 _19728_ (
    .A1(_09531_),
    .A2(_09537_),
    .ZN(_09941_)
  );
  INV_X1 _19729_ (
    .A(_09941_),
    .ZN(_09942_)
  );
  AND2_X1 _19730_ (
    .A1(_09627_),
    .A2(_09634_),
    .ZN(_09943_)
  );
  INV_X1 _19731_ (
    .A(_09943_),
    .ZN(_09944_)
  );
  AND2_X1 _19732_ (
    .A1(_09207_),
    .A2(_09517_),
    .ZN(_09945_)
  );
  INV_X1 _19733_ (
    .A(_09945_),
    .ZN(_09946_)
  );
  AND2_X1 _19734_ (
    .A1(_08674_),
    .A2(_09946_),
    .ZN(_09948_)
  );
  INV_X1 _19735_ (
    .A(_09948_),
    .ZN(_09949_)
  );
  AND2_X1 _19736_ (
    .A1(_08676_),
    .A2(_09945_),
    .ZN(_09950_)
  );
  INV_X1 _19737_ (
    .A(_09950_),
    .ZN(_09951_)
  );
  AND2_X1 _19738_ (
    .A1(_09949_),
    .A2(_09951_),
    .ZN(_09952_)
  );
  INV_X1 _19739_ (
    .A(_09952_),
    .ZN(_09953_)
  );
  AND2_X1 _19740_ (
    .A1(_08998_),
    .A2(_09953_),
    .ZN(_09954_)
  );
  INV_X1 _19741_ (
    .A(_09954_),
    .ZN(_09955_)
  );
  AND2_X1 _19742_ (
    .A1(_08999_),
    .A2(_09952_),
    .ZN(_09956_)
  );
  INV_X1 _19743_ (
    .A(_09956_),
    .ZN(_09957_)
  );
  AND2_X1 _19744_ (
    .A1(_08998_),
    .A2(_09952_),
    .ZN(_09959_)
  );
  INV_X1 _19745_ (
    .A(_09959_),
    .ZN(_09960_)
  );
  AND2_X1 _19746_ (
    .A1(_08999_),
    .A2(_09953_),
    .ZN(_09961_)
  );
  INV_X1 _19747_ (
    .A(_09961_),
    .ZN(_09962_)
  );
  AND2_X1 _19748_ (
    .A1(_09955_),
    .A2(_09957_),
    .ZN(_09963_)
  );
  AND2_X1 _19749_ (
    .A1(_09960_),
    .A2(_09962_),
    .ZN(_09964_)
  );
  AND2_X1 _19750_ (
    .A1(_09944_),
    .A2(_09963_),
    .ZN(_09965_)
  );
  INV_X1 _19751_ (
    .A(_09965_),
    .ZN(_09966_)
  );
  AND2_X1 _19752_ (
    .A1(_09943_),
    .A2(_09964_),
    .ZN(_09967_)
  );
  INV_X1 _19753_ (
    .A(_09967_),
    .ZN(_09968_)
  );
  AND2_X1 _19754_ (
    .A1(_09966_),
    .A2(_09968_),
    .ZN(_09970_)
  );
  INV_X1 _19755_ (
    .A(_09970_),
    .ZN(_09971_)
  );
  AND2_X1 _19756_ (
    .A1(_07082_),
    .A2(_09970_),
    .ZN(_09972_)
  );
  INV_X1 _19757_ (
    .A(_09972_),
    .ZN(_09973_)
  );
  AND2_X1 _19758_ (
    .A1(_07083_),
    .A2(_09971_),
    .ZN(_09974_)
  );
  INV_X1 _19759_ (
    .A(_09974_),
    .ZN(_09975_)
  );
  AND2_X1 _19760_ (
    .A1(_09973_),
    .A2(_09975_),
    .ZN(_09976_)
  );
  INV_X1 _19761_ (
    .A(_09976_),
    .ZN(_09977_)
  );
  AND2_X1 _19762_ (
    .A1(_09942_),
    .A2(_09976_),
    .ZN(_09978_)
  );
  INV_X1 _19763_ (
    .A(_09978_),
    .ZN(_09979_)
  );
  AND2_X1 _19764_ (
    .A1(_09941_),
    .A2(_09977_),
    .ZN(_09981_)
  );
  INV_X1 _19765_ (
    .A(_09981_),
    .ZN(_09982_)
  );
  AND2_X1 _19766_ (
    .A1(_09979_),
    .A2(_09982_),
    .ZN(_09983_)
  );
  INV_X1 _19767_ (
    .A(_09983_),
    .ZN(_09984_)
  );
  AND2_X1 _19768_ (
    .A1(_09940_),
    .A2(_09983_),
    .ZN(_09985_)
  );
  INV_X1 _19769_ (
    .A(_09985_),
    .ZN(_09986_)
  );
  AND2_X1 _19770_ (
    .A1(_09939_),
    .A2(_09984_),
    .ZN(_09987_)
  );
  INV_X1 _19771_ (
    .A(_09987_),
    .ZN(_09988_)
  );
  AND2_X1 _19772_ (
    .A1(_09986_),
    .A2(_09988_),
    .ZN(_09989_)
  );
  INV_X1 _19773_ (
    .A(_09989_),
    .ZN(_09990_)
  );
  AND2_X1 _19774_ (
    .A1(_09937_),
    .A2(_09989_),
    .ZN(_09992_)
  );
  INV_X1 _19775_ (
    .A(_09992_),
    .ZN(_09993_)
  );
  AND2_X1 _19776_ (
    .A1(_09938_),
    .A2(_09990_),
    .ZN(_09994_)
  );
  INV_X1 _19777_ (
    .A(_09994_),
    .ZN(_09995_)
  );
  AND2_X1 _19778_ (
    .A1(_09993_),
    .A2(_09995_),
    .ZN(_09996_)
  );
  INV_X1 _19779_ (
    .A(_09996_),
    .ZN(_09997_)
  );
  AND2_X1 _19780_ (
    .A1(_09770_),
    .A2(_09996_),
    .ZN(_09998_)
  );
  INV_X1 _19781_ (
    .A(_09998_),
    .ZN(_09999_)
  );
  AND2_X1 _19782_ (
    .A1(_09769_),
    .A2(_09997_),
    .ZN(_10000_)
  );
  INV_X1 _19783_ (
    .A(_10000_),
    .ZN(_10001_)
  );
  AND2_X1 _19784_ (
    .A1(_09999_),
    .A2(_10001_),
    .ZN(_10003_)
  );
  INV_X1 _19785_ (
    .A(_10003_),
    .ZN(_10004_)
  );
  AND2_X1 _19786_ (
    .A1(_09654_),
    .A2(_09660_),
    .ZN(_10005_)
  );
  INV_X1 _19787_ (
    .A(_10005_),
    .ZN(_10006_)
  );
  AND2_X1 _19788_ (
    .A1(_07804_),
    .A2(_10006_),
    .ZN(_10007_)
  );
  INV_X1 _19789_ (
    .A(_10007_),
    .ZN(_10008_)
  );
  AND2_X1 _19790_ (
    .A1(_07805_),
    .A2(_10005_),
    .ZN(_10009_)
  );
  INV_X1 _19791_ (
    .A(_10009_),
    .ZN(_10010_)
  );
  AND2_X1 _19792_ (
    .A1(_10008_),
    .A2(_10010_),
    .ZN(_10011_)
  );
  INV_X1 _19793_ (
    .A(_10011_),
    .ZN(_10012_)
  );
  AND2_X1 _19794_ (
    .A1(_08107_),
    .A2(_10011_),
    .ZN(_10014_)
  );
  INV_X1 _19795_ (
    .A(_10014_),
    .ZN(_10015_)
  );
  AND2_X1 _19796_ (
    .A1(_08106_),
    .A2(_10012_),
    .ZN(_10016_)
  );
  INV_X1 _19797_ (
    .A(_10016_),
    .ZN(_10017_)
  );
  AND2_X1 _19798_ (
    .A1(_10015_),
    .A2(_10017_),
    .ZN(_10018_)
  );
  INV_X1 _19799_ (
    .A(_10018_),
    .ZN(_10019_)
  );
  AND2_X1 _19800_ (
    .A1(_10003_),
    .A2(_10018_),
    .ZN(_10020_)
  );
  INV_X1 _19801_ (
    .A(_10020_),
    .ZN(_10021_)
  );
  AND2_X1 _19802_ (
    .A1(_10004_),
    .A2(_10019_),
    .ZN(_10022_)
  );
  INV_X1 _19803_ (
    .A(_10022_),
    .ZN(_10023_)
  );
  AND2_X1 _19804_ (
    .A1(_10021_),
    .A2(_10023_),
    .ZN(_10025_)
  );
  INV_X1 _19805_ (
    .A(_10025_),
    .ZN(_10026_)
  );
  AND2_X1 _19806_ (
    .A1(_09768_),
    .A2(_10025_),
    .ZN(_10027_)
  );
  INV_X1 _19807_ (
    .A(_10027_),
    .ZN(_10028_)
  );
  AND2_X1 _19808_ (
    .A1(_09767_),
    .A2(_10026_),
    .ZN(_10029_)
  );
  INV_X1 _19809_ (
    .A(_10029_),
    .ZN(_10030_)
  );
  AND2_X1 _19810_ (
    .A1(_10028_),
    .A2(_10030_),
    .ZN(_10031_)
  );
  INV_X1 _19811_ (
    .A(_10031_),
    .ZN(_10032_)
  );
  AND2_X1 _19812_ (
    .A1(_09766_),
    .A2(_10031_),
    .ZN(_10033_)
  );
  INV_X1 _19813_ (
    .A(_10033_),
    .ZN(_10034_)
  );
  AND2_X1 _19814_ (
    .A1(_09765_),
    .A2(_10032_),
    .ZN(_10036_)
  );
  INV_X1 _19815_ (
    .A(_10036_),
    .ZN(_10037_)
  );
  AND2_X1 _19816_ (
    .A1(_10034_),
    .A2(_10037_),
    .ZN(_10038_)
  );
  INV_X1 _19817_ (
    .A(_10038_),
    .ZN(_10039_)
  );
  AND2_X1 _19818_ (
    .A1(_09764_),
    .A2(_10038_),
    .ZN(_10040_)
  );
  INV_X1 _19819_ (
    .A(_10040_),
    .ZN(_10041_)
  );
  AND2_X1 _19820_ (
    .A1(_09763_),
    .A2(_10039_),
    .ZN(_10042_)
  );
  INV_X1 _19821_ (
    .A(_10042_),
    .ZN(_10043_)
  );
  AND2_X1 _19822_ (
    .A1(_10041_),
    .A2(_10043_),
    .ZN(_10044_)
  );
  INV_X1 _19823_ (
    .A(_10044_),
    .ZN(_10045_)
  );
  AND2_X1 _19824_ (
    .A1(_09714_),
    .A2(_10044_),
    .ZN(_10047_)
  );
  INV_X1 _19825_ (
    .A(_10047_),
    .ZN(_10048_)
  );
  AND2_X1 _19826_ (
    .A1(_09715_),
    .A2(_10045_),
    .ZN(_10049_)
  );
  INV_X1 _19827_ (
    .A(_10049_),
    .ZN(_10050_)
  );
  AND2_X1 _19828_ (
    .A1(_10048_),
    .A2(_10050_),
    .ZN(_10051_)
  );
  INV_X1 _19829_ (
    .A(_10051_),
    .ZN(_10052_)
  );
  AND2_X1 _19830_ (
    .A1(_09446_),
    .A2(_09722_),
    .ZN(_10053_)
  );
  INV_X1 _19831_ (
    .A(_10053_),
    .ZN(_10054_)
  );
  AND2_X1 _19832_ (
    .A1(_09724_),
    .A2(_10054_),
    .ZN(_10055_)
  );
  AND2_X1 _19833_ (
    .A1(_09722_),
    .A2(_09731_),
    .ZN(_10056_)
  );
  AND2_X1 _19834_ (
    .A1(_10051_),
    .A2(_10055_),
    .ZN(_10058_)
  );
  INV_X1 _19835_ (
    .A(_10058_),
    .ZN(_10059_)
  );
  AND2_X1 _19836_ (
    .A1(_10052_),
    .A2(_10056_),
    .ZN(_10060_)
  );
  INV_X1 _19837_ (
    .A(_10060_),
    .ZN(_10061_)
  );
  AND2_X1 _19838_ (
    .A1(_10059_),
    .A2(_10061_),
    .ZN(_10062_)
  );
  INV_X1 _19839_ (
    .A(_10062_),
    .ZN(_10063_)
  );
  AND2_X1 _19840_ (
    .A1(remainder[65]),
    .A2(_10062_),
    .ZN(_10064_)
  );
  INV_X1 _19841_ (
    .A(_10064_),
    .ZN(_10065_)
  );
  AND2_X1 _19842_ (
    .A1(_04404_),
    .A2(_10063_),
    .ZN(_10066_)
  );
  INV_X1 _19843_ (
    .A(_10066_),
    .ZN(_10067_)
  );
  AND2_X1 _19844_ (
    .A1(_10065_),
    .A2(_10067_),
    .ZN(_10069_)
  );
  INV_X1 _19845_ (
    .A(_10069_),
    .ZN(_10070_)
  );
  AND2_X1 _19846_ (
    .A1(_09762_),
    .A2(_10069_),
    .ZN(_10071_)
  );
  INV_X1 _19847_ (
    .A(_10071_),
    .ZN(_10072_)
  );
  AND2_X1 _19848_ (
    .A1(_09761_),
    .A2(_10070_),
    .ZN(_10073_)
  );
  INV_X1 _19849_ (
    .A(_10073_),
    .ZN(_10074_)
  );
  AND2_X1 _19850_ (
    .A1(_02082_),
    .A2(_10074_),
    .ZN(_10075_)
  );
  AND2_X1 _19851_ (
    .A1(_10072_),
    .A2(_10075_),
    .ZN(_10076_)
  );
  INV_X1 _19852_ (
    .A(_10076_),
    .ZN(_10077_)
  );
  AND2_X1 _19853_ (
    .A1(remainder[59]),
    .A2(_02077_),
    .ZN(_10078_)
  );
  INV_X1 _19854_ (
    .A(_10078_),
    .ZN(_10080_)
  );
  AND2_X1 _19855_ (
    .A1(_04481_),
    .A2(_10451_),
    .ZN(_10081_)
  );
  INV_X1 _19856_ (
    .A(_10081_),
    .ZN(_10082_)
  );
  AND2_X1 _19857_ (
    .A1(_10462_),
    .A2(_01991_),
    .ZN(_10083_)
  );
  INV_X1 _19858_ (
    .A(_10083_),
    .ZN(_10084_)
  );
  AND2_X1 _19859_ (
    .A1(_05983_),
    .A2(_10084_),
    .ZN(_10085_)
  );
  AND2_X1 _19860_ (
    .A1(_10082_),
    .A2(_10085_),
    .ZN(_10086_)
  );
  INV_X1 _19861_ (
    .A(_10086_),
    .ZN(_10087_)
  );
  AND2_X1 _19862_ (
    .A1(_10080_),
    .A2(_10087_),
    .ZN(_10088_)
  );
  AND2_X1 _19863_ (
    .A1(_10077_),
    .A2(_10088_),
    .ZN(_10089_)
  );
  INV_X1 _19864_ (
    .A(_10089_),
    .ZN(_10091_)
  );
  AND2_X1 _19865_ (
    .A1(_06201_),
    .A2(_10091_),
    .ZN(_00080_)
  );
  AND2_X1 _19866_ (
    .A1(_10065_),
    .A2(_10072_),
    .ZN(_10092_)
  );
  INV_X1 _19867_ (
    .A(_10092_),
    .ZN(_10093_)
  );
  AND2_X1 _19868_ (
    .A1(_10048_),
    .A2(_10059_),
    .ZN(_10094_)
  );
  INV_X1 _19869_ (
    .A(_10094_),
    .ZN(_10095_)
  );
  AND2_X1 _19870_ (
    .A1(_10028_),
    .A2(_10034_),
    .ZN(_10096_)
  );
  INV_X1 _19871_ (
    .A(_10096_),
    .ZN(_10097_)
  );
  AND2_X1 _19872_ (
    .A1(_10008_),
    .A2(_10015_),
    .ZN(_10098_)
  );
  INV_X1 _19873_ (
    .A(_10098_),
    .ZN(_10099_)
  );
  AND2_X1 _19874_ (
    .A1(_09999_),
    .A2(_10021_),
    .ZN(_10101_)
  );
  INV_X1 _19875_ (
    .A(_10101_),
    .ZN(_10102_)
  );
  AND2_X1 _19876_ (
    .A1(_09933_),
    .A2(_09993_),
    .ZN(_10103_)
  );
  INV_X1 _19877_ (
    .A(_10103_),
    .ZN(_10104_)
  );
  AND2_X1 _19878_ (
    .A1(_09853_),
    .A2(_09927_),
    .ZN(_10105_)
  );
  INV_X1 _19879_ (
    .A(_10105_),
    .ZN(_10106_)
  );
  AND2_X1 _19880_ (
    .A1(_03249_),
    .A2(_09545_),
    .ZN(_10107_)
  );
  INV_X1 _19881_ (
    .A(_10107_),
    .ZN(_10108_)
  );
  AND2_X1 _19882_ (
    .A1(_03249_),
    .A2(_09547_),
    .ZN(_10109_)
  );
  INV_X1 _19883_ (
    .A(_10109_),
    .ZN(_10110_)
  );
  AND2_X1 _19884_ (
    .A1(_03250_),
    .A2(_09548_),
    .ZN(_10112_)
  );
  INV_X1 _19885_ (
    .A(_10112_),
    .ZN(_10113_)
  );
  AND2_X1 _19886_ (
    .A1(_10110_),
    .A2(_10113_),
    .ZN(_10114_)
  );
  INV_X1 _19887_ (
    .A(_10114_),
    .ZN(_10115_)
  );
  MUX2_X1 _19888_ (
    .A(_05084_),
    .B(_10114_),
    .S(_09780_),
    .Z(_10116_)
  );
  MUX2_X1 _19889_ (
    .A(remainder[1]),
    .B(_10115_),
    .S(_09780_),
    .Z(_10117_)
  );
  AND2_X1 _19890_ (
    .A1(_09807_),
    .A2(_09833_),
    .ZN(_10118_)
  );
  INV_X1 _19891_ (
    .A(_10118_),
    .ZN(_10119_)
  );
  AND2_X1 _19892_ (
    .A1(_09796_),
    .A2(_09800_),
    .ZN(_10120_)
  );
  INV_X1 _19893_ (
    .A(_10120_),
    .ZN(_10121_)
  );
  AND2_X1 _19894_ (
    .A1(divisor[31]),
    .A2(remainder[4]),
    .ZN(_10123_)
  );
  INV_X1 _19895_ (
    .A(_10123_),
    .ZN(_10124_)
  );
  AND2_X1 _19896_ (
    .A1(divisor[32]),
    .A2(remainder[3]),
    .ZN(_10125_)
  );
  INV_X1 _19897_ (
    .A(_10125_),
    .ZN(_10126_)
  );
  AND2_X1 _19898_ (
    .A1(remainder[3]),
    .A2(_09792_),
    .ZN(_10127_)
  );
  INV_X1 _19899_ (
    .A(_10127_),
    .ZN(_10128_)
  );
  MUX2_X1 _19900_ (
    .A(_09792_),
    .B(_05095_),
    .S(_10125_),
    .Z(_10129_)
  );
  MUX2_X1 _19901_ (
    .A(remainder[2]),
    .B(_09794_),
    .S(_10126_),
    .Z(_10130_)
  );
  AND2_X1 _19902_ (
    .A1(_10123_),
    .A2(_10129_),
    .ZN(_10131_)
  );
  INV_X1 _19903_ (
    .A(_10131_),
    .ZN(_10132_)
  );
  AND2_X1 _19904_ (
    .A1(_10124_),
    .A2(_10130_),
    .ZN(_10134_)
  );
  INV_X1 _19905_ (
    .A(_10134_),
    .ZN(_10135_)
  );
  AND2_X1 _19906_ (
    .A1(_10132_),
    .A2(_10135_),
    .ZN(_10136_)
  );
  INV_X1 _19907_ (
    .A(_10136_),
    .ZN(_10137_)
  );
  AND2_X1 _19908_ (
    .A1(_10121_),
    .A2(_10136_),
    .ZN(_10138_)
  );
  INV_X1 _19909_ (
    .A(_10138_),
    .ZN(_10139_)
  );
  AND2_X1 _19910_ (
    .A1(_10120_),
    .A2(_10137_),
    .ZN(_10140_)
  );
  INV_X1 _19911_ (
    .A(_10140_),
    .ZN(_10141_)
  );
  AND2_X1 _19912_ (
    .A1(_10139_),
    .A2(_10141_),
    .ZN(_10142_)
  );
  INV_X1 _19913_ (
    .A(_10142_),
    .ZN(_10143_)
  );
  AND2_X1 _19914_ (
    .A1(divisor[28]),
    .A2(remainder[7]),
    .ZN(_10145_)
  );
  INV_X1 _19915_ (
    .A(_10145_),
    .ZN(_10146_)
  );
  AND2_X1 _19916_ (
    .A1(divisor[29]),
    .A2(remainder[6]),
    .ZN(_10147_)
  );
  INV_X1 _19917_ (
    .A(_10147_),
    .ZN(_10148_)
  );
  AND2_X1 _19918_ (
    .A1(divisor[30]),
    .A2(remainder[6]),
    .ZN(_10149_)
  );
  INV_X1 _19919_ (
    .A(_10149_),
    .ZN(_10150_)
  );
  AND2_X1 _19920_ (
    .A1(_09817_),
    .A2(_10147_),
    .ZN(_10151_)
  );
  INV_X1 _19921_ (
    .A(_10151_),
    .ZN(_10152_)
  );
  AND2_X1 _19922_ (
    .A1(_09818_),
    .A2(_10148_),
    .ZN(_10153_)
  );
  INV_X1 _19923_ (
    .A(_10153_),
    .ZN(_10154_)
  );
  AND2_X1 _19924_ (
    .A1(_10152_),
    .A2(_10154_),
    .ZN(_10156_)
  );
  INV_X1 _19925_ (
    .A(_10156_),
    .ZN(_10157_)
  );
  AND2_X1 _19926_ (
    .A1(_10145_),
    .A2(_10156_),
    .ZN(_10158_)
  );
  INV_X1 _19927_ (
    .A(_10158_),
    .ZN(_10159_)
  );
  AND2_X1 _19928_ (
    .A1(_10146_),
    .A2(_10157_),
    .ZN(_10160_)
  );
  INV_X1 _19929_ (
    .A(_10160_),
    .ZN(_10161_)
  );
  AND2_X1 _19930_ (
    .A1(_10159_),
    .A2(_10161_),
    .ZN(_10162_)
  );
  INV_X1 _19931_ (
    .A(_10162_),
    .ZN(_10163_)
  );
  AND2_X1 _19932_ (
    .A1(_10142_),
    .A2(_10162_),
    .ZN(_10164_)
  );
  INV_X1 _19933_ (
    .A(_10164_),
    .ZN(_10165_)
  );
  AND2_X1 _19934_ (
    .A1(_10143_),
    .A2(_10163_),
    .ZN(_10167_)
  );
  INV_X1 _19935_ (
    .A(_10167_),
    .ZN(_10168_)
  );
  AND2_X1 _19936_ (
    .A1(_10165_),
    .A2(_10168_),
    .ZN(_10169_)
  );
  INV_X1 _19937_ (
    .A(_10169_),
    .ZN(_10170_)
  );
  AND2_X1 _19938_ (
    .A1(_10119_),
    .A2(_10169_),
    .ZN(_10171_)
  );
  INV_X1 _19939_ (
    .A(_10171_),
    .ZN(_10172_)
  );
  AND2_X1 _19940_ (
    .A1(_10118_),
    .A2(_10170_),
    .ZN(_10173_)
  );
  INV_X1 _19941_ (
    .A(_10173_),
    .ZN(_10174_)
  );
  AND2_X1 _19942_ (
    .A1(_10172_),
    .A2(_10174_),
    .ZN(_10175_)
  );
  INV_X1 _19943_ (
    .A(_10175_),
    .ZN(_10176_)
  );
  AND2_X1 _19944_ (
    .A1(_10116_),
    .A2(_10175_),
    .ZN(_10178_)
  );
  INV_X1 _19945_ (
    .A(_10178_),
    .ZN(_10179_)
  );
  AND2_X1 _19946_ (
    .A1(_10117_),
    .A2(_10176_),
    .ZN(_10180_)
  );
  INV_X1 _19947_ (
    .A(_10180_),
    .ZN(_10181_)
  );
  AND2_X1 _19948_ (
    .A1(_10179_),
    .A2(_10181_),
    .ZN(_10182_)
  );
  INV_X1 _19949_ (
    .A(_10182_),
    .ZN(_10183_)
  );
  AND2_X1 _19950_ (
    .A1(_09845_),
    .A2(_10182_),
    .ZN(_10184_)
  );
  INV_X1 _19951_ (
    .A(_10184_),
    .ZN(_10185_)
  );
  AND2_X1 _19952_ (
    .A1(_09846_),
    .A2(_10183_),
    .ZN(_10186_)
  );
  INV_X1 _19953_ (
    .A(_10186_),
    .ZN(_10187_)
  );
  AND2_X1 _19954_ (
    .A1(_10185_),
    .A2(_10187_),
    .ZN(_10189_)
  );
  INV_X1 _19955_ (
    .A(_10189_),
    .ZN(_10190_)
  );
  AND2_X1 _19956_ (
    .A1(_09900_),
    .A2(_09907_),
    .ZN(_10191_)
  );
  INV_X1 _19957_ (
    .A(_10191_),
    .ZN(_10192_)
  );
  AND2_X1 _19958_ (
    .A1(_09887_),
    .A2(_09894_),
    .ZN(_10193_)
  );
  INV_X1 _19959_ (
    .A(_10193_),
    .ZN(_10194_)
  );
  AND2_X1 _19960_ (
    .A1(_09874_),
    .A2(_09880_),
    .ZN(_10195_)
  );
  INV_X1 _19961_ (
    .A(_10195_),
    .ZN(_10196_)
  );
  AND2_X1 _19962_ (
    .A1(_09820_),
    .A2(_09827_),
    .ZN(_10197_)
  );
  INV_X1 _19963_ (
    .A(_10197_),
    .ZN(_10198_)
  );
  MUX2_X1 _19964_ (
    .A(_09868_),
    .B(_05040_),
    .S(_09867_),
    .Z(_10200_)
  );
  AND2_X1 _19965_ (
    .A1(divisor[25]),
    .A2(_10200_),
    .ZN(_10201_)
  );
  INV_X1 _19966_ (
    .A(_10201_),
    .ZN(_10202_)
  );
  MUX2_X1 _19967_ (
    .A(_09472_),
    .B(_05029_),
    .S(_10200_),
    .Z(_10203_)
  );
  MUX2_X1 _19968_ (
    .A(_09473_),
    .B(divisor[25]),
    .S(_10200_),
    .Z(_10204_)
  );
  AND2_X1 _19969_ (
    .A1(_10198_),
    .A2(_10203_),
    .ZN(_10205_)
  );
  INV_X1 _19970_ (
    .A(_10205_),
    .ZN(_10206_)
  );
  AND2_X1 _19971_ (
    .A1(_10197_),
    .A2(_10204_),
    .ZN(_10207_)
  );
  INV_X1 _19972_ (
    .A(_10207_),
    .ZN(_10208_)
  );
  AND2_X1 _19973_ (
    .A1(_10206_),
    .A2(_10208_),
    .ZN(_10209_)
  );
  INV_X1 _19974_ (
    .A(_10209_),
    .ZN(_10211_)
  );
  AND2_X1 _19975_ (
    .A1(_10196_),
    .A2(_10209_),
    .ZN(_10212_)
  );
  INV_X1 _19976_ (
    .A(_10212_),
    .ZN(_10213_)
  );
  AND2_X1 _19977_ (
    .A1(_10195_),
    .A2(_10211_),
    .ZN(_10214_)
  );
  INV_X1 _19978_ (
    .A(_10214_),
    .ZN(_10215_)
  );
  AND2_X1 _19979_ (
    .A1(_10213_),
    .A2(_10215_),
    .ZN(_10216_)
  );
  INV_X1 _19980_ (
    .A(_10216_),
    .ZN(_10217_)
  );
  AND2_X1 _19981_ (
    .A1(_10194_),
    .A2(_10216_),
    .ZN(_10218_)
  );
  INV_X1 _19982_ (
    .A(_10218_),
    .ZN(_10219_)
  );
  AND2_X1 _19983_ (
    .A1(_10193_),
    .A2(_10217_),
    .ZN(_10220_)
  );
  INV_X1 _19984_ (
    .A(_10220_),
    .ZN(_10222_)
  );
  AND2_X1 _19985_ (
    .A1(_10219_),
    .A2(_10222_),
    .ZN(_10223_)
  );
  INV_X1 _19986_ (
    .A(_10223_),
    .ZN(_10224_)
  );
  AND2_X1 _19987_ (
    .A1(_09521_),
    .A2(_10223_),
    .ZN(_10225_)
  );
  INV_X1 _19988_ (
    .A(_10225_),
    .ZN(_10226_)
  );
  AND2_X1 _19989_ (
    .A1(_09522_),
    .A2(_10224_),
    .ZN(_10227_)
  );
  INV_X1 _19990_ (
    .A(_10227_),
    .ZN(_10228_)
  );
  AND2_X1 _19991_ (
    .A1(_10226_),
    .A2(_10228_),
    .ZN(_10229_)
  );
  INV_X1 _19992_ (
    .A(_10229_),
    .ZN(_10230_)
  );
  AND2_X1 _19993_ (
    .A1(_09839_),
    .A2(_10229_),
    .ZN(_10231_)
  );
  INV_X1 _19994_ (
    .A(_10231_),
    .ZN(_10233_)
  );
  AND2_X1 _19995_ (
    .A1(_09840_),
    .A2(_10230_),
    .ZN(_10234_)
  );
  INV_X1 _19996_ (
    .A(_10234_),
    .ZN(_10235_)
  );
  AND2_X1 _19997_ (
    .A1(_10233_),
    .A2(_10235_),
    .ZN(_10236_)
  );
  INV_X1 _19998_ (
    .A(_10236_),
    .ZN(_10237_)
  );
  AND2_X1 _19999_ (
    .A1(_10192_),
    .A2(_10236_),
    .ZN(_10238_)
  );
  INV_X1 _20000_ (
    .A(_10238_),
    .ZN(_10239_)
  );
  AND2_X1 _20001_ (
    .A1(_10191_),
    .A2(_10237_),
    .ZN(_10240_)
  );
  INV_X1 _20002_ (
    .A(_10240_),
    .ZN(_10241_)
  );
  AND2_X1 _20003_ (
    .A1(_10239_),
    .A2(_10241_),
    .ZN(_10242_)
  );
  INV_X1 _20004_ (
    .A(_10242_),
    .ZN(_10244_)
  );
  AND2_X1 _20005_ (
    .A1(_10189_),
    .A2(_10242_),
    .ZN(_10245_)
  );
  INV_X1 _20006_ (
    .A(_10245_),
    .ZN(_10246_)
  );
  AND2_X1 _20007_ (
    .A1(_10190_),
    .A2(_10244_),
    .ZN(_10247_)
  );
  INV_X1 _20008_ (
    .A(_10247_),
    .ZN(_10248_)
  );
  AND2_X1 _20009_ (
    .A1(_10246_),
    .A2(_10248_),
    .ZN(_10249_)
  );
  INV_X1 _20010_ (
    .A(_10249_),
    .ZN(_10250_)
  );
  AND2_X1 _20011_ (
    .A1(_10106_),
    .A2(_10249_),
    .ZN(_10251_)
  );
  INV_X1 _20012_ (
    .A(_10251_),
    .ZN(_10252_)
  );
  AND2_X1 _20013_ (
    .A1(_10105_),
    .A2(_10250_),
    .ZN(_10253_)
  );
  INV_X1 _20014_ (
    .A(_10253_),
    .ZN(_10255_)
  );
  AND2_X1 _20015_ (
    .A1(_10252_),
    .A2(_10255_),
    .ZN(_10256_)
  );
  INV_X1 _20016_ (
    .A(_10256_),
    .ZN(_10257_)
  );
  AND2_X1 _20017_ (
    .A1(_09966_),
    .A2(_09973_),
    .ZN(_10258_)
  );
  INV_X1 _20018_ (
    .A(_10258_),
    .ZN(_10259_)
  );
  AND2_X1 _20019_ (
    .A1(_09913_),
    .A2(_09920_),
    .ZN(_10260_)
  );
  INV_X1 _20020_ (
    .A(_10260_),
    .ZN(_10261_)
  );
  AND2_X1 _20021_ (
    .A1(_08998_),
    .A2(_09950_),
    .ZN(_10262_)
  );
  INV_X1 _20022_ (
    .A(_10262_),
    .ZN(_10263_)
  );
  AND2_X1 _20023_ (
    .A1(_09966_),
    .A2(_10263_),
    .ZN(_10264_)
  );
  INV_X1 _20024_ (
    .A(_10264_),
    .ZN(_10266_)
  );
  AND2_X1 _20025_ (
    .A1(_07082_),
    .A2(_10264_),
    .ZN(_10267_)
  );
  INV_X1 _20026_ (
    .A(_10267_),
    .ZN(_10268_)
  );
  AND2_X1 _20027_ (
    .A1(_07083_),
    .A2(_10266_),
    .ZN(_10269_)
  );
  INV_X1 _20028_ (
    .A(_10269_),
    .ZN(_10270_)
  );
  AND2_X1 _20029_ (
    .A1(_10268_),
    .A2(_10270_),
    .ZN(_10271_)
  );
  INV_X1 _20030_ (
    .A(_10271_),
    .ZN(_10272_)
  );
  AND2_X1 _20031_ (
    .A1(_10261_),
    .A2(_10271_),
    .ZN(_10273_)
  );
  INV_X1 _20032_ (
    .A(_10273_),
    .ZN(_10274_)
  );
  AND2_X1 _20033_ (
    .A1(_10260_),
    .A2(_10272_),
    .ZN(_10275_)
  );
  INV_X1 _20034_ (
    .A(_10275_),
    .ZN(_10277_)
  );
  AND2_X1 _20035_ (
    .A1(_10274_),
    .A2(_10277_),
    .ZN(_10278_)
  );
  INV_X1 _20036_ (
    .A(_10278_),
    .ZN(_10279_)
  );
  AND2_X1 _20037_ (
    .A1(_10259_),
    .A2(_10278_),
    .ZN(_10280_)
  );
  INV_X1 _20038_ (
    .A(_10280_),
    .ZN(_10281_)
  );
  AND2_X1 _20039_ (
    .A1(_10258_),
    .A2(_10279_),
    .ZN(_10282_)
  );
  INV_X1 _20040_ (
    .A(_10282_),
    .ZN(_10283_)
  );
  AND2_X1 _20041_ (
    .A1(_10281_),
    .A2(_10283_),
    .ZN(_10284_)
  );
  INV_X1 _20042_ (
    .A(_10284_),
    .ZN(_10285_)
  );
  AND2_X1 _20043_ (
    .A1(_10256_),
    .A2(_10284_),
    .ZN(_10286_)
  );
  INV_X1 _20044_ (
    .A(_10286_),
    .ZN(_10288_)
  );
  AND2_X1 _20045_ (
    .A1(_10257_),
    .A2(_10285_),
    .ZN(_10289_)
  );
  INV_X1 _20046_ (
    .A(_10289_),
    .ZN(_10290_)
  );
  AND2_X1 _20047_ (
    .A1(_10288_),
    .A2(_10290_),
    .ZN(_10291_)
  );
  INV_X1 _20048_ (
    .A(_10291_),
    .ZN(_10292_)
  );
  AND2_X1 _20049_ (
    .A1(_10104_),
    .A2(_10291_),
    .ZN(_10293_)
  );
  INV_X1 _20050_ (
    .A(_10293_),
    .ZN(_10294_)
  );
  AND2_X1 _20051_ (
    .A1(_10103_),
    .A2(_10292_),
    .ZN(_10295_)
  );
  INV_X1 _20052_ (
    .A(_10295_),
    .ZN(_10296_)
  );
  AND2_X1 _20053_ (
    .A1(_10294_),
    .A2(_10296_),
    .ZN(_10297_)
  );
  INV_X1 _20054_ (
    .A(_10297_),
    .ZN(_10299_)
  );
  AND2_X1 _20055_ (
    .A1(_09979_),
    .A2(_09986_),
    .ZN(_10300_)
  );
  INV_X1 _20056_ (
    .A(_10300_),
    .ZN(_10301_)
  );
  AND2_X1 _20057_ (
    .A1(_07804_),
    .A2(_10301_),
    .ZN(_10302_)
  );
  INV_X1 _20058_ (
    .A(_10302_),
    .ZN(_10303_)
  );
  AND2_X1 _20059_ (
    .A1(_07805_),
    .A2(_10300_),
    .ZN(_10304_)
  );
  INV_X1 _20060_ (
    .A(_10304_),
    .ZN(_10305_)
  );
  AND2_X1 _20061_ (
    .A1(_10303_),
    .A2(_10305_),
    .ZN(_10306_)
  );
  INV_X1 _20062_ (
    .A(_10306_),
    .ZN(_10307_)
  );
  AND2_X1 _20063_ (
    .A1(_08107_),
    .A2(_10306_),
    .ZN(_10308_)
  );
  INV_X1 _20064_ (
    .A(_10308_),
    .ZN(_10310_)
  );
  AND2_X1 _20065_ (
    .A1(_08106_),
    .A2(_10307_),
    .ZN(_10311_)
  );
  INV_X1 _20066_ (
    .A(_10311_),
    .ZN(_10312_)
  );
  AND2_X1 _20067_ (
    .A1(_10310_),
    .A2(_10312_),
    .ZN(_10313_)
  );
  INV_X1 _20068_ (
    .A(_10313_),
    .ZN(_10314_)
  );
  AND2_X1 _20069_ (
    .A1(_10297_),
    .A2(_10313_),
    .ZN(_10315_)
  );
  INV_X1 _20070_ (
    .A(_10315_),
    .ZN(_10316_)
  );
  AND2_X1 _20071_ (
    .A1(_10299_),
    .A2(_10314_),
    .ZN(_10317_)
  );
  INV_X1 _20072_ (
    .A(_10317_),
    .ZN(_10318_)
  );
  AND2_X1 _20073_ (
    .A1(_10316_),
    .A2(_10318_),
    .ZN(_10319_)
  );
  INV_X1 _20074_ (
    .A(_10319_),
    .ZN(_10321_)
  );
  AND2_X1 _20075_ (
    .A1(_10102_),
    .A2(_10319_),
    .ZN(_10322_)
  );
  INV_X1 _20076_ (
    .A(_10322_),
    .ZN(_10323_)
  );
  AND2_X1 _20077_ (
    .A1(_10101_),
    .A2(_10321_),
    .ZN(_10324_)
  );
  INV_X1 _20078_ (
    .A(_10324_),
    .ZN(_10325_)
  );
  AND2_X1 _20079_ (
    .A1(_10323_),
    .A2(_10325_),
    .ZN(_10326_)
  );
  INV_X1 _20080_ (
    .A(_10326_),
    .ZN(_10327_)
  );
  AND2_X1 _20081_ (
    .A1(_10099_),
    .A2(_10326_),
    .ZN(_10328_)
  );
  INV_X1 _20082_ (
    .A(_10328_),
    .ZN(_10329_)
  );
  AND2_X1 _20083_ (
    .A1(_10098_),
    .A2(_10327_),
    .ZN(_10330_)
  );
  INV_X1 _20084_ (
    .A(_10330_),
    .ZN(_10332_)
  );
  AND2_X1 _20085_ (
    .A1(_10329_),
    .A2(_10332_),
    .ZN(_10333_)
  );
  INV_X1 _20086_ (
    .A(_10333_),
    .ZN(_10334_)
  );
  AND2_X1 _20087_ (
    .A1(_10097_),
    .A2(_10333_),
    .ZN(_10335_)
  );
  INV_X1 _20088_ (
    .A(_10335_),
    .ZN(_10336_)
  );
  AND2_X1 _20089_ (
    .A1(_10096_),
    .A2(_10334_),
    .ZN(_10337_)
  );
  INV_X1 _20090_ (
    .A(_10337_),
    .ZN(_10338_)
  );
  AND2_X1 _20091_ (
    .A1(_10336_),
    .A2(_10338_),
    .ZN(_10339_)
  );
  INV_X1 _20092_ (
    .A(_10339_),
    .ZN(_10340_)
  );
  AND2_X1 _20093_ (
    .A1(_10040_),
    .A2(_10339_),
    .ZN(_10341_)
  );
  INV_X1 _20094_ (
    .A(_10341_),
    .ZN(_10343_)
  );
  AND2_X1 _20095_ (
    .A1(_10041_),
    .A2(_10340_),
    .ZN(_10344_)
  );
  INV_X1 _20096_ (
    .A(_10344_),
    .ZN(_10345_)
  );
  AND2_X1 _20097_ (
    .A1(_10343_),
    .A2(_10345_),
    .ZN(_10346_)
  );
  INV_X1 _20098_ (
    .A(_10346_),
    .ZN(_10347_)
  );
  AND2_X1 _20099_ (
    .A1(_10094_),
    .A2(_10347_),
    .ZN(_10348_)
  );
  INV_X1 _20100_ (
    .A(_10348_),
    .ZN(_10349_)
  );
  AND2_X1 _20101_ (
    .A1(_10095_),
    .A2(_10346_),
    .ZN(_10350_)
  );
  INV_X1 _20102_ (
    .A(_10350_),
    .ZN(_10351_)
  );
  AND2_X1 _20103_ (
    .A1(_10349_),
    .A2(_10351_),
    .ZN(_10352_)
  );
  INV_X1 _20104_ (
    .A(_10352_),
    .ZN(_10354_)
  );
  AND2_X1 _20105_ (
    .A1(_04404_),
    .A2(_10354_),
    .ZN(_10355_)
  );
  INV_X1 _20106_ (
    .A(_10355_),
    .ZN(_10356_)
  );
  AND2_X1 _20107_ (
    .A1(remainder[65]),
    .A2(_10352_),
    .ZN(_10357_)
  );
  INV_X1 _20108_ (
    .A(_10357_),
    .ZN(_10358_)
  );
  AND2_X1 _20109_ (
    .A1(_10356_),
    .A2(_10358_),
    .ZN(_10359_)
  );
  INV_X1 _20110_ (
    .A(_10359_),
    .ZN(_10360_)
  );
  AND2_X1 _20111_ (
    .A1(_10092_),
    .A2(_10360_),
    .ZN(_10361_)
  );
  INV_X1 _20112_ (
    .A(_10361_),
    .ZN(_10362_)
  );
  AND2_X1 _20113_ (
    .A1(_10093_),
    .A2(_10359_),
    .ZN(_10363_)
  );
  INV_X1 _20114_ (
    .A(_10363_),
    .ZN(_10365_)
  );
  AND2_X1 _20115_ (
    .A1(_02082_),
    .A2(_10362_),
    .ZN(_10366_)
  );
  AND2_X1 _20116_ (
    .A1(_10365_),
    .A2(_10366_),
    .ZN(_10367_)
  );
  INV_X1 _20117_ (
    .A(_10367_),
    .ZN(_10368_)
  );
  AND2_X1 _20118_ (
    .A1(remainder[60]),
    .A2(_02077_),
    .ZN(_10369_)
  );
  INV_X1 _20119_ (
    .A(_10369_),
    .ZN(_10370_)
  );
  MUX2_X1 _20120_ (
    .A(remainder[59]),
    .B(_02006_),
    .S(_10462_),
    .Z(_10371_)
  );
  AND2_X1 _20121_ (
    .A1(_05983_),
    .A2(_10371_),
    .ZN(_10372_)
  );
  INV_X1 _20122_ (
    .A(_10372_),
    .ZN(_10373_)
  );
  AND2_X1 _20123_ (
    .A1(_10370_),
    .A2(_10373_),
    .ZN(_10374_)
  );
  AND2_X1 _20124_ (
    .A1(_10368_),
    .A2(_10374_),
    .ZN(_10376_)
  );
  INV_X1 _20125_ (
    .A(_10376_),
    .ZN(_10377_)
  );
  AND2_X1 _20126_ (
    .A1(_06201_),
    .A2(_10377_),
    .ZN(_00081_)
  );
  AND2_X1 _20127_ (
    .A1(_09757_),
    .A2(_10069_),
    .ZN(_10378_)
  );
  AND2_X1 _20128_ (
    .A1(_10359_),
    .A2(_10378_),
    .ZN(_10379_)
  );
  INV_X1 _20129_ (
    .A(_10379_),
    .ZN(_10380_)
  );
  AND2_X1 _20130_ (
    .A1(_09759_),
    .A2(_10065_),
    .ZN(_10381_)
  );
  AND2_X1 _20131_ (
    .A1(_10358_),
    .A2(_10381_),
    .ZN(_10382_)
  );
  AND2_X1 _20132_ (
    .A1(_10380_),
    .A2(_10382_),
    .ZN(_10383_)
  );
  INV_X1 _20133_ (
    .A(_10383_),
    .ZN(_10384_)
  );
  AND2_X1 _20134_ (
    .A1(_10323_),
    .A2(_10329_),
    .ZN(_10386_)
  );
  INV_X1 _20135_ (
    .A(_10386_),
    .ZN(_10387_)
  );
  AND2_X1 _20136_ (
    .A1(_10303_),
    .A2(_10310_),
    .ZN(_10388_)
  );
  INV_X1 _20137_ (
    .A(_10388_),
    .ZN(_10389_)
  );
  AND2_X1 _20138_ (
    .A1(_10294_),
    .A2(_10316_),
    .ZN(_10390_)
  );
  INV_X1 _20139_ (
    .A(_10390_),
    .ZN(_10391_)
  );
  AND2_X1 _20140_ (
    .A1(_10252_),
    .A2(_10288_),
    .ZN(_10392_)
  );
  INV_X1 _20141_ (
    .A(_10392_),
    .ZN(_10393_)
  );
  AND2_X1 _20142_ (
    .A1(_10185_),
    .A2(_10246_),
    .ZN(_10394_)
  );
  INV_X1 _20143_ (
    .A(_10394_),
    .ZN(_10395_)
  );
  AND2_X1 _20144_ (
    .A1(_10108_),
    .A2(_10179_),
    .ZN(_10397_)
  );
  INV_X1 _20145_ (
    .A(_10397_),
    .ZN(_10398_)
  );
  AND2_X1 _20146_ (
    .A1(_10139_),
    .A2(_10165_),
    .ZN(_10399_)
  );
  INV_X1 _20147_ (
    .A(_10399_),
    .ZN(_10400_)
  );
  AND2_X1 _20148_ (
    .A1(_10128_),
    .A2(_10132_),
    .ZN(_10401_)
  );
  INV_X1 _20149_ (
    .A(_10401_),
    .ZN(_10402_)
  );
  AND2_X1 _20150_ (
    .A1(divisor[31]),
    .A2(remainder[5]),
    .ZN(_10403_)
  );
  INV_X1 _20151_ (
    .A(_10403_),
    .ZN(_10404_)
  );
  AND2_X1 _20152_ (
    .A1(divisor[32]),
    .A2(remainder[4]),
    .ZN(_10405_)
  );
  INV_X1 _20153_ (
    .A(_10405_),
    .ZN(_10406_)
  );
  AND2_X1 _20154_ (
    .A1(remainder[4]),
    .A2(_10125_),
    .ZN(_10408_)
  );
  INV_X1 _20155_ (
    .A(_10408_),
    .ZN(_10409_)
  );
  MUX2_X1 _20156_ (
    .A(_10125_),
    .B(_05105_),
    .S(_10405_),
    .Z(_10410_)
  );
  MUX2_X1 _20157_ (
    .A(remainder[3]),
    .B(_10126_),
    .S(_10406_),
    .Z(_10411_)
  );
  AND2_X1 _20158_ (
    .A1(_10403_),
    .A2(_10410_),
    .ZN(_10412_)
  );
  INV_X1 _20159_ (
    .A(_10412_),
    .ZN(_10413_)
  );
  AND2_X1 _20160_ (
    .A1(_10404_),
    .A2(_10411_),
    .ZN(_10414_)
  );
  INV_X1 _20161_ (
    .A(_10414_),
    .ZN(_10415_)
  );
  AND2_X1 _20162_ (
    .A1(_10413_),
    .A2(_10415_),
    .ZN(_10416_)
  );
  INV_X1 _20163_ (
    .A(_10416_),
    .ZN(_10417_)
  );
  AND2_X1 _20164_ (
    .A1(_10402_),
    .A2(_10416_),
    .ZN(_10419_)
  );
  INV_X1 _20165_ (
    .A(_10419_),
    .ZN(_10420_)
  );
  AND2_X1 _20166_ (
    .A1(_10401_),
    .A2(_10417_),
    .ZN(_10421_)
  );
  INV_X1 _20167_ (
    .A(_10421_),
    .ZN(_10422_)
  );
  AND2_X1 _20168_ (
    .A1(_10420_),
    .A2(_10422_),
    .ZN(_10423_)
  );
  INV_X1 _20169_ (
    .A(_10423_),
    .ZN(_10424_)
  );
  AND2_X1 _20170_ (
    .A1(divisor[29]),
    .A2(remainder[7]),
    .ZN(_10425_)
  );
  INV_X1 _20171_ (
    .A(_10425_),
    .ZN(_10426_)
  );
  AND2_X1 _20172_ (
    .A1(divisor[30]),
    .A2(remainder[7]),
    .ZN(_10427_)
  );
  INV_X1 _20173_ (
    .A(_10427_),
    .ZN(_10428_)
  );
  AND2_X1 _20174_ (
    .A1(_10147_),
    .A2(_10427_),
    .ZN(_10430_)
  );
  INV_X1 _20175_ (
    .A(_10430_),
    .ZN(_10431_)
  );
  AND2_X1 _20176_ (
    .A1(_10150_),
    .A2(_10426_),
    .ZN(_10432_)
  );
  INV_X1 _20177_ (
    .A(_10432_),
    .ZN(_10433_)
  );
  AND2_X1 _20178_ (
    .A1(_10431_),
    .A2(_10433_),
    .ZN(_10434_)
  );
  INV_X1 _20179_ (
    .A(_10434_),
    .ZN(_10435_)
  );
  AND2_X1 _20180_ (
    .A1(_08005_),
    .A2(_10434_),
    .ZN(_10436_)
  );
  INV_X1 _20181_ (
    .A(_10436_),
    .ZN(_10437_)
  );
  AND2_X1 _20182_ (
    .A1(_08007_),
    .A2(_10435_),
    .ZN(_10438_)
  );
  INV_X1 _20183_ (
    .A(_10438_),
    .ZN(_10439_)
  );
  AND2_X1 _20184_ (
    .A1(_10437_),
    .A2(_10439_),
    .ZN(_10441_)
  );
  INV_X1 _20185_ (
    .A(_10441_),
    .ZN(_10442_)
  );
  AND2_X1 _20186_ (
    .A1(_10423_),
    .A2(_10441_),
    .ZN(_10443_)
  );
  INV_X1 _20187_ (
    .A(_10443_),
    .ZN(_10444_)
  );
  AND2_X1 _20188_ (
    .A1(_10424_),
    .A2(_10442_),
    .ZN(_10445_)
  );
  INV_X1 _20189_ (
    .A(_10445_),
    .ZN(_10446_)
  );
  AND2_X1 _20190_ (
    .A1(_10444_),
    .A2(_10446_),
    .ZN(_10447_)
  );
  INV_X1 _20191_ (
    .A(_10447_),
    .ZN(_10448_)
  );
  AND2_X1 _20192_ (
    .A1(_10400_),
    .A2(_10447_),
    .ZN(_10449_)
  );
  INV_X1 _20193_ (
    .A(_10449_),
    .ZN(_10450_)
  );
  AND2_X1 _20194_ (
    .A1(_10399_),
    .A2(_10448_),
    .ZN(_10452_)
  );
  INV_X1 _20195_ (
    .A(_10452_),
    .ZN(_10453_)
  );
  AND2_X1 _20196_ (
    .A1(_10450_),
    .A2(_10453_),
    .ZN(_10454_)
  );
  INV_X1 _20197_ (
    .A(_10454_),
    .ZN(_10455_)
  );
  AND2_X1 _20198_ (
    .A1(_09545_),
    .A2(_09792_),
    .ZN(_10456_)
  );
  INV_X1 _20199_ (
    .A(_10456_),
    .ZN(_10457_)
  );
  AND2_X1 _20200_ (
    .A1(_09547_),
    .A2(_09792_),
    .ZN(_10458_)
  );
  INV_X1 _20201_ (
    .A(_10458_),
    .ZN(_10459_)
  );
  AND2_X1 _20202_ (
    .A1(_09548_),
    .A2(_09794_),
    .ZN(_10460_)
  );
  INV_X1 _20203_ (
    .A(_10460_),
    .ZN(_10461_)
  );
  AND2_X1 _20204_ (
    .A1(_10459_),
    .A2(_10461_),
    .ZN(_10463_)
  );
  MUX2_X1 _20205_ (
    .A(_09794_),
    .B(_10463_),
    .S(_09546_),
    .Z(_10464_)
  );
  INV_X1 _20206_ (
    .A(_10464_),
    .ZN(_10465_)
  );
  AND2_X1 _20207_ (
    .A1(_03249_),
    .A2(_09548_),
    .ZN(_10466_)
  );
  INV_X1 _20208_ (
    .A(_10466_),
    .ZN(_10467_)
  );
  AND2_X1 _20209_ (
    .A1(_10465_),
    .A2(_10467_),
    .ZN(_10468_)
  );
  INV_X1 _20210_ (
    .A(_10468_),
    .ZN(_10469_)
  );
  AND2_X1 _20211_ (
    .A1(_10464_),
    .A2(_10466_),
    .ZN(_10470_)
  );
  INV_X1 _20212_ (
    .A(_10470_),
    .ZN(_10471_)
  );
  AND2_X1 _20213_ (
    .A1(_10469_),
    .A2(_10471_),
    .ZN(_10472_)
  );
  INV_X1 _20214_ (
    .A(_10472_),
    .ZN(_10474_)
  );
  AND2_X1 _20215_ (
    .A1(_10454_),
    .A2(_10472_),
    .ZN(_10475_)
  );
  INV_X1 _20216_ (
    .A(_10475_),
    .ZN(_10476_)
  );
  AND2_X1 _20217_ (
    .A1(_10455_),
    .A2(_10474_),
    .ZN(_10477_)
  );
  INV_X1 _20218_ (
    .A(_10477_),
    .ZN(_10478_)
  );
  AND2_X1 _20219_ (
    .A1(_10476_),
    .A2(_10478_),
    .ZN(_10479_)
  );
  INV_X1 _20220_ (
    .A(_10479_),
    .ZN(_10480_)
  );
  AND2_X1 _20221_ (
    .A1(_10398_),
    .A2(_10479_),
    .ZN(_10481_)
  );
  INV_X1 _20222_ (
    .A(_10481_),
    .ZN(_10482_)
  );
  AND2_X1 _20223_ (
    .A1(_10397_),
    .A2(_10480_),
    .ZN(_10483_)
  );
  INV_X1 _20224_ (
    .A(_10483_),
    .ZN(_10485_)
  );
  AND2_X1 _20225_ (
    .A1(_10482_),
    .A2(_10485_),
    .ZN(_10486_)
  );
  INV_X1 _20226_ (
    .A(_10486_),
    .ZN(_10487_)
  );
  AND2_X1 _20227_ (
    .A1(_10219_),
    .A2(_10226_),
    .ZN(_10488_)
  );
  INV_X1 _20228_ (
    .A(_10488_),
    .ZN(_10489_)
  );
  AND2_X1 _20229_ (
    .A1(_10206_),
    .A2(_10213_),
    .ZN(_10490_)
  );
  INV_X1 _20230_ (
    .A(_10490_),
    .ZN(_10491_)
  );
  AND2_X1 _20231_ (
    .A1(_09872_),
    .A2(_10202_),
    .ZN(_10492_)
  );
  INV_X1 _20232_ (
    .A(_10492_),
    .ZN(_10493_)
  );
  AND2_X1 _20233_ (
    .A1(_10152_),
    .A2(_10159_),
    .ZN(_10494_)
  );
  INV_X1 _20234_ (
    .A(_10494_),
    .ZN(_10496_)
  );
  AND2_X1 _20235_ (
    .A1(_10203_),
    .A2(_10496_),
    .ZN(_10497_)
  );
  INV_X1 _20236_ (
    .A(_10497_),
    .ZN(_10498_)
  );
  AND2_X1 _20237_ (
    .A1(_10204_),
    .A2(_10494_),
    .ZN(_10499_)
  );
  INV_X1 _20238_ (
    .A(_10499_),
    .ZN(_10500_)
  );
  AND2_X1 _20239_ (
    .A1(_10498_),
    .A2(_10500_),
    .ZN(_10501_)
  );
  INV_X1 _20240_ (
    .A(_10501_),
    .ZN(_10502_)
  );
  AND2_X1 _20241_ (
    .A1(_10493_),
    .A2(_10501_),
    .ZN(_10503_)
  );
  INV_X1 _20242_ (
    .A(_10503_),
    .ZN(_10504_)
  );
  AND2_X1 _20243_ (
    .A1(_10492_),
    .A2(_10502_),
    .ZN(_10505_)
  );
  INV_X1 _20244_ (
    .A(_10505_),
    .ZN(_10507_)
  );
  AND2_X1 _20245_ (
    .A1(_10504_),
    .A2(_10507_),
    .ZN(_10508_)
  );
  INV_X1 _20246_ (
    .A(_10508_),
    .ZN(_10509_)
  );
  AND2_X1 _20247_ (
    .A1(_10491_),
    .A2(_10508_),
    .ZN(_10510_)
  );
  INV_X1 _20248_ (
    .A(_10510_),
    .ZN(_10511_)
  );
  AND2_X1 _20249_ (
    .A1(_10490_),
    .A2(_10509_),
    .ZN(_10512_)
  );
  INV_X1 _20250_ (
    .A(_10512_),
    .ZN(_10513_)
  );
  AND2_X1 _20251_ (
    .A1(_10511_),
    .A2(_10513_),
    .ZN(_10514_)
  );
  INV_X1 _20252_ (
    .A(_10514_),
    .ZN(_10515_)
  );
  AND2_X1 _20253_ (
    .A1(_09521_),
    .A2(_10514_),
    .ZN(_10516_)
  );
  INV_X1 _20254_ (
    .A(_10516_),
    .ZN(_10518_)
  );
  AND2_X1 _20255_ (
    .A1(_09522_),
    .A2(_10515_),
    .ZN(_10519_)
  );
  INV_X1 _20256_ (
    .A(_10519_),
    .ZN(_10520_)
  );
  AND2_X1 _20257_ (
    .A1(_10518_),
    .A2(_10520_),
    .ZN(_10521_)
  );
  INV_X1 _20258_ (
    .A(_10521_),
    .ZN(_10522_)
  );
  AND2_X1 _20259_ (
    .A1(_10171_),
    .A2(_10521_),
    .ZN(_10523_)
  );
  INV_X1 _20260_ (
    .A(_10523_),
    .ZN(_10524_)
  );
  AND2_X1 _20261_ (
    .A1(_10172_),
    .A2(_10522_),
    .ZN(_10525_)
  );
  INV_X1 _20262_ (
    .A(_10525_),
    .ZN(_10526_)
  );
  AND2_X1 _20263_ (
    .A1(_10524_),
    .A2(_10526_),
    .ZN(_10527_)
  );
  INV_X1 _20264_ (
    .A(_10527_),
    .ZN(_10529_)
  );
  AND2_X1 _20265_ (
    .A1(_10489_),
    .A2(_10527_),
    .ZN(_10530_)
  );
  INV_X1 _20266_ (
    .A(_10530_),
    .ZN(_10531_)
  );
  AND2_X1 _20267_ (
    .A1(_10488_),
    .A2(_10529_),
    .ZN(_10532_)
  );
  INV_X1 _20268_ (
    .A(_10532_),
    .ZN(_10533_)
  );
  AND2_X1 _20269_ (
    .A1(_10531_),
    .A2(_10533_),
    .ZN(_10534_)
  );
  INV_X1 _20270_ (
    .A(_10534_),
    .ZN(_10535_)
  );
  AND2_X1 _20271_ (
    .A1(_10486_),
    .A2(_10534_),
    .ZN(_10536_)
  );
  INV_X1 _20272_ (
    .A(_10536_),
    .ZN(_10537_)
  );
  AND2_X1 _20273_ (
    .A1(_10487_),
    .A2(_10535_),
    .ZN(_10538_)
  );
  INV_X1 _20274_ (
    .A(_10538_),
    .ZN(_10540_)
  );
  AND2_X1 _20275_ (
    .A1(_10537_),
    .A2(_10540_),
    .ZN(_10541_)
  );
  INV_X1 _20276_ (
    .A(_10541_),
    .ZN(_10542_)
  );
  AND2_X1 _20277_ (
    .A1(_10395_),
    .A2(_10541_),
    .ZN(_10543_)
  );
  INV_X1 _20278_ (
    .A(_10543_),
    .ZN(_10544_)
  );
  AND2_X1 _20279_ (
    .A1(_10394_),
    .A2(_10542_),
    .ZN(_10545_)
  );
  INV_X1 _20280_ (
    .A(_10545_),
    .ZN(_10546_)
  );
  AND2_X1 _20281_ (
    .A1(_10544_),
    .A2(_10546_),
    .ZN(_10547_)
  );
  INV_X1 _20282_ (
    .A(_10547_),
    .ZN(_10548_)
  );
  AND2_X1 _20283_ (
    .A1(_09966_),
    .A2(_10268_),
    .ZN(_10549_)
  );
  INV_X1 _20284_ (
    .A(_10549_),
    .ZN(_10551_)
  );
  AND2_X1 _20285_ (
    .A1(_10233_),
    .A2(_10239_),
    .ZN(_10552_)
  );
  INV_X1 _20286_ (
    .A(_10552_),
    .ZN(_10553_)
  );
  AND2_X1 _20287_ (
    .A1(_10271_),
    .A2(_10553_),
    .ZN(_10554_)
  );
  INV_X1 _20288_ (
    .A(_10554_),
    .ZN(_10555_)
  );
  AND2_X1 _20289_ (
    .A1(_10272_),
    .A2(_10552_),
    .ZN(_10556_)
  );
  INV_X1 _20290_ (
    .A(_10556_),
    .ZN(_10557_)
  );
  AND2_X1 _20291_ (
    .A1(_10555_),
    .A2(_10557_),
    .ZN(_10558_)
  );
  INV_X1 _20292_ (
    .A(_10558_),
    .ZN(_10559_)
  );
  AND2_X1 _20293_ (
    .A1(_10551_),
    .A2(_10558_),
    .ZN(_10560_)
  );
  INV_X1 _20294_ (
    .A(_10560_),
    .ZN(_10562_)
  );
  AND2_X1 _20295_ (
    .A1(_10549_),
    .A2(_10559_),
    .ZN(_10563_)
  );
  INV_X1 _20296_ (
    .A(_10563_),
    .ZN(_10564_)
  );
  AND2_X1 _20297_ (
    .A1(_10562_),
    .A2(_10564_),
    .ZN(_10565_)
  );
  INV_X1 _20298_ (
    .A(_10565_),
    .ZN(_10566_)
  );
  AND2_X1 _20299_ (
    .A1(_10547_),
    .A2(_10565_),
    .ZN(_10567_)
  );
  INV_X1 _20300_ (
    .A(_10567_),
    .ZN(_10568_)
  );
  AND2_X1 _20301_ (
    .A1(_10548_),
    .A2(_10566_),
    .ZN(_10569_)
  );
  INV_X1 _20302_ (
    .A(_10569_),
    .ZN(_10570_)
  );
  AND2_X1 _20303_ (
    .A1(_10568_),
    .A2(_10570_),
    .ZN(_10571_)
  );
  INV_X1 _20304_ (
    .A(_10571_),
    .ZN(_10573_)
  );
  AND2_X1 _20305_ (
    .A1(_10393_),
    .A2(_10571_),
    .ZN(_10574_)
  );
  INV_X1 _20306_ (
    .A(_10574_),
    .ZN(_10575_)
  );
  AND2_X1 _20307_ (
    .A1(_10392_),
    .A2(_10573_),
    .ZN(_10576_)
  );
  INV_X1 _20308_ (
    .A(_10576_),
    .ZN(_10577_)
  );
  AND2_X1 _20309_ (
    .A1(_10575_),
    .A2(_10577_),
    .ZN(_10578_)
  );
  INV_X1 _20310_ (
    .A(_10578_),
    .ZN(_10579_)
  );
  AND2_X1 _20311_ (
    .A1(_10274_),
    .A2(_10281_),
    .ZN(_10580_)
  );
  INV_X1 _20312_ (
    .A(_10580_),
    .ZN(_10581_)
  );
  AND2_X1 _20313_ (
    .A1(_07804_),
    .A2(_10581_),
    .ZN(_10582_)
  );
  INV_X1 _20314_ (
    .A(_10582_),
    .ZN(_10584_)
  );
  AND2_X1 _20315_ (
    .A1(_07805_),
    .A2(_10580_),
    .ZN(_10585_)
  );
  INV_X1 _20316_ (
    .A(_10585_),
    .ZN(_10586_)
  );
  AND2_X1 _20317_ (
    .A1(_10584_),
    .A2(_10586_),
    .ZN(_10587_)
  );
  INV_X1 _20318_ (
    .A(_10587_),
    .ZN(_10588_)
  );
  AND2_X1 _20319_ (
    .A1(_08107_),
    .A2(_10587_),
    .ZN(_10589_)
  );
  INV_X1 _20320_ (
    .A(_10589_),
    .ZN(_10590_)
  );
  AND2_X1 _20321_ (
    .A1(_08106_),
    .A2(_10588_),
    .ZN(_10591_)
  );
  INV_X1 _20322_ (
    .A(_10591_),
    .ZN(_10592_)
  );
  AND2_X1 _20323_ (
    .A1(_10590_),
    .A2(_10592_),
    .ZN(_10593_)
  );
  INV_X1 _20324_ (
    .A(_10593_),
    .ZN(_10595_)
  );
  AND2_X1 _20325_ (
    .A1(_10578_),
    .A2(_10593_),
    .ZN(_10596_)
  );
  INV_X1 _20326_ (
    .A(_10596_),
    .ZN(_10597_)
  );
  AND2_X1 _20327_ (
    .A1(_10579_),
    .A2(_10595_),
    .ZN(_10598_)
  );
  INV_X1 _20328_ (
    .A(_10598_),
    .ZN(_10599_)
  );
  AND2_X1 _20329_ (
    .A1(_10597_),
    .A2(_10599_),
    .ZN(_10600_)
  );
  INV_X1 _20330_ (
    .A(_10600_),
    .ZN(_10601_)
  );
  AND2_X1 _20331_ (
    .A1(_10391_),
    .A2(_10600_),
    .ZN(_10602_)
  );
  INV_X1 _20332_ (
    .A(_10602_),
    .ZN(_10603_)
  );
  AND2_X1 _20333_ (
    .A1(_10390_),
    .A2(_10601_),
    .ZN(_10604_)
  );
  INV_X1 _20334_ (
    .A(_10604_),
    .ZN(_10606_)
  );
  AND2_X1 _20335_ (
    .A1(_10603_),
    .A2(_10606_),
    .ZN(_10607_)
  );
  INV_X1 _20336_ (
    .A(_10607_),
    .ZN(_10608_)
  );
  AND2_X1 _20337_ (
    .A1(_10389_),
    .A2(_10607_),
    .ZN(_10609_)
  );
  INV_X1 _20338_ (
    .A(_10609_),
    .ZN(_10610_)
  );
  AND2_X1 _20339_ (
    .A1(_10388_),
    .A2(_10608_),
    .ZN(_10611_)
  );
  INV_X1 _20340_ (
    .A(_10611_),
    .ZN(_10612_)
  );
  AND2_X1 _20341_ (
    .A1(_10610_),
    .A2(_10612_),
    .ZN(_10613_)
  );
  INV_X1 _20342_ (
    .A(_10613_),
    .ZN(_10614_)
  );
  AND2_X1 _20343_ (
    .A1(_10387_),
    .A2(_10613_),
    .ZN(_10615_)
  );
  INV_X1 _20344_ (
    .A(_10615_),
    .ZN(_10617_)
  );
  AND2_X1 _20345_ (
    .A1(_10386_),
    .A2(_10614_),
    .ZN(_10618_)
  );
  INV_X1 _20346_ (
    .A(_10618_),
    .ZN(_10619_)
  );
  AND2_X1 _20347_ (
    .A1(_10617_),
    .A2(_10619_),
    .ZN(_10620_)
  );
  INV_X1 _20348_ (
    .A(_10620_),
    .ZN(_10621_)
  );
  AND2_X1 _20349_ (
    .A1(_10335_),
    .A2(_10620_),
    .ZN(_10622_)
  );
  INV_X1 _20350_ (
    .A(_10622_),
    .ZN(_10623_)
  );
  AND2_X1 _20351_ (
    .A1(_10336_),
    .A2(_10621_),
    .ZN(_10624_)
  );
  INV_X1 _20352_ (
    .A(_10624_),
    .ZN(_10625_)
  );
  AND2_X1 _20353_ (
    .A1(_10623_),
    .A2(_10625_),
    .ZN(_10626_)
  );
  INV_X1 _20354_ (
    .A(_10626_),
    .ZN(_10628_)
  );
  AND2_X1 _20355_ (
    .A1(_10094_),
    .A2(_10343_),
    .ZN(_10629_)
  );
  INV_X1 _20356_ (
    .A(_10629_),
    .ZN(_10630_)
  );
  AND2_X1 _20357_ (
    .A1(_10345_),
    .A2(_10630_),
    .ZN(_10631_)
  );
  AND2_X1 _20358_ (
    .A1(_10343_),
    .A2(_10351_),
    .ZN(_10632_)
  );
  AND2_X1 _20359_ (
    .A1(_10626_),
    .A2(_10631_),
    .ZN(_10633_)
  );
  INV_X1 _20360_ (
    .A(_10633_),
    .ZN(_10634_)
  );
  AND2_X1 _20361_ (
    .A1(_10628_),
    .A2(_10632_),
    .ZN(_10635_)
  );
  INV_X1 _20362_ (
    .A(_10635_),
    .ZN(_10636_)
  );
  AND2_X1 _20363_ (
    .A1(_10634_),
    .A2(_10636_),
    .ZN(_10637_)
  );
  INV_X1 _20364_ (
    .A(_10637_),
    .ZN(_10639_)
  );
  AND2_X1 _20365_ (
    .A1(remainder[65]),
    .A2(_10637_),
    .ZN(_10640_)
  );
  INV_X1 _20366_ (
    .A(_10640_),
    .ZN(_10641_)
  );
  AND2_X1 _20367_ (
    .A1(_04404_),
    .A2(_10639_),
    .ZN(_10642_)
  );
  INV_X1 _20368_ (
    .A(_10642_),
    .ZN(_10643_)
  );
  AND2_X1 _20369_ (
    .A1(_10641_),
    .A2(_10643_),
    .ZN(_10644_)
  );
  INV_X1 _20370_ (
    .A(_10644_),
    .ZN(_10645_)
  );
  AND2_X1 _20371_ (
    .A1(_10384_),
    .A2(_10644_),
    .ZN(_10646_)
  );
  INV_X1 _20372_ (
    .A(_10646_),
    .ZN(_10647_)
  );
  AND2_X1 _20373_ (
    .A1(_10383_),
    .A2(_10645_),
    .ZN(_10648_)
  );
  INV_X1 _20374_ (
    .A(_10648_),
    .ZN(_10650_)
  );
  AND2_X1 _20375_ (
    .A1(_02082_),
    .A2(_10650_),
    .ZN(_10651_)
  );
  AND2_X1 _20376_ (
    .A1(_10647_),
    .A2(_10651_),
    .ZN(_10652_)
  );
  INV_X1 _20377_ (
    .A(_10652_),
    .ZN(_10653_)
  );
  AND2_X1 _20378_ (
    .A1(remainder[61]),
    .A2(_02077_),
    .ZN(_10654_)
  );
  INV_X1 _20379_ (
    .A(_10654_),
    .ZN(_10655_)
  );
  AND2_X1 _20380_ (
    .A1(_04459_),
    .A2(_10451_),
    .ZN(_10656_)
  );
  INV_X1 _20381_ (
    .A(_10656_),
    .ZN(_10657_)
  );
  AND2_X1 _20382_ (
    .A1(_10462_),
    .A2(_02018_),
    .ZN(_10658_)
  );
  INV_X1 _20383_ (
    .A(_10658_),
    .ZN(_10659_)
  );
  AND2_X1 _20384_ (
    .A1(_05983_),
    .A2(_10659_),
    .ZN(_10661_)
  );
  AND2_X1 _20385_ (
    .A1(_10657_),
    .A2(_10661_),
    .ZN(_10662_)
  );
  INV_X1 _20386_ (
    .A(_10662_),
    .ZN(_10663_)
  );
  AND2_X1 _20387_ (
    .A1(_10655_),
    .A2(_10663_),
    .ZN(_10664_)
  );
  AND2_X1 _20388_ (
    .A1(_10653_),
    .A2(_10664_),
    .ZN(_10665_)
  );
  INV_X1 _20389_ (
    .A(_10665_),
    .ZN(_10666_)
  );
  AND2_X1 _20390_ (
    .A1(_06201_),
    .A2(_10666_),
    .ZN(_00082_)
  );
  AND2_X1 _20391_ (
    .A1(_10641_),
    .A2(_10647_),
    .ZN(_10667_)
  );
  INV_X1 _20392_ (
    .A(_10667_),
    .ZN(_10668_)
  );
  AND2_X1 _20393_ (
    .A1(_10623_),
    .A2(_10634_),
    .ZN(_10669_)
  );
  INV_X1 _20394_ (
    .A(_10669_),
    .ZN(_10671_)
  );
  AND2_X1 _20395_ (
    .A1(_10603_),
    .A2(_10610_),
    .ZN(_10672_)
  );
  INV_X1 _20396_ (
    .A(_10672_),
    .ZN(_10673_)
  );
  AND2_X1 _20397_ (
    .A1(_10584_),
    .A2(_10590_),
    .ZN(_10674_)
  );
  INV_X1 _20398_ (
    .A(_10674_),
    .ZN(_10675_)
  );
  AND2_X1 _20399_ (
    .A1(_10575_),
    .A2(_10597_),
    .ZN(_10676_)
  );
  INV_X1 _20400_ (
    .A(_10676_),
    .ZN(_10677_)
  );
  AND2_X1 _20401_ (
    .A1(_10544_),
    .A2(_10568_),
    .ZN(_10678_)
  );
  INV_X1 _20402_ (
    .A(_10678_),
    .ZN(_10679_)
  );
  AND2_X1 _20403_ (
    .A1(_10482_),
    .A2(_10537_),
    .ZN(_10680_)
  );
  INV_X1 _20404_ (
    .A(_10680_),
    .ZN(_10682_)
  );
  AND2_X1 _20405_ (
    .A1(_10109_),
    .A2(_10465_),
    .ZN(_10683_)
  );
  INV_X1 _20406_ (
    .A(_10683_),
    .ZN(_10684_)
  );
  AND2_X1 _20407_ (
    .A1(_10476_),
    .A2(_10684_),
    .ZN(_10685_)
  );
  INV_X1 _20408_ (
    .A(_10685_),
    .ZN(_10686_)
  );
  AND2_X1 _20409_ (
    .A1(_03249_),
    .A2(_10464_),
    .ZN(_10687_)
  );
  INV_X1 _20410_ (
    .A(_10687_),
    .ZN(_10688_)
  );
  AND2_X1 _20411_ (
    .A1(_09546_),
    .A2(_10459_),
    .ZN(_10689_)
  );
  INV_X1 _20412_ (
    .A(_10689_),
    .ZN(_10690_)
  );
  AND2_X1 _20413_ (
    .A1(_09797_),
    .A2(_10125_),
    .ZN(_10691_)
  );
  INV_X1 _20414_ (
    .A(_10691_),
    .ZN(_10693_)
  );
  AND2_X1 _20415_ (
    .A1(_09798_),
    .A2(_10126_),
    .ZN(_10694_)
  );
  INV_X1 _20416_ (
    .A(_10694_),
    .ZN(_10695_)
  );
  AND2_X1 _20417_ (
    .A1(_10693_),
    .A2(_10695_),
    .ZN(_10696_)
  );
  INV_X1 _20418_ (
    .A(_10696_),
    .ZN(_10697_)
  );
  AND2_X1 _20419_ (
    .A1(_10690_),
    .A2(_10696_),
    .ZN(_10698_)
  );
  INV_X1 _20420_ (
    .A(_10698_),
    .ZN(_10699_)
  );
  AND2_X1 _20421_ (
    .A1(_10689_),
    .A2(_10697_),
    .ZN(_10700_)
  );
  INV_X1 _20422_ (
    .A(_10700_),
    .ZN(_10701_)
  );
  AND2_X1 _20423_ (
    .A1(_10699_),
    .A2(_10701_),
    .ZN(_10702_)
  );
  INV_X1 _20424_ (
    .A(_10702_),
    .ZN(_10704_)
  );
  AND2_X1 _20425_ (
    .A1(_09784_),
    .A2(_10702_),
    .ZN(_10705_)
  );
  INV_X1 _20426_ (
    .A(_10705_),
    .ZN(_10706_)
  );
  AND2_X1 _20427_ (
    .A1(_09785_),
    .A2(_10704_),
    .ZN(_10707_)
  );
  INV_X1 _20428_ (
    .A(_10707_),
    .ZN(_10708_)
  );
  AND2_X1 _20429_ (
    .A1(_10706_),
    .A2(_10708_),
    .ZN(_10709_)
  );
  INV_X1 _20430_ (
    .A(_10709_),
    .ZN(_10710_)
  );
  AND2_X1 _20431_ (
    .A1(_10687_),
    .A2(_10709_),
    .ZN(_10711_)
  );
  INV_X1 _20432_ (
    .A(_10711_),
    .ZN(_10712_)
  );
  AND2_X1 _20433_ (
    .A1(_10688_),
    .A2(_10710_),
    .ZN(_10713_)
  );
  INV_X1 _20434_ (
    .A(_10713_),
    .ZN(_10714_)
  );
  AND2_X1 _20435_ (
    .A1(_10712_),
    .A2(_10714_),
    .ZN(_10715_)
  );
  INV_X1 _20436_ (
    .A(_10715_),
    .ZN(_10716_)
  );
  AND2_X1 _20437_ (
    .A1(_10420_),
    .A2(_10444_),
    .ZN(_10717_)
  );
  INV_X1 _20438_ (
    .A(_10717_),
    .ZN(_10718_)
  );
  AND2_X1 _20439_ (
    .A1(_10409_),
    .A2(_10413_),
    .ZN(_10719_)
  );
  INV_X1 _20440_ (
    .A(_10719_),
    .ZN(_10720_)
  );
  AND2_X1 _20441_ (
    .A1(divisor[31]),
    .A2(remainder[6]),
    .ZN(_10721_)
  );
  INV_X1 _20442_ (
    .A(_10721_),
    .ZN(_10722_)
  );
  AND2_X1 _20443_ (
    .A1(divisor[32]),
    .A2(remainder[5]),
    .ZN(_10723_)
  );
  INV_X1 _20444_ (
    .A(_10723_),
    .ZN(_10724_)
  );
  AND2_X1 _20445_ (
    .A1(remainder[5]),
    .A2(_10405_),
    .ZN(_10725_)
  );
  INV_X1 _20446_ (
    .A(_10725_),
    .ZN(_10726_)
  );
  MUX2_X1 _20447_ (
    .A(_10405_),
    .B(_05116_),
    .S(_10723_),
    .Z(_10727_)
  );
  MUX2_X1 _20448_ (
    .A(remainder[4]),
    .B(_10406_),
    .S(_10724_),
    .Z(_10728_)
  );
  AND2_X1 _20449_ (
    .A1(_10721_),
    .A2(_10727_),
    .ZN(_10729_)
  );
  INV_X1 _20450_ (
    .A(_10729_),
    .ZN(_10730_)
  );
  AND2_X1 _20451_ (
    .A1(_10722_),
    .A2(_10728_),
    .ZN(_10731_)
  );
  INV_X1 _20452_ (
    .A(_10731_),
    .ZN(_10732_)
  );
  AND2_X1 _20453_ (
    .A1(_10730_),
    .A2(_10732_),
    .ZN(_10733_)
  );
  INV_X1 _20454_ (
    .A(_10733_),
    .ZN(_10734_)
  );
  AND2_X1 _20455_ (
    .A1(_10720_),
    .A2(_10733_),
    .ZN(_10735_)
  );
  INV_X1 _20456_ (
    .A(_10735_),
    .ZN(_10736_)
  );
  AND2_X1 _20457_ (
    .A1(_10719_),
    .A2(_10734_),
    .ZN(_10737_)
  );
  INV_X1 _20458_ (
    .A(_10737_),
    .ZN(_10738_)
  );
  AND2_X1 _20459_ (
    .A1(_10736_),
    .A2(_10738_),
    .ZN(_10739_)
  );
  INV_X1 _20460_ (
    .A(_10739_),
    .ZN(_10740_)
  );
  AND2_X1 _20461_ (
    .A1(remainder[32]),
    .A2(divisor[30]),
    .ZN(_10741_)
  );
  AND2_X1 _20462_ (
    .A1(remainder[32]),
    .A2(divisor[29]),
    .ZN(_10742_)
  );
  INV_X1 _20463_ (
    .A(_10742_),
    .ZN(_10743_)
  );
  AND2_X1 _20464_ (
    .A1(divisor[30]),
    .A2(_10742_),
    .ZN(_10744_)
  );
  INV_X1 _20465_ (
    .A(_10744_),
    .ZN(_10745_)
  );
  AND2_X1 _20466_ (
    .A1(_10427_),
    .A2(_10742_),
    .ZN(_10746_)
  );
  INV_X1 _20467_ (
    .A(_10746_),
    .ZN(_10747_)
  );
  AND2_X1 _20468_ (
    .A1(_10428_),
    .A2(_10743_),
    .ZN(_10748_)
  );
  INV_X1 _20469_ (
    .A(_10748_),
    .ZN(_10749_)
  );
  AND2_X1 _20470_ (
    .A1(_10747_),
    .A2(_10749_),
    .ZN(_10750_)
  );
  INV_X1 _20471_ (
    .A(_10750_),
    .ZN(_10751_)
  );
  AND2_X1 _20472_ (
    .A1(_08005_),
    .A2(_10750_),
    .ZN(_10752_)
  );
  INV_X1 _20473_ (
    .A(_10752_),
    .ZN(_10753_)
  );
  AND2_X1 _20474_ (
    .A1(_08007_),
    .A2(_10751_),
    .ZN(_10754_)
  );
  INV_X1 _20475_ (
    .A(_10754_),
    .ZN(_10755_)
  );
  AND2_X1 _20476_ (
    .A1(_10753_),
    .A2(_10755_),
    .ZN(_10756_)
  );
  INV_X1 _20477_ (
    .A(_10756_),
    .ZN(_10757_)
  );
  AND2_X1 _20478_ (
    .A1(_10739_),
    .A2(_10756_),
    .ZN(_10758_)
  );
  INV_X1 _20479_ (
    .A(_10758_),
    .ZN(_10759_)
  );
  AND2_X1 _20480_ (
    .A1(_10740_),
    .A2(_10757_),
    .ZN(_10760_)
  );
  INV_X1 _20481_ (
    .A(_10760_),
    .ZN(_10761_)
  );
  AND2_X1 _20482_ (
    .A1(_10759_),
    .A2(_10761_),
    .ZN(_10762_)
  );
  INV_X1 _20483_ (
    .A(_10762_),
    .ZN(_10763_)
  );
  AND2_X1 _20484_ (
    .A1(_10456_),
    .A2(_10762_),
    .ZN(_10764_)
  );
  INV_X1 _20485_ (
    .A(_10764_),
    .ZN(_10765_)
  );
  AND2_X1 _20486_ (
    .A1(_10457_),
    .A2(_10763_),
    .ZN(_10766_)
  );
  INV_X1 _20487_ (
    .A(_10766_),
    .ZN(_10767_)
  );
  AND2_X1 _20488_ (
    .A1(_10765_),
    .A2(_10767_),
    .ZN(_10768_)
  );
  INV_X1 _20489_ (
    .A(_10768_),
    .ZN(_10769_)
  );
  AND2_X1 _20490_ (
    .A1(_10718_),
    .A2(_10768_),
    .ZN(_10770_)
  );
  INV_X1 _20491_ (
    .A(_10770_),
    .ZN(_10771_)
  );
  AND2_X1 _20492_ (
    .A1(_10717_),
    .A2(_10769_),
    .ZN(_10772_)
  );
  INV_X1 _20493_ (
    .A(_10772_),
    .ZN(_10773_)
  );
  AND2_X1 _20494_ (
    .A1(_10771_),
    .A2(_10773_),
    .ZN(_10775_)
  );
  INV_X1 _20495_ (
    .A(_10775_),
    .ZN(_10776_)
  );
  AND2_X1 _20496_ (
    .A1(_10715_),
    .A2(_10775_),
    .ZN(_10777_)
  );
  INV_X1 _20497_ (
    .A(_10777_),
    .ZN(_10778_)
  );
  AND2_X1 _20498_ (
    .A1(_10716_),
    .A2(_10776_),
    .ZN(_10779_)
  );
  INV_X1 _20499_ (
    .A(_10779_),
    .ZN(_10780_)
  );
  AND2_X1 _20500_ (
    .A1(_10778_),
    .A2(_10780_),
    .ZN(_10781_)
  );
  INV_X1 _20501_ (
    .A(_10781_),
    .ZN(_10782_)
  );
  AND2_X1 _20502_ (
    .A1(_10686_),
    .A2(_10781_),
    .ZN(_10783_)
  );
  INV_X1 _20503_ (
    .A(_10783_),
    .ZN(_10784_)
  );
  AND2_X1 _20504_ (
    .A1(_10685_),
    .A2(_10782_),
    .ZN(_10786_)
  );
  INV_X1 _20505_ (
    .A(_10786_),
    .ZN(_10787_)
  );
  AND2_X1 _20506_ (
    .A1(_10784_),
    .A2(_10787_),
    .ZN(_10788_)
  );
  INV_X1 _20507_ (
    .A(_10788_),
    .ZN(_10789_)
  );
  AND2_X1 _20508_ (
    .A1(_10511_),
    .A2(_10518_),
    .ZN(_10790_)
  );
  INV_X1 _20509_ (
    .A(_10790_),
    .ZN(_10791_)
  );
  AND2_X1 _20510_ (
    .A1(_10498_),
    .A2(_10504_),
    .ZN(_10792_)
  );
  INV_X1 _20511_ (
    .A(_10792_),
    .ZN(_10793_)
  );
  AND2_X1 _20512_ (
    .A1(_10431_),
    .A2(_10437_),
    .ZN(_10794_)
  );
  INV_X1 _20513_ (
    .A(_10794_),
    .ZN(_10795_)
  );
  AND2_X1 _20514_ (
    .A1(_10203_),
    .A2(_10795_),
    .ZN(_10797_)
  );
  INV_X1 _20515_ (
    .A(_10797_),
    .ZN(_10798_)
  );
  AND2_X1 _20516_ (
    .A1(_10204_),
    .A2(_10794_),
    .ZN(_10799_)
  );
  INV_X1 _20517_ (
    .A(_10799_),
    .ZN(_10800_)
  );
  AND2_X1 _20518_ (
    .A1(_10798_),
    .A2(_10800_),
    .ZN(_10801_)
  );
  INV_X1 _20519_ (
    .A(_10801_),
    .ZN(_10802_)
  );
  AND2_X1 _20520_ (
    .A1(_10493_),
    .A2(_10801_),
    .ZN(_10803_)
  );
  INV_X1 _20521_ (
    .A(_10803_),
    .ZN(_10804_)
  );
  AND2_X1 _20522_ (
    .A1(_10492_),
    .A2(_10802_),
    .ZN(_10805_)
  );
  INV_X1 _20523_ (
    .A(_10805_),
    .ZN(_10806_)
  );
  AND2_X1 _20524_ (
    .A1(_10804_),
    .A2(_10806_),
    .ZN(_10807_)
  );
  INV_X1 _20525_ (
    .A(_10807_),
    .ZN(_10808_)
  );
  AND2_X1 _20526_ (
    .A1(_10793_),
    .A2(_10807_),
    .ZN(_10809_)
  );
  INV_X1 _20527_ (
    .A(_10809_),
    .ZN(_10810_)
  );
  AND2_X1 _20528_ (
    .A1(_10792_),
    .A2(_10808_),
    .ZN(_10811_)
  );
  INV_X1 _20529_ (
    .A(_10811_),
    .ZN(_10812_)
  );
  AND2_X1 _20530_ (
    .A1(_10810_),
    .A2(_10812_),
    .ZN(_10813_)
  );
  INV_X1 _20531_ (
    .A(_10813_),
    .ZN(_10814_)
  );
  AND2_X1 _20532_ (
    .A1(_09521_),
    .A2(_10813_),
    .ZN(_10815_)
  );
  INV_X1 _20533_ (
    .A(_10815_),
    .ZN(_10816_)
  );
  AND2_X1 _20534_ (
    .A1(_09522_),
    .A2(_10814_),
    .ZN(_10818_)
  );
  INV_X1 _20535_ (
    .A(_10818_),
    .ZN(_10819_)
  );
  AND2_X1 _20536_ (
    .A1(_10816_),
    .A2(_10819_),
    .ZN(_10820_)
  );
  INV_X1 _20537_ (
    .A(_10820_),
    .ZN(_10821_)
  );
  AND2_X1 _20538_ (
    .A1(_10449_),
    .A2(_10820_),
    .ZN(_10822_)
  );
  INV_X1 _20539_ (
    .A(_10822_),
    .ZN(_10823_)
  );
  AND2_X1 _20540_ (
    .A1(_10450_),
    .A2(_10821_),
    .ZN(_10824_)
  );
  INV_X1 _20541_ (
    .A(_10824_),
    .ZN(_10825_)
  );
  AND2_X1 _20542_ (
    .A1(_10823_),
    .A2(_10825_),
    .ZN(_10826_)
  );
  INV_X1 _20543_ (
    .A(_10826_),
    .ZN(_10827_)
  );
  AND2_X1 _20544_ (
    .A1(_10791_),
    .A2(_10826_),
    .ZN(_10829_)
  );
  INV_X1 _20545_ (
    .A(_10829_),
    .ZN(_10830_)
  );
  AND2_X1 _20546_ (
    .A1(_10790_),
    .A2(_10827_),
    .ZN(_10831_)
  );
  INV_X1 _20547_ (
    .A(_10831_),
    .ZN(_10832_)
  );
  AND2_X1 _20548_ (
    .A1(_10830_),
    .A2(_10832_),
    .ZN(_10833_)
  );
  INV_X1 _20549_ (
    .A(_10833_),
    .ZN(_10834_)
  );
  AND2_X1 _20550_ (
    .A1(_10788_),
    .A2(_10833_),
    .ZN(_10835_)
  );
  INV_X1 _20551_ (
    .A(_10835_),
    .ZN(_10836_)
  );
  AND2_X1 _20552_ (
    .A1(_10789_),
    .A2(_10834_),
    .ZN(_10837_)
  );
  INV_X1 _20553_ (
    .A(_10837_),
    .ZN(_10838_)
  );
  AND2_X1 _20554_ (
    .A1(_10836_),
    .A2(_10838_),
    .ZN(_10840_)
  );
  INV_X1 _20555_ (
    .A(_10840_),
    .ZN(_10841_)
  );
  AND2_X1 _20556_ (
    .A1(_10682_),
    .A2(_10840_),
    .ZN(_10842_)
  );
  INV_X1 _20557_ (
    .A(_10842_),
    .ZN(_10843_)
  );
  AND2_X1 _20558_ (
    .A1(_10680_),
    .A2(_10841_),
    .ZN(_10844_)
  );
  INV_X1 _20559_ (
    .A(_10844_),
    .ZN(_10845_)
  );
  AND2_X1 _20560_ (
    .A1(_10843_),
    .A2(_10845_),
    .ZN(_10846_)
  );
  INV_X1 _20561_ (
    .A(_10846_),
    .ZN(_10847_)
  );
  AND2_X1 _20562_ (
    .A1(_10524_),
    .A2(_10531_),
    .ZN(_10848_)
  );
  INV_X1 _20563_ (
    .A(_10848_),
    .ZN(_10849_)
  );
  AND2_X1 _20564_ (
    .A1(_10271_),
    .A2(_10849_),
    .ZN(_10851_)
  );
  INV_X1 _20565_ (
    .A(_10851_),
    .ZN(_10852_)
  );
  AND2_X1 _20566_ (
    .A1(_10272_),
    .A2(_10848_),
    .ZN(_10853_)
  );
  INV_X1 _20567_ (
    .A(_10853_),
    .ZN(_10854_)
  );
  AND2_X1 _20568_ (
    .A1(_10852_),
    .A2(_10854_),
    .ZN(_10855_)
  );
  INV_X1 _20569_ (
    .A(_10855_),
    .ZN(_10856_)
  );
  AND2_X1 _20570_ (
    .A1(_10551_),
    .A2(_10855_),
    .ZN(_10857_)
  );
  INV_X1 _20571_ (
    .A(_10857_),
    .ZN(_10858_)
  );
  AND2_X1 _20572_ (
    .A1(_10549_),
    .A2(_10856_),
    .ZN(_10859_)
  );
  INV_X1 _20573_ (
    .A(_10859_),
    .ZN(_10860_)
  );
  AND2_X1 _20574_ (
    .A1(_10858_),
    .A2(_10860_),
    .ZN(_10862_)
  );
  INV_X1 _20575_ (
    .A(_10862_),
    .ZN(_10863_)
  );
  AND2_X1 _20576_ (
    .A1(_10846_),
    .A2(_10862_),
    .ZN(_10864_)
  );
  INV_X1 _20577_ (
    .A(_10864_),
    .ZN(_10865_)
  );
  AND2_X1 _20578_ (
    .A1(_10847_),
    .A2(_10863_),
    .ZN(_10866_)
  );
  INV_X1 _20579_ (
    .A(_10866_),
    .ZN(_10867_)
  );
  AND2_X1 _20580_ (
    .A1(_10865_),
    .A2(_10867_),
    .ZN(_10868_)
  );
  INV_X1 _20581_ (
    .A(_10868_),
    .ZN(_10869_)
  );
  AND2_X1 _20582_ (
    .A1(_10679_),
    .A2(_10868_),
    .ZN(_10870_)
  );
  INV_X1 _20583_ (
    .A(_10870_),
    .ZN(_10871_)
  );
  AND2_X1 _20584_ (
    .A1(_10678_),
    .A2(_10869_),
    .ZN(_10873_)
  );
  INV_X1 _20585_ (
    .A(_10873_),
    .ZN(_10874_)
  );
  AND2_X1 _20586_ (
    .A1(_10871_),
    .A2(_10874_),
    .ZN(_10875_)
  );
  INV_X1 _20587_ (
    .A(_10875_),
    .ZN(_10876_)
  );
  AND2_X1 _20588_ (
    .A1(_10555_),
    .A2(_10562_),
    .ZN(_10877_)
  );
  INV_X1 _20589_ (
    .A(_10877_),
    .ZN(_10878_)
  );
  AND2_X1 _20590_ (
    .A1(_07804_),
    .A2(_10878_),
    .ZN(_10879_)
  );
  INV_X1 _20591_ (
    .A(_10879_),
    .ZN(_10880_)
  );
  AND2_X1 _20592_ (
    .A1(_07805_),
    .A2(_10877_),
    .ZN(_10881_)
  );
  INV_X1 _20593_ (
    .A(_10881_),
    .ZN(_10882_)
  );
  AND2_X1 _20594_ (
    .A1(_10880_),
    .A2(_10882_),
    .ZN(_10884_)
  );
  INV_X1 _20595_ (
    .A(_10884_),
    .ZN(_10885_)
  );
  AND2_X1 _20596_ (
    .A1(_08107_),
    .A2(_10884_),
    .ZN(_10886_)
  );
  INV_X1 _20597_ (
    .A(_10886_),
    .ZN(_10887_)
  );
  AND2_X1 _20598_ (
    .A1(_08106_),
    .A2(_10885_),
    .ZN(_10888_)
  );
  INV_X1 _20599_ (
    .A(_10888_),
    .ZN(_10889_)
  );
  AND2_X1 _20600_ (
    .A1(_10887_),
    .A2(_10889_),
    .ZN(_10890_)
  );
  INV_X1 _20601_ (
    .A(_10890_),
    .ZN(_10891_)
  );
  AND2_X1 _20602_ (
    .A1(_10875_),
    .A2(_10890_),
    .ZN(_10892_)
  );
  INV_X1 _20603_ (
    .A(_10892_),
    .ZN(_10893_)
  );
  AND2_X1 _20604_ (
    .A1(_10876_),
    .A2(_10891_),
    .ZN(_10894_)
  );
  INV_X1 _20605_ (
    .A(_10894_),
    .ZN(_10895_)
  );
  AND2_X1 _20606_ (
    .A1(_10893_),
    .A2(_10895_),
    .ZN(_10896_)
  );
  INV_X1 _20607_ (
    .A(_10896_),
    .ZN(_10897_)
  );
  AND2_X1 _20608_ (
    .A1(_10677_),
    .A2(_10896_),
    .ZN(_10898_)
  );
  INV_X1 _20609_ (
    .A(_10898_),
    .ZN(_10899_)
  );
  AND2_X1 _20610_ (
    .A1(_10676_),
    .A2(_10897_),
    .ZN(_10900_)
  );
  INV_X1 _20611_ (
    .A(_10900_),
    .ZN(_10901_)
  );
  AND2_X1 _20612_ (
    .A1(_10899_),
    .A2(_10901_),
    .ZN(_10902_)
  );
  INV_X1 _20613_ (
    .A(_10902_),
    .ZN(_10903_)
  );
  AND2_X1 _20614_ (
    .A1(_10675_),
    .A2(_10902_),
    .ZN(_10905_)
  );
  INV_X1 _20615_ (
    .A(_10905_),
    .ZN(_10906_)
  );
  AND2_X1 _20616_ (
    .A1(_10674_),
    .A2(_10903_),
    .ZN(_10907_)
  );
  INV_X1 _20617_ (
    .A(_10907_),
    .ZN(_10908_)
  );
  AND2_X1 _20618_ (
    .A1(_10906_),
    .A2(_10908_),
    .ZN(_10909_)
  );
  INV_X1 _20619_ (
    .A(_10909_),
    .ZN(_10910_)
  );
  AND2_X1 _20620_ (
    .A1(_10673_),
    .A2(_10909_),
    .ZN(_10911_)
  );
  INV_X1 _20621_ (
    .A(_10911_),
    .ZN(_10912_)
  );
  AND2_X1 _20622_ (
    .A1(_10672_),
    .A2(_10910_),
    .ZN(_10913_)
  );
  INV_X1 _20623_ (
    .A(_10913_),
    .ZN(_10914_)
  );
  AND2_X1 _20624_ (
    .A1(_10912_),
    .A2(_10914_),
    .ZN(_10916_)
  );
  INV_X1 _20625_ (
    .A(_10916_),
    .ZN(_10917_)
  );
  AND2_X1 _20626_ (
    .A1(_10615_),
    .A2(_10916_),
    .ZN(_10918_)
  );
  INV_X1 _20627_ (
    .A(_10918_),
    .ZN(_10919_)
  );
  AND2_X1 _20628_ (
    .A1(_10617_),
    .A2(_10917_),
    .ZN(_10920_)
  );
  INV_X1 _20629_ (
    .A(_10920_),
    .ZN(_10921_)
  );
  AND2_X1 _20630_ (
    .A1(_10919_),
    .A2(_10921_),
    .ZN(_10922_)
  );
  INV_X1 _20631_ (
    .A(_10922_),
    .ZN(_10923_)
  );
  AND2_X1 _20632_ (
    .A1(_10669_),
    .A2(_10923_),
    .ZN(_10924_)
  );
  INV_X1 _20633_ (
    .A(_10924_),
    .ZN(_10925_)
  );
  AND2_X1 _20634_ (
    .A1(_10671_),
    .A2(_10922_),
    .ZN(_10927_)
  );
  INV_X1 _20635_ (
    .A(_10927_),
    .ZN(_10928_)
  );
  AND2_X1 _20636_ (
    .A1(_10925_),
    .A2(_10928_),
    .ZN(_10929_)
  );
  INV_X1 _20637_ (
    .A(_10929_),
    .ZN(_10930_)
  );
  AND2_X1 _20638_ (
    .A1(_04404_),
    .A2(_10930_),
    .ZN(_10931_)
  );
  INV_X1 _20639_ (
    .A(_10931_),
    .ZN(_10932_)
  );
  AND2_X1 _20640_ (
    .A1(remainder[65]),
    .A2(_10929_),
    .ZN(_10933_)
  );
  INV_X1 _20641_ (
    .A(_10933_),
    .ZN(_10934_)
  );
  AND2_X1 _20642_ (
    .A1(_10932_),
    .A2(_10934_),
    .ZN(_10935_)
  );
  INV_X1 _20643_ (
    .A(_10935_),
    .ZN(_10936_)
  );
  AND2_X1 _20644_ (
    .A1(_10668_),
    .A2(_10935_),
    .ZN(_10938_)
  );
  INV_X1 _20645_ (
    .A(_10938_),
    .ZN(_10939_)
  );
  AND2_X1 _20646_ (
    .A1(_10667_),
    .A2(_10936_),
    .ZN(_10940_)
  );
  INV_X1 _20647_ (
    .A(_10940_),
    .ZN(_10941_)
  );
  AND2_X1 _20648_ (
    .A1(_02082_),
    .A2(_10941_),
    .ZN(_10942_)
  );
  AND2_X1 _20649_ (
    .A1(_10939_),
    .A2(_10942_),
    .ZN(_10943_)
  );
  INV_X1 _20650_ (
    .A(_10943_),
    .ZN(_10944_)
  );
  AND2_X1 _20651_ (
    .A1(remainder[62]),
    .A2(_02077_),
    .ZN(_10945_)
  );
  INV_X1 _20652_ (
    .A(_10945_),
    .ZN(_10946_)
  );
  AND2_X1 _20653_ (
    .A1(_04448_),
    .A2(_10451_),
    .ZN(_10947_)
  );
  INV_X1 _20654_ (
    .A(_10947_),
    .ZN(_10949_)
  );
  AND2_X1 _20655_ (
    .A1(_10462_),
    .A2(_02034_),
    .ZN(_10950_)
  );
  INV_X1 _20656_ (
    .A(_10950_),
    .ZN(_10951_)
  );
  AND2_X1 _20657_ (
    .A1(_05983_),
    .A2(_10951_),
    .ZN(_10952_)
  );
  AND2_X1 _20658_ (
    .A1(_10949_),
    .A2(_10952_),
    .ZN(_10953_)
  );
  INV_X1 _20659_ (
    .A(_10953_),
    .ZN(_10954_)
  );
  AND2_X1 _20660_ (
    .A1(_10946_),
    .A2(_10954_),
    .ZN(_10955_)
  );
  AND2_X1 _20661_ (
    .A1(_10944_),
    .A2(_10955_),
    .ZN(_10956_)
  );
  INV_X1 _20662_ (
    .A(_10956_),
    .ZN(_10957_)
  );
  AND2_X1 _20663_ (
    .A1(_06201_),
    .A2(_10957_),
    .ZN(_00083_)
  );
  AND2_X1 _20664_ (
    .A1(_10646_),
    .A2(_10935_),
    .ZN(_10958_)
  );
  INV_X1 _20665_ (
    .A(_10958_),
    .ZN(_10959_)
  );
  AND2_X1 _20666_ (
    .A1(_10641_),
    .A2(_10934_),
    .ZN(_10960_)
  );
  AND2_X1 _20667_ (
    .A1(_10959_),
    .A2(_10960_),
    .ZN(_10961_)
  );
  INV_X1 _20668_ (
    .A(_10961_),
    .ZN(_10962_)
  );
  AND2_X1 _20669_ (
    .A1(_10899_),
    .A2(_10906_),
    .ZN(_10963_)
  );
  INV_X1 _20670_ (
    .A(_10963_),
    .ZN(_10964_)
  );
  AND2_X1 _20671_ (
    .A1(_10880_),
    .A2(_10887_),
    .ZN(_10965_)
  );
  INV_X1 _20672_ (
    .A(_10965_),
    .ZN(_10966_)
  );
  AND2_X1 _20673_ (
    .A1(_10871_),
    .A2(_10893_),
    .ZN(_10967_)
  );
  INV_X1 _20674_ (
    .A(_10967_),
    .ZN(_10969_)
  );
  AND2_X1 _20675_ (
    .A1(_10843_),
    .A2(_10865_),
    .ZN(_10970_)
  );
  INV_X1 _20676_ (
    .A(_10970_),
    .ZN(_10971_)
  );
  AND2_X1 _20677_ (
    .A1(_10784_),
    .A2(_10836_),
    .ZN(_10972_)
  );
  INV_X1 _20678_ (
    .A(_10972_),
    .ZN(_10973_)
  );
  AND2_X1 _20679_ (
    .A1(_10712_),
    .A2(_10778_),
    .ZN(_10974_)
  );
  INV_X1 _20680_ (
    .A(_10974_),
    .ZN(_10975_)
  );
  AND2_X1 _20681_ (
    .A1(_09796_),
    .A2(_10693_),
    .ZN(_10976_)
  );
  INV_X1 _20682_ (
    .A(_10976_),
    .ZN(_10977_)
  );
  AND2_X1 _20683_ (
    .A1(_10129_),
    .A2(_10405_),
    .ZN(_10978_)
  );
  INV_X1 _20684_ (
    .A(_10978_),
    .ZN(_10980_)
  );
  AND2_X1 _20685_ (
    .A1(_10130_),
    .A2(_10406_),
    .ZN(_10981_)
  );
  INV_X1 _20686_ (
    .A(_10981_),
    .ZN(_10982_)
  );
  AND2_X1 _20687_ (
    .A1(_10980_),
    .A2(_10982_),
    .ZN(_10983_)
  );
  INV_X1 _20688_ (
    .A(_10983_),
    .ZN(_10984_)
  );
  AND2_X1 _20689_ (
    .A1(_10977_),
    .A2(_10983_),
    .ZN(_10985_)
  );
  INV_X1 _20690_ (
    .A(_10985_),
    .ZN(_10986_)
  );
  AND2_X1 _20691_ (
    .A1(_10976_),
    .A2(_10984_),
    .ZN(_10987_)
  );
  INV_X1 _20692_ (
    .A(_10987_),
    .ZN(_10988_)
  );
  AND2_X1 _20693_ (
    .A1(_10986_),
    .A2(_10988_),
    .ZN(_10989_)
  );
  INV_X1 _20694_ (
    .A(_10989_),
    .ZN(_10991_)
  );
  AND2_X1 _20695_ (
    .A1(_10116_),
    .A2(_10989_),
    .ZN(_10992_)
  );
  INV_X1 _20696_ (
    .A(_10992_),
    .ZN(_10993_)
  );
  AND2_X1 _20697_ (
    .A1(_10117_),
    .A2(_10991_),
    .ZN(_10994_)
  );
  INV_X1 _20698_ (
    .A(_10994_),
    .ZN(_10995_)
  );
  AND2_X1 _20699_ (
    .A1(_10993_),
    .A2(_10995_),
    .ZN(_10996_)
  );
  INV_X1 _20700_ (
    .A(_10996_),
    .ZN(_10997_)
  );
  AND2_X1 _20701_ (
    .A1(_10705_),
    .A2(_10996_),
    .ZN(_10998_)
  );
  INV_X1 _20702_ (
    .A(_10998_),
    .ZN(_10999_)
  );
  AND2_X1 _20703_ (
    .A1(_10706_),
    .A2(_10997_),
    .ZN(_11000_)
  );
  INV_X1 _20704_ (
    .A(_11000_),
    .ZN(_11002_)
  );
  AND2_X1 _20705_ (
    .A1(_10999_),
    .A2(_11002_),
    .ZN(_11003_)
  );
  INV_X1 _20706_ (
    .A(_11003_),
    .ZN(_11004_)
  );
  AND2_X1 _20707_ (
    .A1(_10736_),
    .A2(_10759_),
    .ZN(_11005_)
  );
  INV_X1 _20708_ (
    .A(_11005_),
    .ZN(_11006_)
  );
  AND2_X1 _20709_ (
    .A1(_10726_),
    .A2(_10730_),
    .ZN(_11007_)
  );
  INV_X1 _20710_ (
    .A(_11007_),
    .ZN(_11008_)
  );
  AND2_X1 _20711_ (
    .A1(divisor[31]),
    .A2(remainder[7]),
    .ZN(_11009_)
  );
  INV_X1 _20712_ (
    .A(_11009_),
    .ZN(_11010_)
  );
  AND2_X1 _20713_ (
    .A1(divisor[32]),
    .A2(remainder[6]),
    .ZN(_11011_)
  );
  INV_X1 _20714_ (
    .A(_11011_),
    .ZN(_11013_)
  );
  AND2_X1 _20715_ (
    .A1(remainder[5]),
    .A2(_11011_),
    .ZN(_11014_)
  );
  INV_X1 _20716_ (
    .A(_11014_),
    .ZN(_11015_)
  );
  MUX2_X1 _20717_ (
    .A(_11011_),
    .B(_05138_),
    .S(_10723_),
    .Z(_11016_)
  );
  MUX2_X1 _20718_ (
    .A(remainder[6]),
    .B(_11013_),
    .S(_10724_),
    .Z(_11017_)
  );
  AND2_X1 _20719_ (
    .A1(_11009_),
    .A2(_11016_),
    .ZN(_11018_)
  );
  INV_X1 _20720_ (
    .A(_11018_),
    .ZN(_11019_)
  );
  AND2_X1 _20721_ (
    .A1(_11010_),
    .A2(_11017_),
    .ZN(_11020_)
  );
  INV_X1 _20722_ (
    .A(_11020_),
    .ZN(_11021_)
  );
  AND2_X1 _20723_ (
    .A1(_11019_),
    .A2(_11021_),
    .ZN(_11022_)
  );
  INV_X1 _20724_ (
    .A(_11022_),
    .ZN(_11023_)
  );
  AND2_X1 _20725_ (
    .A1(_11008_),
    .A2(_11022_),
    .ZN(_11024_)
  );
  INV_X1 _20726_ (
    .A(_11024_),
    .ZN(_11025_)
  );
  AND2_X1 _20727_ (
    .A1(_11007_),
    .A2(_11023_),
    .ZN(_11026_)
  );
  INV_X1 _20728_ (
    .A(_11026_),
    .ZN(_11027_)
  );
  AND2_X1 _20729_ (
    .A1(_11025_),
    .A2(_11027_),
    .ZN(_11028_)
  );
  INV_X1 _20730_ (
    .A(_11028_),
    .ZN(_11029_)
  );
  MUX2_X1 _20731_ (
    .A(_10742_),
    .B(_05062_),
    .S(_10741_),
    .Z(_11030_)
  );
  AND2_X1 _20732_ (
    .A1(divisor[28]),
    .A2(_11030_),
    .ZN(_11031_)
  );
  INV_X1 _20733_ (
    .A(_11031_),
    .ZN(_11032_)
  );
  MUX2_X1 _20734_ (
    .A(_08005_),
    .B(_05051_),
    .S(_11030_),
    .Z(_11034_)
  );
  MUX2_X1 _20735_ (
    .A(_08007_),
    .B(divisor[28]),
    .S(_11030_),
    .Z(_11035_)
  );
  AND2_X1 _20736_ (
    .A1(_11028_),
    .A2(_11034_),
    .ZN(_11036_)
  );
  INV_X1 _20737_ (
    .A(_11036_),
    .ZN(_11037_)
  );
  AND2_X1 _20738_ (
    .A1(_11029_),
    .A2(_11035_),
    .ZN(_11038_)
  );
  INV_X1 _20739_ (
    .A(_11038_),
    .ZN(_11039_)
  );
  AND2_X1 _20740_ (
    .A1(_11037_),
    .A2(_11039_),
    .ZN(_11040_)
  );
  INV_X1 _20741_ (
    .A(_11040_),
    .ZN(_11041_)
  );
  AND2_X1 _20742_ (
    .A1(_10698_),
    .A2(_11040_),
    .ZN(_11042_)
  );
  INV_X1 _20743_ (
    .A(_11042_),
    .ZN(_11043_)
  );
  AND2_X1 _20744_ (
    .A1(_10699_),
    .A2(_11041_),
    .ZN(_11045_)
  );
  INV_X1 _20745_ (
    .A(_11045_),
    .ZN(_11046_)
  );
  AND2_X1 _20746_ (
    .A1(_11043_),
    .A2(_11046_),
    .ZN(_11047_)
  );
  INV_X1 _20747_ (
    .A(_11047_),
    .ZN(_11048_)
  );
  AND2_X1 _20748_ (
    .A1(_11006_),
    .A2(_11047_),
    .ZN(_11049_)
  );
  INV_X1 _20749_ (
    .A(_11049_),
    .ZN(_11050_)
  );
  AND2_X1 _20750_ (
    .A1(_11005_),
    .A2(_11048_),
    .ZN(_11051_)
  );
  INV_X1 _20751_ (
    .A(_11051_),
    .ZN(_11052_)
  );
  AND2_X1 _20752_ (
    .A1(_11050_),
    .A2(_11052_),
    .ZN(_11053_)
  );
  INV_X1 _20753_ (
    .A(_11053_),
    .ZN(_11054_)
  );
  AND2_X1 _20754_ (
    .A1(_11003_),
    .A2(_11053_),
    .ZN(_11056_)
  );
  INV_X1 _20755_ (
    .A(_11056_),
    .ZN(_11057_)
  );
  AND2_X1 _20756_ (
    .A1(_11004_),
    .A2(_11054_),
    .ZN(_11058_)
  );
  INV_X1 _20757_ (
    .A(_11058_),
    .ZN(_11059_)
  );
  AND2_X1 _20758_ (
    .A1(_11057_),
    .A2(_11059_),
    .ZN(_11060_)
  );
  INV_X1 _20759_ (
    .A(_11060_),
    .ZN(_11061_)
  );
  AND2_X1 _20760_ (
    .A1(_10975_),
    .A2(_11060_),
    .ZN(_11062_)
  );
  INV_X1 _20761_ (
    .A(_11062_),
    .ZN(_11063_)
  );
  AND2_X1 _20762_ (
    .A1(_10974_),
    .A2(_11061_),
    .ZN(_11064_)
  );
  INV_X1 _20763_ (
    .A(_11064_),
    .ZN(_11065_)
  );
  AND2_X1 _20764_ (
    .A1(_11063_),
    .A2(_11065_),
    .ZN(_11067_)
  );
  INV_X1 _20765_ (
    .A(_11067_),
    .ZN(_11068_)
  );
  AND2_X1 _20766_ (
    .A1(_10810_),
    .A2(_10816_),
    .ZN(_11069_)
  );
  INV_X1 _20767_ (
    .A(_11069_),
    .ZN(_11070_)
  );
  AND2_X1 _20768_ (
    .A1(_10765_),
    .A2(_10771_),
    .ZN(_11071_)
  );
  INV_X1 _20769_ (
    .A(_11071_),
    .ZN(_11072_)
  );
  AND2_X1 _20770_ (
    .A1(_10798_),
    .A2(_10804_),
    .ZN(_11073_)
  );
  INV_X1 _20771_ (
    .A(_11073_),
    .ZN(_11074_)
  );
  AND2_X1 _20772_ (
    .A1(_10747_),
    .A2(_10753_),
    .ZN(_11075_)
  );
  INV_X1 _20773_ (
    .A(_11075_),
    .ZN(_11076_)
  );
  AND2_X1 _20774_ (
    .A1(_10203_),
    .A2(_11076_),
    .ZN(_11078_)
  );
  INV_X1 _20775_ (
    .A(_11078_),
    .ZN(_11079_)
  );
  AND2_X1 _20776_ (
    .A1(_10204_),
    .A2(_11075_),
    .ZN(_11080_)
  );
  INV_X1 _20777_ (
    .A(_11080_),
    .ZN(_11081_)
  );
  AND2_X1 _20778_ (
    .A1(_11079_),
    .A2(_11081_),
    .ZN(_11082_)
  );
  INV_X1 _20779_ (
    .A(_11082_),
    .ZN(_11083_)
  );
  AND2_X1 _20780_ (
    .A1(_10493_),
    .A2(_11082_),
    .ZN(_11084_)
  );
  INV_X1 _20781_ (
    .A(_11084_),
    .ZN(_11085_)
  );
  AND2_X1 _20782_ (
    .A1(_10492_),
    .A2(_11083_),
    .ZN(_11086_)
  );
  INV_X1 _20783_ (
    .A(_11086_),
    .ZN(_11087_)
  );
  AND2_X1 _20784_ (
    .A1(_11085_),
    .A2(_11087_),
    .ZN(_11088_)
  );
  INV_X1 _20785_ (
    .A(_11088_),
    .ZN(_11089_)
  );
  AND2_X1 _20786_ (
    .A1(_11074_),
    .A2(_11088_),
    .ZN(_11090_)
  );
  INV_X1 _20787_ (
    .A(_11090_),
    .ZN(_11091_)
  );
  AND2_X1 _20788_ (
    .A1(_11073_),
    .A2(_11089_),
    .ZN(_11092_)
  );
  INV_X1 _20789_ (
    .A(_11092_),
    .ZN(_11093_)
  );
  AND2_X1 _20790_ (
    .A1(_11091_),
    .A2(_11093_),
    .ZN(_11094_)
  );
  INV_X1 _20791_ (
    .A(_11094_),
    .ZN(_11095_)
  );
  AND2_X1 _20792_ (
    .A1(_09521_),
    .A2(_11094_),
    .ZN(_11096_)
  );
  INV_X1 _20793_ (
    .A(_11096_),
    .ZN(_11097_)
  );
  AND2_X1 _20794_ (
    .A1(_09522_),
    .A2(_11095_),
    .ZN(_11099_)
  );
  INV_X1 _20795_ (
    .A(_11099_),
    .ZN(_11100_)
  );
  AND2_X1 _20796_ (
    .A1(_11097_),
    .A2(_11100_),
    .ZN(_11101_)
  );
  INV_X1 _20797_ (
    .A(_11101_),
    .ZN(_11102_)
  );
  AND2_X1 _20798_ (
    .A1(_11072_),
    .A2(_11101_),
    .ZN(_11103_)
  );
  INV_X1 _20799_ (
    .A(_11103_),
    .ZN(_11104_)
  );
  AND2_X1 _20800_ (
    .A1(_11071_),
    .A2(_11102_),
    .ZN(_11105_)
  );
  INV_X1 _20801_ (
    .A(_11105_),
    .ZN(_11106_)
  );
  AND2_X1 _20802_ (
    .A1(_11104_),
    .A2(_11106_),
    .ZN(_11107_)
  );
  INV_X1 _20803_ (
    .A(_11107_),
    .ZN(_11108_)
  );
  AND2_X1 _20804_ (
    .A1(_11070_),
    .A2(_11107_),
    .ZN(_11110_)
  );
  INV_X1 _20805_ (
    .A(_11110_),
    .ZN(_11111_)
  );
  AND2_X1 _20806_ (
    .A1(_11069_),
    .A2(_11108_),
    .ZN(_11112_)
  );
  INV_X1 _20807_ (
    .A(_11112_),
    .ZN(_11113_)
  );
  AND2_X1 _20808_ (
    .A1(_11111_),
    .A2(_11113_),
    .ZN(_11114_)
  );
  INV_X1 _20809_ (
    .A(_11114_),
    .ZN(_11115_)
  );
  AND2_X1 _20810_ (
    .A1(_11067_),
    .A2(_11114_),
    .ZN(_11116_)
  );
  INV_X1 _20811_ (
    .A(_11116_),
    .ZN(_11117_)
  );
  AND2_X1 _20812_ (
    .A1(_11068_),
    .A2(_11115_),
    .ZN(_11118_)
  );
  INV_X1 _20813_ (
    .A(_11118_),
    .ZN(_11119_)
  );
  AND2_X1 _20814_ (
    .A1(_11117_),
    .A2(_11119_),
    .ZN(_11121_)
  );
  INV_X1 _20815_ (
    .A(_11121_),
    .ZN(_11122_)
  );
  AND2_X1 _20816_ (
    .A1(_10973_),
    .A2(_11121_),
    .ZN(_11123_)
  );
  INV_X1 _20817_ (
    .A(_11123_),
    .ZN(_11124_)
  );
  AND2_X1 _20818_ (
    .A1(_10972_),
    .A2(_11122_),
    .ZN(_11125_)
  );
  INV_X1 _20819_ (
    .A(_11125_),
    .ZN(_11126_)
  );
  AND2_X1 _20820_ (
    .A1(_11124_),
    .A2(_11126_),
    .ZN(_11127_)
  );
  INV_X1 _20821_ (
    .A(_11127_),
    .ZN(_11128_)
  );
  AND2_X1 _20822_ (
    .A1(_10823_),
    .A2(_10830_),
    .ZN(_11129_)
  );
  INV_X1 _20823_ (
    .A(_11129_),
    .ZN(_11130_)
  );
  AND2_X1 _20824_ (
    .A1(_10271_),
    .A2(_11130_),
    .ZN(_11132_)
  );
  INV_X1 _20825_ (
    .A(_11132_),
    .ZN(_11133_)
  );
  AND2_X1 _20826_ (
    .A1(_10272_),
    .A2(_11129_),
    .ZN(_11134_)
  );
  INV_X1 _20827_ (
    .A(_11134_),
    .ZN(_11135_)
  );
  AND2_X1 _20828_ (
    .A1(_11133_),
    .A2(_11135_),
    .ZN(_11136_)
  );
  INV_X1 _20829_ (
    .A(_11136_),
    .ZN(_11137_)
  );
  AND2_X1 _20830_ (
    .A1(_10551_),
    .A2(_11136_),
    .ZN(_11138_)
  );
  INV_X1 _20831_ (
    .A(_11138_),
    .ZN(_11139_)
  );
  AND2_X1 _20832_ (
    .A1(_10549_),
    .A2(_11137_),
    .ZN(_11140_)
  );
  INV_X1 _20833_ (
    .A(_11140_),
    .ZN(_11141_)
  );
  AND2_X1 _20834_ (
    .A1(_11139_),
    .A2(_11141_),
    .ZN(_00122_)
  );
  INV_X1 _20835_ (
    .A(_00122_),
    .ZN(_00123_)
  );
  AND2_X1 _20836_ (
    .A1(_11127_),
    .A2(_00122_),
    .ZN(_00124_)
  );
  INV_X1 _20837_ (
    .A(_00124_),
    .ZN(_00125_)
  );
  AND2_X1 _20838_ (
    .A1(_11128_),
    .A2(_00123_),
    .ZN(_00126_)
  );
  INV_X1 _20839_ (
    .A(_00126_),
    .ZN(_00127_)
  );
  AND2_X1 _20840_ (
    .A1(_00125_),
    .A2(_00127_),
    .ZN(_00128_)
  );
  INV_X1 _20841_ (
    .A(_00128_),
    .ZN(_00129_)
  );
  AND2_X1 _20842_ (
    .A1(_10971_),
    .A2(_00128_),
    .ZN(_00130_)
  );
  INV_X1 _20843_ (
    .A(_00130_),
    .ZN(_00131_)
  );
  AND2_X1 _20844_ (
    .A1(_10970_),
    .A2(_00129_),
    .ZN(_00132_)
  );
  INV_X1 _20845_ (
    .A(_00132_),
    .ZN(_00133_)
  );
  AND2_X1 _20846_ (
    .A1(_00131_),
    .A2(_00133_),
    .ZN(_00134_)
  );
  INV_X1 _20847_ (
    .A(_00134_),
    .ZN(_00135_)
  );
  AND2_X1 _20848_ (
    .A1(_10852_),
    .A2(_10858_),
    .ZN(_00136_)
  );
  INV_X1 _20849_ (
    .A(_00136_),
    .ZN(_00137_)
  );
  AND2_X1 _20850_ (
    .A1(_07804_),
    .A2(_00137_),
    .ZN(_00138_)
  );
  INV_X1 _20851_ (
    .A(_00138_),
    .ZN(_00139_)
  );
  AND2_X1 _20852_ (
    .A1(_07805_),
    .A2(_00136_),
    .ZN(_00140_)
  );
  INV_X1 _20853_ (
    .A(_00140_),
    .ZN(_00141_)
  );
  AND2_X1 _20854_ (
    .A1(_00139_),
    .A2(_00141_),
    .ZN(_00143_)
  );
  INV_X1 _20855_ (
    .A(_00143_),
    .ZN(_00144_)
  );
  AND2_X1 _20856_ (
    .A1(_08107_),
    .A2(_00143_),
    .ZN(_00145_)
  );
  INV_X1 _20857_ (
    .A(_00145_),
    .ZN(_00146_)
  );
  AND2_X1 _20858_ (
    .A1(_08106_),
    .A2(_00144_),
    .ZN(_00147_)
  );
  INV_X1 _20859_ (
    .A(_00147_),
    .ZN(_00148_)
  );
  AND2_X1 _20860_ (
    .A1(_00146_),
    .A2(_00148_),
    .ZN(_00149_)
  );
  INV_X1 _20861_ (
    .A(_00149_),
    .ZN(_00150_)
  );
  AND2_X1 _20862_ (
    .A1(_00134_),
    .A2(_00149_),
    .ZN(_00151_)
  );
  INV_X1 _20863_ (
    .A(_00151_),
    .ZN(_00152_)
  );
  AND2_X1 _20864_ (
    .A1(_00135_),
    .A2(_00150_),
    .ZN(_00154_)
  );
  INV_X1 _20865_ (
    .A(_00154_),
    .ZN(_00155_)
  );
  AND2_X1 _20866_ (
    .A1(_00152_),
    .A2(_00155_),
    .ZN(_00156_)
  );
  INV_X1 _20867_ (
    .A(_00156_),
    .ZN(_00157_)
  );
  AND2_X1 _20868_ (
    .A1(_10969_),
    .A2(_00156_),
    .ZN(_00158_)
  );
  INV_X1 _20869_ (
    .A(_00158_),
    .ZN(_00159_)
  );
  AND2_X1 _20870_ (
    .A1(_10967_),
    .A2(_00157_),
    .ZN(_00160_)
  );
  INV_X1 _20871_ (
    .A(_00160_),
    .ZN(_00161_)
  );
  AND2_X1 _20872_ (
    .A1(_00159_),
    .A2(_00161_),
    .ZN(_00162_)
  );
  INV_X1 _20873_ (
    .A(_00162_),
    .ZN(_00163_)
  );
  AND2_X1 _20874_ (
    .A1(_10966_),
    .A2(_00162_),
    .ZN(_00165_)
  );
  INV_X1 _20875_ (
    .A(_00165_),
    .ZN(_00166_)
  );
  AND2_X1 _20876_ (
    .A1(_10965_),
    .A2(_00163_),
    .ZN(_00167_)
  );
  INV_X1 _20877_ (
    .A(_00167_),
    .ZN(_00168_)
  );
  AND2_X1 _20878_ (
    .A1(_00166_),
    .A2(_00168_),
    .ZN(_00169_)
  );
  INV_X1 _20879_ (
    .A(_00169_),
    .ZN(_00170_)
  );
  AND2_X1 _20880_ (
    .A1(_10964_),
    .A2(_00169_),
    .ZN(_00171_)
  );
  INV_X1 _20881_ (
    .A(_00171_),
    .ZN(_00172_)
  );
  AND2_X1 _20882_ (
    .A1(_10963_),
    .A2(_00170_),
    .ZN(_00173_)
  );
  INV_X1 _20883_ (
    .A(_00173_),
    .ZN(_00174_)
  );
  AND2_X1 _20884_ (
    .A1(_00172_),
    .A2(_00174_),
    .ZN(_00176_)
  );
  INV_X1 _20885_ (
    .A(_00176_),
    .ZN(_00177_)
  );
  AND2_X1 _20886_ (
    .A1(_10911_),
    .A2(_00176_),
    .ZN(_00178_)
  );
  INV_X1 _20887_ (
    .A(_00178_),
    .ZN(_00179_)
  );
  AND2_X1 _20888_ (
    .A1(_10912_),
    .A2(_00177_),
    .ZN(_00180_)
  );
  INV_X1 _20889_ (
    .A(_00180_),
    .ZN(_00181_)
  );
  AND2_X1 _20890_ (
    .A1(_00179_),
    .A2(_00181_),
    .ZN(_00182_)
  );
  INV_X1 _20891_ (
    .A(_00182_),
    .ZN(_00183_)
  );
  AND2_X1 _20892_ (
    .A1(_10669_),
    .A2(_10919_),
    .ZN(_00184_)
  );
  INV_X1 _20893_ (
    .A(_00184_),
    .ZN(_00185_)
  );
  AND2_X1 _20894_ (
    .A1(_10921_),
    .A2(_00185_),
    .ZN(_00187_)
  );
  AND2_X1 _20895_ (
    .A1(_10919_),
    .A2(_10928_),
    .ZN(_00188_)
  );
  AND2_X1 _20896_ (
    .A1(_00182_),
    .A2(_00187_),
    .ZN(_00189_)
  );
  INV_X1 _20897_ (
    .A(_00189_),
    .ZN(_00190_)
  );
  AND2_X1 _20898_ (
    .A1(_00183_),
    .A2(_00188_),
    .ZN(_00191_)
  );
  INV_X1 _20899_ (
    .A(_00191_),
    .ZN(_00192_)
  );
  AND2_X1 _20900_ (
    .A1(_00190_),
    .A2(_00192_),
    .ZN(_00193_)
  );
  INV_X1 _20901_ (
    .A(_00193_),
    .ZN(_00194_)
  );
  AND2_X1 _20902_ (
    .A1(remainder[65]),
    .A2(_00193_),
    .ZN(_00195_)
  );
  INV_X1 _20903_ (
    .A(_00195_),
    .ZN(_00196_)
  );
  AND2_X1 _20904_ (
    .A1(_04404_),
    .A2(_00194_),
    .ZN(_00198_)
  );
  INV_X1 _20905_ (
    .A(_00198_),
    .ZN(_00199_)
  );
  AND2_X1 _20906_ (
    .A1(_00196_),
    .A2(_00199_),
    .ZN(_00200_)
  );
  INV_X1 _20907_ (
    .A(_00200_),
    .ZN(_00201_)
  );
  AND2_X1 _20908_ (
    .A1(_10962_),
    .A2(_00200_),
    .ZN(_00202_)
  );
  INV_X1 _20909_ (
    .A(_00202_),
    .ZN(_00203_)
  );
  AND2_X1 _20910_ (
    .A1(_10961_),
    .A2(_00201_),
    .ZN(_00204_)
  );
  INV_X1 _20911_ (
    .A(_00204_),
    .ZN(_00205_)
  );
  AND2_X1 _20912_ (
    .A1(_02082_),
    .A2(_00205_),
    .ZN(_00206_)
  );
  AND2_X1 _20913_ (
    .A1(_00203_),
    .A2(_00206_),
    .ZN(_00207_)
  );
  INV_X1 _20914_ (
    .A(_00207_),
    .ZN(_00209_)
  );
  AND2_X1 _20915_ (
    .A1(remainder[63]),
    .A2(_02077_),
    .ZN(_00210_)
  );
  INV_X1 _20916_ (
    .A(_00210_),
    .ZN(_00211_)
  );
  AND2_X1 _20917_ (
    .A1(_04437_),
    .A2(_10451_),
    .ZN(_00212_)
  );
  INV_X1 _20918_ (
    .A(_00212_),
    .ZN(_00213_)
  );
  AND2_X1 _20919_ (
    .A1(_10462_),
    .A2(_02046_),
    .ZN(_00214_)
  );
  INV_X1 _20920_ (
    .A(_00214_),
    .ZN(_00215_)
  );
  AND2_X1 _20921_ (
    .A1(_05983_),
    .A2(_00215_),
    .ZN(_00216_)
  );
  AND2_X1 _20922_ (
    .A1(_00213_),
    .A2(_00216_),
    .ZN(_00217_)
  );
  INV_X1 _20923_ (
    .A(_00217_),
    .ZN(_00218_)
  );
  AND2_X1 _20924_ (
    .A1(_00211_),
    .A2(_00218_),
    .ZN(_00220_)
  );
  AND2_X1 _20925_ (
    .A1(_00209_),
    .A2(_00220_),
    .ZN(_00221_)
  );
  INV_X1 _20926_ (
    .A(_00221_),
    .ZN(_00222_)
  );
  AND2_X1 _20927_ (
    .A1(_06201_),
    .A2(_00222_),
    .ZN(_00084_)
  );
  AND2_X1 _20928_ (
    .A1(_00196_),
    .A2(_00203_),
    .ZN(_00223_)
  );
  INV_X1 _20929_ (
    .A(_00223_),
    .ZN(_00224_)
  );
  AND2_X1 _20930_ (
    .A1(_00179_),
    .A2(_00190_),
    .ZN(_00225_)
  );
  INV_X1 _20931_ (
    .A(_00225_),
    .ZN(_00226_)
  );
  AND2_X1 _20932_ (
    .A1(_00159_),
    .A2(_00166_),
    .ZN(_00227_)
  );
  INV_X1 _20933_ (
    .A(_00227_),
    .ZN(_00228_)
  );
  AND2_X1 _20934_ (
    .A1(_00139_),
    .A2(_00146_),
    .ZN(_00230_)
  );
  INV_X1 _20935_ (
    .A(_00230_),
    .ZN(_00231_)
  );
  AND2_X1 _20936_ (
    .A1(_00131_),
    .A2(_00152_),
    .ZN(_00232_)
  );
  INV_X1 _20937_ (
    .A(_00232_),
    .ZN(_00233_)
  );
  AND2_X1 _20938_ (
    .A1(_11124_),
    .A2(_00125_),
    .ZN(_00234_)
  );
  INV_X1 _20939_ (
    .A(_00234_),
    .ZN(_00235_)
  );
  AND2_X1 _20940_ (
    .A1(_11063_),
    .A2(_11117_),
    .ZN(_00236_)
  );
  INV_X1 _20941_ (
    .A(_00236_),
    .ZN(_00237_)
  );
  AND2_X1 _20942_ (
    .A1(_10999_),
    .A2(_11057_),
    .ZN(_00238_)
  );
  INV_X1 _20943_ (
    .A(_00238_),
    .ZN(_00239_)
  );
  AND2_X1 _20944_ (
    .A1(_10108_),
    .A2(_10993_),
    .ZN(_00241_)
  );
  INV_X1 _20945_ (
    .A(_00241_),
    .ZN(_00242_)
  );
  AND2_X1 _20946_ (
    .A1(_10109_),
    .A2(_10464_),
    .ZN(_00243_)
  );
  INV_X1 _20947_ (
    .A(_00243_),
    .ZN(_00244_)
  );
  MUX2_X1 _20948_ (
    .A(_10112_),
    .B(_10114_),
    .S(_09794_),
    .Z(_00245_)
  );
  INV_X1 _20949_ (
    .A(_00245_),
    .ZN(_00246_)
  );
  AND2_X1 _20950_ (
    .A1(_00244_),
    .A2(_00246_),
    .ZN(_00247_)
  );
  INV_X1 _20951_ (
    .A(_00247_),
    .ZN(_00248_)
  );
  AND2_X1 _20952_ (
    .A1(_10128_),
    .A2(_10980_),
    .ZN(_00249_)
  );
  INV_X1 _20953_ (
    .A(_00249_),
    .ZN(_00250_)
  );
  AND2_X1 _20954_ (
    .A1(_10410_),
    .A2(_10723_),
    .ZN(_00252_)
  );
  INV_X1 _20955_ (
    .A(_00252_),
    .ZN(_00253_)
  );
  AND2_X1 _20956_ (
    .A1(_10411_),
    .A2(_10724_),
    .ZN(_00254_)
  );
  INV_X1 _20957_ (
    .A(_00254_),
    .ZN(_00255_)
  );
  AND2_X1 _20958_ (
    .A1(_00253_),
    .A2(_00255_),
    .ZN(_00256_)
  );
  INV_X1 _20959_ (
    .A(_00256_),
    .ZN(_00257_)
  );
  AND2_X1 _20960_ (
    .A1(_09545_),
    .A2(_00256_),
    .ZN(_00258_)
  );
  INV_X1 _20961_ (
    .A(_00258_),
    .ZN(_00259_)
  );
  AND2_X1 _20962_ (
    .A1(_09546_),
    .A2(_00257_),
    .ZN(_00260_)
  );
  INV_X1 _20963_ (
    .A(_00260_),
    .ZN(_00261_)
  );
  AND2_X1 _20964_ (
    .A1(_00259_),
    .A2(_00261_),
    .ZN(_00263_)
  );
  INV_X1 _20965_ (
    .A(_00263_),
    .ZN(_00264_)
  );
  AND2_X1 _20966_ (
    .A1(_00250_),
    .A2(_00263_),
    .ZN(_00265_)
  );
  INV_X1 _20967_ (
    .A(_00265_),
    .ZN(_00266_)
  );
  AND2_X1 _20968_ (
    .A1(_00249_),
    .A2(_00264_),
    .ZN(_00267_)
  );
  INV_X1 _20969_ (
    .A(_00267_),
    .ZN(_00268_)
  );
  AND2_X1 _20970_ (
    .A1(_00266_),
    .A2(_00268_),
    .ZN(_00269_)
  );
  INV_X1 _20971_ (
    .A(_00269_),
    .ZN(_00270_)
  );
  AND2_X1 _20972_ (
    .A1(_00248_),
    .A2(_00269_),
    .ZN(_00271_)
  );
  INV_X1 _20973_ (
    .A(_00271_),
    .ZN(_00272_)
  );
  AND2_X1 _20974_ (
    .A1(_00247_),
    .A2(_00270_),
    .ZN(_00274_)
  );
  INV_X1 _20975_ (
    .A(_00274_),
    .ZN(_00275_)
  );
  AND2_X1 _20976_ (
    .A1(_00272_),
    .A2(_00275_),
    .ZN(_00276_)
  );
  INV_X1 _20977_ (
    .A(_00276_),
    .ZN(_00277_)
  );
  AND2_X1 _20978_ (
    .A1(_00242_),
    .A2(_00276_),
    .ZN(_00278_)
  );
  INV_X1 _20979_ (
    .A(_00278_),
    .ZN(_00279_)
  );
  AND2_X1 _20980_ (
    .A1(_00241_),
    .A2(_00277_),
    .ZN(_00280_)
  );
  INV_X1 _20981_ (
    .A(_00280_),
    .ZN(_00281_)
  );
  AND2_X1 _20982_ (
    .A1(_00279_),
    .A2(_00281_),
    .ZN(_00282_)
  );
  INV_X1 _20983_ (
    .A(_00282_),
    .ZN(_00283_)
  );
  AND2_X1 _20984_ (
    .A1(_11025_),
    .A2(_11037_),
    .ZN(_00285_)
  );
  INV_X1 _20985_ (
    .A(_00285_),
    .ZN(_00286_)
  );
  AND2_X1 _20986_ (
    .A1(_11015_),
    .A2(_11019_),
    .ZN(_00287_)
  );
  INV_X1 _20987_ (
    .A(_00287_),
    .ZN(_00288_)
  );
  AND2_X1 _20988_ (
    .A1(remainder[32]),
    .A2(divisor[31]),
    .ZN(_00289_)
  );
  INV_X1 _20989_ (
    .A(_00289_),
    .ZN(_00290_)
  );
  AND2_X1 _20990_ (
    .A1(divisor[32]),
    .A2(remainder[7]),
    .ZN(_00291_)
  );
  AND2_X1 _20991_ (
    .A1(remainder[7]),
    .A2(_11011_),
    .ZN(_00292_)
  );
  INV_X1 _20992_ (
    .A(_00292_),
    .ZN(_00293_)
  );
  MUX2_X1 _20993_ (
    .A(_11011_),
    .B(_05138_),
    .S(_00291_),
    .Z(_00294_)
  );
  MUX2_X1 _20994_ (
    .A(_11013_),
    .B(remainder[6]),
    .S(_00291_),
    .Z(_00296_)
  );
  AND2_X1 _20995_ (
    .A1(_00289_),
    .A2(_00294_),
    .ZN(_00297_)
  );
  INV_X1 _20996_ (
    .A(_00297_),
    .ZN(_00298_)
  );
  AND2_X1 _20997_ (
    .A1(_00290_),
    .A2(_00296_),
    .ZN(_00299_)
  );
  INV_X1 _20998_ (
    .A(_00299_),
    .ZN(_00300_)
  );
  AND2_X1 _20999_ (
    .A1(_00298_),
    .A2(_00300_),
    .ZN(_00301_)
  );
  INV_X1 _21000_ (
    .A(_00301_),
    .ZN(_00302_)
  );
  AND2_X1 _21001_ (
    .A1(_00288_),
    .A2(_00301_),
    .ZN(_00303_)
  );
  INV_X1 _21002_ (
    .A(_00303_),
    .ZN(_00304_)
  );
  AND2_X1 _21003_ (
    .A1(_00287_),
    .A2(_00302_),
    .ZN(_00305_)
  );
  INV_X1 _21004_ (
    .A(_00305_),
    .ZN(_00307_)
  );
  AND2_X1 _21005_ (
    .A1(_00304_),
    .A2(_00307_),
    .ZN(_00308_)
  );
  INV_X1 _21006_ (
    .A(_00308_),
    .ZN(_00309_)
  );
  AND2_X1 _21007_ (
    .A1(_11034_),
    .A2(_00308_),
    .ZN(_00310_)
  );
  INV_X1 _21008_ (
    .A(_00310_),
    .ZN(_00311_)
  );
  AND2_X1 _21009_ (
    .A1(_11035_),
    .A2(_00309_),
    .ZN(_00312_)
  );
  INV_X1 _21010_ (
    .A(_00312_),
    .ZN(_00313_)
  );
  AND2_X1 _21011_ (
    .A1(_00311_),
    .A2(_00313_),
    .ZN(_00314_)
  );
  INV_X1 _21012_ (
    .A(_00314_),
    .ZN(_00315_)
  );
  AND2_X1 _21013_ (
    .A1(_10985_),
    .A2(_00314_),
    .ZN(_00316_)
  );
  INV_X1 _21014_ (
    .A(_00316_),
    .ZN(_00317_)
  );
  AND2_X1 _21015_ (
    .A1(_10986_),
    .A2(_00315_),
    .ZN(_00318_)
  );
  INV_X1 _21016_ (
    .A(_00318_),
    .ZN(_00319_)
  );
  AND2_X1 _21017_ (
    .A1(_00317_),
    .A2(_00319_),
    .ZN(_00320_)
  );
  INV_X1 _21018_ (
    .A(_00320_),
    .ZN(_00321_)
  );
  AND2_X1 _21019_ (
    .A1(_00286_),
    .A2(_00320_),
    .ZN(_00322_)
  );
  INV_X1 _21020_ (
    .A(_00322_),
    .ZN(_00323_)
  );
  AND2_X1 _21021_ (
    .A1(_00285_),
    .A2(_00321_),
    .ZN(_00324_)
  );
  INV_X1 _21022_ (
    .A(_00324_),
    .ZN(_00325_)
  );
  AND2_X1 _21023_ (
    .A1(_00323_),
    .A2(_00325_),
    .ZN(_00326_)
  );
  INV_X1 _21024_ (
    .A(_00326_),
    .ZN(_00328_)
  );
  AND2_X1 _21025_ (
    .A1(_00282_),
    .A2(_00326_),
    .ZN(_00329_)
  );
  INV_X1 _21026_ (
    .A(_00329_),
    .ZN(_00330_)
  );
  AND2_X1 _21027_ (
    .A1(_00283_),
    .A2(_00328_),
    .ZN(_00331_)
  );
  INV_X1 _21028_ (
    .A(_00331_),
    .ZN(_00332_)
  );
  AND2_X1 _21029_ (
    .A1(_00330_),
    .A2(_00332_),
    .ZN(_00333_)
  );
  INV_X1 _21030_ (
    .A(_00333_),
    .ZN(_00334_)
  );
  AND2_X1 _21031_ (
    .A1(_00239_),
    .A2(_00333_),
    .ZN(_00335_)
  );
  INV_X1 _21032_ (
    .A(_00335_),
    .ZN(_00336_)
  );
  AND2_X1 _21033_ (
    .A1(_00238_),
    .A2(_00334_),
    .ZN(_00337_)
  );
  INV_X1 _21034_ (
    .A(_00337_),
    .ZN(_00339_)
  );
  AND2_X1 _21035_ (
    .A1(_00336_),
    .A2(_00339_),
    .ZN(_00340_)
  );
  INV_X1 _21036_ (
    .A(_00340_),
    .ZN(_00341_)
  );
  AND2_X1 _21037_ (
    .A1(_11091_),
    .A2(_11097_),
    .ZN(_00342_)
  );
  INV_X1 _21038_ (
    .A(_00342_),
    .ZN(_00343_)
  );
  AND2_X1 _21039_ (
    .A1(_11043_),
    .A2(_11050_),
    .ZN(_00344_)
  );
  INV_X1 _21040_ (
    .A(_00344_),
    .ZN(_00345_)
  );
  AND2_X1 _21041_ (
    .A1(_11079_),
    .A2(_11085_),
    .ZN(_00346_)
  );
  INV_X1 _21042_ (
    .A(_00346_),
    .ZN(_00347_)
  );
  AND2_X1 _21043_ (
    .A1(_10745_),
    .A2(_11032_),
    .ZN(_00348_)
  );
  INV_X1 _21044_ (
    .A(_00348_),
    .ZN(_00350_)
  );
  AND2_X1 _21045_ (
    .A1(_10203_),
    .A2(_00350_),
    .ZN(_00351_)
  );
  INV_X1 _21046_ (
    .A(_00351_),
    .ZN(_00352_)
  );
  AND2_X1 _21047_ (
    .A1(_10204_),
    .A2(_00348_),
    .ZN(_00353_)
  );
  INV_X1 _21048_ (
    .A(_00353_),
    .ZN(_00354_)
  );
  AND2_X1 _21049_ (
    .A1(_00352_),
    .A2(_00354_),
    .ZN(_00355_)
  );
  INV_X1 _21050_ (
    .A(_00355_),
    .ZN(_00356_)
  );
  AND2_X1 _21051_ (
    .A1(_10492_),
    .A2(_00356_),
    .ZN(_00357_)
  );
  INV_X1 _21052_ (
    .A(_00357_),
    .ZN(_00358_)
  );
  AND2_X1 _21053_ (
    .A1(_10493_),
    .A2(_00355_),
    .ZN(_00359_)
  );
  INV_X1 _21054_ (
    .A(_00359_),
    .ZN(_00361_)
  );
  AND2_X1 _21055_ (
    .A1(_10493_),
    .A2(_00356_),
    .ZN(_00362_)
  );
  INV_X1 _21056_ (
    .A(_00362_),
    .ZN(_00363_)
  );
  AND2_X1 _21057_ (
    .A1(_10492_),
    .A2(_00355_),
    .ZN(_00364_)
  );
  INV_X1 _21058_ (
    .A(_00364_),
    .ZN(_00365_)
  );
  AND2_X1 _21059_ (
    .A1(_00358_),
    .A2(_00361_),
    .ZN(_00366_)
  );
  AND2_X1 _21060_ (
    .A1(_00363_),
    .A2(_00365_),
    .ZN(_00367_)
  );
  AND2_X1 _21061_ (
    .A1(_00347_),
    .A2(_00366_),
    .ZN(_00368_)
  );
  INV_X1 _21062_ (
    .A(_00368_),
    .ZN(_00369_)
  );
  AND2_X1 _21063_ (
    .A1(_00346_),
    .A2(_00367_),
    .ZN(_00370_)
  );
  INV_X1 _21064_ (
    .A(_00370_),
    .ZN(_00372_)
  );
  AND2_X1 _21065_ (
    .A1(_00369_),
    .A2(_00372_),
    .ZN(_00373_)
  );
  INV_X1 _21066_ (
    .A(_00373_),
    .ZN(_00374_)
  );
  AND2_X1 _21067_ (
    .A1(_09521_),
    .A2(_00373_),
    .ZN(_00375_)
  );
  INV_X1 _21068_ (
    .A(_00375_),
    .ZN(_00376_)
  );
  AND2_X1 _21069_ (
    .A1(_09522_),
    .A2(_00374_),
    .ZN(_00377_)
  );
  INV_X1 _21070_ (
    .A(_00377_),
    .ZN(_00378_)
  );
  AND2_X1 _21071_ (
    .A1(_00376_),
    .A2(_00378_),
    .ZN(_00379_)
  );
  INV_X1 _21072_ (
    .A(_00379_),
    .ZN(_00380_)
  );
  AND2_X1 _21073_ (
    .A1(_00345_),
    .A2(_00379_),
    .ZN(_00381_)
  );
  INV_X1 _21074_ (
    .A(_00381_),
    .ZN(_00383_)
  );
  AND2_X1 _21075_ (
    .A1(_00344_),
    .A2(_00380_),
    .ZN(_00384_)
  );
  INV_X1 _21076_ (
    .A(_00384_),
    .ZN(_00385_)
  );
  AND2_X1 _21077_ (
    .A1(_00383_),
    .A2(_00385_),
    .ZN(_00386_)
  );
  INV_X1 _21078_ (
    .A(_00386_),
    .ZN(_00387_)
  );
  AND2_X1 _21079_ (
    .A1(_00343_),
    .A2(_00386_),
    .ZN(_00388_)
  );
  INV_X1 _21080_ (
    .A(_00388_),
    .ZN(_00389_)
  );
  AND2_X1 _21081_ (
    .A1(_00342_),
    .A2(_00387_),
    .ZN(_00390_)
  );
  INV_X1 _21082_ (
    .A(_00390_),
    .ZN(_00391_)
  );
  AND2_X1 _21083_ (
    .A1(_00389_),
    .A2(_00391_),
    .ZN(_00392_)
  );
  INV_X1 _21084_ (
    .A(_00392_),
    .ZN(_00394_)
  );
  AND2_X1 _21085_ (
    .A1(_00340_),
    .A2(_00392_),
    .ZN(_00395_)
  );
  INV_X1 _21086_ (
    .A(_00395_),
    .ZN(_00396_)
  );
  AND2_X1 _21087_ (
    .A1(_00341_),
    .A2(_00394_),
    .ZN(_00397_)
  );
  INV_X1 _21088_ (
    .A(_00397_),
    .ZN(_00398_)
  );
  AND2_X1 _21089_ (
    .A1(_00396_),
    .A2(_00398_),
    .ZN(_00399_)
  );
  INV_X1 _21090_ (
    .A(_00399_),
    .ZN(_00400_)
  );
  AND2_X1 _21091_ (
    .A1(_00237_),
    .A2(_00399_),
    .ZN(_00401_)
  );
  INV_X1 _21092_ (
    .A(_00401_),
    .ZN(_00402_)
  );
  AND2_X1 _21093_ (
    .A1(_00236_),
    .A2(_00400_),
    .ZN(_00403_)
  );
  INV_X1 _21094_ (
    .A(_00403_),
    .ZN(_00405_)
  );
  AND2_X1 _21095_ (
    .A1(_00402_),
    .A2(_00405_),
    .ZN(_00406_)
  );
  INV_X1 _21096_ (
    .A(_00406_),
    .ZN(_00407_)
  );
  AND2_X1 _21097_ (
    .A1(_11104_),
    .A2(_11111_),
    .ZN(_00408_)
  );
  INV_X1 _21098_ (
    .A(_00408_),
    .ZN(_00409_)
  );
  AND2_X1 _21099_ (
    .A1(_10271_),
    .A2(_00409_),
    .ZN(_00410_)
  );
  INV_X1 _21100_ (
    .A(_00410_),
    .ZN(_00411_)
  );
  AND2_X1 _21101_ (
    .A1(_10272_),
    .A2(_00408_),
    .ZN(_00412_)
  );
  INV_X1 _21102_ (
    .A(_00412_),
    .ZN(_00413_)
  );
  AND2_X1 _21103_ (
    .A1(_00411_),
    .A2(_00413_),
    .ZN(_00414_)
  );
  INV_X1 _21104_ (
    .A(_00414_),
    .ZN(_00416_)
  );
  AND2_X1 _21105_ (
    .A1(_10551_),
    .A2(_00414_),
    .ZN(_00417_)
  );
  INV_X1 _21106_ (
    .A(_00417_),
    .ZN(_00418_)
  );
  AND2_X1 _21107_ (
    .A1(_10549_),
    .A2(_00416_),
    .ZN(_00419_)
  );
  INV_X1 _21108_ (
    .A(_00419_),
    .ZN(_00420_)
  );
  AND2_X1 _21109_ (
    .A1(_00418_),
    .A2(_00420_),
    .ZN(_00421_)
  );
  INV_X1 _21110_ (
    .A(_00421_),
    .ZN(_00422_)
  );
  AND2_X1 _21111_ (
    .A1(_00406_),
    .A2(_00421_),
    .ZN(_00423_)
  );
  INV_X1 _21112_ (
    .A(_00423_),
    .ZN(_00424_)
  );
  AND2_X1 _21113_ (
    .A1(_00407_),
    .A2(_00422_),
    .ZN(_00425_)
  );
  INV_X1 _21114_ (
    .A(_00425_),
    .ZN(_00427_)
  );
  AND2_X1 _21115_ (
    .A1(_00424_),
    .A2(_00427_),
    .ZN(_00428_)
  );
  INV_X1 _21116_ (
    .A(_00428_),
    .ZN(_00429_)
  );
  AND2_X1 _21117_ (
    .A1(_00235_),
    .A2(_00428_),
    .ZN(_00430_)
  );
  INV_X1 _21118_ (
    .A(_00430_),
    .ZN(_00431_)
  );
  AND2_X1 _21119_ (
    .A1(_00234_),
    .A2(_00429_),
    .ZN(_00432_)
  );
  INV_X1 _21120_ (
    .A(_00432_),
    .ZN(_00433_)
  );
  AND2_X1 _21121_ (
    .A1(_00431_),
    .A2(_00433_),
    .ZN(_00434_)
  );
  INV_X1 _21122_ (
    .A(_00434_),
    .ZN(_00435_)
  );
  AND2_X1 _21123_ (
    .A1(_11133_),
    .A2(_11139_),
    .ZN(_00436_)
  );
  INV_X1 _21124_ (
    .A(_00436_),
    .ZN(_00438_)
  );
  AND2_X1 _21125_ (
    .A1(_07804_),
    .A2(_00438_),
    .ZN(_00439_)
  );
  INV_X1 _21126_ (
    .A(_00439_),
    .ZN(_00440_)
  );
  AND2_X1 _21127_ (
    .A1(_07805_),
    .A2(_00436_),
    .ZN(_00441_)
  );
  INV_X1 _21128_ (
    .A(_00441_),
    .ZN(_00442_)
  );
  AND2_X1 _21129_ (
    .A1(_00440_),
    .A2(_00442_),
    .ZN(_00443_)
  );
  INV_X1 _21130_ (
    .A(_00443_),
    .ZN(_00444_)
  );
  AND2_X1 _21131_ (
    .A1(_08107_),
    .A2(_00443_),
    .ZN(_00445_)
  );
  INV_X1 _21132_ (
    .A(_00445_),
    .ZN(_00446_)
  );
  AND2_X1 _21133_ (
    .A1(_08106_),
    .A2(_00444_),
    .ZN(_00447_)
  );
  INV_X1 _21134_ (
    .A(_00447_),
    .ZN(_00449_)
  );
  AND2_X1 _21135_ (
    .A1(_00446_),
    .A2(_00449_),
    .ZN(_00450_)
  );
  INV_X1 _21136_ (
    .A(_00450_),
    .ZN(_00451_)
  );
  AND2_X1 _21137_ (
    .A1(_00434_),
    .A2(_00450_),
    .ZN(_00452_)
  );
  INV_X1 _21138_ (
    .A(_00452_),
    .ZN(_00453_)
  );
  AND2_X1 _21139_ (
    .A1(_00435_),
    .A2(_00451_),
    .ZN(_00454_)
  );
  INV_X1 _21140_ (
    .A(_00454_),
    .ZN(_00455_)
  );
  AND2_X1 _21141_ (
    .A1(_00453_),
    .A2(_00455_),
    .ZN(_00456_)
  );
  INV_X1 _21142_ (
    .A(_00456_),
    .ZN(_00457_)
  );
  AND2_X1 _21143_ (
    .A1(_00233_),
    .A2(_00456_),
    .ZN(_00458_)
  );
  INV_X1 _21144_ (
    .A(_00458_),
    .ZN(_00459_)
  );
  AND2_X1 _21145_ (
    .A1(_00232_),
    .A2(_00457_),
    .ZN(_00460_)
  );
  INV_X1 _21146_ (
    .A(_00460_),
    .ZN(_00461_)
  );
  AND2_X1 _21147_ (
    .A1(_00459_),
    .A2(_00461_),
    .ZN(_00462_)
  );
  INV_X1 _21148_ (
    .A(_00462_),
    .ZN(_00463_)
  );
  AND2_X1 _21149_ (
    .A1(_00231_),
    .A2(_00462_),
    .ZN(_00464_)
  );
  INV_X1 _21150_ (
    .A(_00464_),
    .ZN(_00465_)
  );
  AND2_X1 _21151_ (
    .A1(_00230_),
    .A2(_00463_),
    .ZN(_00466_)
  );
  INV_X1 _21152_ (
    .A(_00466_),
    .ZN(_00467_)
  );
  AND2_X1 _21153_ (
    .A1(_00465_),
    .A2(_00467_),
    .ZN(_00468_)
  );
  INV_X1 _21154_ (
    .A(_00468_),
    .ZN(_00470_)
  );
  AND2_X1 _21155_ (
    .A1(_00228_),
    .A2(_00468_),
    .ZN(_00471_)
  );
  INV_X1 _21156_ (
    .A(_00471_),
    .ZN(_00472_)
  );
  AND2_X1 _21157_ (
    .A1(_00227_),
    .A2(_00470_),
    .ZN(_00473_)
  );
  INV_X1 _21158_ (
    .A(_00473_),
    .ZN(_00474_)
  );
  AND2_X1 _21159_ (
    .A1(_00472_),
    .A2(_00474_),
    .ZN(_00475_)
  );
  INV_X1 _21160_ (
    .A(_00475_),
    .ZN(_00476_)
  );
  AND2_X1 _21161_ (
    .A1(_00171_),
    .A2(_00475_),
    .ZN(_00477_)
  );
  INV_X1 _21162_ (
    .A(_00477_),
    .ZN(_00478_)
  );
  AND2_X1 _21163_ (
    .A1(_00172_),
    .A2(_00476_),
    .ZN(_00479_)
  );
  INV_X1 _21164_ (
    .A(_00479_),
    .ZN(_00481_)
  );
  AND2_X1 _21165_ (
    .A1(_00478_),
    .A2(_00481_),
    .ZN(_00482_)
  );
  INV_X1 _21166_ (
    .A(_00482_),
    .ZN(_00483_)
  );
  AND2_X1 _21167_ (
    .A1(_00226_),
    .A2(_00483_),
    .ZN(_00484_)
  );
  INV_X1 _21168_ (
    .A(_00484_),
    .ZN(_00485_)
  );
  AND2_X1 _21169_ (
    .A1(_00225_),
    .A2(_00482_),
    .ZN(_00486_)
  );
  INV_X1 _21170_ (
    .A(_00486_),
    .ZN(_00487_)
  );
  AND2_X1 _21171_ (
    .A1(_00225_),
    .A2(_00483_),
    .ZN(_00488_)
  );
  INV_X1 _21172_ (
    .A(_00488_),
    .ZN(_00489_)
  );
  AND2_X1 _21173_ (
    .A1(_00226_),
    .A2(_00482_),
    .ZN(_00490_)
  );
  INV_X1 _21174_ (
    .A(_00490_),
    .ZN(_00492_)
  );
  AND2_X1 _21175_ (
    .A1(_00485_),
    .A2(_00487_),
    .ZN(_00493_)
  );
  AND2_X1 _21176_ (
    .A1(_00489_),
    .A2(_00492_),
    .ZN(_00494_)
  );
  AND2_X1 _21177_ (
    .A1(_04404_),
    .A2(_00493_),
    .ZN(_00495_)
  );
  INV_X1 _21178_ (
    .A(_00495_),
    .ZN(_00496_)
  );
  AND2_X1 _21179_ (
    .A1(remainder[65]),
    .A2(_00494_),
    .ZN(_00497_)
  );
  INV_X1 _21180_ (
    .A(_00497_),
    .ZN(_00498_)
  );
  AND2_X1 _21181_ (
    .A1(_00496_),
    .A2(_00498_),
    .ZN(_00499_)
  );
  INV_X1 _21182_ (
    .A(_00499_),
    .ZN(_00500_)
  );
  AND2_X1 _21183_ (
    .A1(_00223_),
    .A2(_00500_),
    .ZN(_00501_)
  );
  INV_X1 _21184_ (
    .A(_00501_),
    .ZN(_00503_)
  );
  AND2_X1 _21185_ (
    .A1(_00224_),
    .A2(_00499_),
    .ZN(_00504_)
  );
  INV_X1 _21186_ (
    .A(_00504_),
    .ZN(_00505_)
  );
  AND2_X1 _21187_ (
    .A1(_02082_),
    .A2(_00505_),
    .ZN(_00506_)
  );
  AND2_X1 _21188_ (
    .A1(_00503_),
    .A2(_00506_),
    .ZN(_00507_)
  );
  INV_X1 _21189_ (
    .A(_00507_),
    .ZN(_00508_)
  );
  AND2_X1 _21190_ (
    .A1(remainder[64]),
    .A2(_02077_),
    .ZN(_00509_)
  );
  INV_X1 _21191_ (
    .A(_00509_),
    .ZN(_00510_)
  );
  AND2_X1 _21192_ (
    .A1(_10462_),
    .A2(_02061_),
    .ZN(_00511_)
  );
  INV_X1 _21193_ (
    .A(_00511_),
    .ZN(_00512_)
  );
  AND2_X1 _21194_ (
    .A1(_04426_),
    .A2(_10451_),
    .ZN(_00514_)
  );
  INV_X1 _21195_ (
    .A(_00514_),
    .ZN(_00515_)
  );
  AND2_X1 _21196_ (
    .A1(_05983_),
    .A2(_00512_),
    .ZN(_00516_)
  );
  AND2_X1 _21197_ (
    .A1(_00515_),
    .A2(_00516_),
    .ZN(_00517_)
  );
  INV_X1 _21198_ (
    .A(_00517_),
    .ZN(_00518_)
  );
  AND2_X1 _21199_ (
    .A1(_00510_),
    .A2(_00518_),
    .ZN(_00519_)
  );
  AND2_X1 _21200_ (
    .A1(_00508_),
    .A2(_00519_),
    .ZN(_00520_)
  );
  INV_X1 _21201_ (
    .A(_00520_),
    .ZN(_00521_)
  );
  AND2_X1 _21202_ (
    .A1(_06201_),
    .A2(_00521_),
    .ZN(_00085_)
  );
  AND2_X1 _21203_ (
    .A1(_10958_),
    .A2(_00200_),
    .ZN(_00522_)
  );
  AND2_X1 _21204_ (
    .A1(_00499_),
    .A2(_00522_),
    .ZN(_00524_)
  );
  INV_X1 _21205_ (
    .A(_00524_),
    .ZN(_00525_)
  );
  AND2_X1 _21206_ (
    .A1(_10960_),
    .A2(_00196_),
    .ZN(_00526_)
  );
  AND2_X1 _21207_ (
    .A1(_00498_),
    .A2(_00526_),
    .ZN(_00527_)
  );
  AND2_X1 _21208_ (
    .A1(_00525_),
    .A2(_00527_),
    .ZN(_00528_)
  );
  INV_X1 _21209_ (
    .A(_00528_),
    .ZN(_00529_)
  );
  AND2_X1 _21210_ (
    .A1(_00478_),
    .A2(_00492_),
    .ZN(_00530_)
  );
  INV_X1 _21211_ (
    .A(_00530_),
    .ZN(_00531_)
  );
  AND2_X1 _21212_ (
    .A1(_00459_),
    .A2(_00465_),
    .ZN(_00532_)
  );
  INV_X1 _21213_ (
    .A(_00532_),
    .ZN(_00533_)
  );
  AND2_X1 _21214_ (
    .A1(_00440_),
    .A2(_00446_),
    .ZN(_00535_)
  );
  INV_X1 _21215_ (
    .A(_00535_),
    .ZN(_00536_)
  );
  AND2_X1 _21216_ (
    .A1(_00431_),
    .A2(_00453_),
    .ZN(_00537_)
  );
  INV_X1 _21217_ (
    .A(_00537_),
    .ZN(_00538_)
  );
  AND2_X1 _21218_ (
    .A1(_00336_),
    .A2(_00396_),
    .ZN(_00539_)
  );
  INV_X1 _21219_ (
    .A(_00539_),
    .ZN(_00540_)
  );
  AND2_X1 _21220_ (
    .A1(_00279_),
    .A2(_00330_),
    .ZN(_00541_)
  );
  INV_X1 _21221_ (
    .A(_00541_),
    .ZN(_00542_)
  );
  AND2_X1 _21222_ (
    .A1(_00369_),
    .A2(_00376_),
    .ZN(_00543_)
  );
  INV_X1 _21223_ (
    .A(_00543_),
    .ZN(_00544_)
  );
  AND2_X1 _21224_ (
    .A1(_00542_),
    .A2(_00543_),
    .ZN(_00546_)
  );
  INV_X1 _21225_ (
    .A(_00546_),
    .ZN(_00547_)
  );
  AND2_X1 _21226_ (
    .A1(_00541_),
    .A2(_00544_),
    .ZN(_00548_)
  );
  INV_X1 _21227_ (
    .A(_00548_),
    .ZN(_00549_)
  );
  AND2_X1 _21228_ (
    .A1(_00541_),
    .A2(_00543_),
    .ZN(_00550_)
  );
  INV_X1 _21229_ (
    .A(_00550_),
    .ZN(_00551_)
  );
  AND2_X1 _21230_ (
    .A1(_00542_),
    .A2(_00544_),
    .ZN(_00552_)
  );
  INV_X1 _21231_ (
    .A(_00552_),
    .ZN(_00553_)
  );
  AND2_X1 _21232_ (
    .A1(_00547_),
    .A2(_00549_),
    .ZN(_00554_)
  );
  AND2_X1 _21233_ (
    .A1(_00551_),
    .A2(_00553_),
    .ZN(_00555_)
  );
  AND2_X1 _21234_ (
    .A1(_10684_),
    .A2(_00272_),
    .ZN(_00557_)
  );
  INV_X1 _21235_ (
    .A(_00557_),
    .ZN(_00558_)
  );
  AND2_X1 _21236_ (
    .A1(_00304_),
    .A2(_00311_),
    .ZN(_00559_)
  );
  INV_X1 _21237_ (
    .A(_00559_),
    .ZN(_00560_)
  );
  AND2_X1 _21238_ (
    .A1(_10492_),
    .A2(_00353_),
    .ZN(_00561_)
  );
  INV_X1 _21239_ (
    .A(_00561_),
    .ZN(_00562_)
  );
  AND2_X1 _21240_ (
    .A1(_00369_),
    .A2(_00562_),
    .ZN(_00563_)
  );
  INV_X1 _21241_ (
    .A(_00563_),
    .ZN(_00564_)
  );
  AND2_X1 _21242_ (
    .A1(_09521_),
    .A2(_00559_),
    .ZN(_00565_)
  );
  INV_X1 _21243_ (
    .A(_00565_),
    .ZN(_00566_)
  );
  AND2_X1 _21244_ (
    .A1(_09522_),
    .A2(_00560_),
    .ZN(_00568_)
  );
  INV_X1 _21245_ (
    .A(_00568_),
    .ZN(_00569_)
  );
  AND2_X1 _21246_ (
    .A1(_00566_),
    .A2(_00569_),
    .ZN(_00570_)
  );
  INV_X1 _21247_ (
    .A(_00570_),
    .ZN(_00571_)
  );
  AND2_X1 _21248_ (
    .A1(_00557_),
    .A2(_00571_),
    .ZN(_00572_)
  );
  INV_X1 _21249_ (
    .A(_00572_),
    .ZN(_00573_)
  );
  AND2_X1 _21250_ (
    .A1(_00558_),
    .A2(_00570_),
    .ZN(_00574_)
  );
  INV_X1 _21251_ (
    .A(_00574_),
    .ZN(_00575_)
  );
  AND2_X1 _21252_ (
    .A1(_00573_),
    .A2(_00575_),
    .ZN(_00576_)
  );
  INV_X1 _21253_ (
    .A(_00576_),
    .ZN(_00577_)
  );
  AND2_X1 _21254_ (
    .A1(_00563_),
    .A2(_00577_),
    .ZN(_00579_)
  );
  INV_X1 _21255_ (
    .A(_00579_),
    .ZN(_00580_)
  );
  AND2_X1 _21256_ (
    .A1(_00564_),
    .A2(_00576_),
    .ZN(_00581_)
  );
  INV_X1 _21257_ (
    .A(_00581_),
    .ZN(_00582_)
  );
  AND2_X1 _21258_ (
    .A1(_00580_),
    .A2(_00582_),
    .ZN(_00583_)
  );
  INV_X1 _21259_ (
    .A(_00583_),
    .ZN(_00584_)
  );
  AND2_X1 _21260_ (
    .A1(_00317_),
    .A2(_00323_),
    .ZN(_00585_)
  );
  INV_X1 _21261_ (
    .A(_00585_),
    .ZN(_00586_)
  );
  AND2_X1 _21262_ (
    .A1(_03249_),
    .A2(_10463_),
    .ZN(_00587_)
  );
  INV_X1 _21263_ (
    .A(_00587_),
    .ZN(_00588_)
  );
  AND2_X1 _21264_ (
    .A1(_10409_),
    .A2(_00253_),
    .ZN(_00590_)
  );
  INV_X1 _21265_ (
    .A(_00590_),
    .ZN(_00591_)
  );
  AND2_X1 _21266_ (
    .A1(_00588_),
    .A2(_00590_),
    .ZN(_00592_)
  );
  INV_X1 _21267_ (
    .A(_00592_),
    .ZN(_00593_)
  );
  AND2_X1 _21268_ (
    .A1(_00587_),
    .A2(_00591_),
    .ZN(_00594_)
  );
  INV_X1 _21269_ (
    .A(_00594_),
    .ZN(_00595_)
  );
  AND2_X1 _21270_ (
    .A1(_00588_),
    .A2(_00591_),
    .ZN(_00596_)
  );
  INV_X1 _21271_ (
    .A(_00596_),
    .ZN(_00597_)
  );
  AND2_X1 _21272_ (
    .A1(_00587_),
    .A2(_00590_),
    .ZN(_00598_)
  );
  INV_X1 _21273_ (
    .A(_00598_),
    .ZN(_00599_)
  );
  AND2_X1 _21274_ (
    .A1(_00593_),
    .A2(_00595_),
    .ZN(_00600_)
  );
  AND2_X1 _21275_ (
    .A1(_00597_),
    .A2(_00599_),
    .ZN(_00601_)
  );
  AND2_X1 _21276_ (
    .A1(_00259_),
    .A2(_00266_),
    .ZN(_00602_)
  );
  INV_X1 _21277_ (
    .A(_00602_),
    .ZN(_00603_)
  );
  AND2_X1 _21278_ (
    .A1(_00600_),
    .A2(_00602_),
    .ZN(_00604_)
  );
  INV_X1 _21279_ (
    .A(_00604_),
    .ZN(_00605_)
  );
  AND2_X1 _21280_ (
    .A1(_00601_),
    .A2(_00603_),
    .ZN(_00606_)
  );
  INV_X1 _21281_ (
    .A(_00606_),
    .ZN(_00607_)
  );
  AND2_X1 _21282_ (
    .A1(_00601_),
    .A2(_00602_),
    .ZN(_00608_)
  );
  INV_X1 _21283_ (
    .A(_00608_),
    .ZN(_00609_)
  );
  AND2_X1 _21284_ (
    .A1(_00600_),
    .A2(_00603_),
    .ZN(_00611_)
  );
  INV_X1 _21285_ (
    .A(_00611_),
    .ZN(_00612_)
  );
  AND2_X1 _21286_ (
    .A1(_00605_),
    .A2(_00607_),
    .ZN(_00613_)
  );
  AND2_X1 _21287_ (
    .A1(_00609_),
    .A2(_00612_),
    .ZN(_00614_)
  );
  AND2_X1 _21288_ (
    .A1(_10728_),
    .A2(_11013_),
    .ZN(_00615_)
  );
  INV_X1 _21289_ (
    .A(_00615_),
    .ZN(_00616_)
  );
  AND2_X1 _21290_ (
    .A1(_10727_),
    .A2(_11011_),
    .ZN(_00617_)
  );
  INV_X1 _21291_ (
    .A(_00617_),
    .ZN(_00618_)
  );
  AND2_X1 _21292_ (
    .A1(_10728_),
    .A2(_11011_),
    .ZN(_00619_)
  );
  INV_X1 _21293_ (
    .A(_00619_),
    .ZN(_00620_)
  );
  AND2_X1 _21294_ (
    .A1(_10727_),
    .A2(_11013_),
    .ZN(_00622_)
  );
  INV_X1 _21295_ (
    .A(_00622_),
    .ZN(_00623_)
  );
  AND2_X1 _21296_ (
    .A1(_00616_),
    .A2(_00618_),
    .ZN(_00624_)
  );
  AND2_X1 _21297_ (
    .A1(_00620_),
    .A2(_00623_),
    .ZN(_00625_)
  );
  AND2_X1 _21298_ (
    .A1(_10697_),
    .A2(_00625_),
    .ZN(_00626_)
  );
  INV_X1 _21299_ (
    .A(_00626_),
    .ZN(_00627_)
  );
  AND2_X1 _21300_ (
    .A1(_10696_),
    .A2(_00624_),
    .ZN(_00628_)
  );
  INV_X1 _21301_ (
    .A(_00628_),
    .ZN(_00629_)
  );
  AND2_X1 _21302_ (
    .A1(_10697_),
    .A2(_00624_),
    .ZN(_00630_)
  );
  INV_X1 _21303_ (
    .A(_00630_),
    .ZN(_00631_)
  );
  AND2_X1 _21304_ (
    .A1(_10696_),
    .A2(_00625_),
    .ZN(_00633_)
  );
  INV_X1 _21305_ (
    .A(_00633_),
    .ZN(_00634_)
  );
  AND2_X1 _21306_ (
    .A1(_00627_),
    .A2(_00629_),
    .ZN(_00635_)
  );
  AND2_X1 _21307_ (
    .A1(_00631_),
    .A2(_00634_),
    .ZN(_00636_)
  );
  AND2_X1 _21308_ (
    .A1(_09784_),
    .A2(_10690_),
    .ZN(_00637_)
  );
  INV_X1 _21309_ (
    .A(_00637_),
    .ZN(_00638_)
  );
  AND2_X1 _21310_ (
    .A1(_09785_),
    .A2(_10689_),
    .ZN(_00639_)
  );
  INV_X1 _21311_ (
    .A(_00639_),
    .ZN(_00640_)
  );
  AND2_X1 _21312_ (
    .A1(_09784_),
    .A2(_10689_),
    .ZN(_00641_)
  );
  INV_X1 _21313_ (
    .A(_00641_),
    .ZN(_00642_)
  );
  AND2_X1 _21314_ (
    .A1(_09785_),
    .A2(_10690_),
    .ZN(_00644_)
  );
  INV_X1 _21315_ (
    .A(_00644_),
    .ZN(_00645_)
  );
  AND2_X1 _21316_ (
    .A1(_00638_),
    .A2(_00640_),
    .ZN(_00646_)
  );
  AND2_X1 _21317_ (
    .A1(_00642_),
    .A2(_00645_),
    .ZN(_00647_)
  );
  AND2_X1 _21318_ (
    .A1(_00635_),
    .A2(_00646_),
    .ZN(_00648_)
  );
  INV_X1 _21319_ (
    .A(_00648_),
    .ZN(_00649_)
  );
  AND2_X1 _21320_ (
    .A1(_00636_),
    .A2(_00647_),
    .ZN(_00650_)
  );
  INV_X1 _21321_ (
    .A(_00650_),
    .ZN(_00651_)
  );
  AND2_X1 _21322_ (
    .A1(_00649_),
    .A2(_00651_),
    .ZN(_00652_)
  );
  INV_X1 _21323_ (
    .A(_00652_),
    .ZN(_00653_)
  );
  AND2_X1 _21324_ (
    .A1(_00293_),
    .A2(_00298_),
    .ZN(_00655_)
  );
  INV_X1 _21325_ (
    .A(_00655_),
    .ZN(_00656_)
  );
  AND2_X1 _21326_ (
    .A1(remainder[32]),
    .A2(remainder[7]),
    .ZN(_00657_)
  );
  INV_X1 _21327_ (
    .A(_00657_),
    .ZN(_00658_)
  );
  AND2_X1 _21328_ (
    .A1(_04766_),
    .A2(_05149_),
    .ZN(_00659_)
  );
  INV_X1 _21329_ (
    .A(_00659_),
    .ZN(_00660_)
  );
  AND2_X1 _21330_ (
    .A1(divisor[32]),
    .A2(_00660_),
    .ZN(_00661_)
  );
  AND2_X1 _21331_ (
    .A1(_00658_),
    .A2(_00661_),
    .ZN(_00662_)
  );
  INV_X1 _21332_ (
    .A(_00662_),
    .ZN(_00663_)
  );
  AND2_X1 _21333_ (
    .A1(_00655_),
    .A2(_00662_),
    .ZN(_00664_)
  );
  INV_X1 _21334_ (
    .A(_00664_),
    .ZN(_00666_)
  );
  AND2_X1 _21335_ (
    .A1(_00656_),
    .A2(_00663_),
    .ZN(_00667_)
  );
  INV_X1 _21336_ (
    .A(_00667_),
    .ZN(_00668_)
  );
  AND2_X1 _21337_ (
    .A1(_00656_),
    .A2(_00662_),
    .ZN(_00669_)
  );
  INV_X1 _21338_ (
    .A(_00669_),
    .ZN(_00670_)
  );
  AND2_X1 _21339_ (
    .A1(_00655_),
    .A2(_00663_),
    .ZN(_00671_)
  );
  INV_X1 _21340_ (
    .A(_00671_),
    .ZN(_00672_)
  );
  AND2_X1 _21341_ (
    .A1(_00666_),
    .A2(_00668_),
    .ZN(_00673_)
  );
  AND2_X1 _21342_ (
    .A1(_00670_),
    .A2(_00672_),
    .ZN(_00674_)
  );
  AND2_X1 _21343_ (
    .A1(_11035_),
    .A2(_00290_),
    .ZN(_00675_)
  );
  INV_X1 _21344_ (
    .A(_00675_),
    .ZN(_00677_)
  );
  AND2_X1 _21345_ (
    .A1(_11034_),
    .A2(_00289_),
    .ZN(_00678_)
  );
  INV_X1 _21346_ (
    .A(_00678_),
    .ZN(_00679_)
  );
  AND2_X1 _21347_ (
    .A1(_00677_),
    .A2(_00679_),
    .ZN(_00680_)
  );
  INV_X1 _21348_ (
    .A(_00680_),
    .ZN(_00681_)
  );
  AND2_X1 _21349_ (
    .A1(_00674_),
    .A2(_00680_),
    .ZN(_00682_)
  );
  INV_X1 _21350_ (
    .A(_00682_),
    .ZN(_00683_)
  );
  AND2_X1 _21351_ (
    .A1(_00673_),
    .A2(_00681_),
    .ZN(_00684_)
  );
  INV_X1 _21352_ (
    .A(_00684_),
    .ZN(_00685_)
  );
  AND2_X1 _21353_ (
    .A1(_00673_),
    .A2(_00680_),
    .ZN(_00686_)
  );
  INV_X1 _21354_ (
    .A(_00686_),
    .ZN(_00688_)
  );
  AND2_X1 _21355_ (
    .A1(_00674_),
    .A2(_00681_),
    .ZN(_00689_)
  );
  INV_X1 _21356_ (
    .A(_00689_),
    .ZN(_00690_)
  );
  AND2_X1 _21357_ (
    .A1(_00683_),
    .A2(_00685_),
    .ZN(_00691_)
  );
  AND2_X1 _21358_ (
    .A1(_00688_),
    .A2(_00690_),
    .ZN(_00692_)
  );
  AND2_X1 _21359_ (
    .A1(_00652_),
    .A2(_00692_),
    .ZN(_00693_)
  );
  INV_X1 _21360_ (
    .A(_00693_),
    .ZN(_00694_)
  );
  AND2_X1 _21361_ (
    .A1(_00653_),
    .A2(_00691_),
    .ZN(_00695_)
  );
  INV_X1 _21362_ (
    .A(_00695_),
    .ZN(_00696_)
  );
  AND2_X1 _21363_ (
    .A1(_00653_),
    .A2(_00692_),
    .ZN(_00697_)
  );
  INV_X1 _21364_ (
    .A(_00697_),
    .ZN(_00699_)
  );
  AND2_X1 _21365_ (
    .A1(_00652_),
    .A2(_00691_),
    .ZN(_00700_)
  );
  INV_X1 _21366_ (
    .A(_00700_),
    .ZN(_00701_)
  );
  AND2_X1 _21367_ (
    .A1(_00694_),
    .A2(_00696_),
    .ZN(_00702_)
  );
  AND2_X1 _21368_ (
    .A1(_00699_),
    .A2(_00701_),
    .ZN(_00703_)
  );
  AND2_X1 _21369_ (
    .A1(_00613_),
    .A2(_00703_),
    .ZN(_00704_)
  );
  INV_X1 _21370_ (
    .A(_00704_),
    .ZN(_00705_)
  );
  AND2_X1 _21371_ (
    .A1(_00614_),
    .A2(_00702_),
    .ZN(_00706_)
  );
  INV_X1 _21372_ (
    .A(_00706_),
    .ZN(_00707_)
  );
  AND2_X1 _21373_ (
    .A1(_00614_),
    .A2(_00703_),
    .ZN(_00708_)
  );
  INV_X1 _21374_ (
    .A(_00708_),
    .ZN(_00710_)
  );
  AND2_X1 _21375_ (
    .A1(_00613_),
    .A2(_00702_),
    .ZN(_00711_)
  );
  INV_X1 _21376_ (
    .A(_00711_),
    .ZN(_00712_)
  );
  AND2_X1 _21377_ (
    .A1(_00705_),
    .A2(_00707_),
    .ZN(_00713_)
  );
  AND2_X1 _21378_ (
    .A1(_00710_),
    .A2(_00712_),
    .ZN(_00714_)
  );
  AND2_X1 _21379_ (
    .A1(_00585_),
    .A2(_00713_),
    .ZN(_00715_)
  );
  INV_X1 _21380_ (
    .A(_00715_),
    .ZN(_00716_)
  );
  AND2_X1 _21381_ (
    .A1(_00586_),
    .A2(_00714_),
    .ZN(_00717_)
  );
  INV_X1 _21382_ (
    .A(_00717_),
    .ZN(_00718_)
  );
  AND2_X1 _21383_ (
    .A1(_00585_),
    .A2(_00714_),
    .ZN(_00719_)
  );
  INV_X1 _21384_ (
    .A(_00719_),
    .ZN(_00721_)
  );
  AND2_X1 _21385_ (
    .A1(_00586_),
    .A2(_00713_),
    .ZN(_00722_)
  );
  INV_X1 _21386_ (
    .A(_00722_),
    .ZN(_00723_)
  );
  AND2_X1 _21387_ (
    .A1(_00716_),
    .A2(_00718_),
    .ZN(_00724_)
  );
  AND2_X1 _21388_ (
    .A1(_00721_),
    .A2(_00723_),
    .ZN(_00725_)
  );
  AND2_X1 _21389_ (
    .A1(_00583_),
    .A2(_00724_),
    .ZN(_00726_)
  );
  INV_X1 _21390_ (
    .A(_00726_),
    .ZN(_00727_)
  );
  AND2_X1 _21391_ (
    .A1(_00584_),
    .A2(_00725_),
    .ZN(_00728_)
  );
  INV_X1 _21392_ (
    .A(_00728_),
    .ZN(_00729_)
  );
  AND2_X1 _21393_ (
    .A1(_00583_),
    .A2(_00725_),
    .ZN(_00730_)
  );
  INV_X1 _21394_ (
    .A(_00730_),
    .ZN(_00732_)
  );
  AND2_X1 _21395_ (
    .A1(_00584_),
    .A2(_00724_),
    .ZN(_00733_)
  );
  INV_X1 _21396_ (
    .A(_00733_),
    .ZN(_00734_)
  );
  AND2_X1 _21397_ (
    .A1(_00727_),
    .A2(_00729_),
    .ZN(_00735_)
  );
  AND2_X1 _21398_ (
    .A1(_00732_),
    .A2(_00734_),
    .ZN(_00736_)
  );
  AND2_X1 _21399_ (
    .A1(_00555_),
    .A2(_00736_),
    .ZN(_00737_)
  );
  INV_X1 _21400_ (
    .A(_00737_),
    .ZN(_00738_)
  );
  AND2_X1 _21401_ (
    .A1(_00554_),
    .A2(_00735_),
    .ZN(_00739_)
  );
  INV_X1 _21402_ (
    .A(_00739_),
    .ZN(_00740_)
  );
  AND2_X1 _21403_ (
    .A1(_00554_),
    .A2(_00736_),
    .ZN(_00741_)
  );
  INV_X1 _21404_ (
    .A(_00741_),
    .ZN(_00743_)
  );
  AND2_X1 _21405_ (
    .A1(_00555_),
    .A2(_00735_),
    .ZN(_00744_)
  );
  INV_X1 _21406_ (
    .A(_00744_),
    .ZN(_00745_)
  );
  AND2_X1 _21407_ (
    .A1(_00738_),
    .A2(_00740_),
    .ZN(_00746_)
  );
  AND2_X1 _21408_ (
    .A1(_00743_),
    .A2(_00745_),
    .ZN(_00747_)
  );
  AND2_X1 _21409_ (
    .A1(_00540_),
    .A2(_00746_),
    .ZN(_00748_)
  );
  INV_X1 _21410_ (
    .A(_00748_),
    .ZN(_00749_)
  );
  AND2_X1 _21411_ (
    .A1(_00539_),
    .A2(_00747_),
    .ZN(_00750_)
  );
  INV_X1 _21412_ (
    .A(_00750_),
    .ZN(_00751_)
  );
  AND2_X1 _21413_ (
    .A1(_00749_),
    .A2(_00751_),
    .ZN(_00752_)
  );
  INV_X1 _21414_ (
    .A(_00752_),
    .ZN(_00754_)
  );
  AND2_X1 _21415_ (
    .A1(_00383_),
    .A2(_00389_),
    .ZN(_00755_)
  );
  INV_X1 _21416_ (
    .A(_00755_),
    .ZN(_00756_)
  );
  AND2_X1 _21417_ (
    .A1(_10272_),
    .A2(_00755_),
    .ZN(_00757_)
  );
  INV_X1 _21418_ (
    .A(_00757_),
    .ZN(_00758_)
  );
  AND2_X1 _21419_ (
    .A1(_10271_),
    .A2(_00756_),
    .ZN(_00759_)
  );
  INV_X1 _21420_ (
    .A(_00759_),
    .ZN(_00760_)
  );
  AND2_X1 _21421_ (
    .A1(_10271_),
    .A2(_00755_),
    .ZN(_00761_)
  );
  INV_X1 _21422_ (
    .A(_00761_),
    .ZN(_00762_)
  );
  AND2_X1 _21423_ (
    .A1(_10272_),
    .A2(_00756_),
    .ZN(_00763_)
  );
  INV_X1 _21424_ (
    .A(_00763_),
    .ZN(_00765_)
  );
  AND2_X1 _21425_ (
    .A1(_00758_),
    .A2(_00760_),
    .ZN(_00766_)
  );
  AND2_X1 _21426_ (
    .A1(_00762_),
    .A2(_00765_),
    .ZN(_00767_)
  );
  AND2_X1 _21427_ (
    .A1(_10549_),
    .A2(_00766_),
    .ZN(_00768_)
  );
  INV_X1 _21428_ (
    .A(_00768_),
    .ZN(_00769_)
  );
  AND2_X1 _21429_ (
    .A1(_10551_),
    .A2(_00767_),
    .ZN(_00770_)
  );
  INV_X1 _21430_ (
    .A(_00770_),
    .ZN(_00771_)
  );
  AND2_X1 _21431_ (
    .A1(_00769_),
    .A2(_00771_),
    .ZN(_00772_)
  );
  INV_X1 _21432_ (
    .A(_00772_),
    .ZN(_00773_)
  );
  AND2_X1 _21433_ (
    .A1(_00752_),
    .A2(_00772_),
    .ZN(_00774_)
  );
  INV_X1 _21434_ (
    .A(_00774_),
    .ZN(_00776_)
  );
  AND2_X1 _21435_ (
    .A1(_00754_),
    .A2(_00773_),
    .ZN(_00777_)
  );
  INV_X1 _21436_ (
    .A(_00777_),
    .ZN(_00778_)
  );
  AND2_X1 _21437_ (
    .A1(_00747_),
    .A2(_00767_),
    .ZN(_00779_)
  );
  INV_X1 _21438_ (
    .A(_00779_),
    .ZN(_00780_)
  );
  AND2_X1 _21439_ (
    .A1(_00746_),
    .A2(_00766_),
    .ZN(_00781_)
  );
  INV_X1 _21440_ (
    .A(_00781_),
    .ZN(_00782_)
  );
  AND2_X1 _21441_ (
    .A1(_00780_),
    .A2(_00782_),
    .ZN(_00783_)
  );
  INV_X1 _21442_ (
    .A(_00783_),
    .ZN(_00784_)
  );
  AND2_X1 _21443_ (
    .A1(_10549_),
    .A2(_00539_),
    .ZN(_00785_)
  );
  INV_X1 _21444_ (
    .A(_00785_),
    .ZN(_00787_)
  );
  AND2_X1 _21445_ (
    .A1(_10551_),
    .A2(_00540_),
    .ZN(_00788_)
  );
  INV_X1 _21446_ (
    .A(_00788_),
    .ZN(_00789_)
  );
  AND2_X1 _21447_ (
    .A1(_00787_),
    .A2(_00789_),
    .ZN(_00790_)
  );
  INV_X1 _21448_ (
    .A(_00790_),
    .ZN(_00791_)
  );
  AND2_X1 _21449_ (
    .A1(_00783_),
    .A2(_00790_),
    .ZN(_00792_)
  );
  INV_X1 _21450_ (
    .A(_00792_),
    .ZN(_00793_)
  );
  AND2_X1 _21451_ (
    .A1(_00784_),
    .A2(_00791_),
    .ZN(_00794_)
  );
  INV_X1 _21452_ (
    .A(_00794_),
    .ZN(_00795_)
  );
  AND2_X1 _21453_ (
    .A1(_00776_),
    .A2(_00778_),
    .ZN(_00796_)
  );
  AND2_X1 _21454_ (
    .A1(_00793_),
    .A2(_00795_),
    .ZN(_00798_)
  );
  MUX2_X1 _21455_ (
    .A(_03169_),
    .B(_07803_),
    .S(_07494_),
    .Z(_00799_)
  );
  MUX2_X1 _21456_ (
    .A(_03170_),
    .B(_07802_),
    .S(_07494_),
    .Z(_00800_)
  );
  AND2_X1 _21457_ (
    .A1(_00798_),
    .A2(_00800_),
    .ZN(_00801_)
  );
  INV_X1 _21458_ (
    .A(_00801_),
    .ZN(_00802_)
  );
  AND2_X1 _21459_ (
    .A1(_00796_),
    .A2(_00799_),
    .ZN(_00803_)
  );
  INV_X1 _21460_ (
    .A(_00803_),
    .ZN(_00804_)
  );
  AND2_X1 _21461_ (
    .A1(_00802_),
    .A2(_00804_),
    .ZN(_00805_)
  );
  INV_X1 _21462_ (
    .A(_00805_),
    .ZN(_00806_)
  );
  AND2_X1 _21463_ (
    .A1(_00402_),
    .A2(_00424_),
    .ZN(_00807_)
  );
  INV_X1 _21464_ (
    .A(_00807_),
    .ZN(_00809_)
  );
  AND2_X1 _21465_ (
    .A1(_00411_),
    .A2(_00418_),
    .ZN(_00810_)
  );
  INV_X1 _21466_ (
    .A(_00810_),
    .ZN(_00811_)
  );
  AND2_X1 _21467_ (
    .A1(_00807_),
    .A2(_00810_),
    .ZN(_00812_)
  );
  INV_X1 _21468_ (
    .A(_00812_),
    .ZN(_00813_)
  );
  AND2_X1 _21469_ (
    .A1(_00809_),
    .A2(_00811_),
    .ZN(_00814_)
  );
  INV_X1 _21470_ (
    .A(_00814_),
    .ZN(_00815_)
  );
  AND2_X1 _21471_ (
    .A1(_00813_),
    .A2(_00815_),
    .ZN(_00816_)
  );
  INV_X1 _21472_ (
    .A(_00816_),
    .ZN(_00817_)
  );
  AND2_X1 _21473_ (
    .A1(_00805_),
    .A2(_00816_),
    .ZN(_00818_)
  );
  INV_X1 _21474_ (
    .A(_00818_),
    .ZN(_00820_)
  );
  AND2_X1 _21475_ (
    .A1(_00806_),
    .A2(_00817_),
    .ZN(_00821_)
  );
  INV_X1 _21476_ (
    .A(_00821_),
    .ZN(_00822_)
  );
  AND2_X1 _21477_ (
    .A1(_00820_),
    .A2(_00822_),
    .ZN(_00823_)
  );
  INV_X1 _21478_ (
    .A(_00823_),
    .ZN(_00824_)
  );
  AND2_X1 _21479_ (
    .A1(_00538_),
    .A2(_00823_),
    .ZN(_00825_)
  );
  INV_X1 _21480_ (
    .A(_00825_),
    .ZN(_00826_)
  );
  AND2_X1 _21481_ (
    .A1(_00537_),
    .A2(_00824_),
    .ZN(_00827_)
  );
  INV_X1 _21482_ (
    .A(_00827_),
    .ZN(_00828_)
  );
  AND2_X1 _21483_ (
    .A1(_00538_),
    .A2(_00824_),
    .ZN(_00829_)
  );
  INV_X1 _21484_ (
    .A(_00829_),
    .ZN(_00830_)
  );
  AND2_X1 _21485_ (
    .A1(_00537_),
    .A2(_00823_),
    .ZN(_00831_)
  );
  INV_X1 _21486_ (
    .A(_00831_),
    .ZN(_00832_)
  );
  AND2_X1 _21487_ (
    .A1(_00826_),
    .A2(_00828_),
    .ZN(_00833_)
  );
  AND2_X1 _21488_ (
    .A1(_00830_),
    .A2(_00832_),
    .ZN(_00834_)
  );
  AND2_X1 _21489_ (
    .A1(_00535_),
    .A2(_00833_),
    .ZN(_00835_)
  );
  INV_X1 _21490_ (
    .A(_00835_),
    .ZN(_00836_)
  );
  AND2_X1 _21491_ (
    .A1(_00536_),
    .A2(_00834_),
    .ZN(_00837_)
  );
  INV_X1 _21492_ (
    .A(_00837_),
    .ZN(_00838_)
  );
  AND2_X1 _21493_ (
    .A1(_00535_),
    .A2(_00834_),
    .ZN(_00839_)
  );
  INV_X1 _21494_ (
    .A(_00839_),
    .ZN(_00841_)
  );
  AND2_X1 _21495_ (
    .A1(_00536_),
    .A2(_00833_),
    .ZN(_00842_)
  );
  INV_X1 _21496_ (
    .A(_00842_),
    .ZN(_00843_)
  );
  AND2_X1 _21497_ (
    .A1(_00836_),
    .A2(_00838_),
    .ZN(_00844_)
  );
  AND2_X1 _21498_ (
    .A1(_00841_),
    .A2(_00843_),
    .ZN(_00845_)
  );
  AND2_X1 _21499_ (
    .A1(_00533_),
    .A2(_00844_),
    .ZN(_00846_)
  );
  INV_X1 _21500_ (
    .A(_00846_),
    .ZN(_00847_)
  );
  AND2_X1 _21501_ (
    .A1(_00532_),
    .A2(_00845_),
    .ZN(_00848_)
  );
  INV_X1 _21502_ (
    .A(_00848_),
    .ZN(_00849_)
  );
  AND2_X1 _21503_ (
    .A1(_00533_),
    .A2(_00845_),
    .ZN(_00850_)
  );
  INV_X1 _21504_ (
    .A(_00850_),
    .ZN(_00852_)
  );
  AND2_X1 _21505_ (
    .A1(_00532_),
    .A2(_00844_),
    .ZN(_00853_)
  );
  INV_X1 _21506_ (
    .A(_00853_),
    .ZN(_00854_)
  );
  AND2_X1 _21507_ (
    .A1(_00847_),
    .A2(_00849_),
    .ZN(_00855_)
  );
  AND2_X1 _21508_ (
    .A1(_00852_),
    .A2(_00854_),
    .ZN(_00856_)
  );
  AND2_X1 _21509_ (
    .A1(_04404_),
    .A2(_00472_),
    .ZN(_00857_)
  );
  INV_X1 _21510_ (
    .A(_00857_),
    .ZN(_00858_)
  );
  AND2_X1 _21511_ (
    .A1(remainder[65]),
    .A2(_00471_),
    .ZN(_00859_)
  );
  INV_X1 _21512_ (
    .A(_00859_),
    .ZN(_00860_)
  );
  AND2_X1 _21513_ (
    .A1(_04404_),
    .A2(_00471_),
    .ZN(_00861_)
  );
  INV_X1 _21514_ (
    .A(_00861_),
    .ZN(_00863_)
  );
  AND2_X1 _21515_ (
    .A1(remainder[65]),
    .A2(_00472_),
    .ZN(_00864_)
  );
  INV_X1 _21516_ (
    .A(_00864_),
    .ZN(_00865_)
  );
  AND2_X1 _21517_ (
    .A1(_00858_),
    .A2(_00860_),
    .ZN(_00866_)
  );
  AND2_X1 _21518_ (
    .A1(_00863_),
    .A2(_00865_),
    .ZN(_00867_)
  );
  AND2_X1 _21519_ (
    .A1(_00855_),
    .A2(_00867_),
    .ZN(_00868_)
  );
  INV_X1 _21520_ (
    .A(_00868_),
    .ZN(_00869_)
  );
  AND2_X1 _21521_ (
    .A1(_00856_),
    .A2(_00866_),
    .ZN(_00870_)
  );
  INV_X1 _21522_ (
    .A(_00870_),
    .ZN(_00871_)
  );
  AND2_X1 _21523_ (
    .A1(_00856_),
    .A2(_00867_),
    .ZN(_00872_)
  );
  INV_X1 _21524_ (
    .A(_00872_),
    .ZN(_00874_)
  );
  AND2_X1 _21525_ (
    .A1(_00855_),
    .A2(_00866_),
    .ZN(_00875_)
  );
  INV_X1 _21526_ (
    .A(_00875_),
    .ZN(_00876_)
  );
  AND2_X1 _21527_ (
    .A1(_00869_),
    .A2(_00871_),
    .ZN(_00877_)
  );
  AND2_X1 _21528_ (
    .A1(_00874_),
    .A2(_00876_),
    .ZN(_00878_)
  );
  AND2_X1 _21529_ (
    .A1(_00531_),
    .A2(_00878_),
    .ZN(_00879_)
  );
  INV_X1 _21530_ (
    .A(_00879_),
    .ZN(_00880_)
  );
  AND2_X1 _21531_ (
    .A1(_00530_),
    .A2(_00877_),
    .ZN(_00881_)
  );
  INV_X1 _21532_ (
    .A(_00881_),
    .ZN(_00882_)
  );
  AND2_X1 _21533_ (
    .A1(_00530_),
    .A2(_00878_),
    .ZN(_00883_)
  );
  INV_X1 _21534_ (
    .A(_00883_),
    .ZN(_00885_)
  );
  AND2_X1 _21535_ (
    .A1(_00531_),
    .A2(_00877_),
    .ZN(_00886_)
  );
  INV_X1 _21536_ (
    .A(_00886_),
    .ZN(_00887_)
  );
  AND2_X1 _21537_ (
    .A1(_00880_),
    .A2(_00882_),
    .ZN(_00888_)
  );
  AND2_X1 _21538_ (
    .A1(_00885_),
    .A2(_00887_),
    .ZN(_00889_)
  );
  AND2_X1 _21539_ (
    .A1(_00528_),
    .A2(_00889_),
    .ZN(_00890_)
  );
  INV_X1 _21540_ (
    .A(_00890_),
    .ZN(_00891_)
  );
  AND2_X1 _21541_ (
    .A1(_00529_),
    .A2(_00888_),
    .ZN(_00892_)
  );
  INV_X1 _21542_ (
    .A(_00892_),
    .ZN(_00893_)
  );
  AND2_X1 _21543_ (
    .A1(_06103_),
    .A2(_00893_),
    .ZN(_00894_)
  );
  AND2_X1 _21544_ (
    .A1(_00891_),
    .A2(_00894_),
    .ZN(_00896_)
  );
  INV_X1 _21545_ (
    .A(_00896_),
    .ZN(_00897_)
  );
  AND2_X1 _21546_ (
    .A1(_06114_),
    .A2(_02076_),
    .ZN(_00898_)
  );
  INV_X1 _21547_ (
    .A(_00898_),
    .ZN(_00899_)
  );
  AND2_X1 _21548_ (
    .A1(_05994_),
    .A2(_06201_),
    .ZN(_00900_)
  );
  AND2_X1 _21549_ (
    .A1(_04404_),
    .A2(_06114_),
    .ZN(_00901_)
  );
  INV_X1 _21550_ (
    .A(_00901_),
    .ZN(_00902_)
  );
  AND2_X1 _21551_ (
    .A1(_00900_),
    .A2(_00902_),
    .ZN(_00903_)
  );
  AND2_X1 _21552_ (
    .A1(_00899_),
    .A2(_00903_),
    .ZN(_00904_)
  );
  AND2_X1 _21553_ (
    .A1(_00897_),
    .A2(_00904_),
    .ZN(_00086_)
  );
  AND2_X1 _21554_ (
    .A1(remainder[8]),
    .A2(_06103_),
    .ZN(_00906_)
  );
  INV_X1 _21555_ (
    .A(_00906_),
    .ZN(_00907_)
  );
  MUX2_X1 _21556_ (
    .A(remainder[0]),
    .B(remainder[33]),
    .S(resHi),
    .Z(io_resp_bits_data[0])
  );
  INV_X1 _21557_ (
    .A(io_resp_bits_data[0]),
    .ZN(_00908_)
  );
  AND2_X1 _21558_ (
    .A1(_00898_),
    .A2(io_resp_bits_data[0]),
    .ZN(_00909_)
  );
  INV_X1 _21559_ (
    .A(_00909_),
    .ZN(_00910_)
  );
  AND2_X1 _21560_ (
    .A1(_00907_),
    .A2(_00910_),
    .ZN(_00911_)
  );
  INV_X1 _21561_ (
    .A(_00911_),
    .ZN(_00912_)
  );
  MUX2_X1 _21562_ (
    .A(_10462_),
    .B(_00912_),
    .S(_05994_),
    .Z(_00913_)
  );
  AND2_X1 _21563_ (
    .A1(_06201_),
    .A2(_00913_),
    .ZN(_00914_)
  );
  INV_X1 _21564_ (
    .A(_00914_),
    .ZN(_00916_)
  );
  AND2_X1 _21565_ (
    .A1(io_req_bits_in1[0]),
    .A2(_06190_),
    .ZN(_00917_)
  );
  INV_X1 _21566_ (
    .A(_00917_),
    .ZN(_00918_)
  );
  AND2_X1 _21567_ (
    .A1(_06201_),
    .A2(_02077_),
    .ZN(_00919_)
  );
  AND2_X1 _21568_ (
    .A1(remainder[0]),
    .A2(_00919_),
    .ZN(_00920_)
  );
  INV_X1 _21569_ (
    .A(_00920_),
    .ZN(_00921_)
  );
  AND2_X1 _21570_ (
    .A1(_00918_),
    .A2(_00921_),
    .ZN(_00922_)
  );
  AND2_X1 _21571_ (
    .A1(_00916_),
    .A2(_00922_),
    .ZN(_00923_)
  );
  INV_X1 _21572_ (
    .A(_00923_),
    .ZN(_00087_)
  );
  AND2_X1 _21573_ (
    .A1(remainder[1]),
    .A2(_00919_),
    .ZN(_00924_)
  );
  INV_X1 _21574_ (
    .A(_00924_),
    .ZN(_00926_)
  );
  MUX2_X1 _21575_ (
    .A(remainder[1]),
    .B(remainder[34]),
    .S(resHi),
    .Z(io_resp_bits_data[1])
  );
  INV_X1 _21576_ (
    .A(io_resp_bits_data[1]),
    .ZN(_00927_)
  );
  AND2_X1 _21577_ (
    .A1(_00908_),
    .A2(_00927_),
    .ZN(_00928_)
  );
  INV_X1 _21578_ (
    .A(_00928_),
    .ZN(_00929_)
  );
  AND2_X1 _21579_ (
    .A1(io_resp_bits_data[0]),
    .A2(io_resp_bits_data[1]),
    .ZN(_00930_)
  );
  INV_X1 _21580_ (
    .A(_00930_),
    .ZN(_00931_)
  );
  AND2_X1 _21581_ (
    .A1(_00929_),
    .A2(_00931_),
    .ZN(_00932_)
  );
  AND2_X1 _21582_ (
    .A1(_00898_),
    .A2(_00932_),
    .ZN(_00933_)
  );
  INV_X1 _21583_ (
    .A(_00933_),
    .ZN(_00934_)
  );
  AND2_X1 _21584_ (
    .A1(remainder[9]),
    .A2(_06103_),
    .ZN(_00936_)
  );
  INV_X1 _21585_ (
    .A(_00936_),
    .ZN(_00937_)
  );
  AND2_X1 _21586_ (
    .A1(_00934_),
    .A2(_00937_),
    .ZN(_00938_)
  );
  MUX2_X1 _21587_ (
    .A(_05073_),
    .B(_00938_),
    .S(_05994_),
    .Z(_00939_)
  );
  MUX2_X1 _21588_ (
    .A(_05533_),
    .B(_00939_),
    .S(_06201_),
    .Z(_00940_)
  );
  AND2_X1 _21589_ (
    .A1(_00926_),
    .A2(_00940_),
    .ZN(_00941_)
  );
  INV_X1 _21590_ (
    .A(_00941_),
    .ZN(_00088_)
  );
  AND2_X1 _21591_ (
    .A1(remainder[2]),
    .A2(_00919_),
    .ZN(_00942_)
  );
  INV_X1 _21592_ (
    .A(_00942_),
    .ZN(_00943_)
  );
  AND2_X1 _21593_ (
    .A1(remainder[10]),
    .A2(_06103_),
    .ZN(_00944_)
  );
  INV_X1 _21594_ (
    .A(_00944_),
    .ZN(_00946_)
  );
  AND2_X1 _21595_ (
    .A1(_05994_),
    .A2(_00946_),
    .ZN(_00947_)
  );
  MUX2_X1 _21596_ (
    .A(remainder[2]),
    .B(remainder[35]),
    .S(resHi),
    .Z(io_resp_bits_data[2])
  );
  INV_X1 _21597_ (
    .A(io_resp_bits_data[2]),
    .ZN(_00948_)
  );
  AND2_X1 _21598_ (
    .A1(_00929_),
    .A2(io_resp_bits_data[2]),
    .ZN(_00949_)
  );
  INV_X1 _21599_ (
    .A(_00949_),
    .ZN(_00950_)
  );
  AND2_X1 _21600_ (
    .A1(_00928_),
    .A2(_00948_),
    .ZN(_00951_)
  );
  INV_X1 _21601_ (
    .A(_00951_),
    .ZN(_00952_)
  );
  AND2_X1 _21602_ (
    .A1(_00950_),
    .A2(_00952_),
    .ZN(_00953_)
  );
  AND2_X1 _21603_ (
    .A1(_00898_),
    .A2(_00953_),
    .ZN(_00954_)
  );
  INV_X1 _21604_ (
    .A(_00954_),
    .ZN(_00956_)
  );
  AND2_X1 _21605_ (
    .A1(_00947_),
    .A2(_00956_),
    .ZN(_00957_)
  );
  INV_X1 _21606_ (
    .A(_00957_),
    .ZN(_00958_)
  );
  AND2_X1 _21607_ (
    .A1(_05084_),
    .A2(_05983_),
    .ZN(_00959_)
  );
  INV_X1 _21608_ (
    .A(_00959_),
    .ZN(_00960_)
  );
  AND2_X1 _21609_ (
    .A1(_00958_),
    .A2(_00960_),
    .ZN(_00961_)
  );
  MUX2_X1 _21610_ (
    .A(io_req_bits_in1[2]),
    .B(_00961_),
    .S(_06201_),
    .Z(_00962_)
  );
  INV_X1 _21611_ (
    .A(_00962_),
    .ZN(_00963_)
  );
  AND2_X1 _21612_ (
    .A1(_00943_),
    .A2(_00963_),
    .ZN(_00964_)
  );
  INV_X1 _21613_ (
    .A(_00964_),
    .ZN(_00089_)
  );
  AND2_X1 _21614_ (
    .A1(remainder[3]),
    .A2(_00919_),
    .ZN(_00965_)
  );
  INV_X1 _21615_ (
    .A(_00965_),
    .ZN(_00966_)
  );
  AND2_X1 _21616_ (
    .A1(remainder[11]),
    .A2(_06103_),
    .ZN(_00967_)
  );
  INV_X1 _21617_ (
    .A(_00967_),
    .ZN(_00968_)
  );
  AND2_X1 _21618_ (
    .A1(_05994_),
    .A2(_00968_),
    .ZN(_00969_)
  );
  MUX2_X1 _21619_ (
    .A(remainder[3]),
    .B(remainder[36]),
    .S(resHi),
    .Z(io_resp_bits_data[3])
  );
  INV_X1 _21620_ (
    .A(io_resp_bits_data[3]),
    .ZN(_00970_)
  );
  AND2_X1 _21621_ (
    .A1(_00952_),
    .A2(io_resp_bits_data[3]),
    .ZN(_00971_)
  );
  INV_X1 _21622_ (
    .A(_00971_),
    .ZN(_00972_)
  );
  AND2_X1 _21623_ (
    .A1(_00951_),
    .A2(_00970_),
    .ZN(_00973_)
  );
  INV_X1 _21624_ (
    .A(_00973_),
    .ZN(_00975_)
  );
  AND2_X1 _21625_ (
    .A1(_00972_),
    .A2(_00975_),
    .ZN(_00976_)
  );
  AND2_X1 _21626_ (
    .A1(_00898_),
    .A2(_00976_),
    .ZN(_00977_)
  );
  INV_X1 _21627_ (
    .A(_00977_),
    .ZN(_00978_)
  );
  AND2_X1 _21628_ (
    .A1(_00969_),
    .A2(_00978_),
    .ZN(_00979_)
  );
  INV_X1 _21629_ (
    .A(_00979_),
    .ZN(_00980_)
  );
  AND2_X1 _21630_ (
    .A1(_05095_),
    .A2(_05983_),
    .ZN(_00981_)
  );
  INV_X1 _21631_ (
    .A(_00981_),
    .ZN(_00982_)
  );
  AND2_X1 _21632_ (
    .A1(_00980_),
    .A2(_00982_),
    .ZN(_00983_)
  );
  MUX2_X1 _21633_ (
    .A(io_req_bits_in1[3]),
    .B(_00983_),
    .S(_06201_),
    .Z(_00984_)
  );
  INV_X1 _21634_ (
    .A(_00984_),
    .ZN(_00986_)
  );
  AND2_X1 _21635_ (
    .A1(_00966_),
    .A2(_00986_),
    .ZN(_00987_)
  );
  INV_X1 _21636_ (
    .A(_00987_),
    .ZN(_00090_)
  );
  AND2_X1 _21637_ (
    .A1(remainder[4]),
    .A2(_00919_),
    .ZN(_00988_)
  );
  INV_X1 _21638_ (
    .A(_00988_),
    .ZN(_00989_)
  );
  AND2_X1 _21639_ (
    .A1(remainder[12]),
    .A2(_06103_),
    .ZN(_00990_)
  );
  INV_X1 _21640_ (
    .A(_00990_),
    .ZN(_00991_)
  );
  AND2_X1 _21641_ (
    .A1(_05994_),
    .A2(_00991_),
    .ZN(_00992_)
  );
  MUX2_X1 _21642_ (
    .A(remainder[4]),
    .B(remainder[37]),
    .S(resHi),
    .Z(io_resp_bits_data[4])
  );
  INV_X1 _21643_ (
    .A(io_resp_bits_data[4]),
    .ZN(_00993_)
  );
  AND2_X1 _21644_ (
    .A1(_00975_),
    .A2(io_resp_bits_data[4]),
    .ZN(_00995_)
  );
  INV_X1 _21645_ (
    .A(_00995_),
    .ZN(_00996_)
  );
  AND2_X1 _21646_ (
    .A1(_00973_),
    .A2(_00993_),
    .ZN(_00997_)
  );
  INV_X1 _21647_ (
    .A(_00997_),
    .ZN(_00998_)
  );
  AND2_X1 _21648_ (
    .A1(_00996_),
    .A2(_00998_),
    .ZN(_00999_)
  );
  AND2_X1 _21649_ (
    .A1(_00898_),
    .A2(_00999_),
    .ZN(_01000_)
  );
  INV_X1 _21650_ (
    .A(_01000_),
    .ZN(_01001_)
  );
  AND2_X1 _21651_ (
    .A1(_00992_),
    .A2(_01001_),
    .ZN(_01002_)
  );
  INV_X1 _21652_ (
    .A(_01002_),
    .ZN(_01003_)
  );
  AND2_X1 _21653_ (
    .A1(_05105_),
    .A2(_05983_),
    .ZN(_01004_)
  );
  INV_X1 _21654_ (
    .A(_01004_),
    .ZN(_01006_)
  );
  AND2_X1 _21655_ (
    .A1(_01003_),
    .A2(_01006_),
    .ZN(_01007_)
  );
  MUX2_X1 _21656_ (
    .A(io_req_bits_in1[4]),
    .B(_01007_),
    .S(_06201_),
    .Z(_01008_)
  );
  INV_X1 _21657_ (
    .A(_01008_),
    .ZN(_01009_)
  );
  AND2_X1 _21658_ (
    .A1(_00989_),
    .A2(_01009_),
    .ZN(_01010_)
  );
  INV_X1 _21659_ (
    .A(_01010_),
    .ZN(_00091_)
  );
  AND2_X1 _21660_ (
    .A1(remainder[5]),
    .A2(_00919_),
    .ZN(_01011_)
  );
  INV_X1 _21661_ (
    .A(_01011_),
    .ZN(_01012_)
  );
  AND2_X1 _21662_ (
    .A1(_05116_),
    .A2(_05983_),
    .ZN(_01013_)
  );
  INV_X1 _21663_ (
    .A(_01013_),
    .ZN(_01014_)
  );
  AND2_X1 _21664_ (
    .A1(remainder[13]),
    .A2(_06103_),
    .ZN(_01016_)
  );
  INV_X1 _21665_ (
    .A(_01016_),
    .ZN(_01017_)
  );
  AND2_X1 _21666_ (
    .A1(_05994_),
    .A2(_01017_),
    .ZN(_01018_)
  );
  MUX2_X1 _21667_ (
    .A(remainder[5]),
    .B(remainder[38]),
    .S(resHi),
    .Z(io_resp_bits_data[5])
  );
  INV_X1 _21668_ (
    .A(io_resp_bits_data[5]),
    .ZN(_01019_)
  );
  AND2_X1 _21669_ (
    .A1(_00998_),
    .A2(io_resp_bits_data[5]),
    .ZN(_01020_)
  );
  INV_X1 _21670_ (
    .A(_01020_),
    .ZN(_01021_)
  );
  AND2_X1 _21671_ (
    .A1(_00997_),
    .A2(_01019_),
    .ZN(_01022_)
  );
  INV_X1 _21672_ (
    .A(_01022_),
    .ZN(_01023_)
  );
  AND2_X1 _21673_ (
    .A1(_00898_),
    .A2(_01023_),
    .ZN(_01024_)
  );
  AND2_X1 _21674_ (
    .A1(_01021_),
    .A2(_01024_),
    .ZN(_01026_)
  );
  INV_X1 _21675_ (
    .A(_01026_),
    .ZN(_01027_)
  );
  AND2_X1 _21676_ (
    .A1(_01018_),
    .A2(_01027_),
    .ZN(_01028_)
  );
  INV_X1 _21677_ (
    .A(_01028_),
    .ZN(_01029_)
  );
  AND2_X1 _21678_ (
    .A1(_01014_),
    .A2(_01029_),
    .ZN(_01030_)
  );
  MUX2_X1 _21679_ (
    .A(io_req_bits_in1[5]),
    .B(_01030_),
    .S(_06201_),
    .Z(_01031_)
  );
  INV_X1 _21680_ (
    .A(_01031_),
    .ZN(_01032_)
  );
  AND2_X1 _21681_ (
    .A1(_01012_),
    .A2(_01032_),
    .ZN(_01033_)
  );
  INV_X1 _21682_ (
    .A(_01033_),
    .ZN(_00092_)
  );
  AND2_X1 _21683_ (
    .A1(remainder[6]),
    .A2(_00919_),
    .ZN(_01034_)
  );
  INV_X1 _21684_ (
    .A(_01034_),
    .ZN(_01036_)
  );
  AND2_X1 _21685_ (
    .A1(remainder[14]),
    .A2(_06103_),
    .ZN(_01037_)
  );
  INV_X1 _21686_ (
    .A(_01037_),
    .ZN(_01038_)
  );
  AND2_X1 _21687_ (
    .A1(_05994_),
    .A2(_01038_),
    .ZN(_01039_)
  );
  MUX2_X1 _21688_ (
    .A(remainder[6]),
    .B(remainder[39]),
    .S(resHi),
    .Z(io_resp_bits_data[6])
  );
  INV_X1 _21689_ (
    .A(io_resp_bits_data[6]),
    .ZN(_01040_)
  );
  AND2_X1 _21690_ (
    .A1(_01022_),
    .A2(_01040_),
    .ZN(_01041_)
  );
  INV_X1 _21691_ (
    .A(_01041_),
    .ZN(_01042_)
  );
  AND2_X1 _21692_ (
    .A1(_01023_),
    .A2(io_resp_bits_data[6]),
    .ZN(_01043_)
  );
  INV_X1 _21693_ (
    .A(_01043_),
    .ZN(_01044_)
  );
  AND2_X1 _21694_ (
    .A1(_01042_),
    .A2(_01044_),
    .ZN(_01046_)
  );
  AND2_X1 _21695_ (
    .A1(_00898_),
    .A2(_01046_),
    .ZN(_01047_)
  );
  INV_X1 _21696_ (
    .A(_01047_),
    .ZN(_01048_)
  );
  AND2_X1 _21697_ (
    .A1(_01039_),
    .A2(_01048_),
    .ZN(_01049_)
  );
  INV_X1 _21698_ (
    .A(_01049_),
    .ZN(_01050_)
  );
  AND2_X1 _21699_ (
    .A1(_05127_),
    .A2(_05983_),
    .ZN(_01051_)
  );
  INV_X1 _21700_ (
    .A(_01051_),
    .ZN(_01052_)
  );
  AND2_X1 _21701_ (
    .A1(_01050_),
    .A2(_01052_),
    .ZN(_01053_)
  );
  MUX2_X1 _21702_ (
    .A(io_req_bits_in1[6]),
    .B(_01053_),
    .S(_06201_),
    .Z(_01054_)
  );
  INV_X1 _21703_ (
    .A(_01054_),
    .ZN(_01055_)
  );
  AND2_X1 _21704_ (
    .A1(_01036_),
    .A2(_01055_),
    .ZN(_01057_)
  );
  INV_X1 _21705_ (
    .A(_01057_),
    .ZN(_00093_)
  );
  AND2_X1 _21706_ (
    .A1(remainder[15]),
    .A2(_06103_),
    .ZN(_01058_)
  );
  INV_X1 _21707_ (
    .A(_01058_),
    .ZN(_01059_)
  );
  AND2_X1 _21708_ (
    .A1(_05994_),
    .A2(_01059_),
    .ZN(_01060_)
  );
  MUX2_X1 _21709_ (
    .A(remainder[7]),
    .B(remainder[40]),
    .S(resHi),
    .Z(io_resp_bits_data[7])
  );
  INV_X1 _21710_ (
    .A(io_resp_bits_data[7]),
    .ZN(_01061_)
  );
  AND2_X1 _21711_ (
    .A1(_01042_),
    .A2(io_resp_bits_data[7]),
    .ZN(_01062_)
  );
  INV_X1 _21712_ (
    .A(_01062_),
    .ZN(_01063_)
  );
  AND2_X1 _21713_ (
    .A1(_01041_),
    .A2(_01061_),
    .ZN(_01064_)
  );
  INV_X1 _21714_ (
    .A(_01064_),
    .ZN(_01066_)
  );
  AND2_X1 _21715_ (
    .A1(_00898_),
    .A2(_01066_),
    .ZN(_01067_)
  );
  AND2_X1 _21716_ (
    .A1(_01063_),
    .A2(_01067_),
    .ZN(_01068_)
  );
  INV_X1 _21717_ (
    .A(_01068_),
    .ZN(_01069_)
  );
  AND2_X1 _21718_ (
    .A1(_01060_),
    .A2(_01069_),
    .ZN(_01070_)
  );
  INV_X1 _21719_ (
    .A(_01070_),
    .ZN(_01071_)
  );
  AND2_X1 _21720_ (
    .A1(_05138_),
    .A2(_05983_),
    .ZN(_01072_)
  );
  INV_X1 _21721_ (
    .A(_01072_),
    .ZN(_01073_)
  );
  AND2_X1 _21722_ (
    .A1(_06201_),
    .A2(_01073_),
    .ZN(_01074_)
  );
  AND2_X1 _21723_ (
    .A1(_01071_),
    .A2(_01074_),
    .ZN(_01075_)
  );
  INV_X1 _21724_ (
    .A(_01075_),
    .ZN(_01077_)
  );
  AND2_X1 _21725_ (
    .A1(remainder[7]),
    .A2(_00919_),
    .ZN(_01078_)
  );
  INV_X1 _21726_ (
    .A(_01078_),
    .ZN(_01079_)
  );
  AND2_X1 _21727_ (
    .A1(io_req_bits_in1[7]),
    .A2(_06190_),
    .ZN(_01080_)
  );
  INV_X1 _21728_ (
    .A(_01080_),
    .ZN(_01081_)
  );
  AND2_X1 _21729_ (
    .A1(_01079_),
    .A2(_01081_),
    .ZN(_01082_)
  );
  AND2_X1 _21730_ (
    .A1(_01077_),
    .A2(_01082_),
    .ZN(_01083_)
  );
  INV_X1 _21731_ (
    .A(_01083_),
    .ZN(_00094_)
  );
  AND2_X1 _21732_ (
    .A1(remainder[16]),
    .A2(_06103_),
    .ZN(_01084_)
  );
  INV_X1 _21733_ (
    .A(_01084_),
    .ZN(_01085_)
  );
  AND2_X1 _21734_ (
    .A1(_05994_),
    .A2(_01085_),
    .ZN(_01087_)
  );
  MUX2_X1 _21735_ (
    .A(remainder[8]),
    .B(remainder[41]),
    .S(resHi),
    .Z(io_resp_bits_data[8])
  );
  INV_X1 _21736_ (
    .A(io_resp_bits_data[8]),
    .ZN(_01088_)
  );
  AND2_X1 _21737_ (
    .A1(_01066_),
    .A2(io_resp_bits_data[8]),
    .ZN(_01089_)
  );
  INV_X1 _21738_ (
    .A(_01089_),
    .ZN(_01090_)
  );
  AND2_X1 _21739_ (
    .A1(_01064_),
    .A2(_01088_),
    .ZN(_01091_)
  );
  INV_X1 _21740_ (
    .A(_01091_),
    .ZN(_01092_)
  );
  AND2_X1 _21741_ (
    .A1(_00898_),
    .A2(_01092_),
    .ZN(_01093_)
  );
  AND2_X1 _21742_ (
    .A1(_01090_),
    .A2(_01093_),
    .ZN(_01094_)
  );
  INV_X1 _21743_ (
    .A(_01094_),
    .ZN(_01095_)
  );
  AND2_X1 _21744_ (
    .A1(_01087_),
    .A2(_01095_),
    .ZN(_01096_)
  );
  INV_X1 _21745_ (
    .A(_01096_),
    .ZN(_01097_)
  );
  AND2_X1 _21746_ (
    .A1(_05149_),
    .A2(_05983_),
    .ZN(_01098_)
  );
  INV_X1 _21747_ (
    .A(_01098_),
    .ZN(_01099_)
  );
  AND2_X1 _21748_ (
    .A1(_06201_),
    .A2(_01099_),
    .ZN(_01100_)
  );
  AND2_X1 _21749_ (
    .A1(_01097_),
    .A2(_01100_),
    .ZN(_01101_)
  );
  INV_X1 _21750_ (
    .A(_01101_),
    .ZN(_01102_)
  );
  AND2_X1 _21751_ (
    .A1(remainder[8]),
    .A2(_00919_),
    .ZN(_01103_)
  );
  INV_X1 _21752_ (
    .A(_01103_),
    .ZN(_01104_)
  );
  AND2_X1 _21753_ (
    .A1(io_req_bits_in1[8]),
    .A2(_06190_),
    .ZN(_01105_)
  );
  INV_X1 _21754_ (
    .A(_01105_),
    .ZN(_01107_)
  );
  AND2_X1 _21755_ (
    .A1(_01104_),
    .A2(_01107_),
    .ZN(_01108_)
  );
  AND2_X1 _21756_ (
    .A1(_01102_),
    .A2(_01108_),
    .ZN(_01109_)
  );
  INV_X1 _21757_ (
    .A(_01109_),
    .ZN(_00095_)
  );
  AND2_X1 _21758_ (
    .A1(remainder[17]),
    .A2(_06103_),
    .ZN(_01110_)
  );
  INV_X1 _21759_ (
    .A(_01110_),
    .ZN(_01111_)
  );
  AND2_X1 _21760_ (
    .A1(_05994_),
    .A2(_01111_),
    .ZN(_01112_)
  );
  MUX2_X1 _21761_ (
    .A(remainder[9]),
    .B(remainder[42]),
    .S(resHi),
    .Z(io_resp_bits_data[9])
  );
  INV_X1 _21762_ (
    .A(io_resp_bits_data[9]),
    .ZN(_01113_)
  );
  AND2_X1 _21763_ (
    .A1(_01092_),
    .A2(io_resp_bits_data[9]),
    .ZN(_01114_)
  );
  INV_X1 _21764_ (
    .A(_01114_),
    .ZN(_01116_)
  );
  AND2_X1 _21765_ (
    .A1(_01091_),
    .A2(_01113_),
    .ZN(_01117_)
  );
  INV_X1 _21766_ (
    .A(_01117_),
    .ZN(_01118_)
  );
  AND2_X1 _21767_ (
    .A1(_00898_),
    .A2(_01118_),
    .ZN(_01119_)
  );
  AND2_X1 _21768_ (
    .A1(_01116_),
    .A2(_01119_),
    .ZN(_01120_)
  );
  INV_X1 _21769_ (
    .A(_01120_),
    .ZN(_01121_)
  );
  AND2_X1 _21770_ (
    .A1(_01112_),
    .A2(_01121_),
    .ZN(_01122_)
  );
  INV_X1 _21771_ (
    .A(_01122_),
    .ZN(_01123_)
  );
  AND2_X1 _21772_ (
    .A1(_05160_),
    .A2(_05983_),
    .ZN(_01124_)
  );
  INV_X1 _21773_ (
    .A(_01124_),
    .ZN(_01125_)
  );
  AND2_X1 _21774_ (
    .A1(_06201_),
    .A2(_01125_),
    .ZN(_01127_)
  );
  AND2_X1 _21775_ (
    .A1(_01123_),
    .A2(_01127_),
    .ZN(_01128_)
  );
  INV_X1 _21776_ (
    .A(_01128_),
    .ZN(_01129_)
  );
  AND2_X1 _21777_ (
    .A1(remainder[9]),
    .A2(_00919_),
    .ZN(_01130_)
  );
  INV_X1 _21778_ (
    .A(_01130_),
    .ZN(_01131_)
  );
  AND2_X1 _21779_ (
    .A1(io_req_bits_in1[9]),
    .A2(_06190_),
    .ZN(_01132_)
  );
  INV_X1 _21780_ (
    .A(_01132_),
    .ZN(_01133_)
  );
  AND2_X1 _21781_ (
    .A1(_01131_),
    .A2(_01133_),
    .ZN(_01134_)
  );
  AND2_X1 _21782_ (
    .A1(_01129_),
    .A2(_01134_),
    .ZN(_01135_)
  );
  INV_X1 _21783_ (
    .A(_01135_),
    .ZN(_00096_)
  );
  AND2_X1 _21784_ (
    .A1(remainder[18]),
    .A2(_06103_),
    .ZN(_01137_)
  );
  INV_X1 _21785_ (
    .A(_01137_),
    .ZN(_01138_)
  );
  AND2_X1 _21786_ (
    .A1(_05994_),
    .A2(_01138_),
    .ZN(_01139_)
  );
  MUX2_X1 _21787_ (
    .A(remainder[10]),
    .B(remainder[43]),
    .S(resHi),
    .Z(io_resp_bits_data[10])
  );
  INV_X1 _21788_ (
    .A(io_resp_bits_data[10]),
    .ZN(_01140_)
  );
  AND2_X1 _21789_ (
    .A1(_01118_),
    .A2(io_resp_bits_data[10]),
    .ZN(_01141_)
  );
  INV_X1 _21790_ (
    .A(_01141_),
    .ZN(_01142_)
  );
  AND2_X1 _21791_ (
    .A1(_01117_),
    .A2(_01140_),
    .ZN(_01143_)
  );
  INV_X1 _21792_ (
    .A(_01143_),
    .ZN(_01144_)
  );
  AND2_X1 _21793_ (
    .A1(_00898_),
    .A2(_01144_),
    .ZN(_01145_)
  );
  AND2_X1 _21794_ (
    .A1(_01142_),
    .A2(_01145_),
    .ZN(_01147_)
  );
  INV_X1 _21795_ (
    .A(_01147_),
    .ZN(_01148_)
  );
  AND2_X1 _21796_ (
    .A1(_01139_),
    .A2(_01148_),
    .ZN(_01149_)
  );
  INV_X1 _21797_ (
    .A(_01149_),
    .ZN(_01150_)
  );
  AND2_X1 _21798_ (
    .A1(_05171_),
    .A2(_05983_),
    .ZN(_01151_)
  );
  INV_X1 _21799_ (
    .A(_01151_),
    .ZN(_01152_)
  );
  AND2_X1 _21800_ (
    .A1(_06201_),
    .A2(_01152_),
    .ZN(_01153_)
  );
  AND2_X1 _21801_ (
    .A1(_01150_),
    .A2(_01153_),
    .ZN(_01154_)
  );
  INV_X1 _21802_ (
    .A(_01154_),
    .ZN(_01155_)
  );
  AND2_X1 _21803_ (
    .A1(remainder[10]),
    .A2(_00919_),
    .ZN(_01156_)
  );
  INV_X1 _21804_ (
    .A(_01156_),
    .ZN(_01158_)
  );
  AND2_X1 _21805_ (
    .A1(io_req_bits_in1[10]),
    .A2(_06190_),
    .ZN(_01159_)
  );
  INV_X1 _21806_ (
    .A(_01159_),
    .ZN(_01160_)
  );
  AND2_X1 _21807_ (
    .A1(_01158_),
    .A2(_01160_),
    .ZN(_01161_)
  );
  AND2_X1 _21808_ (
    .A1(_01155_),
    .A2(_01161_),
    .ZN(_01162_)
  );
  INV_X1 _21809_ (
    .A(_01162_),
    .ZN(_00097_)
  );
  AND2_X1 _21810_ (
    .A1(remainder[19]),
    .A2(_06103_),
    .ZN(_01163_)
  );
  INV_X1 _21811_ (
    .A(_01163_),
    .ZN(_01164_)
  );
  AND2_X1 _21812_ (
    .A1(_05994_),
    .A2(_01164_),
    .ZN(_01165_)
  );
  MUX2_X1 _21813_ (
    .A(remainder[11]),
    .B(remainder[44]),
    .S(resHi),
    .Z(io_resp_bits_data[11])
  );
  INV_X1 _21814_ (
    .A(io_resp_bits_data[11]),
    .ZN(_01167_)
  );
  AND2_X1 _21815_ (
    .A1(_01144_),
    .A2(io_resp_bits_data[11]),
    .ZN(_01168_)
  );
  INV_X1 _21816_ (
    .A(_01168_),
    .ZN(_01169_)
  );
  AND2_X1 _21817_ (
    .A1(_01143_),
    .A2(_01167_),
    .ZN(_01170_)
  );
  INV_X1 _21818_ (
    .A(_01170_),
    .ZN(_01171_)
  );
  AND2_X1 _21819_ (
    .A1(_00898_),
    .A2(_01171_),
    .ZN(_01172_)
  );
  AND2_X1 _21820_ (
    .A1(_01169_),
    .A2(_01172_),
    .ZN(_01173_)
  );
  INV_X1 _21821_ (
    .A(_01173_),
    .ZN(_01174_)
  );
  AND2_X1 _21822_ (
    .A1(_01165_),
    .A2(_01174_),
    .ZN(_01175_)
  );
  INV_X1 _21823_ (
    .A(_01175_),
    .ZN(_01176_)
  );
  AND2_X1 _21824_ (
    .A1(_05182_),
    .A2(_05983_),
    .ZN(_01178_)
  );
  INV_X1 _21825_ (
    .A(_01178_),
    .ZN(_01179_)
  );
  AND2_X1 _21826_ (
    .A1(_06201_),
    .A2(_01179_),
    .ZN(_01180_)
  );
  AND2_X1 _21827_ (
    .A1(_01176_),
    .A2(_01180_),
    .ZN(_01181_)
  );
  INV_X1 _21828_ (
    .A(_01181_),
    .ZN(_01182_)
  );
  AND2_X1 _21829_ (
    .A1(remainder[11]),
    .A2(_00919_),
    .ZN(_01183_)
  );
  INV_X1 _21830_ (
    .A(_01183_),
    .ZN(_01184_)
  );
  AND2_X1 _21831_ (
    .A1(io_req_bits_in1[11]),
    .A2(_06190_),
    .ZN(_01185_)
  );
  INV_X1 _21832_ (
    .A(_01185_),
    .ZN(_01186_)
  );
  AND2_X1 _21833_ (
    .A1(_01184_),
    .A2(_01186_),
    .ZN(_01187_)
  );
  AND2_X1 _21834_ (
    .A1(_01182_),
    .A2(_01187_),
    .ZN(_01189_)
  );
  INV_X1 _21835_ (
    .A(_01189_),
    .ZN(_00098_)
  );
  AND2_X1 _21836_ (
    .A1(remainder[20]),
    .A2(_06103_),
    .ZN(_01190_)
  );
  INV_X1 _21837_ (
    .A(_01190_),
    .ZN(_01191_)
  );
  AND2_X1 _21838_ (
    .A1(_05994_),
    .A2(_01191_),
    .ZN(_01192_)
  );
  MUX2_X1 _21839_ (
    .A(remainder[12]),
    .B(remainder[45]),
    .S(resHi),
    .Z(io_resp_bits_data[12])
  );
  INV_X1 _21840_ (
    .A(io_resp_bits_data[12]),
    .ZN(_01193_)
  );
  AND2_X1 _21841_ (
    .A1(_01171_),
    .A2(io_resp_bits_data[12]),
    .ZN(_01194_)
  );
  INV_X1 _21842_ (
    .A(_01194_),
    .ZN(_01195_)
  );
  AND2_X1 _21843_ (
    .A1(_01170_),
    .A2(_01193_),
    .ZN(_01196_)
  );
  INV_X1 _21844_ (
    .A(_01196_),
    .ZN(_01198_)
  );
  AND2_X1 _21845_ (
    .A1(_00898_),
    .A2(_01198_),
    .ZN(_01199_)
  );
  AND2_X1 _21846_ (
    .A1(_01195_),
    .A2(_01199_),
    .ZN(_01200_)
  );
  INV_X1 _21847_ (
    .A(_01200_),
    .ZN(_01201_)
  );
  AND2_X1 _21848_ (
    .A1(_01192_),
    .A2(_01201_),
    .ZN(_01202_)
  );
  INV_X1 _21849_ (
    .A(_01202_),
    .ZN(_01203_)
  );
  AND2_X1 _21850_ (
    .A1(_05193_),
    .A2(_05983_),
    .ZN(_01204_)
  );
  INV_X1 _21851_ (
    .A(_01204_),
    .ZN(_01205_)
  );
  AND2_X1 _21852_ (
    .A1(_06201_),
    .A2(_01205_),
    .ZN(_01206_)
  );
  AND2_X1 _21853_ (
    .A1(_01203_),
    .A2(_01206_),
    .ZN(_01207_)
  );
  INV_X1 _21854_ (
    .A(_01207_),
    .ZN(_01209_)
  );
  AND2_X1 _21855_ (
    .A1(remainder[12]),
    .A2(_00919_),
    .ZN(_01210_)
  );
  INV_X1 _21856_ (
    .A(_01210_),
    .ZN(_01211_)
  );
  AND2_X1 _21857_ (
    .A1(io_req_bits_in1[12]),
    .A2(_06190_),
    .ZN(_01212_)
  );
  INV_X1 _21858_ (
    .A(_01212_),
    .ZN(_01213_)
  );
  AND2_X1 _21859_ (
    .A1(_01211_),
    .A2(_01213_),
    .ZN(_01214_)
  );
  AND2_X1 _21860_ (
    .A1(_01209_),
    .A2(_01214_),
    .ZN(_01215_)
  );
  INV_X1 _21861_ (
    .A(_01215_),
    .ZN(_00099_)
  );
  AND2_X1 _21862_ (
    .A1(remainder[21]),
    .A2(_06103_),
    .ZN(_01216_)
  );
  INV_X1 _21863_ (
    .A(_01216_),
    .ZN(_01217_)
  );
  AND2_X1 _21864_ (
    .A1(_05994_),
    .A2(_01217_),
    .ZN(_01219_)
  );
  MUX2_X1 _21865_ (
    .A(remainder[13]),
    .B(remainder[46]),
    .S(resHi),
    .Z(io_resp_bits_data[13])
  );
  INV_X1 _21866_ (
    .A(io_resp_bits_data[13]),
    .ZN(_01220_)
  );
  AND2_X1 _21867_ (
    .A1(_01198_),
    .A2(io_resp_bits_data[13]),
    .ZN(_01221_)
  );
  INV_X1 _21868_ (
    .A(_01221_),
    .ZN(_01222_)
  );
  AND2_X1 _21869_ (
    .A1(_01196_),
    .A2(_01220_),
    .ZN(_01223_)
  );
  INV_X1 _21870_ (
    .A(_01223_),
    .ZN(_01224_)
  );
  AND2_X1 _21871_ (
    .A1(_00898_),
    .A2(_01224_),
    .ZN(_01225_)
  );
  AND2_X1 _21872_ (
    .A1(_01222_),
    .A2(_01225_),
    .ZN(_01226_)
  );
  INV_X1 _21873_ (
    .A(_01226_),
    .ZN(_01227_)
  );
  AND2_X1 _21874_ (
    .A1(_01219_),
    .A2(_01227_),
    .ZN(_01228_)
  );
  INV_X1 _21875_ (
    .A(_01228_),
    .ZN(_01229_)
  );
  AND2_X1 _21876_ (
    .A1(_05204_),
    .A2(_05983_),
    .ZN(_01230_)
  );
  INV_X1 _21877_ (
    .A(_01230_),
    .ZN(_01231_)
  );
  AND2_X1 _21878_ (
    .A1(_06201_),
    .A2(_01231_),
    .ZN(_01232_)
  );
  AND2_X1 _21879_ (
    .A1(_01229_),
    .A2(_01232_),
    .ZN(_01233_)
  );
  INV_X1 _21880_ (
    .A(_01233_),
    .ZN(_01234_)
  );
  AND2_X1 _21881_ (
    .A1(remainder[13]),
    .A2(_00919_),
    .ZN(_01235_)
  );
  INV_X1 _21882_ (
    .A(_01235_),
    .ZN(_01236_)
  );
  AND2_X1 _21883_ (
    .A1(io_req_bits_in1[13]),
    .A2(_06190_),
    .ZN(_01237_)
  );
  INV_X1 _21884_ (
    .A(_01237_),
    .ZN(_01239_)
  );
  AND2_X1 _21885_ (
    .A1(_01236_),
    .A2(_01239_),
    .ZN(_01240_)
  );
  AND2_X1 _21886_ (
    .A1(_01234_),
    .A2(_01240_),
    .ZN(_01241_)
  );
  INV_X1 _21887_ (
    .A(_01241_),
    .ZN(_00100_)
  );
  AND2_X1 _21888_ (
    .A1(remainder[22]),
    .A2(_06103_),
    .ZN(_01242_)
  );
  INV_X1 _21889_ (
    .A(_01242_),
    .ZN(_01243_)
  );
  AND2_X1 _21890_ (
    .A1(_05994_),
    .A2(_01243_),
    .ZN(_01244_)
  );
  MUX2_X1 _21891_ (
    .A(remainder[14]),
    .B(remainder[47]),
    .S(resHi),
    .Z(io_resp_bits_data[14])
  );
  INV_X1 _21892_ (
    .A(io_resp_bits_data[14]),
    .ZN(_01245_)
  );
  AND2_X1 _21893_ (
    .A1(_01224_),
    .A2(io_resp_bits_data[14]),
    .ZN(_01246_)
  );
  INV_X1 _21894_ (
    .A(_01246_),
    .ZN(_01248_)
  );
  AND2_X1 _21895_ (
    .A1(_01223_),
    .A2(_01245_),
    .ZN(_01249_)
  );
  INV_X1 _21896_ (
    .A(_01249_),
    .ZN(_01250_)
  );
  AND2_X1 _21897_ (
    .A1(_00898_),
    .A2(_01250_),
    .ZN(_01251_)
  );
  AND2_X1 _21898_ (
    .A1(_01248_),
    .A2(_01251_),
    .ZN(_01252_)
  );
  INV_X1 _21899_ (
    .A(_01252_),
    .ZN(_01253_)
  );
  AND2_X1 _21900_ (
    .A1(_01244_),
    .A2(_01253_),
    .ZN(_01254_)
  );
  INV_X1 _21901_ (
    .A(_01254_),
    .ZN(_01255_)
  );
  AND2_X1 _21902_ (
    .A1(_05215_),
    .A2(_05983_),
    .ZN(_01256_)
  );
  INV_X1 _21903_ (
    .A(_01256_),
    .ZN(_01257_)
  );
  AND2_X1 _21904_ (
    .A1(_06201_),
    .A2(_01257_),
    .ZN(_01259_)
  );
  AND2_X1 _21905_ (
    .A1(_01255_),
    .A2(_01259_),
    .ZN(_01260_)
  );
  INV_X1 _21906_ (
    .A(_01260_),
    .ZN(_01261_)
  );
  AND2_X1 _21907_ (
    .A1(remainder[14]),
    .A2(_00919_),
    .ZN(_01262_)
  );
  INV_X1 _21908_ (
    .A(_01262_),
    .ZN(_01263_)
  );
  AND2_X1 _21909_ (
    .A1(io_req_bits_in1[14]),
    .A2(_06190_),
    .ZN(_01264_)
  );
  INV_X1 _21910_ (
    .A(_01264_),
    .ZN(_01265_)
  );
  AND2_X1 _21911_ (
    .A1(_01263_),
    .A2(_01265_),
    .ZN(_01266_)
  );
  AND2_X1 _21912_ (
    .A1(_01261_),
    .A2(_01266_),
    .ZN(_01267_)
  );
  INV_X1 _21913_ (
    .A(_01267_),
    .ZN(_00101_)
  );
  AND2_X1 _21914_ (
    .A1(remainder[23]),
    .A2(_06103_),
    .ZN(_01269_)
  );
  INV_X1 _21915_ (
    .A(_01269_),
    .ZN(_01270_)
  );
  AND2_X1 _21916_ (
    .A1(_05994_),
    .A2(_01270_),
    .ZN(_01271_)
  );
  MUX2_X1 _21917_ (
    .A(remainder[15]),
    .B(remainder[48]),
    .S(resHi),
    .Z(io_resp_bits_data[15])
  );
  INV_X1 _21918_ (
    .A(io_resp_bits_data[15]),
    .ZN(_01272_)
  );
  AND2_X1 _21919_ (
    .A1(_01250_),
    .A2(io_resp_bits_data[15]),
    .ZN(_01273_)
  );
  INV_X1 _21920_ (
    .A(_01273_),
    .ZN(_01274_)
  );
  AND2_X1 _21921_ (
    .A1(_01249_),
    .A2(_01272_),
    .ZN(_01275_)
  );
  INV_X1 _21922_ (
    .A(_01275_),
    .ZN(_01276_)
  );
  AND2_X1 _21923_ (
    .A1(_00898_),
    .A2(_01276_),
    .ZN(_01277_)
  );
  AND2_X1 _21924_ (
    .A1(_01274_),
    .A2(_01277_),
    .ZN(_01279_)
  );
  INV_X1 _21925_ (
    .A(_01279_),
    .ZN(_01280_)
  );
  AND2_X1 _21926_ (
    .A1(_01271_),
    .A2(_01280_),
    .ZN(_01281_)
  );
  INV_X1 _21927_ (
    .A(_01281_),
    .ZN(_01282_)
  );
  AND2_X1 _21928_ (
    .A1(_05226_),
    .A2(_05983_),
    .ZN(_01283_)
  );
  INV_X1 _21929_ (
    .A(_01283_),
    .ZN(_01284_)
  );
  AND2_X1 _21930_ (
    .A1(_06201_),
    .A2(_01284_),
    .ZN(_01285_)
  );
  AND2_X1 _21931_ (
    .A1(_01282_),
    .A2(_01285_),
    .ZN(_01286_)
  );
  INV_X1 _21932_ (
    .A(_01286_),
    .ZN(_01287_)
  );
  AND2_X1 _21933_ (
    .A1(remainder[15]),
    .A2(_00919_),
    .ZN(_01288_)
  );
  INV_X1 _21934_ (
    .A(_01288_),
    .ZN(_01290_)
  );
  AND2_X1 _21935_ (
    .A1(io_req_bits_in1[15]),
    .A2(_06190_),
    .ZN(_01291_)
  );
  INV_X1 _21936_ (
    .A(_01291_),
    .ZN(_01292_)
  );
  AND2_X1 _21937_ (
    .A1(_01290_),
    .A2(_01292_),
    .ZN(_01293_)
  );
  AND2_X1 _21938_ (
    .A1(_01287_),
    .A2(_01293_),
    .ZN(_01294_)
  );
  INV_X1 _21939_ (
    .A(_01294_),
    .ZN(_00102_)
  );
  AND2_X1 _21940_ (
    .A1(remainder[24]),
    .A2(_06103_),
    .ZN(_01295_)
  );
  INV_X1 _21941_ (
    .A(_01295_),
    .ZN(_01296_)
  );
  AND2_X1 _21942_ (
    .A1(_05994_),
    .A2(_01296_),
    .ZN(_01297_)
  );
  MUX2_X1 _21943_ (
    .A(remainder[16]),
    .B(remainder[49]),
    .S(resHi),
    .Z(io_resp_bits_data[16])
  );
  INV_X1 _21944_ (
    .A(io_resp_bits_data[16]),
    .ZN(_01299_)
  );
  AND2_X1 _21945_ (
    .A1(_01276_),
    .A2(io_resp_bits_data[16]),
    .ZN(_01300_)
  );
  INV_X1 _21946_ (
    .A(_01300_),
    .ZN(_01301_)
  );
  AND2_X1 _21947_ (
    .A1(_01275_),
    .A2(_01299_),
    .ZN(_01302_)
  );
  INV_X1 _21948_ (
    .A(_01302_),
    .ZN(_01303_)
  );
  AND2_X1 _21949_ (
    .A1(_00898_),
    .A2(_01303_),
    .ZN(_01304_)
  );
  AND2_X1 _21950_ (
    .A1(_01301_),
    .A2(_01304_),
    .ZN(_01305_)
  );
  INV_X1 _21951_ (
    .A(_01305_),
    .ZN(_01306_)
  );
  AND2_X1 _21952_ (
    .A1(_01297_),
    .A2(_01306_),
    .ZN(_01307_)
  );
  INV_X1 _21953_ (
    .A(_01307_),
    .ZN(_01308_)
  );
  AND2_X1 _21954_ (
    .A1(_05237_),
    .A2(_05983_),
    .ZN(_01310_)
  );
  INV_X1 _21955_ (
    .A(_01310_),
    .ZN(_01311_)
  );
  AND2_X1 _21956_ (
    .A1(_06201_),
    .A2(_01311_),
    .ZN(_01312_)
  );
  AND2_X1 _21957_ (
    .A1(_01308_),
    .A2(_01312_),
    .ZN(_01313_)
  );
  INV_X1 _21958_ (
    .A(_01313_),
    .ZN(_01314_)
  );
  AND2_X1 _21959_ (
    .A1(remainder[16]),
    .A2(_00919_),
    .ZN(_01315_)
  );
  INV_X1 _21960_ (
    .A(_01315_),
    .ZN(_01316_)
  );
  AND2_X1 _21961_ (
    .A1(io_req_bits_in1[16]),
    .A2(_06190_),
    .ZN(_01317_)
  );
  INV_X1 _21962_ (
    .A(_01317_),
    .ZN(_01318_)
  );
  AND2_X1 _21963_ (
    .A1(_01316_),
    .A2(_01318_),
    .ZN(_01319_)
  );
  AND2_X1 _21964_ (
    .A1(_01314_),
    .A2(_01319_),
    .ZN(_01321_)
  );
  INV_X1 _21965_ (
    .A(_01321_),
    .ZN(_00103_)
  );
  AND2_X1 _21966_ (
    .A1(remainder[25]),
    .A2(_06103_),
    .ZN(_01322_)
  );
  INV_X1 _21967_ (
    .A(_01322_),
    .ZN(_01323_)
  );
  AND2_X1 _21968_ (
    .A1(_05994_),
    .A2(_01323_),
    .ZN(_01324_)
  );
  MUX2_X1 _21969_ (
    .A(remainder[17]),
    .B(remainder[50]),
    .S(resHi),
    .Z(io_resp_bits_data[17])
  );
  INV_X1 _21970_ (
    .A(io_resp_bits_data[17]),
    .ZN(_01325_)
  );
  AND2_X1 _21971_ (
    .A1(_01303_),
    .A2(io_resp_bits_data[17]),
    .ZN(_01326_)
  );
  INV_X1 _21972_ (
    .A(_01326_),
    .ZN(_01327_)
  );
  AND2_X1 _21973_ (
    .A1(_01302_),
    .A2(_01325_),
    .ZN(_01328_)
  );
  INV_X1 _21974_ (
    .A(_01328_),
    .ZN(_01330_)
  );
  AND2_X1 _21975_ (
    .A1(_00898_),
    .A2(_01330_),
    .ZN(_01331_)
  );
  AND2_X1 _21976_ (
    .A1(_01327_),
    .A2(_01331_),
    .ZN(_01332_)
  );
  INV_X1 _21977_ (
    .A(_01332_),
    .ZN(_01333_)
  );
  AND2_X1 _21978_ (
    .A1(_01324_),
    .A2(_01333_),
    .ZN(_01334_)
  );
  INV_X1 _21979_ (
    .A(_01334_),
    .ZN(_01335_)
  );
  AND2_X1 _21980_ (
    .A1(_05248_),
    .A2(_05983_),
    .ZN(_01336_)
  );
  INV_X1 _21981_ (
    .A(_01336_),
    .ZN(_01337_)
  );
  AND2_X1 _21982_ (
    .A1(_06201_),
    .A2(_01337_),
    .ZN(_01338_)
  );
  AND2_X1 _21983_ (
    .A1(_01335_),
    .A2(_01338_),
    .ZN(_01339_)
  );
  INV_X1 _21984_ (
    .A(_01339_),
    .ZN(_01341_)
  );
  AND2_X1 _21985_ (
    .A1(remainder[17]),
    .A2(_00919_),
    .ZN(_01342_)
  );
  INV_X1 _21986_ (
    .A(_01342_),
    .ZN(_01343_)
  );
  AND2_X1 _21987_ (
    .A1(io_req_bits_in1[17]),
    .A2(_06190_),
    .ZN(_01344_)
  );
  INV_X1 _21988_ (
    .A(_01344_),
    .ZN(_01345_)
  );
  AND2_X1 _21989_ (
    .A1(_01343_),
    .A2(_01345_),
    .ZN(_01346_)
  );
  AND2_X1 _21990_ (
    .A1(_01341_),
    .A2(_01346_),
    .ZN(_01347_)
  );
  INV_X1 _21991_ (
    .A(_01347_),
    .ZN(_00104_)
  );
  AND2_X1 _21992_ (
    .A1(remainder[26]),
    .A2(_06103_),
    .ZN(_01348_)
  );
  INV_X1 _21993_ (
    .A(_01348_),
    .ZN(_01349_)
  );
  AND2_X1 _21994_ (
    .A1(_05994_),
    .A2(_01349_),
    .ZN(_01351_)
  );
  MUX2_X1 _21995_ (
    .A(remainder[18]),
    .B(remainder[51]),
    .S(resHi),
    .Z(io_resp_bits_data[18])
  );
  INV_X1 _21996_ (
    .A(io_resp_bits_data[18]),
    .ZN(_01352_)
  );
  AND2_X1 _21997_ (
    .A1(_01330_),
    .A2(io_resp_bits_data[18]),
    .ZN(_01353_)
  );
  INV_X1 _21998_ (
    .A(_01353_),
    .ZN(_01354_)
  );
  AND2_X1 _21999_ (
    .A1(_01328_),
    .A2(_01352_),
    .ZN(_01355_)
  );
  INV_X1 _22000_ (
    .A(_01355_),
    .ZN(_01356_)
  );
  AND2_X1 _22001_ (
    .A1(_00898_),
    .A2(_01356_),
    .ZN(_01357_)
  );
  AND2_X1 _22002_ (
    .A1(_01354_),
    .A2(_01357_),
    .ZN(_01358_)
  );
  INV_X1 _22003_ (
    .A(_01358_),
    .ZN(_01359_)
  );
  AND2_X1 _22004_ (
    .A1(_01351_),
    .A2(_01359_),
    .ZN(_01361_)
  );
  INV_X1 _22005_ (
    .A(_01361_),
    .ZN(_01362_)
  );
  AND2_X1 _22006_ (
    .A1(_05259_),
    .A2(_05983_),
    .ZN(_01363_)
  );
  INV_X1 _22007_ (
    .A(_01363_),
    .ZN(_01364_)
  );
  AND2_X1 _22008_ (
    .A1(_06201_),
    .A2(_01364_),
    .ZN(_01365_)
  );
  AND2_X1 _22009_ (
    .A1(_01362_),
    .A2(_01365_),
    .ZN(_01366_)
  );
  INV_X1 _22010_ (
    .A(_01366_),
    .ZN(_01367_)
  );
  AND2_X1 _22011_ (
    .A1(remainder[18]),
    .A2(_00919_),
    .ZN(_01368_)
  );
  INV_X1 _22012_ (
    .A(_01368_),
    .ZN(_01369_)
  );
  AND2_X1 _22013_ (
    .A1(io_req_bits_in1[18]),
    .A2(_06190_),
    .ZN(_01370_)
  );
  INV_X1 _22014_ (
    .A(_01370_),
    .ZN(_01372_)
  );
  AND2_X1 _22015_ (
    .A1(_01369_),
    .A2(_01372_),
    .ZN(_01373_)
  );
  AND2_X1 _22016_ (
    .A1(_01367_),
    .A2(_01373_),
    .ZN(_01374_)
  );
  INV_X1 _22017_ (
    .A(_01374_),
    .ZN(_00105_)
  );
  AND2_X1 _22018_ (
    .A1(remainder[27]),
    .A2(_06103_),
    .ZN(_01375_)
  );
  INV_X1 _22019_ (
    .A(_01375_),
    .ZN(_01376_)
  );
  AND2_X1 _22020_ (
    .A1(_05994_),
    .A2(_01376_),
    .ZN(_01377_)
  );
  MUX2_X1 _22021_ (
    .A(remainder[19]),
    .B(remainder[52]),
    .S(resHi),
    .Z(io_resp_bits_data[19])
  );
  INV_X1 _22022_ (
    .A(io_resp_bits_data[19]),
    .ZN(_01378_)
  );
  AND2_X1 _22023_ (
    .A1(_01356_),
    .A2(io_resp_bits_data[19]),
    .ZN(_01379_)
  );
  INV_X1 _22024_ (
    .A(_01379_),
    .ZN(_01381_)
  );
  AND2_X1 _22025_ (
    .A1(_01355_),
    .A2(_01378_),
    .ZN(_01382_)
  );
  INV_X1 _22026_ (
    .A(_01382_),
    .ZN(_01383_)
  );
  AND2_X1 _22027_ (
    .A1(_00898_),
    .A2(_01383_),
    .ZN(_01384_)
  );
  AND2_X1 _22028_ (
    .A1(_01381_),
    .A2(_01384_),
    .ZN(_01385_)
  );
  INV_X1 _22029_ (
    .A(_01385_),
    .ZN(_01386_)
  );
  AND2_X1 _22030_ (
    .A1(_01377_),
    .A2(_01386_),
    .ZN(_01387_)
  );
  INV_X1 _22031_ (
    .A(_01387_),
    .ZN(_01388_)
  );
  AND2_X1 _22032_ (
    .A1(_05270_),
    .A2(_05983_),
    .ZN(_01389_)
  );
  INV_X1 _22033_ (
    .A(_01389_),
    .ZN(_01390_)
  );
  AND2_X1 _22034_ (
    .A1(_06201_),
    .A2(_01390_),
    .ZN(_01392_)
  );
  AND2_X1 _22035_ (
    .A1(_01388_),
    .A2(_01392_),
    .ZN(_01393_)
  );
  INV_X1 _22036_ (
    .A(_01393_),
    .ZN(_01394_)
  );
  AND2_X1 _22037_ (
    .A1(remainder[19]),
    .A2(_00919_),
    .ZN(_01395_)
  );
  INV_X1 _22038_ (
    .A(_01395_),
    .ZN(_01396_)
  );
  AND2_X1 _22039_ (
    .A1(io_req_bits_in1[19]),
    .A2(_06190_),
    .ZN(_01397_)
  );
  INV_X1 _22040_ (
    .A(_01397_),
    .ZN(_01398_)
  );
  AND2_X1 _22041_ (
    .A1(_01396_),
    .A2(_01398_),
    .ZN(_01399_)
  );
  AND2_X1 _22042_ (
    .A1(_01394_),
    .A2(_01399_),
    .ZN(_01400_)
  );
  INV_X1 _22043_ (
    .A(_01400_),
    .ZN(_00106_)
  );
  AND2_X1 _22044_ (
    .A1(remainder[28]),
    .A2(_06103_),
    .ZN(_01401_)
  );
  INV_X1 _22045_ (
    .A(_01401_),
    .ZN(_01402_)
  );
  AND2_X1 _22046_ (
    .A1(_05994_),
    .A2(_01402_),
    .ZN(_01403_)
  );
  MUX2_X1 _22047_ (
    .A(remainder[20]),
    .B(remainder[53]),
    .S(resHi),
    .Z(io_resp_bits_data[20])
  );
  INV_X1 _22048_ (
    .A(io_resp_bits_data[20]),
    .ZN(_01404_)
  );
  AND2_X1 _22049_ (
    .A1(_01383_),
    .A2(io_resp_bits_data[20]),
    .ZN(_01405_)
  );
  INV_X1 _22050_ (
    .A(_01405_),
    .ZN(_01406_)
  );
  AND2_X1 _22051_ (
    .A1(_01382_),
    .A2(_01404_),
    .ZN(_01407_)
  );
  INV_X1 _22052_ (
    .A(_01407_),
    .ZN(_01408_)
  );
  AND2_X1 _22053_ (
    .A1(_00898_),
    .A2(_01408_),
    .ZN(_01409_)
  );
  AND2_X1 _22054_ (
    .A1(_01406_),
    .A2(_01409_),
    .ZN(_01411_)
  );
  INV_X1 _22055_ (
    .A(_01411_),
    .ZN(_01412_)
  );
  AND2_X1 _22056_ (
    .A1(_01403_),
    .A2(_01412_),
    .ZN(_01413_)
  );
  INV_X1 _22057_ (
    .A(_01413_),
    .ZN(_01414_)
  );
  AND2_X1 _22058_ (
    .A1(_05281_),
    .A2(_05983_),
    .ZN(_01415_)
  );
  INV_X1 _22059_ (
    .A(_01415_),
    .ZN(_01416_)
  );
  AND2_X1 _22060_ (
    .A1(_06201_),
    .A2(_01416_),
    .ZN(_01417_)
  );
  AND2_X1 _22061_ (
    .A1(_01414_),
    .A2(_01417_),
    .ZN(_01418_)
  );
  INV_X1 _22062_ (
    .A(_01418_),
    .ZN(_01419_)
  );
  AND2_X1 _22063_ (
    .A1(remainder[20]),
    .A2(_00919_),
    .ZN(_01420_)
  );
  INV_X1 _22064_ (
    .A(_01420_),
    .ZN(_01422_)
  );
  AND2_X1 _22065_ (
    .A1(io_req_bits_in1[20]),
    .A2(_06190_),
    .ZN(_01423_)
  );
  INV_X1 _22066_ (
    .A(_01423_),
    .ZN(_01424_)
  );
  AND2_X1 _22067_ (
    .A1(_01422_),
    .A2(_01424_),
    .ZN(_01425_)
  );
  AND2_X1 _22068_ (
    .A1(_01419_),
    .A2(_01425_),
    .ZN(_01426_)
  );
  INV_X1 _22069_ (
    .A(_01426_),
    .ZN(_00107_)
  );
  AND2_X1 _22070_ (
    .A1(remainder[29]),
    .A2(_06103_),
    .ZN(_01427_)
  );
  INV_X1 _22071_ (
    .A(_01427_),
    .ZN(_01428_)
  );
  AND2_X1 _22072_ (
    .A1(_05994_),
    .A2(_01428_),
    .ZN(_01429_)
  );
  MUX2_X1 _22073_ (
    .A(remainder[21]),
    .B(remainder[54]),
    .S(resHi),
    .Z(io_resp_bits_data[21])
  );
  INV_X1 _22074_ (
    .A(io_resp_bits_data[21]),
    .ZN(_01431_)
  );
  AND2_X1 _22075_ (
    .A1(_01408_),
    .A2(io_resp_bits_data[21]),
    .ZN(_01432_)
  );
  INV_X1 _22076_ (
    .A(_01432_),
    .ZN(_01433_)
  );
  AND2_X1 _22077_ (
    .A1(_01407_),
    .A2(_01431_),
    .ZN(_01434_)
  );
  INV_X1 _22078_ (
    .A(_01434_),
    .ZN(_01435_)
  );
  AND2_X1 _22079_ (
    .A1(_00898_),
    .A2(_01435_),
    .ZN(_01436_)
  );
  AND2_X1 _22080_ (
    .A1(_01433_),
    .A2(_01436_),
    .ZN(_01437_)
  );
  INV_X1 _22081_ (
    .A(_01437_),
    .ZN(_01438_)
  );
  AND2_X1 _22082_ (
    .A1(_01429_),
    .A2(_01438_),
    .ZN(_01439_)
  );
  INV_X1 _22083_ (
    .A(_01439_),
    .ZN(_01440_)
  );
  AND2_X1 _22084_ (
    .A1(_05292_),
    .A2(_05983_),
    .ZN(_01442_)
  );
  INV_X1 _22085_ (
    .A(_01442_),
    .ZN(_01443_)
  );
  AND2_X1 _22086_ (
    .A1(_06201_),
    .A2(_01443_),
    .ZN(_01444_)
  );
  AND2_X1 _22087_ (
    .A1(_01440_),
    .A2(_01444_),
    .ZN(_01445_)
  );
  INV_X1 _22088_ (
    .A(_01445_),
    .ZN(_01446_)
  );
  AND2_X1 _22089_ (
    .A1(remainder[21]),
    .A2(_00919_),
    .ZN(_01447_)
  );
  INV_X1 _22090_ (
    .A(_01447_),
    .ZN(_01448_)
  );
  AND2_X1 _22091_ (
    .A1(io_req_bits_in1[21]),
    .A2(_06190_),
    .ZN(_01449_)
  );
  INV_X1 _22092_ (
    .A(_01449_),
    .ZN(_01450_)
  );
  AND2_X1 _22093_ (
    .A1(_01448_),
    .A2(_01450_),
    .ZN(_01451_)
  );
  AND2_X1 _22094_ (
    .A1(_01446_),
    .A2(_01451_),
    .ZN(_01453_)
  );
  INV_X1 _22095_ (
    .A(_01453_),
    .ZN(_00108_)
  );
  AND2_X1 _22096_ (
    .A1(remainder[30]),
    .A2(_06103_),
    .ZN(_01454_)
  );
  INV_X1 _22097_ (
    .A(_01454_),
    .ZN(_01455_)
  );
  AND2_X1 _22098_ (
    .A1(_05994_),
    .A2(_01455_),
    .ZN(_01456_)
  );
  MUX2_X1 _22099_ (
    .A(remainder[22]),
    .B(remainder[55]),
    .S(resHi),
    .Z(io_resp_bits_data[22])
  );
  INV_X1 _22100_ (
    .A(io_resp_bits_data[22]),
    .ZN(_01457_)
  );
  AND2_X1 _22101_ (
    .A1(_01435_),
    .A2(io_resp_bits_data[22]),
    .ZN(_01458_)
  );
  INV_X1 _22102_ (
    .A(_01458_),
    .ZN(_01459_)
  );
  AND2_X1 _22103_ (
    .A1(_01434_),
    .A2(_01457_),
    .ZN(_01460_)
  );
  INV_X1 _22104_ (
    .A(_01460_),
    .ZN(_01462_)
  );
  AND2_X1 _22105_ (
    .A1(_00898_),
    .A2(_01462_),
    .ZN(_01463_)
  );
  AND2_X1 _22106_ (
    .A1(_01459_),
    .A2(_01463_),
    .ZN(_01464_)
  );
  INV_X1 _22107_ (
    .A(_01464_),
    .ZN(_01465_)
  );
  AND2_X1 _22108_ (
    .A1(_01456_),
    .A2(_01465_),
    .ZN(_01466_)
  );
  INV_X1 _22109_ (
    .A(_01466_),
    .ZN(_01467_)
  );
  AND2_X1 _22110_ (
    .A1(_05303_),
    .A2(_05983_),
    .ZN(_01468_)
  );
  INV_X1 _22111_ (
    .A(_01468_),
    .ZN(_01469_)
  );
  AND2_X1 _22112_ (
    .A1(_06201_),
    .A2(_01469_),
    .ZN(_01470_)
  );
  AND2_X1 _22113_ (
    .A1(_01467_),
    .A2(_01470_),
    .ZN(_01471_)
  );
  INV_X1 _22114_ (
    .A(_01471_),
    .ZN(_01473_)
  );
  AND2_X1 _22115_ (
    .A1(remainder[22]),
    .A2(_00919_),
    .ZN(_01474_)
  );
  INV_X1 _22116_ (
    .A(_01474_),
    .ZN(_01475_)
  );
  AND2_X1 _22117_ (
    .A1(io_req_bits_in1[22]),
    .A2(_06190_),
    .ZN(_01476_)
  );
  INV_X1 _22118_ (
    .A(_01476_),
    .ZN(_01477_)
  );
  AND2_X1 _22119_ (
    .A1(_01475_),
    .A2(_01477_),
    .ZN(_01478_)
  );
  AND2_X1 _22120_ (
    .A1(_01473_),
    .A2(_01478_),
    .ZN(_01479_)
  );
  INV_X1 _22121_ (
    .A(_01479_),
    .ZN(_00109_)
  );
  AND2_X1 _22122_ (
    .A1(remainder[31]),
    .A2(_06103_),
    .ZN(_01480_)
  );
  INV_X1 _22123_ (
    .A(_01480_),
    .ZN(_01481_)
  );
  AND2_X1 _22124_ (
    .A1(_05994_),
    .A2(_01481_),
    .ZN(_01483_)
  );
  MUX2_X1 _22125_ (
    .A(remainder[23]),
    .B(remainder[56]),
    .S(resHi),
    .Z(io_resp_bits_data[23])
  );
  INV_X1 _22126_ (
    .A(io_resp_bits_data[23]),
    .ZN(_01484_)
  );
  AND2_X1 _22127_ (
    .A1(_01462_),
    .A2(io_resp_bits_data[23]),
    .ZN(_01485_)
  );
  INV_X1 _22128_ (
    .A(_01485_),
    .ZN(_01486_)
  );
  AND2_X1 _22129_ (
    .A1(_01460_),
    .A2(_01484_),
    .ZN(_01487_)
  );
  INV_X1 _22130_ (
    .A(_01487_),
    .ZN(_01488_)
  );
  AND2_X1 _22131_ (
    .A1(_00898_),
    .A2(_01488_),
    .ZN(_01489_)
  );
  AND2_X1 _22132_ (
    .A1(_01486_),
    .A2(_01489_),
    .ZN(_01490_)
  );
  INV_X1 _22133_ (
    .A(_01490_),
    .ZN(_01491_)
  );
  AND2_X1 _22134_ (
    .A1(_01483_),
    .A2(_01491_),
    .ZN(_01493_)
  );
  INV_X1 _22135_ (
    .A(_01493_),
    .ZN(_01494_)
  );
  AND2_X1 _22136_ (
    .A1(_05314_),
    .A2(_05983_),
    .ZN(_01495_)
  );
  INV_X1 _22137_ (
    .A(_01495_),
    .ZN(_01496_)
  );
  AND2_X1 _22138_ (
    .A1(_06201_),
    .A2(_01496_),
    .ZN(_01497_)
  );
  AND2_X1 _22139_ (
    .A1(_01494_),
    .A2(_01497_),
    .ZN(_01498_)
  );
  INV_X1 _22140_ (
    .A(_01498_),
    .ZN(_01499_)
  );
  AND2_X1 _22141_ (
    .A1(remainder[23]),
    .A2(_00919_),
    .ZN(_01500_)
  );
  INV_X1 _22142_ (
    .A(_01500_),
    .ZN(_01501_)
  );
  AND2_X1 _22143_ (
    .A1(io_req_bits_in1[23]),
    .A2(_06190_),
    .ZN(_01502_)
  );
  INV_X1 _22144_ (
    .A(_01502_),
    .ZN(_01504_)
  );
  AND2_X1 _22145_ (
    .A1(_01501_),
    .A2(_01504_),
    .ZN(_01505_)
  );
  AND2_X1 _22146_ (
    .A1(_01499_),
    .A2(_01505_),
    .ZN(_01506_)
  );
  INV_X1 _22147_ (
    .A(_01506_),
    .ZN(_00110_)
  );
  MUX2_X1 _22148_ (
    .A(remainder[24]),
    .B(remainder[57]),
    .S(resHi),
    .Z(io_resp_bits_data[24])
  );
  INV_X1 _22149_ (
    .A(io_resp_bits_data[24]),
    .ZN(_01507_)
  );
  AND2_X1 _22150_ (
    .A1(_01488_),
    .A2(io_resp_bits_data[24]),
    .ZN(_01508_)
  );
  INV_X1 _22151_ (
    .A(_01508_),
    .ZN(_01509_)
  );
  AND2_X1 _22152_ (
    .A1(_01487_),
    .A2(_01507_),
    .ZN(_01510_)
  );
  INV_X1 _22153_ (
    .A(_01510_),
    .ZN(_01511_)
  );
  AND2_X1 _22154_ (
    .A1(_00898_),
    .A2(_01511_),
    .ZN(_01513_)
  );
  AND2_X1 _22155_ (
    .A1(_01509_),
    .A2(_01513_),
    .ZN(_01514_)
  );
  INV_X1 _22156_ (
    .A(_01514_),
    .ZN(_01515_)
  );
  AND2_X1 _22157_ (
    .A1(_04755_),
    .A2(_02468_),
    .ZN(_01516_)
  );
  INV_X1 _22158_ (
    .A(_01516_),
    .ZN(_01517_)
  );
  AND2_X1 _22159_ (
    .A1(_06103_),
    .A2(_02558_),
    .ZN(_01518_)
  );
  AND2_X1 _22160_ (
    .A1(_01517_),
    .A2(_01518_),
    .ZN(_01519_)
  );
  INV_X1 _22161_ (
    .A(_01519_),
    .ZN(_01520_)
  );
  AND2_X1 _22162_ (
    .A1(_05994_),
    .A2(_01520_),
    .ZN(_01521_)
  );
  AND2_X1 _22163_ (
    .A1(_01515_),
    .A2(_01521_),
    .ZN(_01522_)
  );
  INV_X1 _22164_ (
    .A(_01522_),
    .ZN(_01524_)
  );
  AND2_X1 _22165_ (
    .A1(_05325_),
    .A2(_05983_),
    .ZN(_01525_)
  );
  INV_X1 _22166_ (
    .A(_01525_),
    .ZN(_01526_)
  );
  AND2_X1 _22167_ (
    .A1(_06201_),
    .A2(_01526_),
    .ZN(_01527_)
  );
  AND2_X1 _22168_ (
    .A1(_01524_),
    .A2(_01527_),
    .ZN(_01528_)
  );
  INV_X1 _22169_ (
    .A(_01528_),
    .ZN(_01529_)
  );
  AND2_X1 _22170_ (
    .A1(remainder[24]),
    .A2(_00919_),
    .ZN(_01530_)
  );
  INV_X1 _22171_ (
    .A(_01530_),
    .ZN(_01531_)
  );
  AND2_X1 _22172_ (
    .A1(io_req_bits_in1[24]),
    .A2(_06190_),
    .ZN(_01532_)
  );
  INV_X1 _22173_ (
    .A(_01532_),
    .ZN(_01533_)
  );
  AND2_X1 _22174_ (
    .A1(_01531_),
    .A2(_01533_),
    .ZN(_01534_)
  );
  AND2_X1 _22175_ (
    .A1(_01529_),
    .A2(_01534_),
    .ZN(_01535_)
  );
  INV_X1 _22176_ (
    .A(_01535_),
    .ZN(_00111_)
  );
  MUX2_X1 _22177_ (
    .A(remainder[25]),
    .B(remainder[58]),
    .S(resHi),
    .Z(io_resp_bits_data[25])
  );
  INV_X1 _22178_ (
    .A(io_resp_bits_data[25]),
    .ZN(_01536_)
  );
  AND2_X1 _22179_ (
    .A1(_01511_),
    .A2(io_resp_bits_data[25]),
    .ZN(_01537_)
  );
  INV_X1 _22180_ (
    .A(_01537_),
    .ZN(_01538_)
  );
  AND2_X1 _22181_ (
    .A1(_01510_),
    .A2(_01536_),
    .ZN(_01539_)
  );
  INV_X1 _22182_ (
    .A(_01539_),
    .ZN(_01540_)
  );
  AND2_X1 _22183_ (
    .A1(_00898_),
    .A2(_01540_),
    .ZN(_01541_)
  );
  AND2_X1 _22184_ (
    .A1(_01538_),
    .A2(_01541_),
    .ZN(_01543_)
  );
  INV_X1 _22185_ (
    .A(_01543_),
    .ZN(_01544_)
  );
  AND2_X1 _22186_ (
    .A1(_02558_),
    .A2(_02562_),
    .ZN(_01545_)
  );
  INV_X1 _22187_ (
    .A(_01545_),
    .ZN(_01546_)
  );
  AND2_X1 _22188_ (
    .A1(_06103_),
    .A2(_02564_),
    .ZN(_01547_)
  );
  AND2_X1 _22189_ (
    .A1(_01546_),
    .A2(_01547_),
    .ZN(_01548_)
  );
  INV_X1 _22190_ (
    .A(_01548_),
    .ZN(_01549_)
  );
  AND2_X1 _22191_ (
    .A1(_05994_),
    .A2(_01549_),
    .ZN(_01550_)
  );
  AND2_X1 _22192_ (
    .A1(_01544_),
    .A2(_01550_),
    .ZN(_01551_)
  );
  INV_X1 _22193_ (
    .A(_01551_),
    .ZN(_01552_)
  );
  AND2_X1 _22194_ (
    .A1(_05336_),
    .A2(_05983_),
    .ZN(_01554_)
  );
  INV_X1 _22195_ (
    .A(_01554_),
    .ZN(_01555_)
  );
  AND2_X1 _22196_ (
    .A1(_06201_),
    .A2(_01555_),
    .ZN(_01556_)
  );
  AND2_X1 _22197_ (
    .A1(_01552_),
    .A2(_01556_),
    .ZN(_01557_)
  );
  INV_X1 _22198_ (
    .A(_01557_),
    .ZN(_01558_)
  );
  AND2_X1 _22199_ (
    .A1(remainder[25]),
    .A2(_00919_),
    .ZN(_01559_)
  );
  INV_X1 _22200_ (
    .A(_01559_),
    .ZN(_01560_)
  );
  AND2_X1 _22201_ (
    .A1(io_req_bits_in1[25]),
    .A2(_06190_),
    .ZN(_01561_)
  );
  INV_X1 _22202_ (
    .A(_01561_),
    .ZN(_01562_)
  );
  AND2_X1 _22203_ (
    .A1(_01560_),
    .A2(_01562_),
    .ZN(_01563_)
  );
  AND2_X1 _22204_ (
    .A1(_01558_),
    .A2(_01563_),
    .ZN(_01565_)
  );
  INV_X1 _22205_ (
    .A(_01565_),
    .ZN(_00112_)
  );
  MUX2_X1 _22206_ (
    .A(remainder[26]),
    .B(remainder[59]),
    .S(resHi),
    .Z(io_resp_bits_data[26])
  );
  INV_X1 _22207_ (
    .A(io_resp_bits_data[26]),
    .ZN(_01566_)
  );
  AND2_X1 _22208_ (
    .A1(_01540_),
    .A2(io_resp_bits_data[26]),
    .ZN(_01567_)
  );
  INV_X1 _22209_ (
    .A(_01567_),
    .ZN(_01568_)
  );
  AND2_X1 _22210_ (
    .A1(_01539_),
    .A2(_01566_),
    .ZN(_01569_)
  );
  INV_X1 _22211_ (
    .A(_01569_),
    .ZN(_01570_)
  );
  AND2_X1 _22212_ (
    .A1(_00898_),
    .A2(_01570_),
    .ZN(_01571_)
  );
  AND2_X1 _22213_ (
    .A1(_01568_),
    .A2(_01571_),
    .ZN(_01572_)
  );
  INV_X1 _22214_ (
    .A(_01572_),
    .ZN(_01574_)
  );
  AND2_X1 _22215_ (
    .A1(_02565_),
    .A2(_02570_),
    .ZN(_01575_)
  );
  INV_X1 _22216_ (
    .A(_01575_),
    .ZN(_01576_)
  );
  AND2_X1 _22217_ (
    .A1(_06103_),
    .A2(_02572_),
    .ZN(_01577_)
  );
  AND2_X1 _22218_ (
    .A1(_01576_),
    .A2(_01577_),
    .ZN(_01578_)
  );
  INV_X1 _22219_ (
    .A(_01578_),
    .ZN(_01579_)
  );
  AND2_X1 _22220_ (
    .A1(_05994_),
    .A2(_01579_),
    .ZN(_01580_)
  );
  AND2_X1 _22221_ (
    .A1(_01574_),
    .A2(_01580_),
    .ZN(_01581_)
  );
  INV_X1 _22222_ (
    .A(_01581_),
    .ZN(_01582_)
  );
  AND2_X1 _22223_ (
    .A1(_05347_),
    .A2(_05983_),
    .ZN(_01583_)
  );
  INV_X1 _22224_ (
    .A(_01583_),
    .ZN(_01585_)
  );
  AND2_X1 _22225_ (
    .A1(_06201_),
    .A2(_01585_),
    .ZN(_01586_)
  );
  AND2_X1 _22226_ (
    .A1(_01582_),
    .A2(_01586_),
    .ZN(_01587_)
  );
  INV_X1 _22227_ (
    .A(_01587_),
    .ZN(_01588_)
  );
  AND2_X1 _22228_ (
    .A1(remainder[26]),
    .A2(_00919_),
    .ZN(_01589_)
  );
  INV_X1 _22229_ (
    .A(_01589_),
    .ZN(_01590_)
  );
  AND2_X1 _22230_ (
    .A1(io_req_bits_in1[26]),
    .A2(_06190_),
    .ZN(_01591_)
  );
  INV_X1 _22231_ (
    .A(_01591_),
    .ZN(_01592_)
  );
  AND2_X1 _22232_ (
    .A1(_01590_),
    .A2(_01592_),
    .ZN(_01593_)
  );
  AND2_X1 _22233_ (
    .A1(_01588_),
    .A2(_01593_),
    .ZN(_01594_)
  );
  INV_X1 _22234_ (
    .A(_01594_),
    .ZN(_00113_)
  );
  MUX2_X1 _22235_ (
    .A(remainder[27]),
    .B(remainder[60]),
    .S(resHi),
    .Z(io_resp_bits_data[27])
  );
  INV_X1 _22236_ (
    .A(io_resp_bits_data[27]),
    .ZN(_01596_)
  );
  AND2_X1 _22237_ (
    .A1(_01570_),
    .A2(io_resp_bits_data[27]),
    .ZN(_01597_)
  );
  INV_X1 _22238_ (
    .A(_01597_),
    .ZN(_01598_)
  );
  AND2_X1 _22239_ (
    .A1(_01569_),
    .A2(_01596_),
    .ZN(_01599_)
  );
  INV_X1 _22240_ (
    .A(_01599_),
    .ZN(_01600_)
  );
  AND2_X1 _22241_ (
    .A1(_00898_),
    .A2(_01600_),
    .ZN(_01601_)
  );
  AND2_X1 _22242_ (
    .A1(_01598_),
    .A2(_01601_),
    .ZN(_01602_)
  );
  INV_X1 _22243_ (
    .A(_01602_),
    .ZN(_01603_)
  );
  AND2_X1 _22244_ (
    .A1(_02542_),
    .A2(_02544_),
    .ZN(_01605_)
  );
  INV_X1 _22245_ (
    .A(_01605_),
    .ZN(_01606_)
  );
  AND2_X1 _22246_ (
    .A1(_02574_),
    .A2(_01605_),
    .ZN(_01607_)
  );
  INV_X1 _22247_ (
    .A(_01607_),
    .ZN(_01608_)
  );
  AND2_X1 _22248_ (
    .A1(_02573_),
    .A2(_01606_),
    .ZN(_01609_)
  );
  INV_X1 _22249_ (
    .A(_01609_),
    .ZN(_01610_)
  );
  AND2_X1 _22250_ (
    .A1(_06103_),
    .A2(_01608_),
    .ZN(_01611_)
  );
  AND2_X1 _22251_ (
    .A1(_01610_),
    .A2(_01611_),
    .ZN(_01612_)
  );
  INV_X1 _22252_ (
    .A(_01612_),
    .ZN(_01613_)
  );
  AND2_X1 _22253_ (
    .A1(_05994_),
    .A2(_01613_),
    .ZN(_01614_)
  );
  AND2_X1 _22254_ (
    .A1(_01603_),
    .A2(_01614_),
    .ZN(_01616_)
  );
  INV_X1 _22255_ (
    .A(_01616_),
    .ZN(_01617_)
  );
  AND2_X1 _22256_ (
    .A1(_05358_),
    .A2(_05983_),
    .ZN(_01618_)
  );
  INV_X1 _22257_ (
    .A(_01618_),
    .ZN(_01619_)
  );
  AND2_X1 _22258_ (
    .A1(_06201_),
    .A2(_01619_),
    .ZN(_01620_)
  );
  AND2_X1 _22259_ (
    .A1(_01617_),
    .A2(_01620_),
    .ZN(_01621_)
  );
  INV_X1 _22260_ (
    .A(_01621_),
    .ZN(_01622_)
  );
  AND2_X1 _22261_ (
    .A1(remainder[27]),
    .A2(_00919_),
    .ZN(_01623_)
  );
  INV_X1 _22262_ (
    .A(_01623_),
    .ZN(_01624_)
  );
  AND2_X1 _22263_ (
    .A1(io_req_bits_in1[27]),
    .A2(_06190_),
    .ZN(_01625_)
  );
  INV_X1 _22264_ (
    .A(_01625_),
    .ZN(_01627_)
  );
  AND2_X1 _22265_ (
    .A1(_01624_),
    .A2(_01627_),
    .ZN(_01628_)
  );
  AND2_X1 _22266_ (
    .A1(_01622_),
    .A2(_01628_),
    .ZN(_01629_)
  );
  INV_X1 _22267_ (
    .A(_01629_),
    .ZN(_00114_)
  );
  MUX2_X1 _22268_ (
    .A(remainder[28]),
    .B(remainder[61]),
    .S(resHi),
    .Z(io_resp_bits_data[28])
  );
  INV_X1 _22269_ (
    .A(io_resp_bits_data[28]),
    .ZN(_01630_)
  );
  AND2_X1 _22270_ (
    .A1(_01600_),
    .A2(io_resp_bits_data[28]),
    .ZN(_01631_)
  );
  INV_X1 _22271_ (
    .A(_01631_),
    .ZN(_01632_)
  );
  AND2_X1 _22272_ (
    .A1(_01599_),
    .A2(_01630_),
    .ZN(_01633_)
  );
  INV_X1 _22273_ (
    .A(_01633_),
    .ZN(_01634_)
  );
  AND2_X1 _22274_ (
    .A1(_00898_),
    .A2(_01634_),
    .ZN(_01636_)
  );
  AND2_X1 _22275_ (
    .A1(_01632_),
    .A2(_01636_),
    .ZN(_01637_)
  );
  INV_X1 _22276_ (
    .A(_01637_),
    .ZN(_01638_)
  );
  AND2_X1 _22277_ (
    .A1(_02536_),
    .A2(_02579_),
    .ZN(_01639_)
  );
  INV_X1 _22278_ (
    .A(_01639_),
    .ZN(_01640_)
  );
  AND2_X1 _22279_ (
    .A1(_06103_),
    .A2(_02582_),
    .ZN(_01641_)
  );
  AND2_X1 _22280_ (
    .A1(_01640_),
    .A2(_01641_),
    .ZN(_01642_)
  );
  INV_X1 _22281_ (
    .A(_01642_),
    .ZN(_01643_)
  );
  AND2_X1 _22282_ (
    .A1(_05994_),
    .A2(_01643_),
    .ZN(_01644_)
  );
  AND2_X1 _22283_ (
    .A1(_01638_),
    .A2(_01644_),
    .ZN(_01645_)
  );
  INV_X1 _22284_ (
    .A(_01645_),
    .ZN(_01647_)
  );
  AND2_X1 _22285_ (
    .A1(_05369_),
    .A2(_05983_),
    .ZN(_01648_)
  );
  INV_X1 _22286_ (
    .A(_01648_),
    .ZN(_01649_)
  );
  AND2_X1 _22287_ (
    .A1(_06201_),
    .A2(_01649_),
    .ZN(_01650_)
  );
  AND2_X1 _22288_ (
    .A1(_01647_),
    .A2(_01650_),
    .ZN(_01651_)
  );
  INV_X1 _22289_ (
    .A(_01651_),
    .ZN(_01652_)
  );
  AND2_X1 _22290_ (
    .A1(remainder[28]),
    .A2(_00919_),
    .ZN(_01653_)
  );
  INV_X1 _22291_ (
    .A(_01653_),
    .ZN(_01654_)
  );
  AND2_X1 _22292_ (
    .A1(io_req_bits_in1[28]),
    .A2(_06190_),
    .ZN(_01655_)
  );
  INV_X1 _22293_ (
    .A(_01655_),
    .ZN(_01656_)
  );
  AND2_X1 _22294_ (
    .A1(_01654_),
    .A2(_01656_),
    .ZN(_01658_)
  );
  AND2_X1 _22295_ (
    .A1(_01652_),
    .A2(_01658_),
    .ZN(_01659_)
  );
  INV_X1 _22296_ (
    .A(_01659_),
    .ZN(_00115_)
  );
  MUX2_X1 _22297_ (
    .A(remainder[29]),
    .B(remainder[62]),
    .S(resHi),
    .Z(io_resp_bits_data[29])
  );
  INV_X1 _22298_ (
    .A(io_resp_bits_data[29]),
    .ZN(_01660_)
  );
  AND2_X1 _22299_ (
    .A1(_01634_),
    .A2(io_resp_bits_data[29]),
    .ZN(_01661_)
  );
  INV_X1 _22300_ (
    .A(_01661_),
    .ZN(_01662_)
  );
  AND2_X1 _22301_ (
    .A1(_01633_),
    .A2(_01660_),
    .ZN(_01663_)
  );
  INV_X1 _22302_ (
    .A(_01663_),
    .ZN(_01664_)
  );
  AND2_X1 _22303_ (
    .A1(_00898_),
    .A2(_01664_),
    .ZN(_01665_)
  );
  AND2_X1 _22304_ (
    .A1(_01662_),
    .A2(_01665_),
    .ZN(_01667_)
  );
  INV_X1 _22305_ (
    .A(_01667_),
    .ZN(_01668_)
  );
  AND2_X1 _22306_ (
    .A1(_02526_),
    .A2(_02583_),
    .ZN(_01669_)
  );
  INV_X1 _22307_ (
    .A(_01669_),
    .ZN(_01670_)
  );
  AND2_X1 _22308_ (
    .A1(_06103_),
    .A2(_02586_),
    .ZN(_01671_)
  );
  AND2_X1 _22309_ (
    .A1(_01670_),
    .A2(_01671_),
    .ZN(_01672_)
  );
  INV_X1 _22310_ (
    .A(_01672_),
    .ZN(_01673_)
  );
  AND2_X1 _22311_ (
    .A1(_05994_),
    .A2(_01673_),
    .ZN(_01674_)
  );
  AND2_X1 _22312_ (
    .A1(_01668_),
    .A2(_01674_),
    .ZN(_01675_)
  );
  INV_X1 _22313_ (
    .A(_01675_),
    .ZN(_01676_)
  );
  AND2_X1 _22314_ (
    .A1(_05380_),
    .A2(_05983_),
    .ZN(_01678_)
  );
  INV_X1 _22315_ (
    .A(_01678_),
    .ZN(_01679_)
  );
  AND2_X1 _22316_ (
    .A1(_06201_),
    .A2(_01679_),
    .ZN(_01680_)
  );
  AND2_X1 _22317_ (
    .A1(_01676_),
    .A2(_01680_),
    .ZN(_01681_)
  );
  INV_X1 _22318_ (
    .A(_01681_),
    .ZN(_01682_)
  );
  AND2_X1 _22319_ (
    .A1(remainder[29]),
    .A2(_00919_),
    .ZN(_01683_)
  );
  INV_X1 _22320_ (
    .A(_01683_),
    .ZN(_01684_)
  );
  AND2_X1 _22321_ (
    .A1(io_req_bits_in1[29]),
    .A2(_06190_),
    .ZN(_01685_)
  );
  INV_X1 _22322_ (
    .A(_01685_),
    .ZN(_01686_)
  );
  AND2_X1 _22323_ (
    .A1(_01684_),
    .A2(_01686_),
    .ZN(_01687_)
  );
  AND2_X1 _22324_ (
    .A1(_01682_),
    .A2(_01687_),
    .ZN(_01689_)
  );
  INV_X1 _22325_ (
    .A(_01689_),
    .ZN(_00116_)
  );
  MUX2_X1 _22326_ (
    .A(remainder[30]),
    .B(remainder[63]),
    .S(resHi),
    .Z(io_resp_bits_data[30])
  );
  INV_X1 _22327_ (
    .A(io_resp_bits_data[30]),
    .ZN(_01690_)
  );
  AND2_X1 _22328_ (
    .A1(_01664_),
    .A2(io_resp_bits_data[30]),
    .ZN(_01691_)
  );
  INV_X1 _22329_ (
    .A(_01691_),
    .ZN(_01692_)
  );
  AND2_X1 _22330_ (
    .A1(_01663_),
    .A2(_01690_),
    .ZN(_01693_)
  );
  INV_X1 _22331_ (
    .A(_01693_),
    .ZN(_01694_)
  );
  AND2_X1 _22332_ (
    .A1(_00898_),
    .A2(_01694_),
    .ZN(_01695_)
  );
  AND2_X1 _22333_ (
    .A1(_01692_),
    .A2(_01695_),
    .ZN(_01696_)
  );
  INV_X1 _22334_ (
    .A(_01696_),
    .ZN(_01698_)
  );
  AND2_X1 _22335_ (
    .A1(_02587_),
    .A2(_02592_),
    .ZN(_01699_)
  );
  INV_X1 _22336_ (
    .A(_01699_),
    .ZN(_01700_)
  );
  AND2_X1 _22337_ (
    .A1(_06103_),
    .A2(_02594_),
    .ZN(_01701_)
  );
  AND2_X1 _22338_ (
    .A1(_01700_),
    .A2(_01701_),
    .ZN(_01702_)
  );
  INV_X1 _22339_ (
    .A(_01702_),
    .ZN(_01703_)
  );
  AND2_X1 _22340_ (
    .A1(_05994_),
    .A2(_01703_),
    .ZN(_01704_)
  );
  AND2_X1 _22341_ (
    .A1(_01698_),
    .A2(_01704_),
    .ZN(_01705_)
  );
  INV_X1 _22342_ (
    .A(_01705_),
    .ZN(_01706_)
  );
  AND2_X1 _22343_ (
    .A1(_05391_),
    .A2(_05983_),
    .ZN(_01707_)
  );
  INV_X1 _22344_ (
    .A(_01707_),
    .ZN(_01708_)
  );
  AND2_X1 _22345_ (
    .A1(_06201_),
    .A2(_01708_),
    .ZN(_01709_)
  );
  AND2_X1 _22346_ (
    .A1(_01706_),
    .A2(_01709_),
    .ZN(_01710_)
  );
  INV_X1 _22347_ (
    .A(_01710_),
    .ZN(_01711_)
  );
  AND2_X1 _22348_ (
    .A1(remainder[30]),
    .A2(_00919_),
    .ZN(_01712_)
  );
  INV_X1 _22349_ (
    .A(_01712_),
    .ZN(_01713_)
  );
  AND2_X1 _22350_ (
    .A1(io_req_bits_in1[30]),
    .A2(_06190_),
    .ZN(_01714_)
  );
  INV_X1 _22351_ (
    .A(_01714_),
    .ZN(_01715_)
  );
  AND2_X1 _22352_ (
    .A1(_01713_),
    .A2(_01715_),
    .ZN(_01716_)
  );
  AND2_X1 _22353_ (
    .A1(_01711_),
    .A2(_01716_),
    .ZN(_01717_)
  );
  INV_X1 _22354_ (
    .A(_01717_),
    .ZN(_00117_)
  );
  MUX2_X1 _22355_ (
    .A(remainder[31]),
    .B(remainder[64]),
    .S(resHi),
    .Z(io_resp_bits_data[31])
  );
  INV_X1 _22356_ (
    .A(io_resp_bits_data[31]),
    .ZN(_01719_)
  );
  AND2_X1 _22357_ (
    .A1(_01694_),
    .A2(io_resp_bits_data[31]),
    .ZN(_01720_)
  );
  INV_X1 _22358_ (
    .A(_01720_),
    .ZN(_01721_)
  );
  AND2_X1 _22359_ (
    .A1(_01693_),
    .A2(_01719_),
    .ZN(_01722_)
  );
  INV_X1 _22360_ (
    .A(_01722_),
    .ZN(_01723_)
  );
  AND2_X1 _22361_ (
    .A1(_01721_),
    .A2(_01723_),
    .ZN(_01724_)
  );
  AND2_X1 _22362_ (
    .A1(_00898_),
    .A2(_01724_),
    .ZN(_01725_)
  );
  INV_X1 _22363_ (
    .A(_01725_),
    .ZN(_01726_)
  );
  AND2_X1 _22364_ (
    .A1(_02595_),
    .A2(_02600_),
    .ZN(_01728_)
  );
  INV_X1 _22365_ (
    .A(_01728_),
    .ZN(_01729_)
  );
  AND2_X1 _22366_ (
    .A1(_06103_),
    .A2(_01729_),
    .ZN(_01730_)
  );
  AND2_X1 _22367_ (
    .A1(_02602_),
    .A2(_01730_),
    .ZN(_01731_)
  );
  INV_X1 _22368_ (
    .A(_01731_),
    .ZN(_01732_)
  );
  AND2_X1 _22369_ (
    .A1(_05994_),
    .A2(_01732_),
    .ZN(_01733_)
  );
  AND2_X1 _22370_ (
    .A1(_01726_),
    .A2(_01733_),
    .ZN(_01734_)
  );
  INV_X1 _22371_ (
    .A(_01734_),
    .ZN(_01735_)
  );
  AND2_X1 _22372_ (
    .A1(_05402_),
    .A2(_05983_),
    .ZN(_01736_)
  );
  INV_X1 _22373_ (
    .A(_01736_),
    .ZN(_01737_)
  );
  AND2_X1 _22374_ (
    .A1(_06201_),
    .A2(_01737_),
    .ZN(_01739_)
  );
  AND2_X1 _22375_ (
    .A1(_01735_),
    .A2(_01739_),
    .ZN(_01740_)
  );
  INV_X1 _22376_ (
    .A(_01740_),
    .ZN(_01741_)
  );
  AND2_X1 _22377_ (
    .A1(remainder[31]),
    .A2(_00919_),
    .ZN(_01742_)
  );
  INV_X1 _22378_ (
    .A(_01742_),
    .ZN(_01743_)
  );
  AND2_X1 _22379_ (
    .A1(io_req_bits_in1[31]),
    .A2(_06190_),
    .ZN(_01744_)
  );
  INV_X1 _22380_ (
    .A(_01744_),
    .ZN(_01745_)
  );
  AND2_X1 _22381_ (
    .A1(_01743_),
    .A2(_01745_),
    .ZN(_01746_)
  );
  AND2_X1 _22382_ (
    .A1(_01741_),
    .A2(_01746_),
    .ZN(_01747_)
  );
  INV_X1 _22383_ (
    .A(_01747_),
    .ZN(_00118_)
  );
  AND2_X1 _22384_ (
    .A1(_05434_),
    .A2(_06267_),
    .ZN(_01749_)
  );
  INV_X1 _22385_ (
    .A(_01749_),
    .ZN(_01750_)
  );
  AND2_X1 _22386_ (
    .A1(_06462_),
    .A2(_01750_),
    .ZN(_01751_)
  );
  AND2_X1 _22387_ (
    .A1(_04842_),
    .A2(_01751_),
    .ZN(_00119_)
  );
  MUX2_X1 _22388_ (
    .A(isHi),
    .B(_10594_),
    .S(_06190_),
    .Z(_00120_)
  );
  DFF_X1 \count[0]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00014_),
    .Q(count[0]),
    .QN(_count_T_1[0])
  );
  DFF_X1 \count[1]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00015_),
    .Q(count[1]),
    .QN(_00002_)
  );
  DFF_X1 \count[2]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00016_),
    .Q(count[2]),
    .QN(_11210_)
  );
  DFF_X1 \count[3]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00017_),
    .Q(count[3]),
    .QN(_11209_)
  );
  DFF_X1 \count[4]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00018_),
    .Q(count[4]),
    .QN(_11208_)
  );
  DFF_X1 \count[5]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00019_),
    .Q(count[5]),
    .QN(_00001_)
  );
  DFF_X1 \divisor[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00020_),
    .Q(divisor[0]),
    .QN(_11217_[0])
  );
  DFF_X1 \divisor[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00030_),
    .Q(divisor[10]),
    .QN(_11217_[10])
  );
  DFF_X1 \divisor[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00031_),
    .Q(divisor[11]),
    .QN(_11217_[11])
  );
  DFF_X1 \divisor[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00032_),
    .Q(divisor[12]),
    .QN(_11217_[12])
  );
  DFF_X1 \divisor[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00033_),
    .Q(divisor[13]),
    .QN(_11217_[13])
  );
  DFF_X1 \divisor[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00034_),
    .Q(divisor[14]),
    .QN(_11217_[14])
  );
  DFF_X1 \divisor[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00035_),
    .Q(divisor[15]),
    .QN(_11217_[15])
  );
  DFF_X1 \divisor[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00036_),
    .Q(divisor[16]),
    .QN(_11217_[16])
  );
  DFF_X1 \divisor[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00037_),
    .Q(divisor[17]),
    .QN(_11217_[17])
  );
  DFF_X1 \divisor[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00038_),
    .Q(divisor[18]),
    .QN(_11217_[18])
  );
  DFF_X1 \divisor[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00039_),
    .Q(divisor[19]),
    .QN(_11217_[19])
  );
  DFF_X1 \divisor[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00021_),
    .Q(divisor[1]),
    .QN(_11217_[1])
  );
  DFF_X1 \divisor[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00040_),
    .Q(divisor[20]),
    .QN(_11217_[20])
  );
  DFF_X1 \divisor[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00041_),
    .Q(divisor[21]),
    .QN(_11217_[21])
  );
  DFF_X1 \divisor[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00042_),
    .Q(divisor[22]),
    .QN(_11217_[22])
  );
  DFF_X1 \divisor[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00043_),
    .Q(divisor[23]),
    .QN(_11217_[23])
  );
  DFF_X1 \divisor[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00044_),
    .Q(divisor[24]),
    .QN(_11217_[24])
  );
  DFF_X1 \divisor[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00045_),
    .Q(divisor[25]),
    .QN(_11217_[25])
  );
  DFF_X1 \divisor[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00046_),
    .Q(divisor[26]),
    .QN(_11217_[26])
  );
  DFF_X1 \divisor[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00047_),
    .Q(divisor[27]),
    .QN(_11217_[27])
  );
  DFF_X1 \divisor[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00048_),
    .Q(divisor[28]),
    .QN(_11217_[28])
  );
  DFF_X1 \divisor[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00049_),
    .Q(divisor[29]),
    .QN(_11217_[29])
  );
  DFF_X1 \divisor[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00022_),
    .Q(divisor[2]),
    .QN(_11217_[2])
  );
  DFF_X1 \divisor[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00050_),
    .Q(divisor[30]),
    .QN(_11217_[30])
  );
  DFF_X1 \divisor[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00051_),
    .Q(divisor[31]),
    .QN(_11217_[31])
  );
  DFF_X1 \divisor[32]$_DFFE_PP_  (
    .CK(clock),
    .D(_00052_),
    .Q(divisor[32]),
    .QN(_11217_[32])
  );
  DFF_X1 \divisor[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00023_),
    .Q(divisor[3]),
    .QN(_11217_[3])
  );
  DFF_X1 \divisor[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00024_),
    .Q(divisor[4]),
    .QN(_11217_[4])
  );
  DFF_X1 \divisor[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00025_),
    .Q(divisor[5]),
    .QN(_11217_[5])
  );
  DFF_X1 \divisor[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00026_),
    .Q(divisor[6]),
    .QN(_11217_[6])
  );
  DFF_X1 \divisor[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00027_),
    .Q(divisor[7]),
    .QN(_11217_[7])
  );
  DFF_X1 \divisor[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00028_),
    .Q(divisor[8]),
    .QN(_11217_[8])
  );
  DFF_X1 \divisor[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00029_),
    .Q(divisor[9]),
    .QN(_11217_[9])
  );
  DFF_X1 \isHi$_DFFE_PP_  (
    .CK(clock),
    .D(_00120_),
    .Q(isHi),
    .QN(_eOut_T_4)
  );
  DFF_X1 \neg_out$_DFFE_PP_  (
    .CK(clock),
    .D(_00008_),
    .Q(neg_out),
    .QN(_state_T[1])
  );
  DFF_X1 \remainder[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00087_),
    .Q(remainder[0]),
    .QN(_11173_)
  );
  DFF_X1 \remainder[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00097_),
    .Q(remainder[10]),
    .QN(_11163_)
  );
  DFF_X1 \remainder[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00098_),
    .Q(remainder[11]),
    .QN(_11162_)
  );
  DFF_X1 \remainder[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00099_),
    .Q(remainder[12]),
    .QN(_11161_)
  );
  DFF_X1 \remainder[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00100_),
    .Q(remainder[13]),
    .QN(_11160_)
  );
  DFF_X1 \remainder[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00101_),
    .Q(remainder[14]),
    .QN(_11159_)
  );
  DFF_X1 \remainder[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00102_),
    .Q(remainder[15]),
    .QN(_11158_)
  );
  DFF_X1 \remainder[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00103_),
    .Q(remainder[16]),
    .QN(_11157_)
  );
  DFF_X1 \remainder[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00104_),
    .Q(remainder[17]),
    .QN(_11156_)
  );
  DFF_X1 \remainder[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00105_),
    .Q(remainder[18]),
    .QN(_11155_)
  );
  DFF_X1 \remainder[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00106_),
    .Q(remainder[19]),
    .QN(_11154_)
  );
  DFF_X1 \remainder[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00088_),
    .Q(remainder[1]),
    .QN(_11172_)
  );
  DFF_X1 \remainder[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00107_),
    .Q(remainder[20]),
    .QN(_11153_)
  );
  DFF_X1 \remainder[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00108_),
    .Q(remainder[21]),
    .QN(_11152_)
  );
  DFF_X1 \remainder[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00109_),
    .Q(remainder[22]),
    .QN(_11151_)
  );
  DFF_X1 \remainder[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00110_),
    .Q(remainder[23]),
    .QN(_11150_)
  );
  DFF_X1 \remainder[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00111_),
    .Q(remainder[24]),
    .QN(_11149_)
  );
  DFF_X1 \remainder[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00112_),
    .Q(remainder[25]),
    .QN(_11148_)
  );
  DFF_X1 \remainder[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00113_),
    .Q(remainder[26]),
    .QN(_11147_)
  );
  DFF_X1 \remainder[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00114_),
    .Q(remainder[27]),
    .QN(_11146_)
  );
  DFF_X1 \remainder[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00115_),
    .Q(remainder[28]),
    .QN(_11145_)
  );
  DFF_X1 \remainder[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00116_),
    .Q(remainder[29]),
    .QN(_11144_)
  );
  DFF_X1 \remainder[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00089_),
    .Q(remainder[2]),
    .QN(_11171_)
  );
  DFF_X1 \remainder[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00117_),
    .Q(remainder[30]),
    .QN(_11143_)
  );
  DFF_X1 \remainder[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00118_),
    .Q(remainder[31]),
    .QN(_11142_)
  );
  DFF_X1 \remainder[32]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00053_),
    .Q(remainder[32]),
    .QN(_11207_)
  );
  DFF_X1 \remainder[33]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00054_),
    .Q(remainder[33]),
    .QN(_11206_)
  );
  DFF_X1 \remainder[34]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00055_),
    .Q(remainder[34]),
    .QN(_11205_)
  );
  DFF_X1 \remainder[35]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00056_),
    .Q(remainder[35]),
    .QN(_11204_)
  );
  DFF_X1 \remainder[36]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00057_),
    .Q(remainder[36]),
    .QN(_11203_)
  );
  DFF_X1 \remainder[37]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00058_),
    .Q(remainder[37]),
    .QN(_11202_)
  );
  DFF_X1 \remainder[38]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00059_),
    .Q(remainder[38]),
    .QN(_11201_)
  );
  DFF_X1 \remainder[39]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00060_),
    .Q(remainder[39]),
    .QN(_11200_)
  );
  DFF_X1 \remainder[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00090_),
    .Q(remainder[3]),
    .QN(_11170_)
  );
  DFF_X1 \remainder[40]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00061_),
    .Q(remainder[40]),
    .QN(_11199_)
  );
  DFF_X1 \remainder[41]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00062_),
    .Q(remainder[41]),
    .QN(_11198_)
  );
  DFF_X1 \remainder[42]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00063_),
    .Q(remainder[42]),
    .QN(_11197_)
  );
  DFF_X1 \remainder[43]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00064_),
    .Q(remainder[43]),
    .QN(_11196_)
  );
  DFF_X1 \remainder[44]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00065_),
    .Q(remainder[44]),
    .QN(_11195_)
  );
  DFF_X1 \remainder[45]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00066_),
    .Q(remainder[45]),
    .QN(_11194_)
  );
  DFF_X1 \remainder[46]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00067_),
    .Q(remainder[46]),
    .QN(_11193_)
  );
  DFF_X1 \remainder[47]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00068_),
    .Q(remainder[47]),
    .QN(_11192_)
  );
  DFF_X1 \remainder[48]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00069_),
    .Q(remainder[48]),
    .QN(_11191_)
  );
  DFF_X1 \remainder[49]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00070_),
    .Q(remainder[49]),
    .QN(_11190_)
  );
  DFF_X1 \remainder[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00091_),
    .Q(remainder[4]),
    .QN(_11169_)
  );
  DFF_X1 \remainder[50]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00071_),
    .Q(remainder[50]),
    .QN(_11189_)
  );
  DFF_X1 \remainder[51]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00072_),
    .Q(remainder[51]),
    .QN(_11188_)
  );
  DFF_X1 \remainder[52]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00073_),
    .Q(remainder[52]),
    .QN(_11187_)
  );
  DFF_X1 \remainder[53]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00074_),
    .Q(remainder[53]),
    .QN(_11186_)
  );
  DFF_X1 \remainder[54]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00075_),
    .Q(remainder[54]),
    .QN(_11185_)
  );
  DFF_X1 \remainder[55]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00076_),
    .Q(remainder[55]),
    .QN(_11184_)
  );
  DFF_X1 \remainder[56]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00077_),
    .Q(remainder[56]),
    .QN(_11183_)
  );
  DFF_X1 \remainder[57]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00078_),
    .Q(remainder[57]),
    .QN(_11182_)
  );
  DFF_X1 \remainder[58]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00079_),
    .Q(remainder[58]),
    .QN(_11181_)
  );
  DFF_X1 \remainder[59]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00080_),
    .Q(remainder[59]),
    .QN(_11180_)
  );
  DFF_X1 \remainder[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00092_),
    .Q(remainder[5]),
    .QN(_11168_)
  );
  DFF_X1 \remainder[60]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00081_),
    .Q(remainder[60]),
    .QN(_11179_)
  );
  DFF_X1 \remainder[61]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00082_),
    .Q(remainder[61]),
    .QN(_11178_)
  );
  DFF_X1 \remainder[62]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00083_),
    .Q(remainder[62]),
    .QN(_11177_)
  );
  DFF_X1 \remainder[63]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00084_),
    .Q(remainder[63]),
    .QN(_11176_)
  );
  DFF_X1 \remainder[64]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00085_),
    .Q(remainder[64]),
    .QN(_11175_)
  );
  DFF_X1 \remainder[65]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00086_),
    .Q(remainder[65]),
    .QN(_11174_)
  );
  DFF_X1 \remainder[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00093_),
    .Q(remainder[6]),
    .QN(_11167_)
  );
  DFF_X1 \remainder[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00094_),
    .Q(remainder[7]),
    .QN(_11166_)
  );
  DFF_X1 \remainder[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00095_),
    .Q(remainder[8]),
    .QN(_11165_)
  );
  DFF_X1 \remainder[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00096_),
    .Q(remainder[9]),
    .QN(_11164_)
  );
  DFF_X1 \req_tag[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00009_),
    .Q(req_tag[0]),
    .QN(_11215_)
  );
  DFF_X1 \req_tag[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00010_),
    .Q(req_tag[1]),
    .QN(_11214_)
  );
  DFF_X1 \req_tag[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00011_),
    .Q(req_tag[2]),
    .QN(_11213_)
  );
  DFF_X1 \req_tag[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00012_),
    .Q(req_tag[3]),
    .QN(_11212_)
  );
  DFF_X1 \req_tag[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00013_),
    .Q(req_tag[4]),
    .QN(_11211_)
  );
  DFF_X1 \resHi$_SDFF_PP0_  (
    .CK(clock),
    .D(_00005_),
    .Q(resHi),
    .QN(_11216_)
  );
  DFF_X1 \state[0]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00006_),
    .Q(state[0]),
    .QN(_00004_)
  );
  DFF_X1 \state[1]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00007_),
    .Q(state[1]),
    .QN(_00003_)
  );
  DFF_X1 \state[2]$_SDFF_PP0_  (
    .CK(clock),
    .D(_00119_),
    .Q(state[2]),
    .QN(_00000_)
  );
  assign _GEN_0[64:32] = { _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65] };
  assign _GEN_2[64:32] = { _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65] };
  assign _GEN_35 = { remainder[65], remainder[65], remainder[65], remainder[65], remainder[65], remainder[65], remainder[65], remainder[65], remainder[65], remainder[65:33] };
  assign _decoded_T_4[1] = io_req_bits_fn[0];
  assign _decoded_T_6 = io_req_bits_fn[1];
  assign _decoded_T_7[0] = io_req_bits_fn[2];
  assign _decoded_orMatrixOutputs_T_4[0] = io_req_bits_fn[1];
  assign _divisor_T[31:0] = io_req_bits_in2;
  assign _prod_T_2 = { remainder[32], remainder[7:0] };
  assign _remainder_T_2[23:0] = remainder[31:8];
  assign { _state_T[2], _state_T[0] } = 2'h3;
  assign accum = remainder[65:33];
  assign decoded_andMatrixInput_0_3 = io_req_bits_fn[0];
  assign decoded_andMatrixInput_0_4 = io_req_bits_fn[1];
  assign decoded_andMatrixInput_1_2 = io_req_bits_fn[2];
  assign decoded_plaInput = io_req_bits_fn[2:0];
  assign hi = io_req_bits_in1[31:16];
  assign hi_1 = io_req_bits_in2[31:16];
  assign io_resp_bits_tag = req_tag;
  assign lhs_in = io_req_bits_in1;
  assign loOut = io_resp_bits_data[15:0];
  assign mplier = remainder[31:0];
  assign mplierSign = remainder[32];
  assign mulReg = { remainder[65:33], remainder[31:0] };
  assign negated_remainder[0] = io_resp_bits_data[0];
  assign nextMplierSign = _remainder_T_2[32];
  assign nextMulReg[64:0] = { _remainder_T_2[65:33], _remainder_T_2[31:24], remainder[31:8] };
  assign nextMulReg1 = { _remainder_T_2[65:33], _remainder_T_2[31:24], remainder[31:8] };
  assign nextMulReg_hi = { nextMulReg[65], _remainder_T_2[65:33], _remainder_T_2[31:24] };
  assign result = io_resp_bits_data;
  assign rhs_sign = _divisor_T[32];
  assign unrolls_0[32:1] = remainder[31:0];
endmodule
module PlusArgTimeout(clock, reset, io_count);
  input clock;
  wire clock;
  input [31:0] io_count;
  wire [31:0] io_count;
  input reset;
  wire reset;
endmodule
module RVCExpander(io_in, io_out_bits, io_out_rd, io_out_rs1, io_out_rs2, io_rvc);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire [30:0] _GEN_0;
  wire [30:0] _GEN_1;
  wire [31:0] _io_out_T_10_bits;
  wire [4:0] _io_out_T_10_rd;
  wire [4:0] _io_out_T_10_rs1;
  wire [31:0] _io_out_T_12_bits;
  wire [4:0] _io_out_T_12_rd;
  wire [4:0] _io_out_T_12_rs1;
  wire [31:0] _io_out_T_14_bits;
  wire [4:0] _io_out_T_14_rd;
  wire [4:0] _io_out_T_14_rs1;
  wire [31:0] _io_out_T_16_bits;
  wire [4:0] _io_out_T_16_rd;
  wire [4:0] _io_out_T_16_rs1;
  wire [31:0] _io_out_T_18_bits;
  wire [4:0] _io_out_T_18_rd;
  wire [4:0] _io_out_T_18_rs1;
  wire [4:0] _io_out_T_18_rs2;
  wire [4:0] _io_out_T_2;
  wire [31:0] _io_out_T_20_bits;
  wire [4:0] _io_out_T_20_rs2;
  wire [31:0] _io_out_T_22_bits;
  wire [4:0] _io_out_T_22_rs2;
  wire [31:0] _io_out_T_24_bits;
  wire [4:0] _io_out_T_24_rs2;
  wire [31:0] _io_out_T_26_bits;
  wire [4:0] _io_out_T_26_rs2;
  wire [31:0] _io_out_T_28_bits;
  wire [4:0] _io_out_T_28_rs2;
  wire [31:0] _io_out_T_30_bits;
  wire [4:0] _io_out_T_30_rs2;
  wire [31:0] _io_out_T_32_bits;
  wire [4:0] _io_out_T_32_rs2;
  wire [31:0] _io_out_T_34_bits;
  wire [31:0] _io_out_T_36_bits;
  wire [31:0] _io_out_T_38_bits;
  wire [31:0] _io_out_T_40_bits;
  wire [31:0] _io_out_T_42_bits;
  wire [31:0] _io_out_T_44_bits;
  wire [31:0] _io_out_T_46_bits;
  wire [31:0] _io_out_T_48_bits;
  wire [31:0] _io_out_T_4_bits;
  wire [4:0] _io_out_T_4_rd;
  wire [4:0] _io_out_T_4_rs1;
  wire [31:0] _io_out_T_6_bits;
  wire [4:0] _io_out_T_6_rd;
  wire [4:0] _io_out_T_6_rs1;
  wire [31:0] _io_out_T_8_bits;
  wire [4:0] _io_out_T_8_rd;
  wire [4:0] _io_out_T_8_rs1;
  wire [26:0] _io_out_s_T_116;
  wire [26:0] _io_out_s_T_138;
  wire [6:0] _io_out_s_T_148;
  wire [7:0] _io_out_s_T_15;
  wire [11:0] _io_out_s_T_150;
  wire [9:0] _io_out_s_T_161;
  wire [20:0] _io_out_s_T_169;
  wire [4:0] _io_out_s_T_17;
  wire [27:0] _io_out_s_T_20;
  wire [2:0] _io_out_s_T_230;
  wire [25:0] _io_out_s_T_251;
  wire [30:0] _io_out_s_T_260;
  wire [31:0] _io_out_s_T_270;
  wire [24:0] _io_out_s_T_277;
  wire [30:0] _io_out_s_T_278;
  wire [30:0] _io_out_s_T_281;
  wire [31:0] _io_out_s_T_283;
  wire [6:0] _io_out_s_T_31;
  wire [4:0] _io_out_s_T_349;
  wire [12:0] _io_out_s_T_354;
  wire [26:0] _io_out_s_T_36;
  wire [25:0] _io_out_s_T_438;
  wire [28:0] _io_out_s_T_448;
  wire [27:0] _io_out_s_T_457;
  wire [27:0] _io_out_s_T_466;
  wire [8:0] _io_out_s_T_473;
  wire [28:0] _io_out_s_T_480;
  wire [7:0] _io_out_s_T_486;
  wire [27:0] _io_out_s_T_493;
  wire [27:0] _io_out_s_T_506;
  wire [26:0] _io_out_s_T_52;
  wire [4:0] _io_out_s_T_6;
  wire [29:0] _io_out_s_T_7;
  wire [26:0] _io_out_s_T_74;
  wire [27:0] _io_out_s_T_94;
  wire [24:0] _io_out_s_add_T_3;
  wire [24:0] _io_out_s_ebreak_T_1;
  wire [2:0] _io_out_s_funct_T_2;
  wire [2:0] _io_out_s_funct_T_4;
  wire [2:0] _io_out_s_funct_T_6;
  wire [24:0] _io_out_s_jalr_ebreak_T_2;
  wire [24:0] _io_out_s_jr_reserved_T_2;
  wire _io_out_s_load_opc_T_1;
  wire [14:0] _io_out_s_me_T_2;
  wire [31:0] _io_out_s_me_T_4;
  wire [24:0] _io_out_s_mv_T_2;
  input [31:0] io_in;
  wire [31:0] io_in;
  output [31:0] io_out_bits;
  wire [31:0] io_out_bits;
  output [4:0] io_out_rd;
  wire [4:0] io_out_rd;
  output [4:0] io_out_rs1;
  wire [4:0] io_out_rs1;
  output [4:0] io_out_rs2;
  wire [4:0] io_out_rs2;
  wire [31:0] io_out_s_0_bits;
  wire [31:0] io_out_s_10_bits;
  wire [31:0] io_out_s_11_bits;
  wire [4:0] io_out_s_11_rd;
  wire [4:0] io_out_s_11_rs2;
  wire [31:0] io_out_s_12_bits;
  wire [31:0] io_out_s_13_bits;
  wire [31:0] io_out_s_14_bits;
  wire [31:0] io_out_s_15_bits;
  wire [31:0] io_out_s_16_bits;
  wire [31:0] io_out_s_17_bits;
  wire [31:0] io_out_s_18_bits;
  wire [31:0] io_out_s_19_bits;
  wire [31:0] io_out_s_1_bits;
  wire [31:0] io_out_s_20_bits;
  wire [4:0] io_out_s_20_rd;
  wire [4:0] io_out_s_20_rs1;
  wire [4:0] io_out_s_20_rs2;
  wire [31:0] io_out_s_21_bits;
  wire [31:0] io_out_s_22_bits;
  wire [31:0] io_out_s_23_bits;
  wire [4:0] io_out_s_24_rs1;
  wire [4:0] io_out_s_24_rs2;
  wire [31:0] io_out_s_2_bits;
  wire [31:0] io_out_s_3_bits;
  wire [31:0] io_out_s_4_bits;
  wire [31:0] io_out_s_5_bits;
  wire [31:0] io_out_s_6_bits;
  wire [31:0] io_out_s_7_bits;
  wire [31:0] io_out_s_8_bits;
  wire [31:0] io_out_s_9_bits;
  wire [31:0] io_out_s_add_bits;
  wire [24:0] io_out_s_ebreak;
  wire [2:0] io_out_s_funct;
  wire [24:0] io_out_s_jalr;
  wire [31:0] io_out_s_jalr_add_bits;
  wire [4:0] io_out_s_jalr_add_rd;
  wire [4:0] io_out_s_jalr_add_rs1;
  wire [31:0] io_out_s_jalr_ebreak_bits;
  wire [24:0] io_out_s_jr;
  wire [31:0] io_out_s_jr_mv_bits;
  wire [4:0] io_out_s_jr_mv_rd;
  wire [4:0] io_out_s_jr_mv_rs1;
  wire [4:0] io_out_s_jr_mv_rs2;
  wire [31:0] io_out_s_jr_reserved_bits;
  wire [6:0] io_out_s_load_opc;
  wire [31:0] io_out_s_me_bits;
  wire [31:0] io_out_s_mv_bits;
  wire [6:0] io_out_s_opc;
  wire [6:0] io_out_s_opc_1;
  wire [6:0] io_out_s_opc_2;
  wire [6:0] io_out_s_opc_3;
  wire [31:0] io_out_s_res_bits;
  wire [24:0] io_out_s_reserved;
  wire [30:0] io_out_s_sub;
  output io_rvc;
  wire io_rvc;
  INV_X1 _0959_ (
    .A(io_in[6]),
    .ZN(_0769_)
  );
  INV_X1 _0960_ (
    .A(io_in[5]),
    .ZN(_0780_)
  );
  INV_X1 _0961_ (
    .A(io_in[12]),
    .ZN(_0790_)
  );
  INV_X1 _0962_ (
    .A(io_in[8]),
    .ZN(_0801_)
  );
  INV_X1 _0963_ (
    .A(io_in[11]),
    .ZN(_0812_)
  );
  INV_X1 _0964_ (
    .A(io_in[10]),
    .ZN(_0823_)
  );
  INV_X1 _0965_ (
    .A(io_in[0]),
    .ZN(_0833_)
  );
  INV_X1 _0966_ (
    .A(io_in[14]),
    .ZN(_0844_)
  );
  INV_X1 _0967_ (
    .A(io_in[13]),
    .ZN(_0855_)
  );
  INV_X1 _0968_ (
    .A(io_in[1]),
    .ZN(_0865_)
  );
  INV_X1 _0969_ (
    .A(io_in[15]),
    .ZN(_0876_)
  );
  INV_X1 _0970_ (
    .A(io_in[7]),
    .ZN(_0886_)
  );
  INV_X1 _0971_ (
    .A(io_in[9]),
    .ZN(_0896_)
  );
  INV_X1 _0972_ (
    .A(io_in[2]),
    .ZN(_0906_)
  );
  INV_X1 _0973_ (
    .A(io_in[3]),
    .ZN(_0917_)
  );
  INV_X1 _0974_ (
    .A(io_in[4]),
    .ZN(_0928_)
  );
  INV_X1 _0975_ (
    .A(io_in[22]),
    .ZN(_0938_)
  );
  AND2_X1 _0976_ (
    .A1(io_in[0]),
    .A2(io_in[1]),
    .ZN(_0949_)
  );
  INV_X1 _0977_ (
    .A(_0949_),
    .ZN(io_rvc)
  );
  AND2_X1 _0978_ (
    .A1(_0906_),
    .A2(_0949_),
    .ZN(_0010_)
  );
  INV_X1 _0979_ (
    .A(_0010_),
    .ZN(_0020_)
  );
  AND2_X1 _0980_ (
    .A1(_0769_),
    .A2(_0780_),
    .ZN(_0029_)
  );
  INV_X1 _0981_ (
    .A(_0029_),
    .ZN(_0039_)
  );
  AND2_X1 _0982_ (
    .A1(_0906_),
    .A2(_0917_),
    .ZN(_0050_)
  );
  AND2_X1 _0983_ (
    .A1(_0928_),
    .A2(_0050_),
    .ZN(_0059_)
  );
  AND2_X1 _0984_ (
    .A1(_0029_),
    .A2(_0059_),
    .ZN(_0068_)
  );
  INV_X1 _0985_ (
    .A(_0068_),
    .ZN(_0077_)
  );
  AND2_X1 _0986_ (
    .A1(_0790_),
    .A2(_0068_),
    .ZN(_0083_)
  );
  INV_X1 _0987_ (
    .A(_0083_),
    .ZN(_0084_)
  );
  AND2_X1 _0988_ (
    .A1(_0812_),
    .A2(_0823_),
    .ZN(_0085_)
  );
  AND2_X1 _0989_ (
    .A1(_0886_),
    .A2(_0896_),
    .ZN(_0086_)
  );
  AND2_X1 _0990_ (
    .A1(_0085_),
    .A2(_0086_),
    .ZN(_0087_)
  );
  INV_X1 _0991_ (
    .A(_0087_),
    .ZN(_0088_)
  );
  AND2_X1 _0992_ (
    .A1(_0801_),
    .A2(_0087_),
    .ZN(_0089_)
  );
  INV_X1 _0993_ (
    .A(_0089_),
    .ZN(_0090_)
  );
  AND2_X1 _0994_ (
    .A1(_0068_),
    .A2(_0090_),
    .ZN(_0091_)
  );
  INV_X1 _0995_ (
    .A(_0091_),
    .ZN(_0092_)
  );
  AND2_X1 _0996_ (
    .A1(_0844_),
    .A2(_0855_),
    .ZN(_0093_)
  );
  INV_X1 _0997_ (
    .A(_0093_),
    .ZN(_0094_)
  );
  AND2_X1 _0998_ (
    .A1(_0833_),
    .A2(io_in[15]),
    .ZN(_0095_)
  );
  AND2_X1 _0999_ (
    .A1(io_in[1]),
    .A2(_0095_),
    .ZN(_0096_)
  );
  INV_X1 _1000_ (
    .A(_0096_),
    .ZN(_0097_)
  );
  AND2_X1 _1001_ (
    .A1(io_in[1]),
    .A2(_0093_),
    .ZN(_0098_)
  );
  AND2_X1 _1002_ (
    .A1(_0093_),
    .A2(_0096_),
    .ZN(_0099_)
  );
  INV_X1 _1003_ (
    .A(_0099_),
    .ZN(_0100_)
  );
  AND2_X1 _1004_ (
    .A1(_0092_),
    .A2(_0099_),
    .ZN(_0101_)
  );
  INV_X1 _1005_ (
    .A(_0101_),
    .ZN(_0102_)
  );
  AND2_X1 _1006_ (
    .A1(_0084_),
    .A2(_0101_),
    .ZN(_0103_)
  );
  INV_X1 _1007_ (
    .A(_0103_),
    .ZN(_0104_)
  );
  AND2_X1 _1008_ (
    .A1(_0833_),
    .A2(_0876_),
    .ZN(_0105_)
  );
  AND2_X1 _1009_ (
    .A1(io_in[1]),
    .A2(_0105_),
    .ZN(_0106_)
  );
  INV_X1 _1010_ (
    .A(_0106_),
    .ZN(_0107_)
  );
  AND2_X1 _1011_ (
    .A1(io_in[14]),
    .A2(io_in[1]),
    .ZN(_0108_)
  );
  AND2_X1 _1012_ (
    .A1(_0105_),
    .A2(_0108_),
    .ZN(_0109_)
  );
  INV_X1 _1013_ (
    .A(_0109_),
    .ZN(_0110_)
  );
  AND2_X1 _1014_ (
    .A1(io_in[14]),
    .A2(_0855_),
    .ZN(_0111_)
  );
  AND2_X1 _1015_ (
    .A1(_0106_),
    .A2(_0111_),
    .ZN(_0112_)
  );
  INV_X1 _1016_ (
    .A(_0112_),
    .ZN(_0113_)
  );
  AND2_X1 _1017_ (
    .A1(_0865_),
    .A2(_0095_),
    .ZN(_0114_)
  );
  INV_X1 _1018_ (
    .A(_0114_),
    .ZN(_0115_)
  );
  AND2_X1 _1019_ (
    .A1(io_in[14]),
    .A2(_0114_),
    .ZN(_0116_)
  );
  INV_X1 _1020_ (
    .A(_0116_),
    .ZN(_0117_)
  );
  AND2_X1 _1021_ (
    .A1(io_in[14]),
    .A2(io_in[13]),
    .ZN(_0118_)
  );
  AND2_X1 _1022_ (
    .A1(_0114_),
    .A2(_0118_),
    .ZN(_0119_)
  );
  INV_X1 _1023_ (
    .A(_0119_),
    .ZN(_0120_)
  );
  AND2_X1 _1024_ (
    .A1(_0844_),
    .A2(io_in[13]),
    .ZN(_0121_)
  );
  INV_X1 _1025_ (
    .A(_0121_),
    .ZN(_0122_)
  );
  AND2_X1 _1026_ (
    .A1(_0865_),
    .A2(_0121_),
    .ZN(_0123_)
  );
  AND2_X1 _1027_ (
    .A1(_0105_),
    .A2(_0123_),
    .ZN(_0124_)
  );
  INV_X1 _1028_ (
    .A(_0124_),
    .ZN(_0125_)
  );
  AND2_X1 _1029_ (
    .A1(_0790_),
    .A2(_0089_),
    .ZN(_0126_)
  );
  INV_X1 _1030_ (
    .A(_0126_),
    .ZN(_0127_)
  );
  AND2_X1 _1031_ (
    .A1(_0029_),
    .A2(_0126_),
    .ZN(_0128_)
  );
  INV_X1 _1032_ (
    .A(_0128_),
    .ZN(_0129_)
  );
  AND2_X1 _1033_ (
    .A1(_0125_),
    .A2(_0129_),
    .ZN(_0130_)
  );
  INV_X1 _1034_ (
    .A(_0130_),
    .ZN(_0131_)
  );
  AND2_X1 _1035_ (
    .A1(_0865_),
    .A2(_0111_),
    .ZN(_0132_)
  );
  AND2_X1 _1036_ (
    .A1(_0105_),
    .A2(_0132_),
    .ZN(_0133_)
  );
  INV_X1 _1037_ (
    .A(_0133_),
    .ZN(_0134_)
  );
  AND2_X1 _1038_ (
    .A1(_0131_),
    .A2(_0134_),
    .ZN(_0135_)
  );
  INV_X1 _1039_ (
    .A(_0135_),
    .ZN(_0136_)
  );
  AND2_X1 _1040_ (
    .A1(_0105_),
    .A2(_0118_),
    .ZN(_0137_)
  );
  INV_X1 _1041_ (
    .A(_0137_),
    .ZN(_0138_)
  );
  AND2_X1 _1042_ (
    .A1(_0844_),
    .A2(_0095_),
    .ZN(_0139_)
  );
  INV_X1 _1043_ (
    .A(_0139_),
    .ZN(_0140_)
  );
  AND2_X1 _1044_ (
    .A1(_0138_),
    .A2(_0140_),
    .ZN(_0141_)
  );
  INV_X1 _1045_ (
    .A(_0141_),
    .ZN(_0142_)
  );
  AND2_X1 _1046_ (
    .A1(_0865_),
    .A2(_0142_),
    .ZN(_0143_)
  );
  INV_X1 _1047_ (
    .A(_0143_),
    .ZN(_0144_)
  );
  AND2_X1 _1048_ (
    .A1(_0136_),
    .A2(_0144_),
    .ZN(_0145_)
  );
  INV_X1 _1049_ (
    .A(_0145_),
    .ZN(_0146_)
  );
  AND2_X1 _1050_ (
    .A1(_0095_),
    .A2(_0132_),
    .ZN(_0147_)
  );
  INV_X1 _1051_ (
    .A(_0147_),
    .ZN(_0148_)
  );
  MUX2_X1 _1052_ (
    .A(io_in[13]),
    .B(_0146_),
    .S(_0117_),
    .Z(_0149_)
  );
  AND2_X1 _1053_ (
    .A1(_0865_),
    .A2(_0118_),
    .ZN(_0150_)
  );
  AND2_X1 _1054_ (
    .A1(io_in[0]),
    .A2(_0876_),
    .ZN(_0151_)
  );
  AND2_X1 _1055_ (
    .A1(_0150_),
    .A2(_0151_),
    .ZN(_0152_)
  );
  INV_X1 _1056_ (
    .A(_0152_),
    .ZN(_0153_)
  );
  AND2_X1 _1057_ (
    .A1(_0132_),
    .A2(_0151_),
    .ZN(_0154_)
  );
  INV_X1 _1058_ (
    .A(_0154_),
    .ZN(_0155_)
  );
  AND2_X1 _1059_ (
    .A1(_0153_),
    .A2(_0155_),
    .ZN(_0156_)
  );
  AND2_X1 _1060_ (
    .A1(_0865_),
    .A2(_0093_),
    .ZN(_0157_)
  );
  AND2_X1 _1061_ (
    .A1(_0151_),
    .A2(_0157_),
    .ZN(_0158_)
  );
  INV_X1 _1062_ (
    .A(_0158_),
    .ZN(_0159_)
  );
  AND2_X1 _1063_ (
    .A1(_0156_),
    .A2(_0159_),
    .ZN(_0160_)
  );
  INV_X1 _1064_ (
    .A(_0160_),
    .ZN(_0161_)
  );
  AND2_X1 _1065_ (
    .A1(_0149_),
    .A2(_0160_),
    .ZN(_0162_)
  );
  INV_X1 _1066_ (
    .A(_0162_),
    .ZN(_0163_)
  );
  AND2_X1 _1067_ (
    .A1(_0088_),
    .A2(_0152_),
    .ZN(_0164_)
  );
  INV_X1 _1068_ (
    .A(_0164_),
    .ZN(_0165_)
  );
  AND2_X1 _1069_ (
    .A1(_0083_),
    .A2(_0152_),
    .ZN(_0166_)
  );
  INV_X1 _1070_ (
    .A(_0166_),
    .ZN(_0167_)
  );
  AND2_X1 _1071_ (
    .A1(io_in[0]),
    .A2(_0123_),
    .ZN(_0168_)
  );
  INV_X1 _1072_ (
    .A(_0168_),
    .ZN(_0169_)
  );
  AND2_X1 _1073_ (
    .A1(_0123_),
    .A2(_0151_),
    .ZN(_0170_)
  );
  INV_X1 _1074_ (
    .A(_0170_),
    .ZN(_0171_)
  );
  AND2_X1 _1075_ (
    .A1(_0167_),
    .A2(_0171_),
    .ZN(_0172_)
  );
  AND2_X1 _1076_ (
    .A1(_0165_),
    .A2(_0172_),
    .ZN(_0173_)
  );
  AND2_X1 _1077_ (
    .A1(_0163_),
    .A2(_0173_),
    .ZN(_0174_)
  );
  INV_X1 _1078_ (
    .A(_0174_),
    .ZN(_0175_)
  );
  AND2_X1 _1079_ (
    .A1(_0093_),
    .A2(_0106_),
    .ZN(_0176_)
  );
  INV_X1 _1080_ (
    .A(_0176_),
    .ZN(_0177_)
  );
  AND2_X1 _1081_ (
    .A1(io_in[0]),
    .A2(_0865_),
    .ZN(_0178_)
  );
  AND2_X1 _1082_ (
    .A1(io_in[15]),
    .A2(_0178_),
    .ZN(_0179_)
  );
  INV_X1 _1083_ (
    .A(_0179_),
    .ZN(_0180_)
  );
  AND2_X1 _1084_ (
    .A1(io_in[0]),
    .A2(io_in[15]),
    .ZN(_0181_)
  );
  AND2_X1 _1085_ (
    .A1(_0111_),
    .A2(_0179_),
    .ZN(_0182_)
  );
  INV_X1 _1086_ (
    .A(_0182_),
    .ZN(_0183_)
  );
  AND2_X1 _1087_ (
    .A1(_0150_),
    .A2(_0181_),
    .ZN(_0184_)
  );
  INV_X1 _1088_ (
    .A(_0184_),
    .ZN(_0185_)
  );
  AND2_X1 _1089_ (
    .A1(_0183_),
    .A2(_0185_),
    .ZN(_0186_)
  );
  AND2_X1 _1090_ (
    .A1(io_in[14]),
    .A2(_0179_),
    .ZN(_0187_)
  );
  AND2_X1 _1091_ (
    .A1(_0093_),
    .A2(_0179_),
    .ZN(_0188_)
  );
  INV_X1 _1092_ (
    .A(_0188_),
    .ZN(_0189_)
  );
  AND2_X1 _1093_ (
    .A1(_0186_),
    .A2(_0189_),
    .ZN(_0190_)
  );
  AND2_X1 _1094_ (
    .A1(_0177_),
    .A2(_0189_),
    .ZN(_0191_)
  );
  AND2_X1 _1095_ (
    .A1(_0177_),
    .A2(_0186_),
    .ZN(_0192_)
  );
  INV_X1 _1096_ (
    .A(_0192_),
    .ZN(_0193_)
  );
  AND2_X1 _1097_ (
    .A1(_0186_),
    .A2(_0191_),
    .ZN(_0194_)
  );
  INV_X1 _1098_ (
    .A(_0194_),
    .ZN(_0195_)
  );
  AND2_X1 _1099_ (
    .A1(_0175_),
    .A2(_0194_),
    .ZN(_0196_)
  );
  INV_X1 _1100_ (
    .A(_0196_),
    .ZN(_0197_)
  );
  AND2_X1 _1101_ (
    .A1(_0844_),
    .A2(_0106_),
    .ZN(_0198_)
  );
  INV_X1 _1102_ (
    .A(_0198_),
    .ZN(_0199_)
  );
  AND2_X1 _1103_ (
    .A1(_0106_),
    .A2(_0121_),
    .ZN(_0200_)
  );
  INV_X1 _1104_ (
    .A(_0200_),
    .ZN(_0201_)
  );
  AND2_X1 _1105_ (
    .A1(_0121_),
    .A2(_0181_),
    .ZN(_0202_)
  );
  AND2_X1 _1106_ (
    .A1(_0121_),
    .A2(_0179_),
    .ZN(_0203_)
  );
  INV_X1 _1107_ (
    .A(_0203_),
    .ZN(_0204_)
  );
  AND2_X1 _1108_ (
    .A1(_0201_),
    .A2(_0204_),
    .ZN(_0205_)
  );
  AND2_X1 _1109_ (
    .A1(_0197_),
    .A2(_0205_),
    .ZN(_0206_)
  );
  AND2_X1 _1110_ (
    .A1(_0106_),
    .A2(_0118_),
    .ZN(_0207_)
  );
  INV_X1 _1111_ (
    .A(_0207_),
    .ZN(_0208_)
  );
  AND2_X1 _1112_ (
    .A1(_0100_),
    .A2(_0208_),
    .ZN(_0209_)
  );
  AND2_X1 _1113_ (
    .A1(_0089_),
    .A2(_0112_),
    .ZN(_0210_)
  );
  INV_X1 _1114_ (
    .A(_0210_),
    .ZN(_0211_)
  );
  MUX2_X1 _1115_ (
    .A(_0090_),
    .B(_0206_),
    .S(_0113_),
    .Z(_0212_)
  );
  AND2_X1 _1116_ (
    .A1(_0209_),
    .A2(_0212_),
    .ZN(_0213_)
  );
  INV_X1 _1117_ (
    .A(_0213_),
    .ZN(_0214_)
  );
  AND2_X1 _1118_ (
    .A1(_0104_),
    .A2(_0214_),
    .ZN(_0215_)
  );
  INV_X1 _1119_ (
    .A(_0215_),
    .ZN(_0216_)
  );
  AND2_X1 _1120_ (
    .A1(_0095_),
    .A2(_0121_),
    .ZN(_0217_)
  );
  INV_X1 _1121_ (
    .A(_0217_),
    .ZN(_0218_)
  );
  AND2_X1 _1122_ (
    .A1(_0096_),
    .A2(_0121_),
    .ZN(_0219_)
  );
  INV_X1 _1123_ (
    .A(_0219_),
    .ZN(_0220_)
  );
  AND2_X1 _1124_ (
    .A1(_0216_),
    .A2(_0220_),
    .ZN(_0221_)
  );
  INV_X1 _1125_ (
    .A(_0221_),
    .ZN(_0222_)
  );
  AND2_X1 _1126_ (
    .A1(_0096_),
    .A2(_0111_),
    .ZN(_0223_)
  );
  INV_X1 _1127_ (
    .A(_0223_),
    .ZN(_0224_)
  );
  AND2_X1 _1128_ (
    .A1(_0222_),
    .A2(_0224_),
    .ZN(_0225_)
  );
  INV_X1 _1129_ (
    .A(_0225_),
    .ZN(_0226_)
  );
  AND2_X1 _1130_ (
    .A1(_0096_),
    .A2(_0118_),
    .ZN(_0227_)
  );
  INV_X1 _1131_ (
    .A(_0227_),
    .ZN(_0228_)
  );
  AND2_X1 _1132_ (
    .A1(io_rvc),
    .A2(_0228_),
    .ZN(_0229_)
  );
  AND2_X1 _1133_ (
    .A1(_0226_),
    .A2(_0229_),
    .ZN(_0230_)
  );
  INV_X1 _1134_ (
    .A(_0230_),
    .ZN(_0231_)
  );
  AND2_X1 _1135_ (
    .A1(_0020_),
    .A2(_0231_),
    .ZN(io_out_bits[2])
  );
  AND2_X1 _1136_ (
    .A1(io_in[3]),
    .A2(_0949_),
    .ZN(_0232_)
  );
  INV_X1 _1137_ (
    .A(_0232_),
    .ZN(_0233_)
  );
  AND2_X1 _1138_ (
    .A1(_0107_),
    .A2(_0185_),
    .ZN(_0234_)
  );
  AND2_X1 _1139_ (
    .A1(_0183_),
    .A2(_0234_),
    .ZN(_0235_)
  );
  AND2_X1 _1140_ (
    .A1(_0094_),
    .A2(_0105_),
    .ZN(_0236_)
  );
  AND2_X1 _1141_ (
    .A1(_0865_),
    .A2(_0236_),
    .ZN(_0237_)
  );
  INV_X1 _1142_ (
    .A(_0237_),
    .ZN(_0238_)
  );
  AND2_X1 _1143_ (
    .A1(_0128_),
    .A2(_0238_),
    .ZN(_0239_)
  );
  INV_X1 _1144_ (
    .A(_0239_),
    .ZN(_0240_)
  );
  AND2_X1 _1145_ (
    .A1(_0093_),
    .A2(_0114_),
    .ZN(_0241_)
  );
  INV_X1 _1146_ (
    .A(_0241_),
    .ZN(_0242_)
  );
  AND2_X1 _1147_ (
    .A1(_0240_),
    .A2(_0242_),
    .ZN(_0243_)
  );
  INV_X1 _1148_ (
    .A(_0243_),
    .ZN(_0244_)
  );
  AND2_X1 _1149_ (
    .A1(_0865_),
    .A2(_0217_),
    .ZN(_0245_)
  );
  INV_X1 _1150_ (
    .A(_0245_),
    .ZN(_0246_)
  );
  AND2_X1 _1151_ (
    .A1(_0117_),
    .A2(_0246_),
    .ZN(_0247_)
  );
  AND2_X1 _1152_ (
    .A1(_0160_),
    .A2(_0247_),
    .ZN(_0248_)
  );
  AND2_X1 _1153_ (
    .A1(_0117_),
    .A2(_0159_),
    .ZN(_0249_)
  );
  AND2_X1 _1154_ (
    .A1(_0244_),
    .A2(_0248_),
    .ZN(_0250_)
  );
  INV_X1 _1155_ (
    .A(_0250_),
    .ZN(_0251_)
  );
  AND2_X1 _1156_ (
    .A1(_0172_),
    .A2(_0251_),
    .ZN(_0252_)
  );
  INV_X1 _1157_ (
    .A(_0252_),
    .ZN(_0253_)
  );
  AND2_X1 _1158_ (
    .A1(_0189_),
    .A2(_0253_),
    .ZN(_0254_)
  );
  INV_X1 _1159_ (
    .A(_0254_),
    .ZN(_0255_)
  );
  AND2_X1 _1160_ (
    .A1(io_in[11]),
    .A2(io_in[10]),
    .ZN(_0256_)
  );
  INV_X1 _1161_ (
    .A(_0256_),
    .ZN(_0257_)
  );
  AND2_X1 _1162_ (
    .A1(_0188_),
    .A2(_0256_),
    .ZN(_0258_)
  );
  INV_X1 _1163_ (
    .A(_0258_),
    .ZN(_0259_)
  );
  AND2_X1 _1164_ (
    .A1(io_in[12]),
    .A2(_0258_),
    .ZN(_0260_)
  );
  INV_X1 _1165_ (
    .A(_0260_),
    .ZN(_0261_)
  );
  AND2_X1 _1166_ (
    .A1(_0204_),
    .A2(_0261_),
    .ZN(_0262_)
  );
  AND2_X1 _1167_ (
    .A1(_0255_),
    .A2(_0262_),
    .ZN(_0263_)
  );
  INV_X1 _1168_ (
    .A(_0263_),
    .ZN(_0264_)
  );
  AND2_X1 _1169_ (
    .A1(_0235_),
    .A2(_0264_),
    .ZN(_0265_)
  );
  INV_X1 _1170_ (
    .A(_0265_),
    .ZN(_0266_)
  );
  AND2_X1 _1171_ (
    .A1(_0100_),
    .A2(_0211_),
    .ZN(_0267_)
  );
  AND2_X1 _1172_ (
    .A1(_0266_),
    .A2(_0267_),
    .ZN(_0268_)
  );
  INV_X1 _1173_ (
    .A(_0268_),
    .ZN(_0269_)
  );
  AND2_X1 _1174_ (
    .A1(_0089_),
    .A2(_0093_),
    .ZN(_0270_)
  );
  AND2_X1 _1175_ (
    .A1(_0068_),
    .A2(_0089_),
    .ZN(_0271_)
  );
  AND2_X1 _1176_ (
    .A1(_0083_),
    .A2(_0270_),
    .ZN(_0272_)
  );
  INV_X1 _1177_ (
    .A(_0272_),
    .ZN(_0273_)
  );
  AND2_X1 _1178_ (
    .A1(_0096_),
    .A2(_0273_),
    .ZN(_0274_)
  );
  INV_X1 _1179_ (
    .A(_0274_),
    .ZN(_0275_)
  );
  AND2_X1 _1180_ (
    .A1(io_rvc),
    .A2(_0275_),
    .ZN(_0276_)
  );
  AND2_X1 _1181_ (
    .A1(_0269_),
    .A2(_0276_),
    .ZN(_0277_)
  );
  INV_X1 _1182_ (
    .A(_0277_),
    .ZN(_0278_)
  );
  AND2_X1 _1183_ (
    .A1(_0233_),
    .A2(_0278_),
    .ZN(_0279_)
  );
  INV_X1 _1184_ (
    .A(_0279_),
    .ZN(io_out_bits[3])
  );
  AND2_X1 _1185_ (
    .A1(io_in[4]),
    .A2(_0949_),
    .ZN(_0280_)
  );
  INV_X1 _1186_ (
    .A(_0280_),
    .ZN(_0281_)
  );
  AND2_X1 _1187_ (
    .A1(io_in[1]),
    .A2(_0094_),
    .ZN(_0282_)
  );
  AND2_X1 _1188_ (
    .A1(_0094_),
    .A2(_0096_),
    .ZN(_0283_)
  );
  INV_X1 _1189_ (
    .A(_0283_),
    .ZN(_0284_)
  );
  AND2_X1 _1190_ (
    .A1(io_in[1]),
    .A2(_0202_),
    .ZN(_0285_)
  );
  INV_X1 _1191_ (
    .A(_0285_),
    .ZN(_0286_)
  );
  AND2_X1 _1192_ (
    .A1(_0098_),
    .A2(_0181_),
    .ZN(_0287_)
  );
  INV_X1 _1193_ (
    .A(_0287_),
    .ZN(_0288_)
  );
  AND2_X1 _1194_ (
    .A1(_0286_),
    .A2(_0288_),
    .ZN(_0289_)
  );
  AND2_X1 _1195_ (
    .A1(_0108_),
    .A2(_0181_),
    .ZN(_0290_)
  );
  AND2_X1 _1196_ (
    .A1(io_in[15]),
    .A2(_0949_),
    .ZN(_0291_)
  );
  INV_X1 _1197_ (
    .A(_0291_),
    .ZN(_0292_)
  );
  AND2_X1 _1198_ (
    .A1(_0098_),
    .A2(_0151_),
    .ZN(_0293_)
  );
  INV_X1 _1199_ (
    .A(_0293_),
    .ZN(_0294_)
  );
  AND2_X1 _1200_ (
    .A1(_0876_),
    .A2(_0949_),
    .ZN(_0295_)
  );
  INV_X1 _1201_ (
    .A(_0295_),
    .ZN(_0296_)
  );
  AND2_X1 _1202_ (
    .A1(io_rvc),
    .A2(_0284_),
    .ZN(_0297_)
  );
  INV_X1 _1203_ (
    .A(_0297_),
    .ZN(_0298_)
  );
  AND2_X1 _1204_ (
    .A1(_0115_),
    .A2(_0238_),
    .ZN(_0299_)
  );
  INV_X1 _1205_ (
    .A(_0299_),
    .ZN(_0300_)
  );
  AND2_X1 _1206_ (
    .A1(_0148_),
    .A2(_0238_),
    .ZN(_0301_)
  );
  AND2_X1 _1207_ (
    .A1(_0246_),
    .A2(_0301_),
    .ZN(_0302_)
  );
  AND2_X1 _1208_ (
    .A1(_0120_),
    .A2(_0302_),
    .ZN(_0303_)
  );
  AND2_X1 _1209_ (
    .A1(_0183_),
    .A2(_0204_),
    .ZN(_0304_)
  );
  AND2_X1 _1210_ (
    .A1(_0186_),
    .A2(_0204_),
    .ZN(_0305_)
  );
  INV_X1 _1211_ (
    .A(_0305_),
    .ZN(_0306_)
  );
  AND2_X1 _1212_ (
    .A1(_0169_),
    .A2(_0186_),
    .ZN(_0307_)
  );
  AND2_X1 _1213_ (
    .A1(_0094_),
    .A2(_0106_),
    .ZN(_0308_)
  );
  INV_X1 _1214_ (
    .A(_0308_),
    .ZN(_0309_)
  );
  AND2_X1 _1215_ (
    .A1(_0113_),
    .A2(_0303_),
    .ZN(_0310_)
  );
  AND2_X1 _1216_ (
    .A1(_0307_),
    .A2(_0310_),
    .ZN(_0311_)
  );
  AND2_X1 _1217_ (
    .A1(_0201_),
    .A2(_0311_),
    .ZN(_0312_)
  );
  INV_X1 _1218_ (
    .A(_0312_),
    .ZN(_0313_)
  );
  AND2_X1 _1219_ (
    .A1(_0211_),
    .A2(_0313_),
    .ZN(_0314_)
  );
  INV_X1 _1220_ (
    .A(_0314_),
    .ZN(_0315_)
  );
  AND2_X1 _1221_ (
    .A1(_0209_),
    .A2(_0315_),
    .ZN(_0316_)
  );
  INV_X1 _1222_ (
    .A(_0316_),
    .ZN(_0317_)
  );
  AND2_X1 _1223_ (
    .A1(_0102_),
    .A2(_0317_),
    .ZN(_0318_)
  );
  INV_X1 _1224_ (
    .A(_0318_),
    .ZN(_0319_)
  );
  AND2_X1 _1225_ (
    .A1(_0297_),
    .A2(_0319_),
    .ZN(_0320_)
  );
  INV_X1 _1226_ (
    .A(_0320_),
    .ZN(_0321_)
  );
  AND2_X1 _1227_ (
    .A1(_0281_),
    .A2(_0321_),
    .ZN(_0322_)
  );
  INV_X1 _1228_ (
    .A(_0322_),
    .ZN(io_out_bits[4])
  );
  AND2_X1 _1229_ (
    .A1(_0259_),
    .A2(_0307_),
    .ZN(_0323_)
  );
  AND2_X1 _1230_ (
    .A1(io_in[5]),
    .A2(_0949_),
    .ZN(_0324_)
  );
  INV_X1 _1231_ (
    .A(_0324_),
    .ZN(_0325_)
  );
  AND2_X1 _1232_ (
    .A1(_0115_),
    .A2(_0325_),
    .ZN(_0326_)
  );
  AND2_X1 _1233_ (
    .A1(_0165_),
    .A2(_0326_),
    .ZN(_0327_)
  );
  AND2_X1 _1234_ (
    .A1(_0323_),
    .A2(_0327_),
    .ZN(_0328_)
  );
  AND2_X1 _1235_ (
    .A1(_0275_),
    .A2(_0328_),
    .ZN(_0329_)
  );
  INV_X1 _1236_ (
    .A(_0329_),
    .ZN(io_out_bits[5])
  );
  AND2_X1 _1237_ (
    .A1(_0068_),
    .A2(_0099_),
    .ZN(_0330_)
  );
  INV_X1 _1238_ (
    .A(_0330_),
    .ZN(_0331_)
  );
  AND2_X1 _1239_ (
    .A1(_0127_),
    .A2(_0330_),
    .ZN(_0332_)
  );
  INV_X1 _1240_ (
    .A(_0332_),
    .ZN(_0333_)
  );
  AND2_X1 _1241_ (
    .A1(io_in[6]),
    .A2(_0949_),
    .ZN(_0334_)
  );
  INV_X1 _1242_ (
    .A(_0334_),
    .ZN(_0335_)
  );
  AND2_X1 _1243_ (
    .A1(_0307_),
    .A2(_0335_),
    .ZN(_0336_)
  );
  AND2_X1 _1244_ (
    .A1(_0333_),
    .A2(_0336_),
    .ZN(_0337_)
  );
  INV_X1 _1245_ (
    .A(_0337_),
    .ZN(io_out_bits[6])
  );
  AND2_X1 _1246_ (
    .A1(io_in[7]),
    .A2(_0949_),
    .ZN(_0338_)
  );
  INV_X1 _1247_ (
    .A(_0338_),
    .ZN(_0339_)
  );
  AND2_X1 _1248_ (
    .A1(io_in[7]),
    .A2(_0158_),
    .ZN(_0340_)
  );
  INV_X1 _1249_ (
    .A(_0340_),
    .ZN(_0341_)
  );
  AND2_X1 _1250_ (
    .A1(_0171_),
    .A2(_0341_),
    .ZN(_0342_)
  );
  AND2_X1 _1251_ (
    .A1(_0115_),
    .A2(_0159_),
    .ZN(_0343_)
  );
  AND2_X1 _1252_ (
    .A1(io_in[2]),
    .A2(_0343_),
    .ZN(_0344_)
  );
  INV_X1 _1253_ (
    .A(_0344_),
    .ZN(_0345_)
  );
  AND2_X1 _1254_ (
    .A1(_0342_),
    .A2(_0345_),
    .ZN(_0346_)
  );
  INV_X1 _1255_ (
    .A(_0346_),
    .ZN(_0347_)
  );
  AND2_X1 _1256_ (
    .A1(_0156_),
    .A2(_0189_),
    .ZN(_0348_)
  );
  INV_X1 _1257_ (
    .A(_0348_),
    .ZN(_0349_)
  );
  MUX2_X1 _1258_ (
    .A(io_in[7]),
    .B(_0347_),
    .S(_0348_),
    .Z(_0350_)
  );
  AND2_X1 _1259_ (
    .A1(_0305_),
    .A2(_0350_),
    .ZN(_0351_)
  );
  INV_X1 _1260_ (
    .A(_0351_),
    .ZN(_0352_)
  );
  AND2_X1 _1261_ (
    .A1(io_in[12]),
    .A2(_0187_),
    .ZN(_0353_)
  );
  INV_X1 _1262_ (
    .A(_0353_),
    .ZN(_0354_)
  );
  AND2_X1 _1263_ (
    .A1(_0352_),
    .A2(_0354_),
    .ZN(_0355_)
  );
  INV_X1 _1264_ (
    .A(_0355_),
    .ZN(_0356_)
  );
  AND2_X1 _1265_ (
    .A1(_0107_),
    .A2(_0356_),
    .ZN(_0357_)
  );
  INV_X1 _1266_ (
    .A(_0357_),
    .ZN(_0358_)
  );
  AND2_X1 _1267_ (
    .A1(io_in[7]),
    .A2(_0106_),
    .ZN(_0359_)
  );
  INV_X1 _1268_ (
    .A(_0359_),
    .ZN(_0360_)
  );
  AND2_X1 _1269_ (
    .A1(_0100_),
    .A2(_0360_),
    .ZN(_0361_)
  );
  AND2_X1 _1270_ (
    .A1(_0358_),
    .A2(_0361_),
    .ZN(_0362_)
  );
  INV_X1 _1271_ (
    .A(_0362_),
    .ZN(_0363_)
  );
  AND2_X1 _1272_ (
    .A1(io_in[12]),
    .A2(_0091_),
    .ZN(_0364_)
  );
  INV_X1 _1273_ (
    .A(_0364_),
    .ZN(_0365_)
  );
  AND2_X1 _1274_ (
    .A1(io_in[7]),
    .A2(_0077_),
    .ZN(_0366_)
  );
  INV_X1 _1275_ (
    .A(_0366_),
    .ZN(_0367_)
  );
  AND2_X1 _1276_ (
    .A1(_0099_),
    .A2(_0367_),
    .ZN(_0368_)
  );
  AND2_X1 _1277_ (
    .A1(_0365_),
    .A2(_0368_),
    .ZN(_0369_)
  );
  INV_X1 _1278_ (
    .A(_0369_),
    .ZN(_0370_)
  );
  AND2_X1 _1279_ (
    .A1(_0297_),
    .A2(_0370_),
    .ZN(_0371_)
  );
  AND2_X1 _1280_ (
    .A1(_0363_),
    .A2(_0371_),
    .ZN(_0372_)
  );
  INV_X1 _1281_ (
    .A(_0372_),
    .ZN(_0373_)
  );
  AND2_X1 _1282_ (
    .A1(_0339_),
    .A2(_0373_),
    .ZN(_0374_)
  );
  INV_X1 _1283_ (
    .A(_0374_),
    .ZN(io_out_bits[7])
  );
  AND2_X1 _1284_ (
    .A1(io_in[8]),
    .A2(_0949_),
    .ZN(_0375_)
  );
  INV_X1 _1285_ (
    .A(_0375_),
    .ZN(_0376_)
  );
  AND2_X1 _1286_ (
    .A1(_0077_),
    .A2(_0099_),
    .ZN(_0377_)
  );
  INV_X1 _1287_ (
    .A(_0377_),
    .ZN(_0378_)
  );
  AND2_X1 _1288_ (
    .A1(io_in[8]),
    .A2(_0377_),
    .ZN(_0379_)
  );
  INV_X1 _1289_ (
    .A(_0379_),
    .ZN(_0380_)
  );
  AND2_X1 _1290_ (
    .A1(io_in[8]),
    .A2(_0106_),
    .ZN(_0381_)
  );
  INV_X1 _1291_ (
    .A(_0381_),
    .ZN(_0382_)
  );
  AND2_X1 _1292_ (
    .A1(io_in[8]),
    .A2(_0349_),
    .ZN(_0383_)
  );
  INV_X1 _1293_ (
    .A(_0383_),
    .ZN(_0384_)
  );
  AND2_X1 _1294_ (
    .A1(io_in[8]),
    .A2(_0158_),
    .ZN(_0385_)
  );
  INV_X1 _1295_ (
    .A(_0385_),
    .ZN(_0386_)
  );
  AND2_X1 _1296_ (
    .A1(io_in[3]),
    .A2(_0343_),
    .ZN(_0387_)
  );
  INV_X1 _1297_ (
    .A(_0387_),
    .ZN(_0388_)
  );
  AND2_X1 _1298_ (
    .A1(_0386_),
    .A2(_0388_),
    .ZN(_0389_)
  );
  INV_X1 _1299_ (
    .A(_0389_),
    .ZN(_0390_)
  );
  AND2_X1 _1300_ (
    .A1(_0171_),
    .A2(_0348_),
    .ZN(_0391_)
  );
  AND2_X1 _1301_ (
    .A1(_0153_),
    .A2(_0171_),
    .ZN(_0392_)
  );
  INV_X1 _1302_ (
    .A(_0392_),
    .ZN(_0393_)
  );
  AND2_X1 _1303_ (
    .A1(_0390_),
    .A2(_0391_),
    .ZN(_0394_)
  );
  INV_X1 _1304_ (
    .A(_0394_),
    .ZN(_0395_)
  );
  AND2_X1 _1305_ (
    .A1(_0384_),
    .A2(_0395_),
    .ZN(_0396_)
  );
  INV_X1 _1306_ (
    .A(_0396_),
    .ZN(_0397_)
  );
  AND2_X1 _1307_ (
    .A1(_0107_),
    .A2(_0204_),
    .ZN(_0398_)
  );
  AND2_X1 _1308_ (
    .A1(_0397_),
    .A2(_0398_),
    .ZN(_0399_)
  );
  INV_X1 _1309_ (
    .A(_0399_),
    .ZN(_0400_)
  );
  AND2_X1 _1310_ (
    .A1(_0382_),
    .A2(_0400_),
    .ZN(_0401_)
  );
  INV_X1 _1311_ (
    .A(_0401_),
    .ZN(_0402_)
  );
  AND2_X1 _1312_ (
    .A1(_0100_),
    .A2(_0402_),
    .ZN(_0403_)
  );
  INV_X1 _1313_ (
    .A(_0403_),
    .ZN(_0404_)
  );
  AND2_X1 _1314_ (
    .A1(_0380_),
    .A2(_0404_),
    .ZN(_0405_)
  );
  INV_X1 _1315_ (
    .A(_0405_),
    .ZN(_0406_)
  );
  AND2_X1 _1316_ (
    .A1(_0297_),
    .A2(_0406_),
    .ZN(_0407_)
  );
  INV_X1 _1317_ (
    .A(_0407_),
    .ZN(_0408_)
  );
  AND2_X1 _1318_ (
    .A1(_0376_),
    .A2(_0408_),
    .ZN(_0409_)
  );
  INV_X1 _1319_ (
    .A(_0409_),
    .ZN(io_out_bits[8])
  );
  AND2_X1 _1320_ (
    .A1(io_in[9]),
    .A2(_0106_),
    .ZN(_0410_)
  );
  INV_X1 _1321_ (
    .A(_0410_),
    .ZN(_0411_)
  );
  AND2_X1 _1322_ (
    .A1(io_in[9]),
    .A2(_0349_),
    .ZN(_0412_)
  );
  INV_X1 _1323_ (
    .A(_0412_),
    .ZN(_0413_)
  );
  AND2_X1 _1324_ (
    .A1(_0769_),
    .A2(_0122_),
    .ZN(_0414_)
  );
  INV_X1 _1325_ (
    .A(_0414_),
    .ZN(_0415_)
  );
  MUX2_X1 _1326_ (
    .A(io_in[4]),
    .B(_0415_),
    .S(_0114_),
    .Z(_0416_)
  );
  AND2_X1 _1327_ (
    .A1(_0246_),
    .A2(_0416_),
    .ZN(_0417_)
  );
  MUX2_X1 _1328_ (
    .A(io_in[9]),
    .B(_0417_),
    .S(_0159_),
    .Z(_0418_)
  );
  AND2_X1 _1329_ (
    .A1(_0391_),
    .A2(_0418_),
    .ZN(_0419_)
  );
  INV_X1 _1330_ (
    .A(_0419_),
    .ZN(_0420_)
  );
  AND2_X1 _1331_ (
    .A1(_0413_),
    .A2(_0420_),
    .ZN(_0421_)
  );
  INV_X1 _1332_ (
    .A(_0421_),
    .ZN(_0422_)
  );
  AND2_X1 _1333_ (
    .A1(_0398_),
    .A2(_0422_),
    .ZN(_0423_)
  );
  INV_X1 _1334_ (
    .A(_0423_),
    .ZN(_0424_)
  );
  AND2_X1 _1335_ (
    .A1(_0411_),
    .A2(_0424_),
    .ZN(_0425_)
  );
  INV_X1 _1336_ (
    .A(_0425_),
    .ZN(_0426_)
  );
  AND2_X1 _1337_ (
    .A1(io_rvc),
    .A2(_0097_),
    .ZN(_0427_)
  );
  AND2_X1 _1338_ (
    .A1(_0426_),
    .A2(_0427_),
    .ZN(_0428_)
  );
  INV_X1 _1339_ (
    .A(_0428_),
    .ZN(_0429_)
  );
  AND2_X1 _1340_ (
    .A1(io_in[15]),
    .A2(_0108_),
    .ZN(_0430_)
  );
  INV_X1 _1341_ (
    .A(_0430_),
    .ZN(_0431_)
  );
  AND2_X1 _1342_ (
    .A1(io_rvc),
    .A2(_0431_),
    .ZN(_0432_)
  );
  AND2_X1 _1343_ (
    .A1(_0378_),
    .A2(_0432_),
    .ZN(_0433_)
  );
  INV_X1 _1344_ (
    .A(_0433_),
    .ZN(_0434_)
  );
  AND2_X1 _1345_ (
    .A1(io_in[9]),
    .A2(_0434_),
    .ZN(_0435_)
  );
  INV_X1 _1346_ (
    .A(_0435_),
    .ZN(_0436_)
  );
  AND2_X1 _1347_ (
    .A1(_0429_),
    .A2(_0436_),
    .ZN(_0437_)
  );
  INV_X1 _1348_ (
    .A(_0437_),
    .ZN(io_out_bits[9])
  );
  AND2_X1 _1349_ (
    .A1(_0155_),
    .A2(_0343_),
    .ZN(_0438_)
  );
  AND2_X1 _1350_ (
    .A1(_0235_),
    .A2(_0438_),
    .ZN(_0439_)
  );
  AND2_X1 _1351_ (
    .A1(_0297_),
    .A2(_0439_),
    .ZN(_0440_)
  );
  INV_X1 _1352_ (
    .A(_0440_),
    .ZN(_0441_)
  );
  AND2_X1 _1353_ (
    .A1(_0823_),
    .A2(_0441_),
    .ZN(_0442_)
  );
  INV_X1 _1354_ (
    .A(_0442_),
    .ZN(_0443_)
  );
  MUX2_X1 _1355_ (
    .A(io_in[10]),
    .B(_0171_),
    .S(_0153_),
    .Z(_0444_)
  );
  AND2_X1 _1356_ (
    .A1(_0204_),
    .A2(_0444_),
    .ZN(_0445_)
  );
  AND2_X1 _1357_ (
    .A1(_0100_),
    .A2(_0445_),
    .ZN(_0446_)
  );
  INV_X1 _1358_ (
    .A(_0446_),
    .ZN(_0447_)
  );
  AND2_X1 _1359_ (
    .A1(io_in[10]),
    .A2(_0377_),
    .ZN(_0448_)
  );
  INV_X1 _1360_ (
    .A(_0448_),
    .ZN(_0449_)
  );
  AND2_X1 _1361_ (
    .A1(_0447_),
    .A2(_0449_),
    .ZN(_0450_)
  );
  INV_X1 _1362_ (
    .A(_0450_),
    .ZN(_0451_)
  );
  AND2_X1 _1363_ (
    .A1(_0443_),
    .A2(_0451_),
    .ZN(io_out_bits[10])
  );
  AND2_X1 _1364_ (
    .A1(_0156_),
    .A2(_0343_),
    .ZN(_0452_)
  );
  AND2_X1 _1365_ (
    .A1(_0297_),
    .A2(_0378_),
    .ZN(_0453_)
  );
  INV_X1 _1366_ (
    .A(_0453_),
    .ZN(_0454_)
  );
  AND2_X1 _1367_ (
    .A1(_0235_),
    .A2(_0453_),
    .ZN(_0455_)
  );
  AND2_X1 _1368_ (
    .A1(_0452_),
    .A2(_0455_),
    .ZN(_0456_)
  );
  INV_X1 _1369_ (
    .A(_0456_),
    .ZN(_0457_)
  );
  AND2_X1 _1370_ (
    .A1(io_in[11]),
    .A2(_0457_),
    .ZN(io_out_bits[11])
  );
  AND2_X1 _1371_ (
    .A1(io_in[6]),
    .A2(io_in[5]),
    .ZN(_0458_)
  );
  INV_X1 _1372_ (
    .A(_0458_),
    .ZN(_0459_)
  );
  AND2_X1 _1373_ (
    .A1(_0256_),
    .A2(_0459_),
    .ZN(_0460_)
  );
  INV_X1 _1374_ (
    .A(_0460_),
    .ZN(_0461_)
  );
  AND2_X1 _1375_ (
    .A1(_0188_),
    .A2(_0461_),
    .ZN(_0462_)
  );
  INV_X1 _1376_ (
    .A(_0462_),
    .ZN(_0463_)
  );
  AND2_X1 _1377_ (
    .A1(_0125_),
    .A2(_0218_),
    .ZN(_0464_)
  );
  AND2_X1 _1378_ (
    .A1(_0185_),
    .A2(_0199_),
    .ZN(_0465_)
  );
  AND2_X1 _1379_ (
    .A1(_0464_),
    .A2(_0465_),
    .ZN(_0466_)
  );
  AND2_X1 _1380_ (
    .A1(io_in[2]),
    .A2(_0164_),
    .ZN(_0467_)
  );
  INV_X1 _1381_ (
    .A(_0467_),
    .ZN(_0468_)
  );
  AND2_X1 _1382_ (
    .A1(_0466_),
    .A2(_0468_),
    .ZN(_0469_)
  );
  AND2_X1 _1383_ (
    .A1(io_in[12]),
    .A2(_0949_),
    .ZN(_0470_)
  );
  INV_X1 _1384_ (
    .A(_0470_),
    .ZN(_0471_)
  );
  AND2_X1 _1385_ (
    .A1(io_in[12]),
    .A2(_0170_),
    .ZN(_0472_)
  );
  INV_X1 _1386_ (
    .A(_0472_),
    .ZN(_0473_)
  );
  AND2_X1 _1387_ (
    .A1(io_in[12]),
    .A2(_0203_),
    .ZN(_0474_)
  );
  INV_X1 _1388_ (
    .A(_0474_),
    .ZN(_0475_)
  );
  AND2_X1 _1389_ (
    .A1(_0473_),
    .A2(_0475_),
    .ZN(_0476_)
  );
  AND2_X1 _1390_ (
    .A1(_0463_),
    .A2(_0476_),
    .ZN(_0477_)
  );
  AND2_X1 _1391_ (
    .A1(_0471_),
    .A2(_0477_),
    .ZN(_0478_)
  );
  AND2_X1 _1392_ (
    .A1(_0469_),
    .A2(_0478_),
    .ZN(_0479_)
  );
  INV_X1 _1393_ (
    .A(_0479_),
    .ZN(io_out_bits[12])
  );
  AND2_X1 _1394_ (
    .A1(io_in[3]),
    .A2(_0164_),
    .ZN(_0480_)
  );
  INV_X1 _1395_ (
    .A(_0480_),
    .ZN(_0481_)
  );
  AND2_X1 _1396_ (
    .A1(_0299_),
    .A2(_0476_),
    .ZN(_0482_)
  );
  AND2_X1 _1397_ (
    .A1(io_in[11]),
    .A2(_0823_),
    .ZN(_0483_)
  );
  INV_X1 _1398_ (
    .A(_0483_),
    .ZN(_0484_)
  );
  AND2_X1 _1399_ (
    .A1(io_in[6]),
    .A2(io_in[11]),
    .ZN(_0485_)
  );
  INV_X1 _1400_ (
    .A(_0485_),
    .ZN(_0486_)
  );
  AND2_X1 _1401_ (
    .A1(_0484_),
    .A2(_0486_),
    .ZN(_0487_)
  );
  INV_X1 _1402_ (
    .A(_0487_),
    .ZN(_0488_)
  );
  AND2_X1 _1403_ (
    .A1(_0188_),
    .A2(_0488_),
    .ZN(_0489_)
  );
  INV_X1 _1404_ (
    .A(_0489_),
    .ZN(_0490_)
  );
  AND2_X1 _1405_ (
    .A1(io_in[0]),
    .A2(_0855_),
    .ZN(_0491_)
  );
  INV_X1 _1406_ (
    .A(_0491_),
    .ZN(_0492_)
  );
  AND2_X1 _1407_ (
    .A1(_0282_),
    .A2(_0492_),
    .ZN(_0493_)
  );
  INV_X1 _1408_ (
    .A(_0493_),
    .ZN(_0494_)
  );
  AND2_X1 _1409_ (
    .A1(_0490_),
    .A2(_0494_),
    .ZN(_0495_)
  );
  AND2_X1 _1410_ (
    .A1(_0481_),
    .A2(_0495_),
    .ZN(_0496_)
  );
  AND2_X1 _1411_ (
    .A1(_0482_),
    .A2(_0496_),
    .ZN(_0497_)
  );
  INV_X1 _1412_ (
    .A(_0497_),
    .ZN(io_out_bits[13])
  );
  AND2_X1 _1413_ (
    .A1(io_in[4]),
    .A2(_0164_),
    .ZN(_0498_)
  );
  INV_X1 _1414_ (
    .A(_0498_),
    .ZN(_0499_)
  );
  AND2_X1 _1415_ (
    .A1(_0790_),
    .A2(_0039_),
    .ZN(_0500_)
  );
  INV_X1 _1416_ (
    .A(_0500_),
    .ZN(_0501_)
  );
  AND2_X1 _1417_ (
    .A1(_0256_),
    .A2(_0501_),
    .ZN(_0502_)
  );
  INV_X1 _1418_ (
    .A(_0502_),
    .ZN(_0503_)
  );
  AND2_X1 _1419_ (
    .A1(_0188_),
    .A2(_0503_),
    .ZN(_0504_)
  );
  INV_X1 _1420_ (
    .A(_0504_),
    .ZN(_0505_)
  );
  AND2_X1 _1421_ (
    .A1(io_in[14]),
    .A2(_0949_),
    .ZN(_0506_)
  );
  INV_X1 _1422_ (
    .A(_0506_),
    .ZN(_0507_)
  );
  AND2_X1 _1423_ (
    .A1(_0476_),
    .A2(_0507_),
    .ZN(_0508_)
  );
  AND2_X1 _1424_ (
    .A1(_0505_),
    .A2(_0508_),
    .ZN(_0509_)
  );
  AND2_X1 _1425_ (
    .A1(_0499_),
    .A2(_0509_),
    .ZN(_0510_)
  );
  INV_X1 _1426_ (
    .A(_0510_),
    .ZN(io_out_bits[14])
  );
  AND2_X1 _1427_ (
    .A1(_0238_),
    .A2(_0343_),
    .ZN(_0511_)
  );
  INV_X1 _1428_ (
    .A(_0511_),
    .ZN(_0512_)
  );
  AND2_X1 _1429_ (
    .A1(io_in[7]),
    .A2(_0512_),
    .ZN(_0513_)
  );
  INV_X1 _1430_ (
    .A(_0513_),
    .ZN(_0514_)
  );
  AND2_X1 _1431_ (
    .A1(_0790_),
    .A2(_0077_),
    .ZN(_0515_)
  );
  INV_X1 _1432_ (
    .A(_0515_),
    .ZN(_0516_)
  );
  AND2_X1 _1433_ (
    .A1(io_in[7]),
    .A2(_0099_),
    .ZN(_0517_)
  );
  INV_X1 _1434_ (
    .A(_0517_),
    .ZN(_0518_)
  );
  AND2_X1 _1435_ (
    .A1(_0516_),
    .A2(_0517_),
    .ZN(_0519_)
  );
  INV_X1 _1436_ (
    .A(_0519_),
    .ZN(_0520_)
  );
  AND2_X1 _1437_ (
    .A1(_0292_),
    .A2(_0520_),
    .ZN(_0521_)
  );
  AND2_X1 _1438_ (
    .A1(_0514_),
    .A2(_0521_),
    .ZN(_0522_)
  );
  AND2_X1 _1439_ (
    .A1(io_in[7]),
    .A2(_0195_),
    .ZN(_0523_)
  );
  INV_X1 _1440_ (
    .A(_0523_),
    .ZN(_0524_)
  );
  AND2_X1 _1441_ (
    .A1(io_in[5]),
    .A2(_0164_),
    .ZN(_0525_)
  );
  INV_X1 _1442_ (
    .A(_0525_),
    .ZN(_0526_)
  );
  AND2_X1 _1443_ (
    .A1(_0476_),
    .A2(_0526_),
    .ZN(_0527_)
  );
  AND2_X1 _1444_ (
    .A1(_0524_),
    .A2(_0527_),
    .ZN(_0528_)
  );
  AND2_X1 _1445_ (
    .A1(_0522_),
    .A2(_0528_),
    .ZN(_0529_)
  );
  INV_X1 _1446_ (
    .A(_0529_),
    .ZN(io_out_bits[15])
  );
  AND2_X1 _1447_ (
    .A1(_0099_),
    .A2(_0516_),
    .ZN(_0530_)
  );
  INV_X1 _1448_ (
    .A(_0530_),
    .ZN(_0531_)
  );
  AND2_X1 _1449_ (
    .A1(io_in[8]),
    .A2(_0530_),
    .ZN(_0532_)
  );
  INV_X1 _1450_ (
    .A(_0532_),
    .ZN(_0533_)
  );
  AND2_X1 _1451_ (
    .A1(_0769_),
    .A2(_0088_),
    .ZN(_0534_)
  );
  INV_X1 _1452_ (
    .A(_0534_),
    .ZN(_0535_)
  );
  AND2_X1 _1453_ (
    .A1(_0090_),
    .A2(_0152_),
    .ZN(_0536_)
  );
  AND2_X1 _1454_ (
    .A1(_0535_),
    .A2(_0536_),
    .ZN(_0537_)
  );
  INV_X1 _1455_ (
    .A(_0537_),
    .ZN(_0538_)
  );
  AND2_X1 _1456_ (
    .A1(io_in[8]),
    .A2(_0188_),
    .ZN(_0539_)
  );
  INV_X1 _1457_ (
    .A(_0539_),
    .ZN(_0540_)
  );
  AND2_X1 _1458_ (
    .A1(_0801_),
    .A2(_0512_),
    .ZN(_0541_)
  );
  INV_X1 _1459_ (
    .A(_0541_),
    .ZN(_0542_)
  );
  MUX2_X1 _1460_ (
    .A(io_in[12]),
    .B(_0542_),
    .S(_0171_),
    .Z(_0543_)
  );
  AND2_X1 _1461_ (
    .A1(_0348_),
    .A2(_0543_),
    .ZN(_0544_)
  );
  INV_X1 _1462_ (
    .A(_0544_),
    .ZN(_0545_)
  );
  AND2_X1 _1463_ (
    .A1(_0540_),
    .A2(_0545_),
    .ZN(_0546_)
  );
  AND2_X1 _1464_ (
    .A1(_0538_),
    .A2(_0546_),
    .ZN(_0547_)
  );
  INV_X1 _1465_ (
    .A(_0547_),
    .ZN(_0548_)
  );
  AND2_X1 _1466_ (
    .A1(_0801_),
    .A2(_0193_),
    .ZN(_0549_)
  );
  INV_X1 _1467_ (
    .A(_0549_),
    .ZN(_0550_)
  );
  AND2_X1 _1468_ (
    .A1(io_rvc),
    .A2(_0100_),
    .ZN(_0551_)
  );
  AND2_X1 _1469_ (
    .A1(_0100_),
    .A2(_0550_),
    .ZN(_0552_)
  );
  MUX2_X1 _1470_ (
    .A(io_in[12]),
    .B(_0548_),
    .S(_0204_),
    .Z(_0553_)
  );
  AND2_X1 _1471_ (
    .A1(_0552_),
    .A2(_0553_),
    .ZN(_0554_)
  );
  INV_X1 _1472_ (
    .A(_0554_),
    .ZN(_0555_)
  );
  AND2_X1 _1473_ (
    .A1(_0533_),
    .A2(_0555_),
    .ZN(_0556_)
  );
  INV_X1 _1474_ (
    .A(_0556_),
    .ZN(_0557_)
  );
  MUX2_X1 _1475_ (
    .A(io_in[16]),
    .B(_0557_),
    .S(io_rvc),
    .Z(io_out_bits[16])
  );
  AND2_X1 _1476_ (
    .A1(_0511_),
    .A2(_0531_),
    .ZN(_0558_)
  );
  INV_X1 _1477_ (
    .A(_0558_),
    .ZN(_0559_)
  );
  AND2_X1 _1478_ (
    .A1(io_in[9]),
    .A2(_0559_),
    .ZN(_0560_)
  );
  INV_X1 _1479_ (
    .A(_0560_),
    .ZN(_0561_)
  );
  AND2_X1 _1480_ (
    .A1(io_in[17]),
    .A2(_0949_),
    .ZN(_0562_)
  );
  INV_X1 _1481_ (
    .A(_0562_),
    .ZN(_0563_)
  );
  AND2_X1 _1482_ (
    .A1(_0561_),
    .A2(_0563_),
    .ZN(_0564_)
  );
  AND2_X1 _1483_ (
    .A1(io_in[9]),
    .A2(_0195_),
    .ZN(_0565_)
  );
  INV_X1 _1484_ (
    .A(_0565_),
    .ZN(_0566_)
  );
  AND2_X1 _1485_ (
    .A1(io_in[12]),
    .A2(_0152_),
    .ZN(_0567_)
  );
  INV_X1 _1486_ (
    .A(_0567_),
    .ZN(_0568_)
  );
  AND2_X1 _1487_ (
    .A1(_0790_),
    .A2(_0088_),
    .ZN(_0569_)
  );
  INV_X1 _1488_ (
    .A(_0569_),
    .ZN(_0570_)
  );
  AND2_X1 _1489_ (
    .A1(_0152_),
    .A2(_0570_),
    .ZN(_0571_)
  );
  INV_X1 _1490_ (
    .A(_0571_),
    .ZN(_0572_)
  );
  AND2_X1 _1491_ (
    .A1(_0088_),
    .A2(_0567_),
    .ZN(_0573_)
  );
  INV_X1 _1492_ (
    .A(_0573_),
    .ZN(_0574_)
  );
  AND2_X1 _1493_ (
    .A1(_0476_),
    .A2(_0574_),
    .ZN(_0575_)
  );
  AND2_X1 _1494_ (
    .A1(_0566_),
    .A2(_0575_),
    .ZN(_0576_)
  );
  AND2_X1 _1495_ (
    .A1(_0564_),
    .A2(_0576_),
    .ZN(_0577_)
  );
  INV_X1 _1496_ (
    .A(_0577_),
    .ZN(io_out_bits[17])
  );
  AND2_X1 _1497_ (
    .A1(io_in[10]),
    .A2(_0176_),
    .ZN(_0578_)
  );
  INV_X1 _1498_ (
    .A(_0578_),
    .ZN(_0579_)
  );
  AND2_X1 _1499_ (
    .A1(_0289_),
    .A2(_0296_),
    .ZN(_0580_)
  );
  INV_X1 _1500_ (
    .A(_0580_),
    .ZN(_0581_)
  );
  AND2_X1 _1501_ (
    .A1(io_in[18]),
    .A2(_0581_),
    .ZN(_0582_)
  );
  INV_X1 _1502_ (
    .A(_0582_),
    .ZN(_0583_)
  );
  AND2_X1 _1503_ (
    .A1(_0579_),
    .A2(_0583_),
    .ZN(_0584_)
  );
  AND2_X1 _1504_ (
    .A1(io_in[10]),
    .A2(_0530_),
    .ZN(_0585_)
  );
  INV_X1 _1505_ (
    .A(_0585_),
    .ZN(_0586_)
  );
  AND2_X1 _1506_ (
    .A1(_0190_),
    .A2(_0586_),
    .ZN(_0587_)
  );
  AND2_X1 _1507_ (
    .A1(io_in[10]),
    .A2(_0158_),
    .ZN(_0588_)
  );
  INV_X1 _1508_ (
    .A(_0588_),
    .ZN(_0589_)
  );
  AND2_X1 _1509_ (
    .A1(io_in[18]),
    .A2(_0290_),
    .ZN(_0590_)
  );
  INV_X1 _1510_ (
    .A(_0590_),
    .ZN(_0591_)
  );
  AND2_X1 _1511_ (
    .A1(_0589_),
    .A2(_0591_),
    .ZN(_0592_)
  );
  AND2_X1 _1512_ (
    .A1(_0482_),
    .A2(_0592_),
    .ZN(_0593_)
  );
  AND2_X1 _1513_ (
    .A1(_0574_),
    .A2(_0593_),
    .ZN(_0594_)
  );
  AND2_X1 _1514_ (
    .A1(_0587_),
    .A2(_0594_),
    .ZN(_0595_)
  );
  AND2_X1 _1515_ (
    .A1(_0584_),
    .A2(_0595_),
    .ZN(_0596_)
  );
  INV_X1 _1516_ (
    .A(_0596_),
    .ZN(io_out_bits[18])
  );
  AND2_X1 _1517_ (
    .A1(io_in[11]),
    .A2(_0158_),
    .ZN(_0597_)
  );
  INV_X1 _1518_ (
    .A(_0597_),
    .ZN(_0598_)
  );
  AND2_X1 _1519_ (
    .A1(io_in[19]),
    .A2(_0290_),
    .ZN(_0599_)
  );
  INV_X1 _1520_ (
    .A(_0599_),
    .ZN(_0600_)
  );
  AND2_X1 _1521_ (
    .A1(_0598_),
    .A2(_0600_),
    .ZN(_0601_)
  );
  AND2_X1 _1522_ (
    .A1(io_in[11]),
    .A2(_0176_),
    .ZN(_0602_)
  );
  INV_X1 _1523_ (
    .A(_0602_),
    .ZN(_0603_)
  );
  AND2_X1 _1524_ (
    .A1(io_in[19]),
    .A2(_0581_),
    .ZN(_0604_)
  );
  INV_X1 _1525_ (
    .A(_0604_),
    .ZN(_0605_)
  );
  AND2_X1 _1526_ (
    .A1(_0603_),
    .A2(_0605_),
    .ZN(_0606_)
  );
  AND2_X1 _1527_ (
    .A1(io_in[11]),
    .A2(_0530_),
    .ZN(_0607_)
  );
  INV_X1 _1528_ (
    .A(_0607_),
    .ZN(_0608_)
  );
  AND2_X1 _1529_ (
    .A1(_0575_),
    .A2(_0608_),
    .ZN(_0609_)
  );
  AND2_X1 _1530_ (
    .A1(_0606_),
    .A2(_0609_),
    .ZN(_0610_)
  );
  AND2_X1 _1531_ (
    .A1(_0601_),
    .A2(_0610_),
    .ZN(_0611_)
  );
  INV_X1 _1532_ (
    .A(_0611_),
    .ZN(io_out_bits[19])
  );
  AND2_X1 _1533_ (
    .A1(_0191_),
    .A2(_0284_),
    .ZN(_0612_)
  );
  AND2_X1 _1534_ (
    .A1(_0438_),
    .A2(_0612_),
    .ZN(_0613_)
  );
  INV_X1 _1535_ (
    .A(_0613_),
    .ZN(_0614_)
  );
  AND2_X1 _1536_ (
    .A1(io_in[2]),
    .A2(_0614_),
    .ZN(_0615_)
  );
  INV_X1 _1537_ (
    .A(_0615_),
    .ZN(_0616_)
  );
  AND2_X1 _1538_ (
    .A1(io_in[12]),
    .A2(_0271_),
    .ZN(_0617_)
  );
  INV_X1 _1539_ (
    .A(_0617_),
    .ZN(_0618_)
  );
  AND2_X1 _1540_ (
    .A1(_0906_),
    .A2(_0618_),
    .ZN(_0619_)
  );
  INV_X1 _1541_ (
    .A(_0619_),
    .ZN(_0620_)
  );
  AND2_X1 _1542_ (
    .A1(_0099_),
    .A2(_0620_),
    .ZN(_0621_)
  );
  INV_X1 _1543_ (
    .A(_0621_),
    .ZN(_0622_)
  );
  AND2_X1 _1544_ (
    .A1(io_in[20]),
    .A2(_0949_),
    .ZN(_0623_)
  );
  INV_X1 _1545_ (
    .A(_0623_),
    .ZN(_0624_)
  );
  AND2_X1 _1546_ (
    .A1(_0575_),
    .A2(_0624_),
    .ZN(_0625_)
  );
  AND2_X1 _1547_ (
    .A1(_0622_),
    .A2(_0625_),
    .ZN(_0626_)
  );
  AND2_X1 _1548_ (
    .A1(_0616_),
    .A2(_0626_),
    .ZN(_0627_)
  );
  INV_X1 _1549_ (
    .A(_0627_),
    .ZN(io_out_bits[20])
  );
  AND2_X1 _1550_ (
    .A1(_0171_),
    .A2(_0438_),
    .ZN(_0628_)
  );
  AND2_X1 _1551_ (
    .A1(_0189_),
    .A2(_0204_),
    .ZN(_0629_)
  );
  AND2_X1 _1552_ (
    .A1(_0097_),
    .A2(_0177_),
    .ZN(_0630_)
  );
  AND2_X1 _1553_ (
    .A1(_0629_),
    .A2(_0630_),
    .ZN(_0631_)
  );
  AND2_X1 _1554_ (
    .A1(_0628_),
    .A2(_0631_),
    .ZN(_0632_)
  );
  INV_X1 _1555_ (
    .A(_0632_),
    .ZN(_0633_)
  );
  AND2_X1 _1556_ (
    .A1(io_in[3]),
    .A2(_0633_),
    .ZN(_0634_)
  );
  INV_X1 _1557_ (
    .A(_0634_),
    .ZN(_0635_)
  );
  AND2_X1 _1558_ (
    .A1(io_in[21]),
    .A2(_0949_),
    .ZN(_0636_)
  );
  INV_X1 _1559_ (
    .A(_0636_),
    .ZN(_0637_)
  );
  AND2_X1 _1560_ (
    .A1(_0574_),
    .A2(_0637_),
    .ZN(_0638_)
  );
  AND2_X1 _1561_ (
    .A1(_0635_),
    .A2(_0638_),
    .ZN(_0639_)
  );
  INV_X1 _1562_ (
    .A(_0639_),
    .ZN(io_out_bits[21])
  );
  AND2_X1 _1563_ (
    .A1(_0094_),
    .A2(_0295_),
    .ZN(_0640_)
  );
  INV_X1 _1564_ (
    .A(_0640_),
    .ZN(_0641_)
  );
  AND2_X1 _1565_ (
    .A1(_0292_),
    .A2(_0641_),
    .ZN(_0642_)
  );
  INV_X1 _1566_ (
    .A(_0642_),
    .ZN(_0643_)
  );
  AND2_X1 _1567_ (
    .A1(io_in[22]),
    .A2(_0949_),
    .ZN(_0644_)
  );
  INV_X1 _1568_ (
    .A(_0644_),
    .ZN(_0645_)
  );
  AND2_X1 _1569_ (
    .A1(_0833_),
    .A2(io_in[1]),
    .ZN(_0646_)
  );
  AND2_X1 _1570_ (
    .A1(_0097_),
    .A2(_0110_),
    .ZN(_0647_)
  );
  INV_X1 _1571_ (
    .A(_0647_),
    .ZN(_0648_)
  );
  AND2_X1 _1572_ (
    .A1(io_in[4]),
    .A2(_0648_),
    .ZN(_0649_)
  );
  INV_X1 _1573_ (
    .A(_0649_),
    .ZN(_0650_)
  );
  AND2_X1 _1574_ (
    .A1(io_in[4]),
    .A2(_0176_),
    .ZN(_0651_)
  );
  INV_X1 _1575_ (
    .A(_0651_),
    .ZN(_0652_)
  );
  AND2_X1 _1576_ (
    .A1(io_in[6]),
    .A2(_0125_),
    .ZN(_0653_)
  );
  MUX2_X1 _1577_ (
    .A(io_in[4]),
    .B(_0653_),
    .S(_0628_),
    .Z(_0654_)
  );
  AND2_X1 _1578_ (
    .A1(_0153_),
    .A2(_0654_),
    .ZN(_0655_)
  );
  INV_X1 _1579_ (
    .A(_0655_),
    .ZN(_0656_)
  );
  AND2_X1 _1580_ (
    .A1(_0574_),
    .A2(_0629_),
    .ZN(_0657_)
  );
  AND2_X1 _1581_ (
    .A1(_0656_),
    .A2(_0657_),
    .ZN(_0658_)
  );
  INV_X1 _1582_ (
    .A(_0658_),
    .ZN(_0659_)
  );
  AND2_X1 _1583_ (
    .A1(_0177_),
    .A2(_0180_),
    .ZN(_0660_)
  );
  INV_X1 _1584_ (
    .A(_0660_),
    .ZN(_0661_)
  );
  AND2_X1 _1585_ (
    .A1(io_in[4]),
    .A2(_0192_),
    .ZN(_0662_)
  );
  INV_X1 _1586_ (
    .A(_0662_),
    .ZN(_0663_)
  );
  AND2_X1 _1587_ (
    .A1(_0661_),
    .A2(_0663_),
    .ZN(_0664_)
  );
  INV_X1 _1588_ (
    .A(_0664_),
    .ZN(_0665_)
  );
  AND2_X1 _1589_ (
    .A1(_0659_),
    .A2(_0665_),
    .ZN(_0666_)
  );
  INV_X1 _1590_ (
    .A(_0666_),
    .ZN(_0667_)
  );
  AND2_X1 _1591_ (
    .A1(_0652_),
    .A2(_0667_),
    .ZN(_0668_)
  );
  INV_X1 _1592_ (
    .A(_0668_),
    .ZN(_0669_)
  );
  AND2_X1 _1593_ (
    .A1(_0097_),
    .A2(_0309_),
    .ZN(_0670_)
  );
  AND2_X1 _1594_ (
    .A1(_0669_),
    .A2(_0670_),
    .ZN(_0671_)
  );
  INV_X1 _1595_ (
    .A(_0671_),
    .ZN(_0672_)
  );
  AND2_X1 _1596_ (
    .A1(_0650_),
    .A2(_0672_),
    .ZN(_0673_)
  );
  INV_X1 _1597_ (
    .A(_0673_),
    .ZN(_0674_)
  );
  MUX2_X1 _1598_ (
    .A(io_in[22]),
    .B(_0674_),
    .S(io_rvc),
    .Z(io_out_bits[22])
  );
  AND2_X1 _1599_ (
    .A1(io_rvc),
    .A2(_0186_),
    .ZN(_0675_)
  );
  AND2_X1 _1600_ (
    .A1(_0153_),
    .A2(_0238_),
    .ZN(_0676_)
  );
  AND2_X1 _1601_ (
    .A1(io_in[5]),
    .A2(_0676_),
    .ZN(_0677_)
  );
  INV_X1 _1602_ (
    .A(_0677_),
    .ZN(_0678_)
  );
  AND2_X1 _1603_ (
    .A1(_0188_),
    .A2(_0257_),
    .ZN(_0679_)
  );
  INV_X1 _1604_ (
    .A(_0679_),
    .ZN(_0680_)
  );
  AND2_X1 _1605_ (
    .A1(_0823_),
    .A2(_0115_),
    .ZN(_0681_)
  );
  INV_X1 _1606_ (
    .A(_0681_),
    .ZN(_0682_)
  );
  AND2_X1 _1607_ (
    .A1(_0300_),
    .A2(_0682_),
    .ZN(_0683_)
  );
  INV_X1 _1608_ (
    .A(_0683_),
    .ZN(_0684_)
  );
  AND2_X1 _1609_ (
    .A1(_0189_),
    .A2(_0574_),
    .ZN(_0685_)
  );
  AND2_X1 _1610_ (
    .A1(_0684_),
    .A2(_0685_),
    .ZN(_0686_)
  );
  INV_X1 _1611_ (
    .A(_0686_),
    .ZN(_0687_)
  );
  AND2_X1 _1612_ (
    .A1(_0680_),
    .A2(_0687_),
    .ZN(_0688_)
  );
  INV_X1 _1613_ (
    .A(_0688_),
    .ZN(_0689_)
  );
  AND2_X1 _1614_ (
    .A1(_0678_),
    .A2(_0689_),
    .ZN(_0690_)
  );
  INV_X1 _1615_ (
    .A(_0690_),
    .ZN(_0691_)
  );
  AND2_X1 _1616_ (
    .A1(_0675_),
    .A2(_0691_),
    .ZN(_0692_)
  );
  INV_X1 _1617_ (
    .A(_0692_),
    .ZN(_0693_)
  );
  AND2_X1 _1618_ (
    .A1(io_in[23]),
    .A2(_0949_),
    .ZN(_0694_)
  );
  INV_X1 _1619_ (
    .A(_0694_),
    .ZN(_0695_)
  );
  AND2_X1 _1620_ (
    .A1(_0693_),
    .A2(_0695_),
    .ZN(_0696_)
  );
  INV_X1 _1621_ (
    .A(_0696_),
    .ZN(io_out_bits[23])
  );
  AND2_X1 _1622_ (
    .A1(io_in[24]),
    .A2(_0949_),
    .ZN(_0697_)
  );
  INV_X1 _1623_ (
    .A(_0697_),
    .ZN(_0698_)
  );
  AND2_X1 _1624_ (
    .A1(io_in[11]),
    .A2(_0452_),
    .ZN(_0699_)
  );
  INV_X1 _1625_ (
    .A(_0699_),
    .ZN(_0700_)
  );
  AND2_X1 _1626_ (
    .A1(_0574_),
    .A2(_0700_),
    .ZN(_0701_)
  );
  INV_X1 _1627_ (
    .A(_0701_),
    .ZN(_0702_)
  );
  AND2_X1 _1628_ (
    .A1(_0189_),
    .A2(_0702_),
    .ZN(_0703_)
  );
  INV_X1 _1629_ (
    .A(_0703_),
    .ZN(_0704_)
  );
  AND2_X1 _1630_ (
    .A1(_0161_),
    .A2(_0165_),
    .ZN(_0705_)
  );
  INV_X1 _1631_ (
    .A(_0705_),
    .ZN(_0706_)
  );
  AND2_X1 _1632_ (
    .A1(_0189_),
    .A2(_0706_),
    .ZN(_0707_)
  );
  INV_X1 _1633_ (
    .A(_0707_),
    .ZN(_0708_)
  );
  AND2_X1 _1634_ (
    .A1(io_in[6]),
    .A2(_0708_),
    .ZN(_0709_)
  );
  INV_X1 _1635_ (
    .A(_0709_),
    .ZN(_0710_)
  );
  AND2_X1 _1636_ (
    .A1(_0704_),
    .A2(_0710_),
    .ZN(_0711_)
  );
  INV_X1 _1637_ (
    .A(_0711_),
    .ZN(_0712_)
  );
  AND2_X1 _1638_ (
    .A1(_0097_),
    .A2(_0235_),
    .ZN(_0713_)
  );
  AND2_X1 _1639_ (
    .A1(_0259_),
    .A2(_0713_),
    .ZN(_0714_)
  );
  AND2_X1 _1640_ (
    .A1(_0712_),
    .A2(_0714_),
    .ZN(_0715_)
  );
  INV_X1 _1641_ (
    .A(_0715_),
    .ZN(_0716_)
  );
  AND2_X1 _1642_ (
    .A1(io_in[6]),
    .A2(_0646_),
    .ZN(_0717_)
  );
  INV_X1 _1643_ (
    .A(_0717_),
    .ZN(_0718_)
  );
  AND2_X1 _1644_ (
    .A1(_0716_),
    .A2(_0718_),
    .ZN(_0719_)
  );
  INV_X1 _1645_ (
    .A(_0719_),
    .ZN(_0720_)
  );
  AND2_X1 _1646_ (
    .A1(_0698_),
    .A2(_0718_),
    .ZN(_0721_)
  );
  INV_X1 _1647_ (
    .A(_0721_),
    .ZN(io_out_rs2[4])
  );
  MUX2_X1 _1648_ (
    .A(io_in[24]),
    .B(_0720_),
    .S(io_rvc),
    .Z(io_out_bits[24])
  );
  AND2_X1 _1649_ (
    .A1(io_in[25]),
    .A2(_0949_),
    .ZN(_0722_)
  );
  INV_X1 _1650_ (
    .A(_0722_),
    .ZN(_0723_)
  );
  MUX2_X1 _1651_ (
    .A(_0257_),
    .B(_0392_),
    .S(_0189_),
    .Z(_0724_)
  );
  AND2_X1 _1652_ (
    .A1(io_in[12]),
    .A2(_0724_),
    .ZN(_0725_)
  );
  INV_X1 _1653_ (
    .A(_0725_),
    .ZN(_0726_)
  );
  AND2_X1 _1654_ (
    .A1(_0574_),
    .A2(_0726_),
    .ZN(_0727_)
  );
  INV_X1 _1655_ (
    .A(_0727_),
    .ZN(_0728_)
  );
  AND2_X1 _1656_ (
    .A1(_0305_),
    .A2(_0728_),
    .ZN(_0729_)
  );
  INV_X1 _1657_ (
    .A(_0729_),
    .ZN(_0730_)
  );
  AND2_X1 _1658_ (
    .A1(_0171_),
    .A2(_0572_),
    .ZN(_0731_)
  );
  AND2_X1 _1659_ (
    .A1(_0305_),
    .A2(_0731_),
    .ZN(_0732_)
  );
  INV_X1 _1660_ (
    .A(_0732_),
    .ZN(_0733_)
  );
  AND2_X1 _1661_ (
    .A1(io_in[2]),
    .A2(_0733_),
    .ZN(_0734_)
  );
  INV_X1 _1662_ (
    .A(_0734_),
    .ZN(_0735_)
  );
  AND2_X1 _1663_ (
    .A1(_0730_),
    .A2(_0735_),
    .ZN(_0736_)
  );
  INV_X1 _1664_ (
    .A(_0736_),
    .ZN(_0737_)
  );
  AND2_X1 _1665_ (
    .A1(_0551_),
    .A2(_0737_),
    .ZN(_0738_)
  );
  INV_X1 _1666_ (
    .A(_0738_),
    .ZN(_0739_)
  );
  AND2_X1 _1667_ (
    .A1(_0723_),
    .A2(_0739_),
    .ZN(_0740_)
  );
  INV_X1 _1668_ (
    .A(_0740_),
    .ZN(io_out_bits[25])
  );
  AND2_X1 _1669_ (
    .A1(io_in[26]),
    .A2(_0949_),
    .ZN(_0741_)
  );
  INV_X1 _1670_ (
    .A(_0741_),
    .ZN(_0742_)
  );
  AND2_X1 _1671_ (
    .A1(io_in[2]),
    .A2(_0308_),
    .ZN(_0743_)
  );
  INV_X1 _1672_ (
    .A(_0743_),
    .ZN(_0744_)
  );
  AND2_X1 _1673_ (
    .A1(_0238_),
    .A2(_0438_),
    .ZN(_0745_)
  );
  AND2_X1 _1674_ (
    .A1(io_in[7]),
    .A2(_0745_),
    .ZN(_0746_)
  );
  INV_X1 _1675_ (
    .A(_0746_),
    .ZN(_0747_)
  );
  AND2_X1 _1676_ (
    .A1(io_in[12]),
    .A2(_0154_),
    .ZN(_0748_)
  );
  INV_X1 _1677_ (
    .A(_0748_),
    .ZN(_0749_)
  );
  AND2_X1 _1678_ (
    .A1(io_in[12]),
    .A2(_0158_),
    .ZN(_0750_)
  );
  INV_X1 _1679_ (
    .A(_0750_),
    .ZN(_0751_)
  );
  AND2_X1 _1680_ (
    .A1(_0749_),
    .A2(_0751_),
    .ZN(_0752_)
  );
  AND2_X1 _1681_ (
    .A1(_0747_),
    .A2(_0752_),
    .ZN(_0753_)
  );
  INV_X1 _1682_ (
    .A(_0753_),
    .ZN(_0754_)
  );
  AND2_X1 _1683_ (
    .A1(_0153_),
    .A2(_0754_),
    .ZN(_0755_)
  );
  INV_X1 _1684_ (
    .A(_0755_),
    .ZN(_0756_)
  );
  AND2_X1 _1685_ (
    .A1(_0153_),
    .A2(_0299_),
    .ZN(_0757_)
  );
  INV_X1 _1686_ (
    .A(_0757_),
    .ZN(_0758_)
  );
  AND2_X1 _1687_ (
    .A1(io_in[5]),
    .A2(_0758_),
    .ZN(_0759_)
  );
  MUX2_X1 _1688_ (
    .A(io_in[12]),
    .B(_0759_),
    .S(_0165_),
    .Z(_0760_)
  );
  INV_X1 _1689_ (
    .A(_0760_),
    .ZN(_0761_)
  );
  AND2_X1 _1690_ (
    .A1(_0756_),
    .A2(_0761_),
    .ZN(_0762_)
  );
  INV_X1 _1691_ (
    .A(_0762_),
    .ZN(_0763_)
  );
  AND2_X1 _1692_ (
    .A1(_0190_),
    .A2(_0763_),
    .ZN(_0764_)
  );
  INV_X1 _1693_ (
    .A(_0764_),
    .ZN(_0765_)
  );
  AND2_X1 _1694_ (
    .A1(io_in[5]),
    .A2(_0187_),
    .ZN(_0766_)
  );
  INV_X1 _1695_ (
    .A(_0766_),
    .ZN(_0767_)
  );
  AND2_X1 _1696_ (
    .A1(io_in[12]),
    .A2(_0483_),
    .ZN(_0768_)
  );
  AND2_X1 _1697_ (
    .A1(_0188_),
    .A2(_0768_),
    .ZN(_0770_)
  );
  INV_X1 _1698_ (
    .A(_0770_),
    .ZN(_0771_)
  );
  AND2_X1 _1699_ (
    .A1(_0767_),
    .A2(_0771_),
    .ZN(_0772_)
  );
  AND2_X1 _1700_ (
    .A1(_0765_),
    .A2(_0772_),
    .ZN(_0773_)
  );
  INV_X1 _1701_ (
    .A(_0773_),
    .ZN(_0774_)
  );
  AND2_X1 _1702_ (
    .A1(_0107_),
    .A2(_0774_),
    .ZN(_0775_)
  );
  INV_X1 _1703_ (
    .A(_0775_),
    .ZN(_0776_)
  );
  AND2_X1 _1704_ (
    .A1(_0744_),
    .A2(_0776_),
    .ZN(_0777_)
  );
  INV_X1 _1705_ (
    .A(_0777_),
    .ZN(_0778_)
  );
  AND2_X1 _1706_ (
    .A1(_0551_),
    .A2(_0778_),
    .ZN(_0779_)
  );
  INV_X1 _1707_ (
    .A(_0779_),
    .ZN(_0781_)
  );
  AND2_X1 _1708_ (
    .A1(_0742_),
    .A2(_0781_),
    .ZN(_0782_)
  );
  INV_X1 _1709_ (
    .A(_0782_),
    .ZN(io_out_bits[26])
  );
  AND2_X1 _1710_ (
    .A1(io_in[27]),
    .A2(_0949_),
    .ZN(_0783_)
  );
  INV_X1 _1711_ (
    .A(_0783_),
    .ZN(_0784_)
  );
  AND2_X1 _1712_ (
    .A1(io_in[3]),
    .A2(_0308_),
    .ZN(_0785_)
  );
  INV_X1 _1713_ (
    .A(_0785_),
    .ZN(_0786_)
  );
  AND2_X1 _1714_ (
    .A1(_0917_),
    .A2(_0087_),
    .ZN(_0787_)
  );
  INV_X1 _1715_ (
    .A(_0787_),
    .ZN(_0788_)
  );
  AND2_X1 _1716_ (
    .A1(_0571_),
    .A2(_0788_),
    .ZN(_0789_)
  );
  INV_X1 _1717_ (
    .A(_0789_),
    .ZN(_0791_)
  );
  AND2_X1 _1718_ (
    .A1(io_in[6]),
    .A2(_0245_),
    .ZN(_0792_)
  );
  INV_X1 _1719_ (
    .A(_0792_),
    .ZN(_0793_)
  );
  MUX2_X1 _1720_ (
    .A(io_in[8]),
    .B(io_in[6]),
    .S(_0124_),
    .Z(_0794_)
  );
  AND2_X1 _1721_ (
    .A1(_0144_),
    .A2(_0794_),
    .ZN(_0795_)
  );
  AND2_X1 _1722_ (
    .A1(_0134_),
    .A2(_0795_),
    .ZN(_0796_)
  );
  INV_X1 _1723_ (
    .A(_0796_),
    .ZN(_0797_)
  );
  AND2_X1 _1724_ (
    .A1(_0793_),
    .A2(_0797_),
    .ZN(_0798_)
  );
  INV_X1 _1725_ (
    .A(_0798_),
    .ZN(_0799_)
  );
  AND2_X1 _1726_ (
    .A1(_0249_),
    .A2(_0799_),
    .ZN(_0800_)
  );
  INV_X1 _1727_ (
    .A(_0800_),
    .ZN(_0802_)
  );
  AND2_X1 _1728_ (
    .A1(_0171_),
    .A2(_0751_),
    .ZN(_0803_)
  );
  AND2_X1 _1729_ (
    .A1(_0802_),
    .A2(_0803_),
    .ZN(_0804_)
  );
  INV_X1 _1730_ (
    .A(_0804_),
    .ZN(_0805_)
  );
  AND2_X1 _1731_ (
    .A1(_0769_),
    .A2(_0170_),
    .ZN(_0806_)
  );
  INV_X1 _1732_ (
    .A(_0806_),
    .ZN(_0807_)
  );
  AND2_X1 _1733_ (
    .A1(_0805_),
    .A2(_0807_),
    .ZN(_0808_)
  );
  MUX2_X1 _1734_ (
    .A(io_in[12]),
    .B(_0808_),
    .S(_0155_),
    .Z(_0809_)
  );
  AND2_X1 _1735_ (
    .A1(_0153_),
    .A2(_0809_),
    .ZN(_0810_)
  );
  INV_X1 _1736_ (
    .A(_0810_),
    .ZN(_0811_)
  );
  AND2_X1 _1737_ (
    .A1(_0791_),
    .A2(_0811_),
    .ZN(_0813_)
  );
  MUX2_X1 _1738_ (
    .A(_0093_),
    .B(_0813_),
    .S(_0180_),
    .Z(_0814_)
  );
  AND2_X1 _1739_ (
    .A1(_0771_),
    .A2(_0814_),
    .ZN(_0815_)
  );
  INV_X1 _1740_ (
    .A(_0815_),
    .ZN(_0816_)
  );
  AND2_X1 _1741_ (
    .A1(_0769_),
    .A2(_0306_),
    .ZN(_0817_)
  );
  INV_X1 _1742_ (
    .A(_0817_),
    .ZN(_0818_)
  );
  AND2_X1 _1743_ (
    .A1(_0107_),
    .A2(_0818_),
    .ZN(_0819_)
  );
  AND2_X1 _1744_ (
    .A1(_0816_),
    .A2(_0819_),
    .ZN(_0820_)
  );
  INV_X1 _1745_ (
    .A(_0820_),
    .ZN(_0821_)
  );
  AND2_X1 _1746_ (
    .A1(_0786_),
    .A2(_0821_),
    .ZN(_0822_)
  );
  INV_X1 _1747_ (
    .A(_0822_),
    .ZN(_0824_)
  );
  AND2_X1 _1748_ (
    .A1(_0551_),
    .A2(_0824_),
    .ZN(_0825_)
  );
  INV_X1 _1749_ (
    .A(_0825_),
    .ZN(_0826_)
  );
  AND2_X1 _1750_ (
    .A1(_0784_),
    .A2(_0826_),
    .ZN(_0827_)
  );
  INV_X1 _1751_ (
    .A(_0827_),
    .ZN(io_out_bits[27])
  );
  AND2_X1 _1752_ (
    .A1(io_in[28]),
    .A2(_0949_),
    .ZN(_0828_)
  );
  INV_X1 _1753_ (
    .A(_0828_),
    .ZN(_0829_)
  );
  AND2_X1 _1754_ (
    .A1(io_in[4]),
    .A2(_0200_),
    .ZN(_0830_)
  );
  INV_X1 _1755_ (
    .A(_0830_),
    .ZN(_0831_)
  );
  AND2_X1 _1756_ (
    .A1(io_in[9]),
    .A2(_0745_),
    .ZN(_0832_)
  );
  INV_X1 _1757_ (
    .A(_0832_),
    .ZN(_0834_)
  );
  AND2_X1 _1758_ (
    .A1(_0752_),
    .A2(_0834_),
    .ZN(_0835_)
  );
  INV_X1 _1759_ (
    .A(_0835_),
    .ZN(_0836_)
  );
  AND2_X1 _1760_ (
    .A1(_0153_),
    .A2(_0836_),
    .ZN(_0837_)
  );
  INV_X1 _1761_ (
    .A(_0837_),
    .ZN(_0838_)
  );
  AND2_X1 _1762_ (
    .A1(_0928_),
    .A2(_0087_),
    .ZN(_0839_)
  );
  INV_X1 _1763_ (
    .A(_0839_),
    .ZN(_0840_)
  );
  AND2_X1 _1764_ (
    .A1(_0571_),
    .A2(_0840_),
    .ZN(_0841_)
  );
  INV_X1 _1765_ (
    .A(_0841_),
    .ZN(_0842_)
  );
  AND2_X1 _1766_ (
    .A1(_0838_),
    .A2(_0842_),
    .ZN(_0843_)
  );
  INV_X1 _1767_ (
    .A(_0843_),
    .ZN(_0845_)
  );
  AND2_X1 _1768_ (
    .A1(_0190_),
    .A2(_0845_),
    .ZN(_0846_)
  );
  INV_X1 _1769_ (
    .A(_0846_),
    .ZN(_0847_)
  );
  AND2_X1 _1770_ (
    .A1(_0354_),
    .A2(_0771_),
    .ZN(_0848_)
  );
  AND2_X1 _1771_ (
    .A1(_0847_),
    .A2(_0848_),
    .ZN(_0849_)
  );
  INV_X1 _1772_ (
    .A(_0849_),
    .ZN(_0850_)
  );
  AND2_X1 _1773_ (
    .A1(_0199_),
    .A2(_0850_),
    .ZN(_0851_)
  );
  INV_X1 _1774_ (
    .A(_0851_),
    .ZN(_0852_)
  );
  AND2_X1 _1775_ (
    .A1(_0831_),
    .A2(_0852_),
    .ZN(_0853_)
  );
  INV_X1 _1776_ (
    .A(_0853_),
    .ZN(_0854_)
  );
  AND2_X1 _1777_ (
    .A1(_0113_),
    .A2(_0432_),
    .ZN(_0856_)
  );
  AND2_X1 _1778_ (
    .A1(_0209_),
    .A2(_0856_),
    .ZN(_0857_)
  );
  AND2_X1 _1779_ (
    .A1(_0854_),
    .A2(_0857_),
    .ZN(_0858_)
  );
  INV_X1 _1780_ (
    .A(_0858_),
    .ZN(_0859_)
  );
  AND2_X1 _1781_ (
    .A1(_0829_),
    .A2(_0859_),
    .ZN(_0860_)
  );
  INV_X1 _1782_ (
    .A(_0860_),
    .ZN(io_out_bits[28])
  );
  AND2_X1 _1783_ (
    .A1(io_in[29]),
    .A2(_0949_),
    .ZN(_0861_)
  );
  INV_X1 _1784_ (
    .A(_0861_),
    .ZN(_0862_)
  );
  AND2_X1 _1785_ (
    .A1(io_in[10]),
    .A2(_0745_),
    .ZN(_0863_)
  );
  INV_X1 _1786_ (
    .A(_0863_),
    .ZN(_0864_)
  );
  AND2_X1 _1787_ (
    .A1(_0568_),
    .A2(_0752_),
    .ZN(_0866_)
  );
  AND2_X1 _1788_ (
    .A1(_0771_),
    .A2(_0866_),
    .ZN(_0867_)
  );
  AND2_X1 _1789_ (
    .A1(_0864_),
    .A2(_0867_),
    .ZN(_0868_)
  );
  INV_X1 _1790_ (
    .A(_0868_),
    .ZN(_0869_)
  );
  MUX2_X1 _1791_ (
    .A(_0186_),
    .B(_0768_),
    .S(_0188_),
    .Z(_0870_)
  );
  AND2_X1 _1792_ (
    .A1(_0790_),
    .A2(_0152_),
    .ZN(_0871_)
  );
  INV_X1 _1793_ (
    .A(_0871_),
    .ZN(_0872_)
  );
  AND2_X1 _1794_ (
    .A1(_0870_),
    .A2(_0872_),
    .ZN(_0873_)
  );
  AND2_X1 _1795_ (
    .A1(_0869_),
    .A2(_0873_),
    .ZN(_0874_)
  );
  INV_X1 _1796_ (
    .A(_0874_),
    .ZN(_0875_)
  );
  AND2_X1 _1797_ (
    .A1(_0354_),
    .A2(_0875_),
    .ZN(_0877_)
  );
  INV_X1 _1798_ (
    .A(_0877_),
    .ZN(_0878_)
  );
  AND2_X1 _1799_ (
    .A1(_0865_),
    .A2(_0878_),
    .ZN(_0879_)
  );
  INV_X1 _1800_ (
    .A(_0879_),
    .ZN(_0880_)
  );
  AND2_X1 _1801_ (
    .A1(_0862_),
    .A2(_0880_),
    .ZN(_0881_)
  );
  INV_X1 _1802_ (
    .A(_0881_),
    .ZN(io_out_bits[29])
  );
  AND2_X1 _1803_ (
    .A1(io_in[30]),
    .A2(_0949_),
    .ZN(_0882_)
  );
  INV_X1 _1804_ (
    .A(_0882_),
    .ZN(_0883_)
  );
  AND2_X1 _1805_ (
    .A1(_0354_),
    .A2(_0883_),
    .ZN(_0884_)
  );
  AND2_X1 _1806_ (
    .A1(io_in[11]),
    .A2(_0039_),
    .ZN(_0885_)
  );
  INV_X1 _1807_ (
    .A(_0885_),
    .ZN(_0887_)
  );
  AND2_X1 _1808_ (
    .A1(_0188_),
    .A2(_0887_),
    .ZN(_0888_)
  );
  AND2_X1 _1809_ (
    .A1(io_in[10]),
    .A2(_0888_),
    .ZN(_0889_)
  );
  INV_X1 _1810_ (
    .A(_0889_),
    .ZN(_0890_)
  );
  AND2_X1 _1811_ (
    .A1(io_in[8]),
    .A2(_0168_),
    .ZN(_0891_)
  );
  INV_X1 _1812_ (
    .A(_0891_),
    .ZN(_0892_)
  );
  AND2_X1 _1813_ (
    .A1(_0890_),
    .A2(_0892_),
    .ZN(_0893_)
  );
  AND2_X1 _1814_ (
    .A1(_0884_),
    .A2(_0893_),
    .ZN(_0894_)
  );
  AND2_X1 _1815_ (
    .A1(_0867_),
    .A2(_0894_),
    .ZN(_0895_)
  );
  INV_X1 _1816_ (
    .A(_0895_),
    .ZN(io_out_bits[30])
  );
  AND2_X1 _1817_ (
    .A1(io_in[31]),
    .A2(_0949_),
    .ZN(_0897_)
  );
  INV_X1 _1818_ (
    .A(_0897_),
    .ZN(_0898_)
  );
  AND2_X1 _1819_ (
    .A1(_0476_),
    .A2(_0898_),
    .ZN(_0899_)
  );
  AND2_X1 _1820_ (
    .A1(_0848_),
    .A2(_0899_),
    .ZN(_0900_)
  );
  AND2_X1 _1821_ (
    .A1(_0866_),
    .A2(_0900_),
    .ZN(_0901_)
  );
  INV_X1 _1822_ (
    .A(_0901_),
    .ZN(io_out_bits[31])
  );
  AND2_X1 _1823_ (
    .A1(_0886_),
    .A2(_0298_),
    .ZN(_0902_)
  );
  INV_X1 _1824_ (
    .A(_0902_),
    .ZN(_0903_)
  );
  AND2_X1 _1825_ (
    .A1(io_in[7]),
    .A2(_0182_),
    .ZN(_0904_)
  );
  INV_X1 _1826_ (
    .A(_0904_),
    .ZN(_0905_)
  );
  AND2_X1 _1827_ (
    .A1(io_in[2]),
    .A2(_0159_),
    .ZN(_0907_)
  );
  INV_X1 _1828_ (
    .A(_0907_),
    .ZN(_0908_)
  );
  AND2_X1 _1829_ (
    .A1(_0342_),
    .A2(_0908_),
    .ZN(_0909_)
  );
  INV_X1 _1830_ (
    .A(_0909_),
    .ZN(_0910_)
  );
  MUX2_X1 _1831_ (
    .A(io_in[7]),
    .B(_0910_),
    .S(_0348_),
    .Z(_0911_)
  );
  AND2_X1 _1832_ (
    .A1(_0304_),
    .A2(_0911_),
    .ZN(_0912_)
  );
  INV_X1 _1833_ (
    .A(_0912_),
    .ZN(_0913_)
  );
  AND2_X1 _1834_ (
    .A1(_0905_),
    .A2(_0913_),
    .ZN(_0914_)
  );
  INV_X1 _1835_ (
    .A(_0914_),
    .ZN(_0915_)
  );
  AND2_X1 _1836_ (
    .A1(_0234_),
    .A2(_0915_),
    .ZN(_0916_)
  );
  INV_X1 _1837_ (
    .A(_0916_),
    .ZN(_0918_)
  );
  AND2_X1 _1838_ (
    .A1(_0360_),
    .A2(_0918_),
    .ZN(_0919_)
  );
  INV_X1 _1839_ (
    .A(_0919_),
    .ZN(_0920_)
  );
  AND2_X1 _1840_ (
    .A1(_0100_),
    .A2(_0920_),
    .ZN(_0921_)
  );
  INV_X1 _1841_ (
    .A(_0921_),
    .ZN(_0922_)
  );
  AND2_X1 _1842_ (
    .A1(_0331_),
    .A2(_0518_),
    .ZN(_0923_)
  );
  INV_X1 _1843_ (
    .A(_0923_),
    .ZN(_0924_)
  );
  AND2_X1 _1844_ (
    .A1(_0084_),
    .A2(_0924_),
    .ZN(_0925_)
  );
  INV_X1 _1845_ (
    .A(_0925_),
    .ZN(_0926_)
  );
  AND2_X1 _1846_ (
    .A1(_0297_),
    .A2(_0926_),
    .ZN(_0927_)
  );
  AND2_X1 _1847_ (
    .A1(_0922_),
    .A2(_0927_),
    .ZN(_0929_)
  );
  INV_X1 _1848_ (
    .A(_0929_),
    .ZN(_0930_)
  );
  AND2_X1 _1849_ (
    .A1(_0903_),
    .A2(_0930_),
    .ZN(io_out_rd[0])
  );
  AND2_X1 _1850_ (
    .A1(io_in[8]),
    .A2(_0454_),
    .ZN(_0931_)
  );
  INV_X1 _1851_ (
    .A(_0931_),
    .ZN(_0932_)
  );
  AND2_X1 _1852_ (
    .A1(io_in[8]),
    .A2(_0182_),
    .ZN(_0933_)
  );
  INV_X1 _1853_ (
    .A(_0933_),
    .ZN(_0934_)
  );
  MUX2_X1 _1854_ (
    .A(io_in[3]),
    .B(io_in[8]),
    .S(_0158_),
    .Z(_0935_)
  );
  AND2_X1 _1855_ (
    .A1(_0391_),
    .A2(_0935_),
    .ZN(_0936_)
  );
  INV_X1 _1856_ (
    .A(_0936_),
    .ZN(_0937_)
  );
  AND2_X1 _1857_ (
    .A1(_0384_),
    .A2(_0937_),
    .ZN(_0939_)
  );
  INV_X1 _1858_ (
    .A(_0939_),
    .ZN(_0940_)
  );
  AND2_X1 _1859_ (
    .A1(_0304_),
    .A2(_0940_),
    .ZN(_0941_)
  );
  INV_X1 _1860_ (
    .A(_0941_),
    .ZN(_0942_)
  );
  AND2_X1 _1861_ (
    .A1(_0934_),
    .A2(_0942_),
    .ZN(_0943_)
  );
  INV_X1 _1862_ (
    .A(_0943_),
    .ZN(_0944_)
  );
  AND2_X1 _1863_ (
    .A1(_0234_),
    .A2(_0944_),
    .ZN(_0945_)
  );
  INV_X1 _1864_ (
    .A(_0945_),
    .ZN(_0946_)
  );
  AND2_X1 _1865_ (
    .A1(_0382_),
    .A2(_0946_),
    .ZN(_0947_)
  );
  INV_X1 _1866_ (
    .A(_0947_),
    .ZN(_0948_)
  );
  AND2_X1 _1867_ (
    .A1(_0427_),
    .A2(_0948_),
    .ZN(_0950_)
  );
  INV_X1 _1868_ (
    .A(_0950_),
    .ZN(_0951_)
  );
  AND2_X1 _1869_ (
    .A1(_0932_),
    .A2(_0951_),
    .ZN(_0952_)
  );
  INV_X1 _1870_ (
    .A(_0952_),
    .ZN(io_out_rd[1])
  );
  AND2_X1 _1871_ (
    .A1(io_in[9]),
    .A2(_0454_),
    .ZN(_0953_)
  );
  INV_X1 _1872_ (
    .A(_0953_),
    .ZN(_0954_)
  );
  AND2_X1 _1873_ (
    .A1(io_in[9]),
    .A2(_0182_),
    .ZN(_0955_)
  );
  INV_X1 _1874_ (
    .A(_0955_),
    .ZN(_0956_)
  );
  MUX2_X1 _1875_ (
    .A(io_in[4]),
    .B(io_in[9]),
    .S(_0158_),
    .Z(_0957_)
  );
  AND2_X1 _1876_ (
    .A1(_0391_),
    .A2(_0957_),
    .ZN(_0958_)
  );
  INV_X1 _1877_ (
    .A(_0958_),
    .ZN(_0000_)
  );
  AND2_X1 _1878_ (
    .A1(_0413_),
    .A2(_0000_),
    .ZN(_0001_)
  );
  INV_X1 _1879_ (
    .A(_0001_),
    .ZN(_0002_)
  );
  AND2_X1 _1880_ (
    .A1(_0304_),
    .A2(_0002_),
    .ZN(_0003_)
  );
  INV_X1 _1881_ (
    .A(_0003_),
    .ZN(_0004_)
  );
  AND2_X1 _1882_ (
    .A1(_0956_),
    .A2(_0004_),
    .ZN(_0005_)
  );
  INV_X1 _1883_ (
    .A(_0005_),
    .ZN(_0006_)
  );
  AND2_X1 _1884_ (
    .A1(_0234_),
    .A2(_0006_),
    .ZN(_0007_)
  );
  INV_X1 _1885_ (
    .A(_0007_),
    .ZN(_0008_)
  );
  AND2_X1 _1886_ (
    .A1(_0411_),
    .A2(_0008_),
    .ZN(_0009_)
  );
  INV_X1 _1887_ (
    .A(_0009_),
    .ZN(_0011_)
  );
  AND2_X1 _1888_ (
    .A1(_0427_),
    .A2(_0011_),
    .ZN(_0012_)
  );
  INV_X1 _1889_ (
    .A(_0012_),
    .ZN(_0013_)
  );
  AND2_X1 _1890_ (
    .A1(_0954_),
    .A2(_0013_),
    .ZN(_0014_)
  );
  INV_X1 _1891_ (
    .A(_0014_),
    .ZN(io_out_rd[2])
  );
  AND2_X1 _1892_ (
    .A1(_0169_),
    .A2(_0185_),
    .ZN(_0015_)
  );
  AND2_X1 _1893_ (
    .A1(_0100_),
    .A2(_0015_),
    .ZN(_0016_)
  );
  INV_X1 _1894_ (
    .A(_0016_),
    .ZN(_0017_)
  );
  AND2_X1 _1895_ (
    .A1(_0449_),
    .A2(_0017_),
    .ZN(_0018_)
  );
  INV_X1 _1896_ (
    .A(_0018_),
    .ZN(_0019_)
  );
  AND2_X1 _1897_ (
    .A1(_0107_),
    .A2(_0160_),
    .ZN(_0021_)
  );
  AND2_X1 _1898_ (
    .A1(_0297_),
    .A2(_0021_),
    .ZN(_0022_)
  );
  INV_X1 _1899_ (
    .A(_0022_),
    .ZN(_0023_)
  );
  AND2_X1 _1900_ (
    .A1(_0823_),
    .A2(_0023_),
    .ZN(_0024_)
  );
  INV_X1 _1901_ (
    .A(_0024_),
    .ZN(_0025_)
  );
  AND2_X1 _1902_ (
    .A1(_0019_),
    .A2(_0025_),
    .ZN(io_out_rd[3])
  );
  AND2_X1 _1903_ (
    .A1(_0453_),
    .A2(_0021_),
    .ZN(_0026_)
  );
  INV_X1 _1904_ (
    .A(_0026_),
    .ZN(_0027_)
  );
  AND2_X1 _1905_ (
    .A1(io_in[11]),
    .A2(_0027_),
    .ZN(io_out_rd[4])
  );
  AND2_X1 _1906_ (
    .A1(_0153_),
    .A2(_0660_),
    .ZN(_0028_)
  );
  INV_X1 _1907_ (
    .A(_0028_),
    .ZN(_0030_)
  );
  AND2_X1 _1908_ (
    .A1(_0392_),
    .A2(_0660_),
    .ZN(_0031_)
  );
  INV_X1 _1909_ (
    .A(_0031_),
    .ZN(_0032_)
  );
  AND2_X1 _1910_ (
    .A1(io_in[7]),
    .A2(_0032_),
    .ZN(_0033_)
  );
  INV_X1 _1911_ (
    .A(_0033_),
    .ZN(_0034_)
  );
  AND2_X1 _1912_ (
    .A1(_0522_),
    .A2(_0034_),
    .ZN(_0035_)
  );
  INV_X1 _1913_ (
    .A(_0035_),
    .ZN(io_out_rs1[0])
  );
  MUX2_X1 _1914_ (
    .A(_0801_),
    .B(_0541_),
    .S(_0171_),
    .Z(_0036_)
  );
  INV_X1 _1915_ (
    .A(_0036_),
    .ZN(_0037_)
  );
  AND2_X1 _1916_ (
    .A1(io_in[8]),
    .A2(_0030_),
    .ZN(_0038_)
  );
  INV_X1 _1917_ (
    .A(_0038_),
    .ZN(_0040_)
  );
  AND2_X1 _1918_ (
    .A1(_0156_),
    .A2(_0660_),
    .ZN(_0041_)
  );
  INV_X1 _1919_ (
    .A(_0041_),
    .ZN(_0042_)
  );
  AND2_X1 _1920_ (
    .A1(_0040_),
    .A2(_0042_),
    .ZN(_0043_)
  );
  INV_X1 _1921_ (
    .A(_0043_),
    .ZN(_0044_)
  );
  AND2_X1 _1922_ (
    .A1(_0037_),
    .A2(_0044_),
    .ZN(_0045_)
  );
  AND2_X1 _1923_ (
    .A1(_0100_),
    .A2(_0045_),
    .ZN(_0046_)
  );
  INV_X1 _1924_ (
    .A(_0046_),
    .ZN(_0047_)
  );
  AND2_X1 _1925_ (
    .A1(_0533_),
    .A2(_0047_),
    .ZN(_0048_)
  );
  INV_X1 _1926_ (
    .A(_0048_),
    .ZN(_0049_)
  );
  MUX2_X1 _1927_ (
    .A(io_in[16]),
    .B(_0049_),
    .S(io_rvc),
    .Z(io_out_rs1[1])
  );
  AND2_X1 _1928_ (
    .A1(io_in[9]),
    .A2(_0032_),
    .ZN(_0051_)
  );
  INV_X1 _1929_ (
    .A(_0051_),
    .ZN(_0052_)
  );
  AND2_X1 _1930_ (
    .A1(_0564_),
    .A2(_0052_),
    .ZN(_0053_)
  );
  INV_X1 _1931_ (
    .A(_0053_),
    .ZN(io_out_rs1[2])
  );
  AND2_X1 _1932_ (
    .A1(io_in[10]),
    .A2(_0393_),
    .ZN(_0054_)
  );
  INV_X1 _1933_ (
    .A(_0054_),
    .ZN(_0055_)
  );
  AND2_X1 _1934_ (
    .A1(_0204_),
    .A2(_0299_),
    .ZN(_0056_)
  );
  AND2_X1 _1935_ (
    .A1(_0592_),
    .A2(_0056_),
    .ZN(_0057_)
  );
  AND2_X1 _1936_ (
    .A1(_0055_),
    .A2(_0057_),
    .ZN(_0058_)
  );
  AND2_X1 _1937_ (
    .A1(_0587_),
    .A2(_0058_),
    .ZN(_0060_)
  );
  AND2_X1 _1938_ (
    .A1(_0584_),
    .A2(_0060_),
    .ZN(_0061_)
  );
  INV_X1 _1939_ (
    .A(_0061_),
    .ZN(io_out_rs1[3])
  );
  AND2_X1 _1940_ (
    .A1(_0601_),
    .A2(_0606_),
    .ZN(_0062_)
  );
  AND2_X1 _1941_ (
    .A1(io_in[11]),
    .A2(_0393_),
    .ZN(_0063_)
  );
  INV_X1 _1942_ (
    .A(_0063_),
    .ZN(_0064_)
  );
  AND2_X1 _1943_ (
    .A1(_0608_),
    .A2(_0064_),
    .ZN(_0065_)
  );
  AND2_X1 _1944_ (
    .A1(_0062_),
    .A2(_0065_),
    .ZN(_0066_)
  );
  INV_X1 _1945_ (
    .A(_0066_),
    .ZN(io_out_rs1[4])
  );
  AND2_X1 _1946_ (
    .A1(io_in[2]),
    .A2(_0675_),
    .ZN(_0067_)
  );
  INV_X1 _1947_ (
    .A(_0067_),
    .ZN(_0069_)
  );
  AND2_X1 _1948_ (
    .A1(_0624_),
    .A2(_0069_),
    .ZN(_0070_)
  );
  INV_X1 _1949_ (
    .A(_0070_),
    .ZN(io_out_rs2[0])
  );
  AND2_X1 _1950_ (
    .A1(io_in[3]),
    .A2(_0675_),
    .ZN(_0071_)
  );
  INV_X1 _1951_ (
    .A(_0071_),
    .ZN(_0072_)
  );
  AND2_X1 _1952_ (
    .A1(_0637_),
    .A2(_0072_),
    .ZN(_0073_)
  );
  INV_X1 _1953_ (
    .A(_0073_),
    .ZN(io_out_rs2[1])
  );
  AND2_X1 _1954_ (
    .A1(_0938_),
    .A2(_0643_),
    .ZN(_0074_)
  );
  INV_X1 _1955_ (
    .A(_0074_),
    .ZN(_0075_)
  );
  AND2_X1 _1956_ (
    .A1(io_in[4]),
    .A2(_0294_),
    .ZN(_0076_)
  );
  AND2_X1 _1957_ (
    .A1(_0186_),
    .A2(_0076_),
    .ZN(_0078_)
  );
  INV_X1 _1958_ (
    .A(_0078_),
    .ZN(_0079_)
  );
  AND2_X1 _1959_ (
    .A1(_0645_),
    .A2(_0079_),
    .ZN(_0080_)
  );
  INV_X1 _1960_ (
    .A(_0080_),
    .ZN(_0081_)
  );
  AND2_X1 _1961_ (
    .A1(_0075_),
    .A2(_0081_),
    .ZN(io_out_rs2[2])
  );
  MUX2_X1 _1962_ (
    .A(_0186_),
    .B(io_in[5]),
    .S(_0646_),
    .Z(_0082_)
  );
  MUX2_X1 _1963_ (
    .A(io_in[23]),
    .B(_0082_),
    .S(io_rvc),
    .Z(io_out_rs2[3])
  );
  assign _GEN_0 = { 5'h00, io_in[12], io_in[6:2], 2'h1, io_in[9:7], 5'h15, io_in[9:7], 7'h13 };
  assign { _GEN_1[30:15], _GEN_1[11:0] } = { 8'h01, io_in[4:2], 2'h1, io_in[9:7], 2'h1, io_in[9:7], 3'h3, io_in[12], 3'h3 };
  assign { _io_out_T_10_bits[31:30], _io_out_T_10_bits[25], _io_out_T_10_bits[19], _io_out_T_10_bits[14:13], _io_out_T_10_bits[6], _io_out_T_10_bits[1:0] } = { 2'h0, io_in[12], 2'h0, _io_out_T_10_bits[18], 3'h3 };
  assign _io_out_T_10_rd = { 2'h1, io_in[4:2] };
  assign _io_out_T_10_rs1 = { 1'h0, _io_out_T_10_bits[18:15] };
  assign { _io_out_T_12_bits[31:30], _io_out_T_12_bits[25], _io_out_T_12_bits[19], _io_out_T_12_bits[14:13], _io_out_T_12_bits[6], _io_out_T_12_bits[1:0] } = { 2'h0, io_in[12], 2'h0, _io_out_T_12_bits[18], 3'h3 };
  assign _io_out_T_12_rd = { 2'h1, io_in[4:2] };
  assign _io_out_T_12_rs1 = { 1'h0, _io_out_T_12_bits[18:15] };
  assign { _io_out_T_14_bits[31:30], _io_out_T_14_bits[25], _io_out_T_14_bits[19], _io_out_T_14_bits[14:13], _io_out_T_14_bits[6], _io_out_T_14_bits[1:0] } = { 2'h0, io_in[12], 2'h0, _io_out_T_14_bits[18], 3'h3 };
  assign _io_out_T_14_rd = { 2'h1, io_in[4:2] };
  assign _io_out_T_14_rs1 = { 1'h0, _io_out_T_14_bits[18:15] };
  assign { _io_out_T_16_bits[31:30], _io_out_T_16_bits[25], _io_out_T_16_bits[19], _io_out_T_16_bits[14:13], _io_out_T_16_bits[6], _io_out_T_16_bits[1:0] } = { 2'h0, io_in[12], 2'h0, _io_out_T_16_bits[18], 3'h3 };
  assign _io_out_T_16_rd = { 2'h1, io_in[4:2] };
  assign _io_out_T_16_rs1 = { 1'h0, _io_out_T_16_bits[18:15] };
  assign { _io_out_T_18_bits[30], _io_out_T_18_bits[25], _io_out_T_18_bits[14], _io_out_T_18_bits[6], _io_out_T_18_bits[1:0] } = { _io_out_T_18_bits[31], io_in[12], 4'h3 };
  assign _io_out_T_18_rd[4] = _io_out_T_18_bits[19];
  assign _io_out_T_18_rs1 = _io_out_T_18_bits[19:15];
  assign _io_out_T_18_rs2 = { 2'h1, io_in[4:2] };
  assign _io_out_T_2 = { io_in[1:0], io_in[15:13] };
  assign _io_out_T_20_bits[1:0] = 2'h3;
  assign _io_out_T_20_rs2 = { 2'h1, io_in[4:2] };
  assign _io_out_T_22_bits[1:0] = 2'h3;
  assign _io_out_T_22_rs2 = { 2'h1, io_in[4:2] };
  assign _io_out_T_24_bits[1:0] = 2'h3;
  assign _io_out_T_24_rs2 = { 2'h1, io_in[4:2] };
  assign _io_out_T_26_bits[1:0] = 2'h3;
  assign _io_out_T_26_rs2 = { 2'h1, io_in[4:2] };
  assign _io_out_T_28_bits[1:0] = 2'h3;
  assign _io_out_T_28_rs2 = { 2'h1, io_in[4:2] };
  assign _io_out_T_30_bits[1:0] = 2'h3;
  assign _io_out_T_30_rs2[4] = 1'h0;
  assign _io_out_T_32_bits[1:0] = 2'h3;
  assign _io_out_T_32_rs2[4] = 1'h0;
  assign _io_out_T_34_bits[1:0] = 2'h3;
  assign _io_out_T_36_bits[1:0] = 2'h3;
  assign _io_out_T_38_bits[1:0] = 2'h3;
  assign _io_out_T_40_bits[1:0] = 2'h3;
  assign _io_out_T_42_bits[1:0] = 2'h3;
  assign _io_out_T_44_bits[1:0] = 2'h3;
  assign _io_out_T_46_bits[1:0] = 2'h3;
  assign _io_out_T_48_bits[1:0] = 2'h3;
  assign { _io_out_T_4_bits[31:30], _io_out_T_4_bits[25:24], _io_out_T_4_bits[21:19], _io_out_T_4_bits[14:5], _io_out_T_4_bits[1:0] } = { 2'h0, io_in[12:11], 4'h0, _io_out_T_4_bits[18], _io_out_T_4_bits[18], 2'h1, io_in[4:2], 4'h3 };
  assign _io_out_T_4_rd = { 2'h1, io_in[4:2] };
  assign _io_out_T_4_rs1 = { 1'h0, _io_out_T_4_bits[18:15] };
  assign { _io_out_T_6_bits[31:30], _io_out_T_6_bits[25:24], _io_out_T_6_bits[21:19], _io_out_T_6_bits[14:13], _io_out_T_6_bits[11:5], _io_out_T_6_bits[1:0] } = { 2'h0, io_in[12:11], 4'h0, _io_out_T_6_bits[18], 2'h1, io_in[4:2], 4'h3 };
  assign _io_out_T_6_rd = { 2'h1, io_in[4:2] };
  assign _io_out_T_6_rs1 = { 1'h0, _io_out_T_6_bits[18:15] };
  assign { _io_out_T_8_bits[31:30], _io_out_T_8_bits[25:24], _io_out_T_8_bits[21:19], _io_out_T_8_bits[14:13], _io_out_T_8_bits[11:5], _io_out_T_8_bits[1:0] } = { 2'h0, io_in[12:11], 4'h0, _io_out_T_8_bits[18], 2'h1, io_in[4:2], 4'h3 };
  assign _io_out_T_8_rd = { 2'h1, io_in[4:2] };
  assign _io_out_T_8_rs1 = { 1'h0, _io_out_T_8_bits[18:15] };
  assign _io_out_s_T_116 = { io_in[5], io_in[12], 2'h1, io_in[4:2], 2'h1, io_in[9:7], 3'h2, io_in[11:10], io_in[6], 9'h023 };
  assign _io_out_s_T_138 = { io_in[5], io_in[12], 2'h1, io_in[4:2], 2'h1, io_in[9:7], 3'h2, io_in[11:10], io_in[6], 9'h027 };
  assign _io_out_s_T_148 = { io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12] };
  assign _io_out_s_T_15 = { io_in[6:5], io_in[12:10], 3'h0 };
  assign _io_out_s_T_150 = { io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[6:2] };
  assign _io_out_s_T_161 = { io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12] };
  assign _io_out_s_T_169 = { io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[8], io_in[10:9], io_in[6], io_in[7], io_in[2], io_in[11], io_in[5:3], 1'h0 };
  assign _io_out_s_T_17 = { 2'h1, io_in[9:7] };
  assign _io_out_s_T_20 = { io_in[6:5], io_in[12:10], 5'h01, io_in[9:7], 5'h0d, io_in[4:2], 7'h07 };
  assign _io_out_s_T_230 = { io_in[12], io_in[12], io_in[12] };
  assign _io_out_s_T_251 = { io_in[12], io_in[6:2], 2'h1, io_in[9:7], 5'h15, io_in[9:7], 7'h13 };
  assign _io_out_s_T_260 = { 5'h10, io_in[12], io_in[6:2], 2'h1, io_in[9:7], 5'h15, io_in[9:7], 7'h13 };
  assign _io_out_s_T_270 = { io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[6:2], 2'h1, io_in[9:7], 5'h1d, io_in[9:7], 7'h13 };
  assign _io_out_s_T_277 = { 2'h1, io_in[4:2], 2'h1, io_in[9:7], _GEN_1[14:12], 2'h1, io_in[9:7], 3'h3, io_in[12], 3'h3 };
  assign _io_out_s_T_278[29:0] = { 7'h01, io_in[4:2], 2'h1, io_in[9:7], _GEN_1[14:12], 2'h1, io_in[9:7], 3'h3, io_in[12], 3'h3 };
  assign _io_out_s_T_281[29:0] = { 4'h0, io_in[12], io_in[6:2], 2'h1, io_in[9:7], 5'h15, io_in[9:7], 7'h13 };
  assign { _io_out_s_T_283[29:14], _io_out_s_T_283[12:0] } = { _io_out_s_T_283[31], _io_out_s_T_283[31], _io_out_s_T_283[31], _io_out_s_T_283[31], io_in[12], io_in[6:2], 2'h1, io_in[9:7], 4'hd, io_in[9:7], 7'h13 };
  assign _io_out_s_T_31 = { io_in[5], io_in[12:10], io_in[6], 2'h0 };
  assign _io_out_s_T_349 = { io_in[12], io_in[12], io_in[12], io_in[12], io_in[12] };
  assign _io_out_s_T_354 = { io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[6:5], io_in[2], io_in[11:10], io_in[4:3], 1'h0 };
  assign _io_out_s_T_36 = { io_in[5], io_in[12:10], io_in[6], 4'h1, io_in[9:7], 5'h09, io_in[4:2], 7'h03 };
  assign _io_out_s_T_438 = { io_in[12], io_in[6:2], io_in[11:7], 3'h1, io_in[11:7], 7'h13 };
  assign _io_out_s_T_448 = { io_in[4:2], io_in[12], io_in[6:5], 11'h013, io_in[11:7], 7'h07 };
  assign { _io_out_s_T_457[27:5], _io_out_s_T_457[3:0] } = { io_in[3:2], io_in[12], io_in[6:4], 10'h012, io_in[11:7], 2'h0, _io_out_s_T_457[4], _io_out_s_T_457[4], 2'h3 };
  assign _io_out_s_T_466 = { io_in[3:2], io_in[12], io_in[6:4], 10'h012, io_in[11:7], 7'h07 };
  assign _io_out_s_T_473 = { io_in[9:7], io_in[12:10], 3'h0 };
  assign _io_out_s_T_480 = { io_in[9:7], io_in[12], io_in[6:2], 8'h13, io_in[11:10], 10'h027 };
  assign _io_out_s_T_486 = { io_in[8:7], io_in[12:9], 2'h0 };
  assign _io_out_s_T_493 = { io_in[8:7], io_in[12], io_in[6:2], 8'h12, io_in[11:9], 9'h023 };
  assign _io_out_s_T_506 = { io_in[8:7], io_in[12], io_in[6:2], 8'h12, io_in[11:9], 9'h027 };
  assign _io_out_s_T_52 = { io_in[5], io_in[12:10], io_in[6], 4'h1, io_in[9:7], 5'h09, io_in[4:2], 7'h07 };
  assign _io_out_s_T_6 = { 2'h1, io_in[4:2] };
  assign { _io_out_s_T_7[29:4], _io_out_s_T_7[2:0] } = { io_in[10:7], io_in[12:11], io_in[5], io_in[6], 12'h041, io_in[4:2], 3'h1, _io_out_s_T_7[3], 2'h3 };
  assign _io_out_s_T_74 = { io_in[5], io_in[12], 2'h1, io_in[4:2], 2'h1, io_in[9:7], 3'h2, io_in[11:10], io_in[6], 9'h03f };
  assign _io_out_s_T_94 = { io_in[6:5], io_in[12], 2'h1, io_in[4:2], 2'h1, io_in[9:7], 3'h3, io_in[11:10], 10'h027 };
  assign _io_out_s_add_T_3 = { io_in[6:2], io_in[11:7], 3'h0, io_in[11:7], 7'h33 };
  assign _io_out_s_ebreak_T_1 = { io_in[6:2], io_in[11:7], 15'h0073 };
  assign _io_out_s_funct_T_2 = { io_in[12], io_in[6:5] };
  assign _io_out_s_funct_T_4[1:0] = 2'h0;
  assign _io_out_s_funct_T_6[0] = 1'h0;
  assign { _io_out_s_jalr_ebreak_T_2[24:21], _io_out_s_jalr_ebreak_T_2[19:8], _io_out_s_jalr_ebreak_T_2[6:0] } = { io_in[6:3], io_in[11:7], 9'h003, _io_out_s_T_457[4], 1'h0, _io_out_s_jalr_ebreak_T_2[7], 2'h3 };
  assign _io_out_s_jr_reserved_T_2 = { io_in[6:2], io_in[11:7], 8'h00, _io_out_s_jalr_ebreak_T_2[7], _io_out_s_jalr_ebreak_T_2[7], _io_out_s_T_457[4], _io_out_s_T_457[4], 3'h7 };
  assign _io_out_s_load_opc_T_1 = _io_out_s_jalr_ebreak_T_2[7];
  assign _io_out_s_me_T_2 = { io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12] };
  assign _io_out_s_me_T_4 = { io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[6:2], 12'h000 };
  assign _io_out_s_mv_T_2 = { io_in[6:2], 8'h00, io_in[11:7], 7'h33 };
  assign io_out_bits[1:0] = 2'h3;
  assign io_out_s_0_bits = { 2'h0, io_in[10:7], io_in[12:11], io_in[5], io_in[6], 12'h041, io_in[4:2], 3'h1, _io_out_s_T_7[3], _io_out_s_T_7[3], 2'h3 };
  assign io_out_s_10_bits = { io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[6:2], 8'h00, io_in[11:7], 7'h13 };
  assign { io_out_s_11_bits[31:29], io_out_s_11_bits[22:20], io_out_s_11_bits[11:6], io_out_s_11_bits[4], io_out_s_11_bits[1:0] } = { io_in[12], io_in[12], io_in[12], io_out_s_11_bits[23], io_out_s_11_bits[23], io_out_s_11_bits[23], io_in[11:7], 4'h7 };
  assign io_out_s_11_rd = io_in[11:7];
  assign io_out_s_11_rs2 = { 2'h1, io_in[4:2] };
  assign { io_out_s_12_bits[29:26], io_out_s_12_bits[22:15], io_out_s_12_bits[11:6], io_out_s_12_bits[4], io_out_s_12_bits[2:0] } = { io_out_s_12_bits[31], io_out_s_12_bits[31], io_out_s_12_bits[31], io_out_s_12_bits[31], io_in[4:2], 2'h1, io_in[9:7], 2'h1, io_in[9:7], 5'h0b };
  assign io_out_s_13_bits = { io_in[12], io_in[8], io_in[10:9], io_in[6], io_in[7], io_in[2], io_in[11], io_in[5:3], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], 12'h06f };
  assign io_out_s_14_bits = { io_in[12], io_in[12], io_in[12], io_in[12], io_in[6:5], io_in[2], 7'h01, io_in[9:7], 3'h0, io_in[11:10], io_in[4:3], io_in[12], 7'h63 };
  assign io_out_s_15_bits = { io_in[12], io_in[12], io_in[12], io_in[12], io_in[6:5], io_in[2], 7'h01, io_in[9:7], 3'h1, io_in[11:10], io_in[4:3], io_in[12], 7'h63 };
  assign io_out_s_16_bits = { 6'h00, io_in[12], io_in[6:2], io_in[11:7], 3'h1, io_in[11:7], 7'h13 };
  assign io_out_s_17_bits = { 3'h0, io_in[4:2], io_in[12], io_in[6:5], 11'h013, io_in[11:7], 7'h07 };
  assign io_out_s_18_bits = { 4'h0, io_in[3:2], io_in[12], io_in[6:4], 10'h012, io_in[11:7], 2'h0, _io_out_s_T_457[4], _io_out_s_T_457[4], _io_out_s_T_457[4], 2'h3 };
  assign io_out_s_19_bits = { 4'h0, io_in[3:2], io_in[12], io_in[6:4], 10'h012, io_in[11:7], 7'h07 };
  assign io_out_s_1_bits = { 4'h0, io_in[6:5], io_in[12:10], 5'h01, io_in[9:7], 5'h0d, io_in[4:2], 7'h07 };
  assign { io_out_s_20_bits[31:21], io_out_s_20_bits[14:12], io_out_s_20_bits[1:0] } = { 7'h00, io_in[6:3], 5'h03 };
  assign io_out_s_20_rd[4:1] = io_out_s_20_bits[11:8];
  assign io_out_s_20_rs1 = io_out_s_20_bits[19:15];
  assign io_out_s_20_rs2 = io_in[6:2];
  assign io_out_s_21_bits = { 3'h0, io_in[9:7], io_in[12], io_in[6:2], 8'h13, io_in[11:10], 10'h027 };
  assign io_out_s_22_bits = { 4'h0, io_in[8:7], io_in[12], io_in[6:2], 8'h12, io_in[11:9], 9'h023 };
  assign io_out_s_23_bits = { 4'h0, io_in[8:7], io_in[12], io_in[6:2], 8'h12, io_in[11:9], 9'h027 };
  assign io_out_s_24_rs1 = io_in[19:15];
  assign io_out_s_24_rs2 = io_in[24:20];
  assign io_out_s_2_bits = { 5'h00, io_in[5], io_in[12:10], io_in[6], 4'h1, io_in[9:7], 5'h09, io_in[4:2], 7'h03 };
  assign io_out_s_3_bits = { 5'h00, io_in[5], io_in[12:10], io_in[6], 4'h1, io_in[9:7], 5'h09, io_in[4:2], 7'h07 };
  assign io_out_s_4_bits = { 5'h00, io_in[5], io_in[12], 2'h1, io_in[4:2], 2'h1, io_in[9:7], 3'h2, io_in[11:10], io_in[6], 9'h03f };
  assign io_out_s_5_bits = { 4'h0, io_in[6:5], io_in[12], 2'h1, io_in[4:2], 2'h1, io_in[9:7], 3'h3, io_in[11:10], 10'h027 };
  assign io_out_s_6_bits = { 5'h00, io_in[5], io_in[12], 2'h1, io_in[4:2], 2'h1, io_in[9:7], 3'h2, io_in[11:10], io_in[6], 9'h023 };
  assign io_out_s_7_bits = { 5'h00, io_in[5], io_in[12], 2'h1, io_in[4:2], 2'h1, io_in[9:7], 3'h2, io_in[11:10], io_in[6], 9'h027 };
  assign io_out_s_8_bits = { io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[6:2], io_in[11:7], 3'h0, io_in[11:7], 7'h13 };
  assign io_out_s_9_bits = { io_in[12], io_in[8], io_in[10:9], io_in[6], io_in[7], io_in[2], io_in[11], io_in[5:3], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], 12'h0ef };
  assign io_out_s_add_bits = { 7'h00, io_in[6:2], io_in[11:7], 3'h0, io_in[11:7], 7'h33 };
  assign io_out_s_ebreak = { io_in[6:3], 1'h1, io_in[11:7], 15'h0073 };
  assign io_out_s_funct = _GEN_1[14:12];
  assign io_out_s_jalr = { io_in[6:2], io_in[11:7], 15'h00e7 };
  assign { io_out_s_jalr_add_bits[31:21], io_out_s_jalr_add_bits[19:8], io_out_s_jalr_add_bits[5:3], io_out_s_jalr_add_bits[1:0] } = { 7'h00, io_in[6:3], io_in[11:7], 3'h0, io_out_s_20_bits[11:8], 1'h1, io_out_s_20_bits[4], 3'h3 };
  assign io_out_s_jalr_add_rd[4:1] = io_out_s_20_bits[11:8];
  assign io_out_s_jalr_add_rs1 = io_in[11:7];
  assign io_out_s_jalr_ebreak_bits = { 7'h00, io_in[6:3], _io_out_s_jalr_ebreak_T_2[20], io_in[11:7], 7'h00, _io_out_s_jalr_ebreak_T_2[7], 2'h3, _io_out_s_T_457[4], 1'h0, _io_out_s_jalr_ebreak_T_2[7], 2'h3 };
  assign io_out_s_jr = { io_in[6:2], io_in[11:7], 15'h0067 };
  assign { io_out_s_jr_mv_bits[31:20], io_out_s_jr_mv_bits[14:8], io_out_s_jr_mv_bits[6], io_out_s_jr_mv_bits[4], io_out_s_jr_mv_bits[2:0] } = { 7'h00, io_in[6:2], 3'h0, io_out_s_20_bits[11:8], io_out_s_jalr_add_bits[2], io_out_s_20_bits[4], io_out_s_jalr_add_bits[6], 2'h3 };
  assign io_out_s_jr_mv_rd = { io_out_s_20_bits[11:8], io_out_s_jr_mv_bits[7] };
  assign io_out_s_jr_mv_rs1 = io_out_s_jr_mv_bits[19:15];
  assign io_out_s_jr_mv_rs2 = io_in[6:2];
  assign io_out_s_jr_reserved_bits = { 7'h00, io_in[6:2], io_in[11:7], 8'h00, _io_out_s_jalr_ebreak_T_2[7], _io_out_s_jalr_ebreak_T_2[7], _io_out_s_T_457[4], _io_out_s_T_457[4], 3'h7 };
  assign io_out_s_load_opc = { 2'h0, _io_out_s_T_457[4], _io_out_s_T_457[4], _io_out_s_T_457[4], 2'h3 };
  assign io_out_s_me_bits = { io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[6:2], io_in[11:7], 3'h3, io_out_s_11_bits[3], 3'h7 };
  assign io_out_s_mv_bits = { 7'h00, io_in[6:2], 8'h00, io_in[11:7], 7'h33 };
  assign io_out_s_opc = { 3'h1, _io_out_s_T_7[3], _io_out_s_T_7[3], 2'h3 };
  assign io_out_s_opc_1 = { 3'h3, io_out_s_11_bits[3], 3'h7 };
  assign io_out_s_opc_2 = { 3'h1, io_out_s_11_bits[3], io_out_s_11_bits[3], 2'h3 };
  assign io_out_s_opc_3 = { 3'h3, io_in[12], 3'h3 };
  assign io_out_s_res_bits = { io_in[12], io_in[12], io_in[12], io_in[4:3], io_in[5], io_in[2], io_in[6], 4'h0, io_in[11:7], 3'h0, io_in[11:7], 3'h1, io_out_s_11_bits[3], io_out_s_11_bits[3], 2'h3 };
  assign io_out_s_reserved = { io_in[6:2], io_in[11:7], 15'h001f };
  assign io_out_s_sub = { _io_out_s_T_278[30], 30'h00000000 };
endmodule
module Rocket(clock, reset, io_hartid, io_interrupts_debug, io_interrupts_mtip, io_interrupts_msip, io_interrupts_meip, io_imem_might_request, io_imem_req_valid, io_imem_req_bits_pc, io_imem_req_bits_speculative, io_imem_resp_ready, io_imem_resp_valid, io_imem_resp_bits_pc, io_imem_resp_bits_data, io_imem_resp_bits_xcpt_ae_inst, io_imem_resp_bits_replay, io_imem_btb_update_valid, io_imem_bht_update_valid, io_imem_flush_icache, io_dmem_req_ready
, io_dmem_req_valid, io_dmem_req_bits_addr, io_dmem_req_bits_tag, io_dmem_req_bits_cmd, io_dmem_req_bits_size, io_dmem_req_bits_signed, io_dmem_req_bits_dv, io_dmem_s1_kill, io_dmem_s1_data_data, io_dmem_s2_nack, io_dmem_resp_valid, io_dmem_resp_bits_tag, io_dmem_resp_bits_data, io_dmem_resp_bits_replay, io_dmem_resp_bits_has_data, io_dmem_resp_bits_data_word_bypass, io_dmem_replay_next, io_dmem_s2_xcpt_ma_ld, io_dmem_s2_xcpt_ma_st, io_dmem_s2_xcpt_pf_ld, io_dmem_s2_xcpt_pf_st
, io_dmem_s2_xcpt_ae_ld, io_dmem_s2_xcpt_ae_st, io_dmem_ordered, io_dmem_perf_grant, io_ptw_status_debug, io_ptw_pmp_0_cfg_l, io_ptw_pmp_0_cfg_a, io_ptw_pmp_0_cfg_x, io_ptw_pmp_0_cfg_w, io_ptw_pmp_0_cfg_r, io_ptw_pmp_0_addr, io_ptw_pmp_0_mask, io_ptw_pmp_1_cfg_l, io_ptw_pmp_1_cfg_a, io_ptw_pmp_1_cfg_x, io_ptw_pmp_1_cfg_w, io_ptw_pmp_1_cfg_r, io_ptw_pmp_1_addr, io_ptw_pmp_1_mask, io_ptw_pmp_2_cfg_l, io_ptw_pmp_2_cfg_a
, io_ptw_pmp_2_cfg_x, io_ptw_pmp_2_cfg_w, io_ptw_pmp_2_cfg_r, io_ptw_pmp_2_addr, io_ptw_pmp_2_mask, io_ptw_pmp_3_cfg_l, io_ptw_pmp_3_cfg_a, io_ptw_pmp_3_cfg_x, io_ptw_pmp_3_cfg_w, io_ptw_pmp_3_cfg_r, io_ptw_pmp_3_addr, io_ptw_pmp_3_mask, io_ptw_pmp_4_cfg_l, io_ptw_pmp_4_cfg_a, io_ptw_pmp_4_cfg_x, io_ptw_pmp_4_cfg_w, io_ptw_pmp_4_cfg_r, io_ptw_pmp_4_addr, io_ptw_pmp_4_mask, io_ptw_pmp_5_cfg_l, io_ptw_pmp_5_cfg_a
, io_ptw_pmp_5_cfg_x, io_ptw_pmp_5_cfg_w, io_ptw_pmp_5_cfg_r, io_ptw_pmp_5_addr, io_ptw_pmp_5_mask, io_ptw_pmp_6_cfg_l, io_ptw_pmp_6_cfg_a, io_ptw_pmp_6_cfg_x, io_ptw_pmp_6_cfg_w, io_ptw_pmp_6_cfg_r, io_ptw_pmp_6_addr, io_ptw_pmp_6_mask, io_ptw_pmp_7_cfg_l, io_ptw_pmp_7_cfg_a, io_ptw_pmp_7_cfg_x, io_ptw_pmp_7_cfg_w, io_ptw_pmp_7_cfg_r, io_ptw_pmp_7_addr, io_ptw_pmp_7_mask, io_ptw_customCSRs_csrs_0_value, io_rocc_cmd_valid
, io_wfi);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire [1:0] _15563_;
  wire [1:0] _15564_;
  wire PlusArgTimeout_clock;
  wire [31:0] PlusArgTimeout_io_count;
  wire PlusArgTimeout_reset;
  wire [4:0] _T_11;
  wire [2:0] _T_113;
  wire [2:0] _T_114;
  wire [2:0] _T_115;
  wire [4:0] _T_116;
  wire [4:0] _T_118;
  wire [4:0] _T_119;
  wire [4:0] _T_12;
  wire [4:0] _T_13;
  wire [31:0] _T_143;
  wire [2:0] _T_35;
  wire [2:0] _T_37;
  wire _T_40;
  wire _T_41;
  wire _T_42;
  wire [3:0] _T_74;
  wire _T_93;
  wire [1:0] _bypass_src_T;
  wire [1:0] _bypass_src_T_2;
  wire [15:0] _csr_io_inst_0_T_3;
  wire [2:0] _csr_io_rw_cmd_T;
  wire [2:0] _csr_io_rw_cmd_T_1;
  wire _ctrl_stalld_T_15;
  wire _ex_imm_b11_T_5;
  wire _ex_imm_b11_T_8;
  wire [7:0] _ex_imm_b19_12_T_4;
  wire [10:0] _ex_imm_b30_20_T_2;
  wire _ex_imm_sign_T_2;
  wire [31:0] _ex_op1_T;
  wire [31:0] _ex_op2_T;
  wire [3:0] _ex_op2_T_1;
  wire _ex_reg_valid_T;
  wire [31:0] _ex_rs_T_13;
  wire [31:0] _ex_rs_T_6;
  wire [7:0] _id_ctrl_decoder_decoded_T;
  wire [8:0] _id_ctrl_decoder_decoded_T_10;
  wire [8:0] _id_ctrl_decoder_decoded_T_100;
  wire [8:0] _id_ctrl_decoder_decoded_T_102;
  wire [9:0] _id_ctrl_decoder_decoded_T_104;
  wire [13:0] _id_ctrl_decoder_decoded_T_106;
  wire [14:0] _id_ctrl_decoder_decoded_T_108;
  wire [14:0] _id_ctrl_decoder_decoded_T_110;
  wire [13:0] _id_ctrl_decoder_decoded_T_112;
  wire [16:0] _id_ctrl_decoder_decoded_T_114;
  wire [19:0] _id_ctrl_decoder_decoded_T_116;
  wire [27:0] _id_ctrl_decoder_decoded_T_118;
  wire [5:0] _id_ctrl_decoder_decoded_T_12;
  wire [30:0] _id_ctrl_decoder_decoded_T_120;
  wire [14:0] _id_ctrl_decoder_decoded_T_122;
  wire [12:0] _id_ctrl_decoder_decoded_T_124;
  wire [27:0] _id_ctrl_decoder_decoded_T_126;
  wire [31:0] _id_ctrl_decoder_decoded_T_128;
  wire [16:0] _id_ctrl_decoder_decoded_T_130;
  wire [12:0] _id_ctrl_decoder_decoded_T_132;
  wire [15:0] _id_ctrl_decoder_decoded_T_134;
  wire [27:0] _id_ctrl_decoder_decoded_T_136;
  wire [31:0] _id_ctrl_decoder_decoded_T_138;
  wire [6:0] _id_ctrl_decoder_decoded_T_14;
  wire [12:0] _id_ctrl_decoder_decoded_T_140;
  wire [8:0] _id_ctrl_decoder_decoded_T_16;
  wire [7:0] _id_ctrl_decoder_decoded_T_18;
  wire [7:0] _id_ctrl_decoder_decoded_T_2;
  wire [8:0] _id_ctrl_decoder_decoded_T_20;
  wire [15:0] _id_ctrl_decoder_decoded_T_22;
  wire [12:0] _id_ctrl_decoder_decoded_T_24;
  wire [7:0] _id_ctrl_decoder_decoded_T_26;
  wire [8:0] _id_ctrl_decoder_decoded_T_28;
  wire [8:0] _id_ctrl_decoder_decoded_T_30;
  wire [9:0] _id_ctrl_decoder_decoded_T_32;
  wire [6:0] _id_ctrl_decoder_decoded_T_34;
  wire [27:0] _id_ctrl_decoder_decoded_T_36;
  wire [30:0] _id_ctrl_decoder_decoded_T_38;
  wire [7:0] _id_ctrl_decoder_decoded_T_4;
  wire [9:0] _id_ctrl_decoder_decoded_T_40;
  wire [14:0] _id_ctrl_decoder_decoded_T_42;
  wire [15:0] _id_ctrl_decoder_decoded_T_44;
  wire [7:0] _id_ctrl_decoder_decoded_T_46;
  wire [8:0] _id_ctrl_decoder_decoded_T_48;
  wire [8:0] _id_ctrl_decoder_decoded_T_50;
  wire [7:0] _id_ctrl_decoder_decoded_T_52;
  wire [7:0] _id_ctrl_decoder_decoded_T_54;
  wire [8:0] _id_ctrl_decoder_decoded_T_56;
  wire [11:0] _id_ctrl_decoder_decoded_T_58;
  wire [7:0] _id_ctrl_decoder_decoded_T_6;
  wire [14:0] _id_ctrl_decoder_decoded_T_60;
  wire [15:0] _id_ctrl_decoder_decoded_T_62;
  wire [7:0] _id_ctrl_decoder_decoded_T_64;
  wire [8:0] _id_ctrl_decoder_decoded_T_66;
  wire [8:0] _id_ctrl_decoder_decoded_T_68;
  wire [14:0] _id_ctrl_decoder_decoded_T_70;
  wire [8:0] _id_ctrl_decoder_decoded_T_72;
  wire [13:0] _id_ctrl_decoder_decoded_T_74;
  wire [7:0] _id_ctrl_decoder_decoded_T_76;
  wire [14:0] _id_ctrl_decoder_decoded_T_78;
  wire [7:0] _id_ctrl_decoder_decoded_T_8;
  wire [15:0] _id_ctrl_decoder_decoded_T_80;
  wire [15:0] _id_ctrl_decoder_decoded_T_82;
  wire [15:0] _id_ctrl_decoder_decoded_T_84;
  wire [14:0] _id_ctrl_decoder_decoded_T_86;
  wire [7:0] _id_ctrl_decoder_decoded_T_88;
  wire [8:0] _id_ctrl_decoder_decoded_T_90;
  wire [8:0] _id_ctrl_decoder_decoded_T_92;
  wire [8:0] _id_ctrl_decoder_decoded_T_94;
  wire [14:0] _id_ctrl_decoder_decoded_T_96;
  wire [7:0] _id_ctrl_decoder_decoded_T_98;
  wire _id_illegal_insn_T_11;
  wire _id_illegal_insn_T_15;
  wire _id_illegal_insn_T_33;
  wire [31:0] _io_fpu_time_T;
  wire [31:0] _mem_br_target_T_3;
  wire [31:0] _mem_br_target_T_5;
  wire [3:0] _mem_br_target_T_6;
  wire [31:0] _mem_br_target_T_7;
  wire [31:0] _mem_br_target_T_8;
  wire _mem_reg_load_T_1;
  wire [31:0] _mem_reg_rs2_T_3;
  wire [31:0] _mem_reg_rs2_T_6;
  wire [31:0] _mem_reg_rs2_T_7;
  wire _mem_reg_valid_T;
  wire [31:0] _mem_reg_wdata_T;
  wire [31:0] _r;
  wire _take_pc_mem_T;
  wire _wb_reg_replay_T;
  wire _wb_reg_valid_T;
  wire [31:0] alu_io_adder_out;
  wire alu_io_cmp_out;
  wire [3:0] alu_io_fn;
  wire [31:0] alu_io_in1;
  wire [31:0] alu_io_in2;
  wire [31:0] alu_io_out;
  wire blocked;
  wire [31:0] bpu_io_bp_0_address;
  wire bpu_io_bp_0_control_action;
  wire bpu_io_bp_0_control_r;
  wire [1:0] bpu_io_bp_0_control_tmatch;
  wire bpu_io_bp_0_control_w;
  wire bpu_io_bp_0_control_x;
  wire bpu_io_debug_if;
  wire bpu_io_debug_ld;
  wire bpu_io_debug_st;
  wire [31:0] bpu_io_ea;
  wire [31:0] bpu_io_pc;
  wire bpu_io_status_debug;
  wire bpu_io_xcpt_if;
  wire bpu_io_xcpt_ld;
  wire bpu_io_xcpt_st;
  input clock;
  wire clock;
  wire [31:0] coreMonitorBundle_inst;
  wire [31:0] coreMonitorBundle_pc;
  wire csr_clock;
  wire [31:0] csr_io_bp_0_address;
  wire csr_io_bp_0_control_action;
  wire csr_io_bp_0_control_r;
  wire [1:0] csr_io_bp_0_control_tmatch;
  wire csr_io_bp_0_control_w;
  wire csr_io_bp_0_control_x;
  wire [31:0] csr_io_cause;
  wire csr_io_csr_stall;
  wire [31:0] csr_io_customCSRs_0_value;
  wire csr_io_decode_0_fp_csr;
  wire csr_io_decode_0_fp_illegal;
  wire [31:0] csr_io_decode_0_inst;
  wire csr_io_decode_0_read_illegal;
  wire csr_io_decode_0_rocc_illegal;
  wire csr_io_decode_0_system_illegal;
  wire csr_io_decode_0_write_flush;
  wire csr_io_decode_0_write_illegal;
  wire csr_io_eret;
  wire [31:0] csr_io_evec;
  wire csr_io_exception;
  wire csr_io_gva;
  wire csr_io_hartid;
  wire csr_io_inhibit_cycle;
  wire [31:0] csr_io_inst_0;
  wire csr_io_interrupt;
  wire [31:0] csr_io_interrupt_cause;
  wire csr_io_interrupts_debug;
  wire csr_io_interrupts_meip;
  wire csr_io_interrupts_msip;
  wire csr_io_interrupts_mtip;
  wire [31:0] csr_io_pc;
  wire [29:0] csr_io_pmp_0_addr;
  wire [1:0] csr_io_pmp_0_cfg_a;
  wire csr_io_pmp_0_cfg_l;
  wire csr_io_pmp_0_cfg_r;
  wire csr_io_pmp_0_cfg_w;
  wire csr_io_pmp_0_cfg_x;
  wire [31:0] csr_io_pmp_0_mask;
  wire [29:0] csr_io_pmp_1_addr;
  wire [1:0] csr_io_pmp_1_cfg_a;
  wire csr_io_pmp_1_cfg_l;
  wire csr_io_pmp_1_cfg_r;
  wire csr_io_pmp_1_cfg_w;
  wire csr_io_pmp_1_cfg_x;
  wire [31:0] csr_io_pmp_1_mask;
  wire [29:0] csr_io_pmp_2_addr;
  wire [1:0] csr_io_pmp_2_cfg_a;
  wire csr_io_pmp_2_cfg_l;
  wire csr_io_pmp_2_cfg_r;
  wire csr_io_pmp_2_cfg_w;
  wire csr_io_pmp_2_cfg_x;
  wire [31:0] csr_io_pmp_2_mask;
  wire [29:0] csr_io_pmp_3_addr;
  wire [1:0] csr_io_pmp_3_cfg_a;
  wire csr_io_pmp_3_cfg_l;
  wire csr_io_pmp_3_cfg_r;
  wire csr_io_pmp_3_cfg_w;
  wire csr_io_pmp_3_cfg_x;
  wire [31:0] csr_io_pmp_3_mask;
  wire [29:0] csr_io_pmp_4_addr;
  wire [1:0] csr_io_pmp_4_cfg_a;
  wire csr_io_pmp_4_cfg_l;
  wire csr_io_pmp_4_cfg_r;
  wire csr_io_pmp_4_cfg_w;
  wire csr_io_pmp_4_cfg_x;
  wire [31:0] csr_io_pmp_4_mask;
  wire [29:0] csr_io_pmp_5_addr;
  wire [1:0] csr_io_pmp_5_cfg_a;
  wire csr_io_pmp_5_cfg_l;
  wire csr_io_pmp_5_cfg_r;
  wire csr_io_pmp_5_cfg_w;
  wire csr_io_pmp_5_cfg_x;
  wire [31:0] csr_io_pmp_5_mask;
  wire [29:0] csr_io_pmp_6_addr;
  wire [1:0] csr_io_pmp_6_cfg_a;
  wire csr_io_pmp_6_cfg_l;
  wire csr_io_pmp_6_cfg_r;
  wire csr_io_pmp_6_cfg_w;
  wire csr_io_pmp_6_cfg_x;
  wire [31:0] csr_io_pmp_6_mask;
  wire [29:0] csr_io_pmp_7_addr;
  wire [1:0] csr_io_pmp_7_cfg_a;
  wire csr_io_pmp_7_cfg_l;
  wire csr_io_pmp_7_cfg_r;
  wire csr_io_pmp_7_cfg_w;
  wire csr_io_pmp_7_cfg_x;
  wire [31:0] csr_io_pmp_7_mask;
  wire csr_io_retire;
  wire [11:0] csr_io_rw_addr;
  wire [2:0] csr_io_rw_cmd;
  wire [31:0] csr_io_rw_rdata;
  wire [31:0] csr_io_rw_wdata;
  wire csr_io_singleStep;
  wire csr_io_status_cease;
  wire csr_io_status_debug;
  wire [1:0] csr_io_status_dprv;
  wire csr_io_status_dv;
  wire [1:0] csr_io_status_fs;
  wire csr_io_status_gva;
  wire csr_io_status_hie;
  wire [31:0] csr_io_status_isa;
  wire csr_io_status_mbe;
  wire csr_io_status_mie;
  wire csr_io_status_mpie;
  wire [1:0] csr_io_status_mpp;
  wire csr_io_status_mprv;
  wire csr_io_status_mpv;
  wire csr_io_status_mxr;
  wire [1:0] csr_io_status_prv;
  wire csr_io_status_sbe;
  wire csr_io_status_sd;
  wire csr_io_status_sd_rv32;
  wire csr_io_status_sie;
  wire csr_io_status_spie;
  wire csr_io_status_spp;
  wire csr_io_status_sum;
  wire [1:0] csr_io_status_sxl;
  wire csr_io_status_tsr;
  wire csr_io_status_tvm;
  wire csr_io_status_tw;
  wire csr_io_status_ube;
  wire csr_io_status_uie;
  wire csr_io_status_upie;
  wire [1:0] csr_io_status_uxl;
  wire csr_io_status_v;
  wire [1:0] csr_io_status_vs;
  wire csr_io_status_wfi;
  wire [1:0] csr_io_status_xs;
  wire [7:0] csr_io_status_zero1;
  wire [22:0] csr_io_status_zero2;
  wire [31:0] csr_io_time;
  wire csr_io_trace_0_exception;
  wire [31:0] csr_io_trace_0_iaddr;
  wire [31:0] csr_io_trace_0_insn;
  wire csr_io_trace_0_valid;
  wire [31:0] csr_io_tval;
  wire csr_io_ungated_clock;
  wire csr_reset;
  wire div_clock;
  wire div_io_kill;
  wire div_io_kill_REG;
  wire [3:0] div_io_req_bits_fn;
  wire [31:0] div_io_req_bits_in1;
  wire [31:0] div_io_req_bits_in2;
  wire [4:0] div_io_req_bits_tag;
  wire div_io_req_ready;
  wire div_io_req_valid;
  wire [31:0] div_io_resp_bits_data;
  wire [4:0] div_io_resp_bits_tag;
  wire div_io_resp_ready;
  wire div_io_resp_valid;
  wire div_reset;
  wire [4:0] dmem_resp_waddr;
  wire [3:0] ex_ctrl_alu_fn;
  wire ex_ctrl_branch;
  wire [2:0] ex_ctrl_csr;
  wire ex_ctrl_div;
  wire ex_ctrl_fence_i;
  wire ex_ctrl_fp;
  wire ex_ctrl_jal;
  wire ex_ctrl_jalr;
  wire ex_ctrl_mem;
  wire [4:0] ex_ctrl_mem_cmd;
  wire ex_ctrl_mul;
  wire ex_ctrl_rfs1;
  wire ex_ctrl_rfs2;
  wire ex_ctrl_rocc;
  wire ex_ctrl_rxs2;
  wire [1:0] ex_ctrl_sel_alu1;
  wire [1:0] ex_ctrl_sel_alu2;
  wire [2:0] ex_ctrl_sel_imm;
  wire ex_ctrl_wfd;
  wire ex_ctrl_wxd;
  wire [5:0] ex_dcache_tag;
  wire [31:0] ex_reg_cause;
  wire ex_reg_flush_pipe;
  wire [31:0] ex_reg_inst;
  wire ex_reg_load_use;
  wire [1:0] ex_reg_mem_size;
  wire [31:0] ex_reg_pc;
  wire [31:0] ex_reg_raw_inst;
  wire ex_reg_replay;
  wire ex_reg_rs_bypass_0;
  wire ex_reg_rs_bypass_1;
  wire [1:0] ex_reg_rs_lsb_0;
  wire [1:0] ex_reg_rs_lsb_1;
  wire [29:0] ex_reg_rs_msb_0;
  wire [29:0] ex_reg_rs_msb_1;
  wire ex_reg_rvc;
  wire ex_reg_valid;
  wire ex_reg_xcpt;
  wire ex_reg_xcpt_interrupt;
  wire [31:0] ex_rs_1;
  wire [4:0] ex_waddr;
  wire ibuf_clock;
  wire [31:0] ibuf_io_imem_bits_data;
  wire [31:0] ibuf_io_imem_bits_pc;
  wire ibuf_io_imem_bits_replay;
  wire ibuf_io_imem_bits_xcpt_ae_inst;
  wire ibuf_io_imem_ready;
  wire ibuf_io_imem_valid;
  wire [31:0] ibuf_io_inst_0_bits_inst_bits;
  wire [4:0] ibuf_io_inst_0_bits_inst_rd;
  wire [4:0] ibuf_io_inst_0_bits_inst_rs1;
  wire [4:0] ibuf_io_inst_0_bits_inst_rs2;
  wire [31:0] ibuf_io_inst_0_bits_raw;
  wire ibuf_io_inst_0_bits_replay;
  wire ibuf_io_inst_0_bits_rvc;
  wire ibuf_io_inst_0_bits_xcpt0_ae_inst;
  wire ibuf_io_inst_0_bits_xcpt1_ae_inst;
  wire ibuf_io_inst_0_bits_xcpt1_gf_inst;
  wire ibuf_io_inst_0_bits_xcpt1_pf_inst;
  wire ibuf_io_inst_0_ready;
  wire ibuf_io_inst_0_valid;
  wire ibuf_io_kill;
  wire [31:0] ibuf_io_pc;
  wire ibuf_reset;
  wire id_amo_aq;
  wire id_amo_rl;
  wire id_ctrl_decoder_1;
  wire [4:0] id_ctrl_decoder_15;
  wire id_ctrl_decoder_16;
  wire id_ctrl_decoder_17;
  wire id_ctrl_decoder_19;
  wire id_ctrl_decoder_2;
  wire id_ctrl_decoder_20;
  wire id_ctrl_decoder_27;
  wire id_ctrl_decoder_8;
  wire id_ctrl_decoder_decoded_andMatrixInput_0;
  wire id_ctrl_decoder_decoded_andMatrixInput_1;
  wire id_ctrl_decoder_decoded_andMatrixInput_10;
  wire id_ctrl_decoder_decoded_andMatrixInput_10_20;
  wire id_ctrl_decoder_decoded_andMatrixInput_11;
  wire id_ctrl_decoder_decoded_andMatrixInput_11_1;
  wire id_ctrl_decoder_decoded_andMatrixInput_12;
  wire id_ctrl_decoder_decoded_andMatrixInput_12_2;
  wire id_ctrl_decoder_decoded_andMatrixInput_12_25;
  wire id_ctrl_decoder_decoded_andMatrixInput_12_33;
  wire id_ctrl_decoder_decoded_andMatrixInput_13;
  wire id_ctrl_decoder_decoded_andMatrixInput_13_1;
  wire id_ctrl_decoder_decoded_andMatrixInput_13_19;
  wire id_ctrl_decoder_decoded_andMatrixInput_14;
  wire id_ctrl_decoder_decoded_andMatrixInput_14_1;
  wire id_ctrl_decoder_decoded_andMatrixInput_15;
  wire id_ctrl_decoder_decoded_andMatrixInput_15_1;
  wire id_ctrl_decoder_decoded_andMatrixInput_15_14;
  wire id_ctrl_decoder_decoded_andMatrixInput_16;
  wire id_ctrl_decoder_decoded_andMatrixInput_17;
  wire id_ctrl_decoder_decoded_andMatrixInput_17_3;
  wire id_ctrl_decoder_decoded_andMatrixInput_17_5;
  wire id_ctrl_decoder_decoded_andMatrixInput_18;
  wire id_ctrl_decoder_decoded_andMatrixInput_19;
  wire id_ctrl_decoder_decoded_andMatrixInput_19_3;
  wire id_ctrl_decoder_decoded_andMatrixInput_2;
  wire id_ctrl_decoder_decoded_andMatrixInput_20;
  wire id_ctrl_decoder_decoded_andMatrixInput_20_6;
  wire id_ctrl_decoder_decoded_andMatrixInput_2_5;
  wire id_ctrl_decoder_decoded_andMatrixInput_3;
  wire id_ctrl_decoder_decoded_andMatrixInput_3_5;
  wire id_ctrl_decoder_decoded_andMatrixInput_4;
  wire id_ctrl_decoder_decoded_andMatrixInput_4_18;
  wire id_ctrl_decoder_decoded_andMatrixInput_4_6;
  wire id_ctrl_decoder_decoded_andMatrixInput_5;
  wire id_ctrl_decoder_decoded_andMatrixInput_5_18;
  wire id_ctrl_decoder_decoded_andMatrixInput_5_8;
  wire id_ctrl_decoder_decoded_andMatrixInput_6;
  wire id_ctrl_decoder_decoded_andMatrixInput_6_1;
  wire id_ctrl_decoder_decoded_andMatrixInput_6_12;
  wire id_ctrl_decoder_decoded_andMatrixInput_6_17;
  wire id_ctrl_decoder_decoded_andMatrixInput_7;
  wire id_ctrl_decoder_decoded_andMatrixInput_7_15;
  wire id_ctrl_decoder_decoded_andMatrixInput_7_17;
  wire id_ctrl_decoder_decoded_andMatrixInput_7_2;
  wire id_ctrl_decoder_decoded_andMatrixInput_7_24;
  wire id_ctrl_decoder_decoded_andMatrixInput_7_50;
  wire id_ctrl_decoder_decoded_andMatrixInput_7_54;
  wire id_ctrl_decoder_decoded_andMatrixInput_8_22;
  wire id_ctrl_decoder_decoded_andMatrixInput_8_8;
  wire [9:0] id_ctrl_decoder_decoded_hi_58;
  wire [6:0] id_ctrl_decoder_decoded_hi_lo_17;
  wire [7:0] id_ctrl_decoder_decoded_hi_lo_18;
  wire [6:0] id_ctrl_decoder_decoded_hi_lo_62;
  wire [31:0] id_ctrl_decoder_decoded_invInputs;
  wire [40:0] id_ctrl_decoder_decoded_invMatrixOutputs;
  wire [4:0] id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_lo;
  wire [9:0] id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi;
  wire [9:0] id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo;
  wire [7:0] id_ctrl_decoder_decoded_lo_11;
  wire [5:0] id_ctrl_decoder_decoded_lo_12;
  wire [13:0] id_ctrl_decoder_decoded_lo_18;
  wire [14:0] id_ctrl_decoder_decoded_lo_19;
  wire [7:0] id_ctrl_decoder_decoded_lo_22;
  wire [5:0] id_ctrl_decoder_decoded_lo_29;
  wire [7:0] id_ctrl_decoder_decoded_lo_31;
  wire [6:0] id_ctrl_decoder_decoded_lo_35;
  wire [6:0] id_ctrl_decoder_decoded_lo_37;
  wire [6:0] id_ctrl_decoder_decoded_lo_39;
  wire [7:0] id_ctrl_decoder_decoded_lo_40;
  wire [7:0] id_ctrl_decoder_decoded_lo_41;
  wire [6:0] id_ctrl_decoder_decoded_lo_53;
  wire [6:0] id_ctrl_decoder_decoded_lo_56;
  wire [7:0] id_ctrl_decoder_decoded_lo_57;
  wire [9:0] id_ctrl_decoder_decoded_lo_58;
  wire [13:0] id_ctrl_decoder_decoded_lo_59;
  wire [14:0] id_ctrl_decoder_decoded_lo_60;
  wire [6:0] id_ctrl_decoder_decoded_lo_61;
  wire [5:0] id_ctrl_decoder_decoded_lo_62;
  wire [13:0] id_ctrl_decoder_decoded_lo_63;
  wire [15:0] id_ctrl_decoder_decoded_lo_64;
  wire [7:0] id_ctrl_decoder_decoded_lo_65;
  wire [5:0] id_ctrl_decoder_decoded_lo_66;
  wire [7:0] id_ctrl_decoder_decoded_lo_67;
  wire [13:0] id_ctrl_decoder_decoded_lo_68;
  wire [15:0] id_ctrl_decoder_decoded_lo_69;
  wire [5:0] id_ctrl_decoder_decoded_lo_70;
  wire [6:0] id_ctrl_decoder_decoded_lo_lo_15;
  wire [6:0] id_ctrl_decoder_decoded_lo_lo_56;
  wire [6:0] id_ctrl_decoder_decoded_lo_lo_60;
  wire [7:0] id_ctrl_decoder_decoded_lo_lo_61;
  wire [6:0] id_ctrl_decoder_decoded_lo_lo_65;
  wire [7:0] id_ctrl_decoder_decoded_lo_lo_66;
  wire [40:0] id_ctrl_decoder_decoded_orMatrixOutputs;
  wire [4:0] id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_6;
  wire [19:0] id_ctrl_decoder_decoded_orMatrixOutputs_lo_17;
  wire [9:0] id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_10;
  wire [31:0] id_ctrl_decoder_decoded_plaInput;
  wire [3:0] id_fence_succ;
  wire [4:0] id_raddr1;
  wire [4:0] id_raddr2;
  wire id_reg_fence;
  wire id_reg_pause;
  wire [4:0] id_waddr;
  wire imem_might_request_reg;
  wire [31:0] inst;
  input io_dmem_ordered;
  wire io_dmem_ordered;
  input io_dmem_perf_grant;
  wire io_dmem_perf_grant;
  input io_dmem_replay_next;
  wire io_dmem_replay_next;
  output [31:0] io_dmem_req_bits_addr;
  wire [31:0] io_dmem_req_bits_addr;
  output [4:0] io_dmem_req_bits_cmd;
  wire [4:0] io_dmem_req_bits_cmd;
  output io_dmem_req_bits_dv;
  wire io_dmem_req_bits_dv;
  output io_dmem_req_bits_signed;
  wire io_dmem_req_bits_signed;
  output [1:0] io_dmem_req_bits_size;
  wire [1:0] io_dmem_req_bits_size;
  output [6:0] io_dmem_req_bits_tag;
  wire [6:0] io_dmem_req_bits_tag;
  input io_dmem_req_ready;
  wire io_dmem_req_ready;
  output io_dmem_req_valid;
  wire io_dmem_req_valid;
  input [31:0] io_dmem_resp_bits_data;
  wire [31:0] io_dmem_resp_bits_data;
  input [31:0] io_dmem_resp_bits_data_word_bypass;
  wire [31:0] io_dmem_resp_bits_data_word_bypass;
  input io_dmem_resp_bits_has_data;
  wire io_dmem_resp_bits_has_data;
  input io_dmem_resp_bits_replay;
  wire io_dmem_resp_bits_replay;
  input [6:0] io_dmem_resp_bits_tag;
  wire [6:0] io_dmem_resp_bits_tag;
  input io_dmem_resp_valid;
  wire io_dmem_resp_valid;
  output [31:0] io_dmem_s1_data_data;
  wire [31:0] io_dmem_s1_data_data;
  output io_dmem_s1_kill;
  wire io_dmem_s1_kill;
  input io_dmem_s2_nack;
  wire io_dmem_s2_nack;
  input io_dmem_s2_xcpt_ae_ld;
  wire io_dmem_s2_xcpt_ae_ld;
  input io_dmem_s2_xcpt_ae_st;
  wire io_dmem_s2_xcpt_ae_st;
  input io_dmem_s2_xcpt_ma_ld;
  wire io_dmem_s2_xcpt_ma_ld;
  input io_dmem_s2_xcpt_ma_st;
  wire io_dmem_s2_xcpt_ma_st;
  input io_dmem_s2_xcpt_pf_ld;
  wire io_dmem_s2_xcpt_pf_ld;
  input io_dmem_s2_xcpt_pf_st;
  wire io_dmem_s2_xcpt_pf_st;
  input io_hartid;
  wire io_hartid;
  output io_imem_bht_update_valid;
  wire io_imem_bht_update_valid;
  output io_imem_btb_update_valid;
  wire io_imem_btb_update_valid;
  output io_imem_flush_icache;
  wire io_imem_flush_icache;
  output io_imem_might_request;
  wire io_imem_might_request;
  output [31:0] io_imem_req_bits_pc;
  wire [31:0] io_imem_req_bits_pc;
  output io_imem_req_bits_speculative;
  wire io_imem_req_bits_speculative;
  output io_imem_req_valid;
  wire io_imem_req_valid;
  input [31:0] io_imem_resp_bits_data;
  wire [31:0] io_imem_resp_bits_data;
  input [31:0] io_imem_resp_bits_pc;
  wire [31:0] io_imem_resp_bits_pc;
  input io_imem_resp_bits_replay;
  wire io_imem_resp_bits_replay;
  input io_imem_resp_bits_xcpt_ae_inst;
  wire io_imem_resp_bits_xcpt_ae_inst;
  output io_imem_resp_ready;
  wire io_imem_resp_ready;
  input io_imem_resp_valid;
  wire io_imem_resp_valid;
  input io_interrupts_debug;
  wire io_interrupts_debug;
  input io_interrupts_meip;
  wire io_interrupts_meip;
  input io_interrupts_msip;
  wire io_interrupts_msip;
  input io_interrupts_mtip;
  wire io_interrupts_mtip;
  output [31:0] io_ptw_customCSRs_csrs_0_value;
  wire [31:0] io_ptw_customCSRs_csrs_0_value;
  output [29:0] io_ptw_pmp_0_addr;
  wire [29:0] io_ptw_pmp_0_addr;
  output [1:0] io_ptw_pmp_0_cfg_a;
  wire [1:0] io_ptw_pmp_0_cfg_a;
  output io_ptw_pmp_0_cfg_l;
  wire io_ptw_pmp_0_cfg_l;
  output io_ptw_pmp_0_cfg_r;
  wire io_ptw_pmp_0_cfg_r;
  output io_ptw_pmp_0_cfg_w;
  wire io_ptw_pmp_0_cfg_w;
  output io_ptw_pmp_0_cfg_x;
  wire io_ptw_pmp_0_cfg_x;
  output [31:0] io_ptw_pmp_0_mask;
  wire [31:0] io_ptw_pmp_0_mask;
  output [29:0] io_ptw_pmp_1_addr;
  wire [29:0] io_ptw_pmp_1_addr;
  output [1:0] io_ptw_pmp_1_cfg_a;
  wire [1:0] io_ptw_pmp_1_cfg_a;
  output io_ptw_pmp_1_cfg_l;
  wire io_ptw_pmp_1_cfg_l;
  output io_ptw_pmp_1_cfg_r;
  wire io_ptw_pmp_1_cfg_r;
  output io_ptw_pmp_1_cfg_w;
  wire io_ptw_pmp_1_cfg_w;
  output io_ptw_pmp_1_cfg_x;
  wire io_ptw_pmp_1_cfg_x;
  output [31:0] io_ptw_pmp_1_mask;
  wire [31:0] io_ptw_pmp_1_mask;
  output [29:0] io_ptw_pmp_2_addr;
  wire [29:0] io_ptw_pmp_2_addr;
  output [1:0] io_ptw_pmp_2_cfg_a;
  wire [1:0] io_ptw_pmp_2_cfg_a;
  output io_ptw_pmp_2_cfg_l;
  wire io_ptw_pmp_2_cfg_l;
  output io_ptw_pmp_2_cfg_r;
  wire io_ptw_pmp_2_cfg_r;
  output io_ptw_pmp_2_cfg_w;
  wire io_ptw_pmp_2_cfg_w;
  output io_ptw_pmp_2_cfg_x;
  wire io_ptw_pmp_2_cfg_x;
  output [31:0] io_ptw_pmp_2_mask;
  wire [31:0] io_ptw_pmp_2_mask;
  output [29:0] io_ptw_pmp_3_addr;
  wire [29:0] io_ptw_pmp_3_addr;
  output [1:0] io_ptw_pmp_3_cfg_a;
  wire [1:0] io_ptw_pmp_3_cfg_a;
  output io_ptw_pmp_3_cfg_l;
  wire io_ptw_pmp_3_cfg_l;
  output io_ptw_pmp_3_cfg_r;
  wire io_ptw_pmp_3_cfg_r;
  output io_ptw_pmp_3_cfg_w;
  wire io_ptw_pmp_3_cfg_w;
  output io_ptw_pmp_3_cfg_x;
  wire io_ptw_pmp_3_cfg_x;
  output [31:0] io_ptw_pmp_3_mask;
  wire [31:0] io_ptw_pmp_3_mask;
  output [29:0] io_ptw_pmp_4_addr;
  wire [29:0] io_ptw_pmp_4_addr;
  output [1:0] io_ptw_pmp_4_cfg_a;
  wire [1:0] io_ptw_pmp_4_cfg_a;
  output io_ptw_pmp_4_cfg_l;
  wire io_ptw_pmp_4_cfg_l;
  output io_ptw_pmp_4_cfg_r;
  wire io_ptw_pmp_4_cfg_r;
  output io_ptw_pmp_4_cfg_w;
  wire io_ptw_pmp_4_cfg_w;
  output io_ptw_pmp_4_cfg_x;
  wire io_ptw_pmp_4_cfg_x;
  output [31:0] io_ptw_pmp_4_mask;
  wire [31:0] io_ptw_pmp_4_mask;
  output [29:0] io_ptw_pmp_5_addr;
  wire [29:0] io_ptw_pmp_5_addr;
  output [1:0] io_ptw_pmp_5_cfg_a;
  wire [1:0] io_ptw_pmp_5_cfg_a;
  output io_ptw_pmp_5_cfg_l;
  wire io_ptw_pmp_5_cfg_l;
  output io_ptw_pmp_5_cfg_r;
  wire io_ptw_pmp_5_cfg_r;
  output io_ptw_pmp_5_cfg_w;
  wire io_ptw_pmp_5_cfg_w;
  output io_ptw_pmp_5_cfg_x;
  wire io_ptw_pmp_5_cfg_x;
  output [31:0] io_ptw_pmp_5_mask;
  wire [31:0] io_ptw_pmp_5_mask;
  output [29:0] io_ptw_pmp_6_addr;
  wire [29:0] io_ptw_pmp_6_addr;
  output [1:0] io_ptw_pmp_6_cfg_a;
  wire [1:0] io_ptw_pmp_6_cfg_a;
  output io_ptw_pmp_6_cfg_l;
  wire io_ptw_pmp_6_cfg_l;
  output io_ptw_pmp_6_cfg_r;
  wire io_ptw_pmp_6_cfg_r;
  output io_ptw_pmp_6_cfg_w;
  wire io_ptw_pmp_6_cfg_w;
  output io_ptw_pmp_6_cfg_x;
  wire io_ptw_pmp_6_cfg_x;
  output [31:0] io_ptw_pmp_6_mask;
  wire [31:0] io_ptw_pmp_6_mask;
  output [29:0] io_ptw_pmp_7_addr;
  wire [29:0] io_ptw_pmp_7_addr;
  output [1:0] io_ptw_pmp_7_cfg_a;
  wire [1:0] io_ptw_pmp_7_cfg_a;
  output io_ptw_pmp_7_cfg_l;
  wire io_ptw_pmp_7_cfg_l;
  output io_ptw_pmp_7_cfg_r;
  wire io_ptw_pmp_7_cfg_r;
  output io_ptw_pmp_7_cfg_w;
  wire io_ptw_pmp_7_cfg_w;
  output io_ptw_pmp_7_cfg_x;
  wire io_ptw_pmp_7_cfg_x;
  output [31:0] io_ptw_pmp_7_mask;
  wire [31:0] io_ptw_pmp_7_mask;
  output io_ptw_status_debug;
  wire io_ptw_status_debug;
  output io_rocc_cmd_valid;
  wire io_rocc_cmd_valid;
  output io_wfi;
  wire io_wfi;
  wire [31:0] ll_wdata;
  wire mem_br_taken;
  wire [31:0] mem_br_target;
  wire [5:0] mem_br_target_b10_5;
  wire [3:0] mem_br_target_b4_1;
  wire mem_br_target_hi_hi_hi;
  wire [10:0] mem_br_target_hi_hi_lo;
  wire [7:0] mem_br_target_hi_lo_hi;
  wire [7:0] mem_br_target_hi_lo_hi_1;
  wire mem_br_target_hi_lo_lo;
  wire mem_br_target_hi_lo_lo_1;
  wire mem_br_target_sign;
  wire mem_ctrl_branch;
  wire [2:0] mem_ctrl_csr;
  wire mem_ctrl_div;
  wire mem_ctrl_fence_i;
  wire mem_ctrl_fp;
  wire mem_ctrl_jal;
  wire mem_ctrl_jalr;
  wire mem_ctrl_mem;
  wire mem_ctrl_mul;
  wire mem_ctrl_rocc;
  wire mem_ctrl_wxd;
  wire [3:0] mem_ldst_cause;
  wire [31:0] mem_npc;
  wire [31:0] mem_reg_cause;
  wire mem_reg_flush_pipe;
  wire mem_reg_hls_or_dv;
  wire [31:0] mem_reg_inst;
  wire mem_reg_load;
  wire [31:0] mem_reg_pc;
  wire [31:0] mem_reg_raw_inst;
  wire mem_reg_replay;
  wire [31:0] mem_reg_rs2;
  wire mem_reg_rvc;
  wire mem_reg_slow_bypass;
  wire mem_reg_store;
  wire mem_reg_valid;
  wire [31:0] mem_reg_wdata;
  wire mem_reg_xcpt;
  wire mem_reg_xcpt_interrupt;
  wire [4:0] mem_waddr;
  wire [31:0] r;
  wire replay_wb_rocc;
  input reset;
  wire reset;
  wire [31:0] \rf[0] ;
  wire [31:0] \rf[10] ;
  wire [31:0] \rf[11] ;
  wire [31:0] \rf[12] ;
  wire [31:0] \rf[13] ;
  wire [31:0] \rf[14] ;
  wire [31:0] \rf[15] ;
  wire [31:0] \rf[16] ;
  wire [31:0] \rf[17] ;
  wire [31:0] \rf[18] ;
  wire [31:0] \rf[19] ;
  wire [31:0] \rf[1] ;
  wire [31:0] \rf[20] ;
  wire [31:0] \rf[21] ;
  wire [31:0] \rf[22] ;
  wire [31:0] \rf[23] ;
  wire [31:0] \rf[24] ;
  wire [31:0] \rf[25] ;
  wire [31:0] \rf[26] ;
  wire [31:0] \rf[27] ;
  wire [31:0] \rf[28] ;
  wire [31:0] \rf[29] ;
  wire [31:0] \rf[2] ;
  wire [31:0] \rf[30] ;
  wire [31:0] \rf[3] ;
  wire [31:0] \rf[4] ;
  wire [31:0] \rf[5] ;
  wire [31:0] \rf[6] ;
  wire [31:0] \rf[7] ;
  wire [31:0] \rf[8] ;
  wire [31:0] \rf[9] ;
  wire rf_MPORT_mask;
  wire rf_id_rs_MPORT_1_en;
  wire rf_id_rs_MPORT_en;
  wire [1:0] size;
  wire take_pc_mem_wb;
  wire tval_dmem_addr;
  wire [2:0] wb_ctrl_csr;
  wire wb_ctrl_div;
  wire wb_ctrl_fence_i;
  wire wb_ctrl_mem;
  wire wb_ctrl_rocc;
  wire wb_ctrl_wxd;
  wire [31:0] wb_reg_cause;
  wire wb_reg_flush_pipe;
  wire wb_reg_hls_or_dv;
  wire [31:0] wb_reg_inst;
  wire [31:0] wb_reg_pc;
  wire [31:0] wb_reg_raw_inst;
  wire wb_reg_replay;
  wire wb_reg_valid;
  wire [31:0] wb_reg_wdata;
  wire wb_reg_xcpt;
  wire wb_valid;
  wire [4:0] wb_waddr;
  wire wb_xcpt;
  INV_X1 _15565_ (
    .A(id_reg_pause),
    .ZN(_07940_)
  );
  INV_X1 _15566_ (
    .A(csr_io_interrupt),
    .ZN(_07941_)
  );
  INV_X1 _15567_ (
    .A(_r[31]),
    .ZN(_07942_)
  );
  INV_X1 _15568_ (
    .A(_r[29]),
    .ZN(_07943_)
  );
  INV_X1 _15569_ (
    .A(_r[27]),
    .ZN(_07944_)
  );
  INV_X1 _15570_ (
    .A(_r[25]),
    .ZN(_07945_)
  );
  INV_X1 _15571_ (
    .A(_r[15]),
    .ZN(_07946_)
  );
  INV_X1 _15572_ (
    .A(_r[13]),
    .ZN(_07947_)
  );
  INV_X1 _15573_ (
    .A(_r[11]),
    .ZN(_07948_)
  );
  INV_X1 _15574_ (
    .A(_r[9]),
    .ZN(_07949_)
  );
  INV_X1 _15575_ (
    .A(_r[7]),
    .ZN(_07950_)
  );
  INV_X1 _15576_ (
    .A(_r[5]),
    .ZN(_07951_)
  );
  INV_X1 _15577_ (
    .A(_r[3]),
    .ZN(_07952_)
  );
  INV_X1 _15578_ (
    .A(_r[1]),
    .ZN(_07953_)
  );
  INV_X1 _15579_ (
    .A(reset),
    .ZN(_07954_)
  );
  INV_X1 _15580_ (
    .A(ex_reg_rs_lsb_0[0]),
    .ZN(_07955_)
  );
  INV_X1 _15581_ (
    .A(ex_reg_rs_lsb_0[1]),
    .ZN(_07956_)
  );
  INV_X1 _15582_ (
    .A(wb_reg_cause[4]),
    .ZN(_07957_)
  );
  INV_X1 _15583_ (
    .A(wb_reg_cause[5]),
    .ZN(_07958_)
  );
  INV_X1 _15584_ (
    .A(wb_reg_cause[6]),
    .ZN(_07959_)
  );
  INV_X1 _15585_ (
    .A(wb_reg_cause[7]),
    .ZN(_07960_)
  );
  INV_X1 _15586_ (
    .A(wb_reg_cause[8]),
    .ZN(_07961_)
  );
  INV_X1 _15587_ (
    .A(wb_reg_cause[9]),
    .ZN(_07962_)
  );
  INV_X1 _15588_ (
    .A(wb_reg_cause[10]),
    .ZN(_07963_)
  );
  INV_X1 _15589_ (
    .A(wb_reg_cause[11]),
    .ZN(_07964_)
  );
  INV_X1 _15590_ (
    .A(wb_reg_cause[12]),
    .ZN(_07965_)
  );
  INV_X1 _15591_ (
    .A(wb_reg_cause[13]),
    .ZN(_07966_)
  );
  INV_X1 _15592_ (
    .A(wb_reg_cause[14]),
    .ZN(_07967_)
  );
  INV_X1 _15593_ (
    .A(wb_reg_cause[15]),
    .ZN(_07968_)
  );
  INV_X1 _15594_ (
    .A(wb_reg_cause[16]),
    .ZN(_07969_)
  );
  INV_X1 _15595_ (
    .A(wb_reg_cause[17]),
    .ZN(_07970_)
  );
  INV_X1 _15596_ (
    .A(wb_reg_cause[18]),
    .ZN(_07971_)
  );
  INV_X1 _15597_ (
    .A(wb_reg_cause[19]),
    .ZN(_07972_)
  );
  INV_X1 _15598_ (
    .A(wb_reg_cause[20]),
    .ZN(_07973_)
  );
  INV_X1 _15599_ (
    .A(wb_reg_cause[21]),
    .ZN(_07974_)
  );
  INV_X1 _15600_ (
    .A(wb_reg_cause[22]),
    .ZN(_07975_)
  );
  INV_X1 _15601_ (
    .A(wb_reg_cause[23]),
    .ZN(_07976_)
  );
  INV_X1 _15602_ (
    .A(wb_reg_cause[24]),
    .ZN(_07977_)
  );
  INV_X1 _15603_ (
    .A(wb_reg_cause[25]),
    .ZN(_07978_)
  );
  INV_X1 _15604_ (
    .A(wb_reg_cause[26]),
    .ZN(_07979_)
  );
  INV_X1 _15605_ (
    .A(wb_reg_cause[27]),
    .ZN(_07980_)
  );
  INV_X1 _15606_ (
    .A(wb_reg_cause[28]),
    .ZN(_07981_)
  );
  INV_X1 _15607_ (
    .A(wb_reg_cause[29]),
    .ZN(_07982_)
  );
  INV_X1 _15608_ (
    .A(wb_reg_cause[30]),
    .ZN(_07983_)
  );
  INV_X1 _15609_ (
    .A(wb_reg_cause[31]),
    .ZN(_07984_)
  );
  INV_X1 _15610_ (
    .A(mem_reg_pc[1]),
    .ZN(_07985_)
  );
  INV_X1 _15611_ (
    .A(mem_reg_pc[2]),
    .ZN(_07986_)
  );
  INV_X1 _15612_ (
    .A(mem_reg_pc[3]),
    .ZN(_07987_)
  );
  INV_X1 _15613_ (
    .A(mem_reg_pc[4]),
    .ZN(_07988_)
  );
  INV_X1 _15614_ (
    .A(wb_reg_pc[5]),
    .ZN(_07989_)
  );
  INV_X1 _15615_ (
    .A(mem_reg_pc[5]),
    .ZN(_07990_)
  );
  INV_X1 _15616_ (
    .A(wb_reg_pc[6]),
    .ZN(_07991_)
  );
  INV_X1 _15617_ (
    .A(mem_reg_pc[6]),
    .ZN(_07992_)
  );
  INV_X1 _15618_ (
    .A(wb_reg_pc[7]),
    .ZN(_07993_)
  );
  INV_X1 _15619_ (
    .A(mem_reg_pc[7]),
    .ZN(_07994_)
  );
  INV_X1 _15620_ (
    .A(wb_reg_pc[8]),
    .ZN(_07995_)
  );
  INV_X1 _15621_ (
    .A(mem_reg_pc[8]),
    .ZN(_07996_)
  );
  INV_X1 _15622_ (
    .A(wb_reg_pc[9]),
    .ZN(_07997_)
  );
  INV_X1 _15623_ (
    .A(mem_reg_pc[9]),
    .ZN(_07998_)
  );
  INV_X1 _15624_ (
    .A(wb_reg_pc[10]),
    .ZN(_07999_)
  );
  INV_X1 _15625_ (
    .A(mem_reg_pc[10]),
    .ZN(_08000_)
  );
  INV_X1 _15626_ (
    .A(wb_reg_pc[11]),
    .ZN(_08001_)
  );
  INV_X1 _15627_ (
    .A(mem_reg_pc[11]),
    .ZN(_08002_)
  );
  INV_X1 _15628_ (
    .A(wb_reg_pc[12]),
    .ZN(_08003_)
  );
  INV_X1 _15629_ (
    .A(mem_reg_pc[12]),
    .ZN(_08004_)
  );
  INV_X1 _15630_ (
    .A(wb_reg_pc[13]),
    .ZN(_08005_)
  );
  INV_X1 _15631_ (
    .A(mem_reg_pc[13]),
    .ZN(_08006_)
  );
  INV_X1 _15632_ (
    .A(wb_reg_pc[14]),
    .ZN(_08007_)
  );
  INV_X1 _15633_ (
    .A(mem_reg_pc[14]),
    .ZN(_08008_)
  );
  INV_X1 _15634_ (
    .A(wb_reg_pc[15]),
    .ZN(_08009_)
  );
  INV_X1 _15635_ (
    .A(mem_reg_pc[15]),
    .ZN(_08010_)
  );
  INV_X1 _15636_ (
    .A(wb_reg_pc[16]),
    .ZN(_08011_)
  );
  INV_X1 _15637_ (
    .A(mem_reg_pc[16]),
    .ZN(_08012_)
  );
  INV_X1 _15638_ (
    .A(wb_reg_pc[17]),
    .ZN(_08013_)
  );
  INV_X1 _15639_ (
    .A(mem_reg_pc[17]),
    .ZN(_08014_)
  );
  INV_X1 _15640_ (
    .A(wb_reg_pc[18]),
    .ZN(_08015_)
  );
  INV_X1 _15641_ (
    .A(mem_reg_pc[18]),
    .ZN(_08016_)
  );
  INV_X1 _15642_ (
    .A(wb_reg_pc[19]),
    .ZN(_08017_)
  );
  INV_X1 _15643_ (
    .A(mem_reg_pc[19]),
    .ZN(_08018_)
  );
  INV_X1 _15644_ (
    .A(wb_reg_pc[20]),
    .ZN(_08019_)
  );
  INV_X1 _15645_ (
    .A(mem_reg_pc[20]),
    .ZN(_08020_)
  );
  INV_X1 _15646_ (
    .A(wb_reg_pc[21]),
    .ZN(_08021_)
  );
  INV_X1 _15647_ (
    .A(mem_reg_pc[21]),
    .ZN(_08022_)
  );
  INV_X1 _15648_ (
    .A(wb_reg_pc[22]),
    .ZN(_08023_)
  );
  INV_X1 _15649_ (
    .A(mem_reg_pc[22]),
    .ZN(_08024_)
  );
  INV_X1 _15650_ (
    .A(wb_reg_pc[23]),
    .ZN(_08025_)
  );
  INV_X1 _15651_ (
    .A(mem_reg_pc[23]),
    .ZN(_08026_)
  );
  INV_X1 _15652_ (
    .A(wb_reg_pc[24]),
    .ZN(_08027_)
  );
  INV_X1 _15653_ (
    .A(mem_reg_pc[24]),
    .ZN(_08028_)
  );
  INV_X1 _15654_ (
    .A(wb_reg_pc[25]),
    .ZN(_08029_)
  );
  INV_X1 _15655_ (
    .A(mem_reg_pc[25]),
    .ZN(_08030_)
  );
  INV_X1 _15656_ (
    .A(wb_reg_pc[26]),
    .ZN(_08031_)
  );
  INV_X1 _15657_ (
    .A(mem_reg_pc[26]),
    .ZN(_08032_)
  );
  INV_X1 _15658_ (
    .A(wb_reg_pc[27]),
    .ZN(_08033_)
  );
  INV_X1 _15659_ (
    .A(mem_reg_pc[27]),
    .ZN(_08034_)
  );
  INV_X1 _15660_ (
    .A(wb_reg_pc[28]),
    .ZN(_08035_)
  );
  INV_X1 _15661_ (
    .A(mem_reg_pc[28]),
    .ZN(_08036_)
  );
  INV_X1 _15662_ (
    .A(wb_reg_pc[29]),
    .ZN(_08037_)
  );
  INV_X1 _15663_ (
    .A(mem_reg_pc[29]),
    .ZN(_08038_)
  );
  INV_X1 _15664_ (
    .A(wb_reg_pc[30]),
    .ZN(_08039_)
  );
  INV_X1 _15665_ (
    .A(mem_reg_pc[30]),
    .ZN(_08040_)
  );
  INV_X1 _15666_ (
    .A(wb_reg_pc[31]),
    .ZN(_08041_)
  );
  INV_X1 _15667_ (
    .A(mem_reg_pc[31]),
    .ZN(_08042_)
  );
  INV_X1 _15668_ (
    .A(mem_reg_rs2[8]),
    .ZN(_08043_)
  );
  INV_X1 _15669_ (
    .A(mem_reg_rs2[9]),
    .ZN(_08044_)
  );
  INV_X1 _15670_ (
    .A(mem_reg_rs2[10]),
    .ZN(_08045_)
  );
  INV_X1 _15671_ (
    .A(mem_reg_rs2[11]),
    .ZN(_08046_)
  );
  INV_X1 _15672_ (
    .A(mem_reg_rs2[12]),
    .ZN(_08047_)
  );
  INV_X1 _15673_ (
    .A(mem_reg_rs2[13]),
    .ZN(_08048_)
  );
  INV_X1 _15674_ (
    .A(mem_reg_rs2[24]),
    .ZN(_08049_)
  );
  INV_X1 _15675_ (
    .A(mem_reg_rs2[25]),
    .ZN(_08050_)
  );
  INV_X1 _15676_ (
    .A(mem_reg_rs2[26]),
    .ZN(_08051_)
  );
  INV_X1 _15677_ (
    .A(mem_reg_rs2[27]),
    .ZN(_08052_)
  );
  INV_X1 _15678_ (
    .A(mem_reg_rs2[28]),
    .ZN(_08053_)
  );
  INV_X1 _15679_ (
    .A(mem_reg_rs2[29]),
    .ZN(_08054_)
  );
  INV_X1 _15680_ (
    .A(mem_reg_rs2[30]),
    .ZN(_08055_)
  );
  INV_X1 _15681_ (
    .A(mem_reg_rs2[31]),
    .ZN(_08056_)
  );
  INV_X1 _15682_ (
    .A(mem_reg_wdata[5]),
    .ZN(_08057_)
  );
  INV_X1 _15683_ (
    .A(mem_reg_wdata[6]),
    .ZN(_08058_)
  );
  INV_X1 _15684_ (
    .A(mem_reg_wdata[7]),
    .ZN(_08059_)
  );
  INV_X1 _15685_ (
    .A(mem_reg_wdata[8]),
    .ZN(_08060_)
  );
  INV_X1 _15686_ (
    .A(mem_reg_wdata[9]),
    .ZN(_08061_)
  );
  INV_X1 _15687_ (
    .A(mem_reg_wdata[10]),
    .ZN(_08062_)
  );
  INV_X1 _15688_ (
    .A(mem_reg_wdata[11]),
    .ZN(_08063_)
  );
  INV_X1 _15689_ (
    .A(mem_reg_wdata[12]),
    .ZN(_08064_)
  );
  INV_X1 _15690_ (
    .A(mem_reg_wdata[13]),
    .ZN(_08065_)
  );
  INV_X1 _15691_ (
    .A(mem_reg_wdata[14]),
    .ZN(_08066_)
  );
  INV_X1 _15692_ (
    .A(mem_reg_wdata[15]),
    .ZN(_08067_)
  );
  INV_X1 _15693_ (
    .A(mem_reg_wdata[16]),
    .ZN(_08068_)
  );
  INV_X1 _15694_ (
    .A(mem_reg_wdata[17]),
    .ZN(_08069_)
  );
  INV_X1 _15695_ (
    .A(mem_reg_wdata[18]),
    .ZN(_08070_)
  );
  INV_X1 _15696_ (
    .A(mem_reg_wdata[19]),
    .ZN(_08071_)
  );
  INV_X1 _15697_ (
    .A(mem_reg_wdata[20]),
    .ZN(_08072_)
  );
  INV_X1 _15698_ (
    .A(mem_reg_wdata[21]),
    .ZN(_08073_)
  );
  INV_X1 _15699_ (
    .A(mem_reg_wdata[22]),
    .ZN(_08074_)
  );
  INV_X1 _15700_ (
    .A(mem_reg_wdata[23]),
    .ZN(_08075_)
  );
  INV_X1 _15701_ (
    .A(mem_reg_wdata[24]),
    .ZN(_08076_)
  );
  INV_X1 _15702_ (
    .A(mem_reg_wdata[25]),
    .ZN(_08077_)
  );
  INV_X1 _15703_ (
    .A(mem_reg_wdata[26]),
    .ZN(_08078_)
  );
  INV_X1 _15704_ (
    .A(mem_reg_wdata[27]),
    .ZN(_08079_)
  );
  INV_X1 _15705_ (
    .A(mem_reg_wdata[28]),
    .ZN(_08080_)
  );
  INV_X1 _15706_ (
    .A(mem_reg_wdata[29]),
    .ZN(_08081_)
  );
  INV_X1 _15707_ (
    .A(mem_reg_wdata[30]),
    .ZN(_08082_)
  );
  INV_X1 _15708_ (
    .A(mem_reg_wdata[31]),
    .ZN(_08083_)
  );
  INV_X1 _15709_ (
    .A(mem_reg_inst[7]),
    .ZN(_08084_)
  );
  INV_X1 _15710_ (
    .A(ex_reg_inst[7]),
    .ZN(_08085_)
  );
  INV_X1 _15711_ (
    .A(mem_reg_inst[8]),
    .ZN(_08086_)
  );
  INV_X1 _15712_ (
    .A(ex_reg_inst[8]),
    .ZN(_08087_)
  );
  INV_X1 _15713_ (
    .A(mem_reg_inst[9]),
    .ZN(_08088_)
  );
  INV_X1 _15714_ (
    .A(ex_reg_inst[9]),
    .ZN(_08089_)
  );
  INV_X1 _15715_ (
    .A(mem_reg_inst[10]),
    .ZN(_08090_)
  );
  INV_X1 _15716_ (
    .A(ex_reg_inst[10]),
    .ZN(_08091_)
  );
  INV_X1 _15717_ (
    .A(mem_reg_inst[11]),
    .ZN(_08092_)
  );
  INV_X1 _15718_ (
    .A(ex_reg_inst[11]),
    .ZN(_08093_)
  );
  INV_X1 _15719_ (
    .A(ex_reg_inst[20]),
    .ZN(_08094_)
  );
  INV_X1 _15720_ (
    .A(ex_reg_pc[0]),
    .ZN(_08095_)
  );
  INV_X1 _15721_ (
    .A(ex_reg_pc[1]),
    .ZN(_08096_)
  );
  INV_X1 _15722_ (
    .A(ex_reg_pc[2]),
    .ZN(_08097_)
  );
  INV_X1 _15723_ (
    .A(ex_reg_pc[3]),
    .ZN(_08098_)
  );
  INV_X1 _15724_ (
    .A(ex_reg_pc[4]),
    .ZN(_08099_)
  );
  INV_X1 _15725_ (
    .A(ex_reg_pc[5]),
    .ZN(_08100_)
  );
  INV_X1 _15726_ (
    .A(ex_reg_pc[6]),
    .ZN(_08101_)
  );
  INV_X1 _15727_ (
    .A(ex_reg_pc[7]),
    .ZN(_08102_)
  );
  INV_X1 _15728_ (
    .A(ex_reg_pc[8]),
    .ZN(_08103_)
  );
  INV_X1 _15729_ (
    .A(ex_reg_pc[9]),
    .ZN(_08104_)
  );
  INV_X1 _15730_ (
    .A(ex_reg_pc[10]),
    .ZN(_08105_)
  );
  INV_X1 _15731_ (
    .A(ex_reg_pc[11]),
    .ZN(_08106_)
  );
  INV_X1 _15732_ (
    .A(ex_reg_pc[12]),
    .ZN(_08107_)
  );
  INV_X1 _15733_ (
    .A(ex_reg_pc[13]),
    .ZN(_08108_)
  );
  INV_X1 _15734_ (
    .A(ex_reg_pc[14]),
    .ZN(_08109_)
  );
  INV_X1 _15735_ (
    .A(ex_reg_pc[15]),
    .ZN(_08110_)
  );
  INV_X1 _15736_ (
    .A(ex_reg_pc[16]),
    .ZN(_08111_)
  );
  INV_X1 _15737_ (
    .A(ex_reg_pc[17]),
    .ZN(_08112_)
  );
  INV_X1 _15738_ (
    .A(ex_reg_pc[18]),
    .ZN(_08113_)
  );
  INV_X1 _15739_ (
    .A(ex_reg_pc[19]),
    .ZN(_08114_)
  );
  INV_X1 _15740_ (
    .A(ex_reg_pc[20]),
    .ZN(_08115_)
  );
  INV_X1 _15741_ (
    .A(ex_reg_pc[21]),
    .ZN(_08116_)
  );
  INV_X1 _15742_ (
    .A(ex_reg_pc[22]),
    .ZN(_08117_)
  );
  INV_X1 _15743_ (
    .A(ex_reg_pc[23]),
    .ZN(_08118_)
  );
  INV_X1 _15744_ (
    .A(ex_reg_pc[24]),
    .ZN(_08119_)
  );
  INV_X1 _15745_ (
    .A(ex_reg_pc[25]),
    .ZN(_08120_)
  );
  INV_X1 _15746_ (
    .A(ex_reg_pc[26]),
    .ZN(_08121_)
  );
  INV_X1 _15747_ (
    .A(ex_reg_pc[27]),
    .ZN(_08122_)
  );
  INV_X1 _15748_ (
    .A(ex_reg_pc[28]),
    .ZN(_08123_)
  );
  INV_X1 _15749_ (
    .A(ex_reg_pc[29]),
    .ZN(_08124_)
  );
  INV_X1 _15750_ (
    .A(ex_reg_pc[30]),
    .ZN(_08125_)
  );
  INV_X1 _15751_ (
    .A(ex_reg_pc[31]),
    .ZN(_08126_)
  );
  INV_X1 _15752_ (
    .A(ibuf_io_inst_0_bits_raw[0]),
    .ZN(_08127_)
  );
  INV_X1 _15753_ (
    .A(csr_io_decode_0_inst[7]),
    .ZN(_08128_)
  );
  INV_X1 _15754_ (
    .A(csr_io_decode_0_inst[8]),
    .ZN(_08129_)
  );
  INV_X1 _15755_ (
    .A(csr_io_decode_0_inst[9]),
    .ZN(_08130_)
  );
  INV_X1 _15756_ (
    .A(csr_io_decode_0_inst[10]),
    .ZN(_08131_)
  );
  INV_X1 _15757_ (
    .A(csr_io_decode_0_inst[11]),
    .ZN(_08132_)
  );
  INV_X1 _15758_ (
    .A(csr_io_decode_0_inst[12]),
    .ZN(_08133_)
  );
  INV_X1 _15759_ (
    .A(csr_io_decode_0_inst[13]),
    .ZN(_08134_)
  );
  INV_X1 _15760_ (
    .A(csr_io_decode_0_inst[14]),
    .ZN(_08135_)
  );
  INV_X1 _15761_ (
    .A(csr_io_decode_0_inst[15]),
    .ZN(_08136_)
  );
  INV_X1 _15762_ (
    .A(csr_io_decode_0_inst[16]),
    .ZN(_08137_)
  );
  INV_X1 _15763_ (
    .A(csr_io_decode_0_inst[17]),
    .ZN(_08138_)
  );
  INV_X1 _15764_ (
    .A(csr_io_decode_0_inst[18]),
    .ZN(_08139_)
  );
  INV_X1 _15765_ (
    .A(csr_io_decode_0_inst[19]),
    .ZN(_08140_)
  );
  INV_X1 _15766_ (
    .A(csr_io_decode_0_inst[20]),
    .ZN(_08141_)
  );
  INV_X1 _15767_ (
    .A(csr_io_decode_0_inst[21]),
    .ZN(_08142_)
  );
  INV_X1 _15768_ (
    .A(csr_io_decode_0_inst[22]),
    .ZN(_08143_)
  );
  INV_X1 _15769_ (
    .A(csr_io_decode_0_inst[23]),
    .ZN(_08144_)
  );
  INV_X1 _15770_ (
    .A(csr_io_decode_0_inst[24]),
    .ZN(_08145_)
  );
  INV_X1 _15771_ (
    .A(csr_io_decode_0_inst[25]),
    .ZN(_08146_)
  );
  INV_X1 _15772_ (
    .A(csr_io_decode_0_inst[26]),
    .ZN(_08147_)
  );
  INV_X1 _15773_ (
    .A(csr_io_decode_0_inst[27]),
    .ZN(_08148_)
  );
  INV_X1 _15774_ (
    .A(csr_io_decode_0_inst[28]),
    .ZN(_08149_)
  );
  INV_X1 _15775_ (
    .A(csr_io_decode_0_inst[29]),
    .ZN(_08150_)
  );
  INV_X1 _15776_ (
    .A(csr_io_decode_0_inst[30]),
    .ZN(_08151_)
  );
  INV_X1 _15777_ (
    .A(csr_io_decode_0_inst[31]),
    .ZN(_08152_)
  );
  INV_X1 _15778_ (
    .A(ex_reg_mem_size[0]),
    .ZN(_08153_)
  );
  INV_X1 _15779_ (
    .A(ex_reg_mem_size[1]),
    .ZN(_08154_)
  );
  INV_X1 _15780_ (
    .A(bpu_io_pc[0]),
    .ZN(_08155_)
  );
  INV_X1 _15781_ (
    .A(bpu_io_pc[1]),
    .ZN(_08156_)
  );
  INV_X1 _15782_ (
    .A(bpu_io_pc[2]),
    .ZN(_08157_)
  );
  INV_X1 _15783_ (
    .A(bpu_io_pc[3]),
    .ZN(_08158_)
  );
  INV_X1 _15784_ (
    .A(bpu_io_pc[4]),
    .ZN(_08159_)
  );
  INV_X1 _15785_ (
    .A(bpu_io_pc[5]),
    .ZN(_08160_)
  );
  INV_X1 _15786_ (
    .A(bpu_io_pc[6]),
    .ZN(_08161_)
  );
  INV_X1 _15787_ (
    .A(bpu_io_pc[7]),
    .ZN(_08162_)
  );
  INV_X1 _15788_ (
    .A(bpu_io_pc[8]),
    .ZN(_08163_)
  );
  INV_X1 _15789_ (
    .A(bpu_io_pc[9]),
    .ZN(_08164_)
  );
  INV_X1 _15790_ (
    .A(bpu_io_pc[10]),
    .ZN(_08165_)
  );
  INV_X1 _15791_ (
    .A(bpu_io_pc[11]),
    .ZN(_08166_)
  );
  INV_X1 _15792_ (
    .A(bpu_io_pc[12]),
    .ZN(_08167_)
  );
  INV_X1 _15793_ (
    .A(bpu_io_pc[13]),
    .ZN(_08168_)
  );
  INV_X1 _15794_ (
    .A(bpu_io_pc[14]),
    .ZN(_08169_)
  );
  INV_X1 _15795_ (
    .A(bpu_io_pc[15]),
    .ZN(_08170_)
  );
  INV_X1 _15796_ (
    .A(bpu_io_pc[16]),
    .ZN(_08171_)
  );
  INV_X1 _15797_ (
    .A(bpu_io_pc[17]),
    .ZN(_08172_)
  );
  INV_X1 _15798_ (
    .A(bpu_io_pc[18]),
    .ZN(_08173_)
  );
  INV_X1 _15799_ (
    .A(bpu_io_pc[19]),
    .ZN(_08174_)
  );
  INV_X1 _15800_ (
    .A(bpu_io_pc[20]),
    .ZN(_08175_)
  );
  INV_X1 _15801_ (
    .A(bpu_io_pc[21]),
    .ZN(_08176_)
  );
  INV_X1 _15802_ (
    .A(bpu_io_pc[22]),
    .ZN(_08177_)
  );
  INV_X1 _15803_ (
    .A(bpu_io_pc[23]),
    .ZN(_08178_)
  );
  INV_X1 _15804_ (
    .A(bpu_io_pc[24]),
    .ZN(_08179_)
  );
  INV_X1 _15805_ (
    .A(bpu_io_pc[25]),
    .ZN(_08180_)
  );
  INV_X1 _15806_ (
    .A(bpu_io_pc[26]),
    .ZN(_08181_)
  );
  INV_X1 _15807_ (
    .A(bpu_io_pc[27]),
    .ZN(_08182_)
  );
  INV_X1 _15808_ (
    .A(bpu_io_pc[28]),
    .ZN(_08183_)
  );
  INV_X1 _15809_ (
    .A(bpu_io_pc[29]),
    .ZN(_08184_)
  );
  INV_X1 _15810_ (
    .A(bpu_io_pc[30]),
    .ZN(_08185_)
  );
  INV_X1 _15811_ (
    .A(bpu_io_pc[31]),
    .ZN(_08186_)
  );
  INV_X1 _15812_ (
    .A(ex_reg_flush_pipe),
    .ZN(_08187_)
  );
  INV_X1 _15813_ (
    .A(wb_ctrl_csr[0]),
    .ZN(_08188_)
  );
  INV_X1 _15814_ (
    .A(mem_ctrl_csr[0]),
    .ZN(_08189_)
  );
  INV_X1 _15815_ (
    .A(wb_ctrl_csr[1]),
    .ZN(_08190_)
  );
  INV_X1 _15816_ (
    .A(mem_ctrl_csr[1]),
    .ZN(_08191_)
  );
  INV_X1 _15817_ (
    .A(wb_ctrl_csr[2]),
    .ZN(_08192_)
  );
  INV_X1 _15818_ (
    .A(mem_ctrl_csr[2]),
    .ZN(_08193_)
  );
  INV_X1 _15819_ (
    .A(wb_ctrl_div),
    .ZN(_08194_)
  );
  INV_X1 _15820_ (
    .A(mem_ctrl_div),
    .ZN(_08195_)
  );
  INV_X1 _15821_ (
    .A(wb_reg_inst[7]),
    .ZN(_08196_)
  );
  INV_X1 _15822_ (
    .A(wb_reg_inst[8]),
    .ZN(_08197_)
  );
  INV_X1 _15823_ (
    .A(wb_reg_inst[9]),
    .ZN(_08198_)
  );
  INV_X1 _15824_ (
    .A(wb_reg_inst[10]),
    .ZN(_08199_)
  );
  INV_X1 _15825_ (
    .A(wb_reg_inst[11]),
    .ZN(_08200_)
  );
  INV_X1 _15826_ (
    .A(ex_ctrl_csr[0]),
    .ZN(_08201_)
  );
  INV_X1 _15827_ (
    .A(ex_ctrl_csr[1]),
    .ZN(_08202_)
  );
  INV_X1 _15828_ (
    .A(ex_ctrl_csr[2]),
    .ZN(_08203_)
  );
  INV_X1 _15829_ (
    .A(ex_ctrl_div),
    .ZN(_08204_)
  );
  INV_X1 _15830_ (
    .A(ex_ctrl_mem),
    .ZN(_08205_)
  );
  INV_X1 _15831_ (
    .A(mem_ctrl_jalr),
    .ZN(_08206_)
  );
  INV_X1 _15832_ (
    .A(ex_ctrl_jalr),
    .ZN(_08207_)
  );
  INV_X1 _15833_ (
    .A(mem_ctrl_jal),
    .ZN(_08208_)
  );
  INV_X1 _15834_ (
    .A(ex_ctrl_fence_i),
    .ZN(_08209_)
  );
  INV_X1 _15835_ (
    .A(ex_ctrl_mem_cmd[0]),
    .ZN(_08210_)
  );
  INV_X1 _15836_ (
    .A(ex_ctrl_mem_cmd[1]),
    .ZN(_08211_)
  );
  INV_X1 _15837_ (
    .A(ex_ctrl_mem_cmd[2]),
    .ZN(_08212_)
  );
  INV_X1 _15838_ (
    .A(ex_ctrl_mem_cmd[3]),
    .ZN(_08213_)
  );
  INV_X1 _15839_ (
    .A(ex_ctrl_sel_imm[0]),
    .ZN(_08214_)
  );
  INV_X1 _15840_ (
    .A(ex_ctrl_sel_imm[1]),
    .ZN(_08215_)
  );
  INV_X1 _15841_ (
    .A(ex_ctrl_sel_imm[2]),
    .ZN(_08216_)
  );
  INV_X1 _15842_ (
    .A(ex_ctrl_sel_alu1[0]),
    .ZN(_08217_)
  );
  INV_X1 _15843_ (
    .A(ex_ctrl_sel_alu1[1]),
    .ZN(_08218_)
  );
  INV_X1 _15844_ (
    .A(ex_ctrl_sel_alu2[0]),
    .ZN(_08219_)
  );
  INV_X1 _15845_ (
    .A(ex_reg_rs_lsb_1[0]),
    .ZN(_08220_)
  );
  INV_X1 _15846_ (
    .A(ex_reg_rs_lsb_1[1]),
    .ZN(_08221_)
  );
  INV_X1 _15847_ (
    .A(wb_reg_cause[0]),
    .ZN(_08222_)
  );
  INV_X1 _15848_ (
    .A(wb_reg_cause[1]),
    .ZN(_08223_)
  );
  INV_X1 _15849_ (
    .A(wb_reg_cause[2]),
    .ZN(_08224_)
  );
  INV_X1 _15850_ (
    .A(wb_reg_cause[3]),
    .ZN(_08225_)
  );
  INV_X1 _15851_ (
    .A(\rf[8] [31]),
    .ZN(_08226_)
  );
  INV_X1 _15852_ (
    .A(\rf[28] [31]),
    .ZN(_08227_)
  );
  INV_X1 _15853_ (
    .A(\rf[24] [31]),
    .ZN(_08228_)
  );
  INV_X1 _15854_ (
    .A(\rf[21] [31]),
    .ZN(_08229_)
  );
  INV_X1 _15855_ (
    .A(\rf[20] [31]),
    .ZN(_08230_)
  );
  INV_X1 _15856_ (
    .A(\rf[17] [31]),
    .ZN(_08231_)
  );
  INV_X1 _15857_ (
    .A(\rf[16] [31]),
    .ZN(_08232_)
  );
  INV_X1 _15858_ (
    .A(\rf[14] [31]),
    .ZN(_08233_)
  );
  INV_X1 _15859_ (
    .A(\rf[12] [31]),
    .ZN(_08234_)
  );
  INV_X1 _15860_ (
    .A(\rf[10] [31]),
    .ZN(_08235_)
  );
  INV_X1 _15861_ (
    .A(\rf[25] [4]),
    .ZN(_08236_)
  );
  INV_X1 _15862_ (
    .A(\rf[25] [6]),
    .ZN(_08237_)
  );
  INV_X1 _15863_ (
    .A(\rf[25] [7]),
    .ZN(_08238_)
  );
  INV_X1 _15864_ (
    .A(\rf[25] [8]),
    .ZN(_08239_)
  );
  INV_X1 _15865_ (
    .A(\rf[25] [9]),
    .ZN(_08240_)
  );
  INV_X1 _15866_ (
    .A(\rf[25] [11]),
    .ZN(_08241_)
  );
  INV_X1 _15867_ (
    .A(\rf[25] [12]),
    .ZN(_08242_)
  );
  INV_X1 _15868_ (
    .A(\rf[25] [13]),
    .ZN(_08243_)
  );
  INV_X1 _15869_ (
    .A(\rf[6] [0]),
    .ZN(_08244_)
  );
  INV_X1 _15870_ (
    .A(\rf[6] [1]),
    .ZN(_08245_)
  );
  INV_X1 _15871_ (
    .A(\rf[6] [20]),
    .ZN(_08246_)
  );
  INV_X1 _15872_ (
    .A(\rf[6] [29]),
    .ZN(_08247_)
  );
  INV_X1 _15873_ (
    .A(\rf[4] [0]),
    .ZN(_08248_)
  );
  INV_X1 _15874_ (
    .A(\rf[4] [1]),
    .ZN(_08249_)
  );
  INV_X1 _15875_ (
    .A(\rf[4] [20]),
    .ZN(_08250_)
  );
  INV_X1 _15876_ (
    .A(ex_ctrl_sel_alu2[1]),
    .ZN(_08251_)
  );
  INV_X1 _15877_ (
    .A(\rf[4] [29]),
    .ZN(_08252_)
  );
  INV_X1 _15878_ (
    .A(\rf[0] [0]),
    .ZN(_08253_)
  );
  INV_X1 _15879_ (
    .A(\rf[0] [1]),
    .ZN(_08254_)
  );
  INV_X1 _15880_ (
    .A(\rf[0] [20]),
    .ZN(_08255_)
  );
  INV_X1 _15881_ (
    .A(\rf[0] [29]),
    .ZN(_08256_)
  );
  INV_X1 _15882_ (
    .A(\rf[8] [0]),
    .ZN(_08257_)
  );
  INV_X1 _15883_ (
    .A(\rf[8] [1]),
    .ZN(_08258_)
  );
  INV_X1 _15884_ (
    .A(\rf[8] [6]),
    .ZN(_08259_)
  );
  INV_X1 _15885_ (
    .A(\rf[8] [8]),
    .ZN(_08260_)
  );
  INV_X1 _15886_ (
    .A(\rf[8] [9]),
    .ZN(_08261_)
  );
  INV_X1 _15887_ (
    .A(\rf[8] [11]),
    .ZN(_08262_)
  );
  INV_X1 _15888_ (
    .A(\rf[8] [14]),
    .ZN(_08263_)
  );
  INV_X1 _15889_ (
    .A(\rf[8] [18]),
    .ZN(_08264_)
  );
  INV_X1 _15890_ (
    .A(\rf[8] [20]),
    .ZN(_08265_)
  );
  INV_X1 _15891_ (
    .A(\rf[8] [21]),
    .ZN(_08266_)
  );
  INV_X1 _15892_ (
    .A(\rf[8] [22]),
    .ZN(_08267_)
  );
  INV_X1 _15893_ (
    .A(\rf[8] [24]),
    .ZN(_08268_)
  );
  INV_X1 _15894_ (
    .A(\rf[8] [25]),
    .ZN(_08269_)
  );
  INV_X1 _15895_ (
    .A(\rf[8] [27]),
    .ZN(_08270_)
  );
  INV_X1 _15896_ (
    .A(\rf[8] [28]),
    .ZN(_08271_)
  );
  INV_X1 _15897_ (
    .A(\rf[8] [29]),
    .ZN(_08272_)
  );
  INV_X1 _15898_ (
    .A(\rf[8] [30]),
    .ZN(_08273_)
  );
  INV_X1 _15899_ (
    .A(\rf[16] [0]),
    .ZN(_08274_)
  );
  INV_X1 _15900_ (
    .A(\rf[16] [1]),
    .ZN(_08275_)
  );
  INV_X1 _15901_ (
    .A(\rf[16] [2]),
    .ZN(_08276_)
  );
  INV_X1 _15902_ (
    .A(\rf[16] [3]),
    .ZN(_08277_)
  );
  INV_X1 _15903_ (
    .A(\rf[16] [4]),
    .ZN(_08278_)
  );
  INV_X1 _15904_ (
    .A(\rf[16] [5]),
    .ZN(_08279_)
  );
  INV_X1 _15905_ (
    .A(\rf[16] [6]),
    .ZN(_08280_)
  );
  INV_X1 _15906_ (
    .A(\rf[16] [7]),
    .ZN(_08281_)
  );
  INV_X1 _15907_ (
    .A(\rf[16] [8]),
    .ZN(_08282_)
  );
  INV_X1 _15908_ (
    .A(\rf[16] [9]),
    .ZN(_08283_)
  );
  INV_X1 _15909_ (
    .A(\rf[16] [10]),
    .ZN(_08284_)
  );
  INV_X1 _15910_ (
    .A(\rf[16] [11]),
    .ZN(_08285_)
  );
  INV_X1 _15911_ (
    .A(\rf[16] [12]),
    .ZN(_08286_)
  );
  INV_X1 _15912_ (
    .A(\rf[16] [13]),
    .ZN(_08287_)
  );
  INV_X1 _15913_ (
    .A(\rf[16] [14]),
    .ZN(_08288_)
  );
  INV_X1 _15914_ (
    .A(\rf[16] [15]),
    .ZN(_08289_)
  );
  INV_X1 _15915_ (
    .A(\rf[16] [16]),
    .ZN(_08290_)
  );
  INV_X1 _15916_ (
    .A(\rf[16] [17]),
    .ZN(_08291_)
  );
  INV_X1 _15917_ (
    .A(\rf[16] [18]),
    .ZN(_08292_)
  );
  INV_X1 _15918_ (
    .A(\rf[16] [19]),
    .ZN(_08293_)
  );
  INV_X1 _15919_ (
    .A(\rf[16] [20]),
    .ZN(_08294_)
  );
  INV_X1 _15920_ (
    .A(\rf[16] [21]),
    .ZN(_08295_)
  );
  INV_X1 _15921_ (
    .A(\rf[16] [22]),
    .ZN(_08296_)
  );
  INV_X1 _15922_ (
    .A(\rf[16] [23]),
    .ZN(_08297_)
  );
  INV_X1 _15923_ (
    .A(\rf[16] [24]),
    .ZN(_08298_)
  );
  INV_X1 _15924_ (
    .A(\rf[16] [25]),
    .ZN(_08299_)
  );
  INV_X1 _15925_ (
    .A(\rf[16] [26]),
    .ZN(_08300_)
  );
  INV_X1 _15926_ (
    .A(\rf[16] [27]),
    .ZN(_08301_)
  );
  INV_X1 _15927_ (
    .A(\rf[16] [28]),
    .ZN(_08302_)
  );
  INV_X1 _15928_ (
    .A(\rf[16] [29]),
    .ZN(_08303_)
  );
  INV_X1 _15929_ (
    .A(\rf[16] [30]),
    .ZN(_08304_)
  );
  INV_X1 _15930_ (
    .A(\rf[17] [0]),
    .ZN(_08305_)
  );
  INV_X1 _15931_ (
    .A(\rf[17] [2]),
    .ZN(_08306_)
  );
  INV_X1 _15932_ (
    .A(\rf[17] [3]),
    .ZN(_08307_)
  );
  INV_X1 _15933_ (
    .A(\rf[17] [4]),
    .ZN(_08308_)
  );
  INV_X1 _15934_ (
    .A(\rf[17] [5]),
    .ZN(_08309_)
  );
  INV_X1 _15935_ (
    .A(\rf[17] [6]),
    .ZN(_08310_)
  );
  INV_X1 _15936_ (
    .A(\rf[17] [7]),
    .ZN(_08311_)
  );
  INV_X1 _15937_ (
    .A(\rf[17] [8]),
    .ZN(_08312_)
  );
  INV_X1 _15938_ (
    .A(\rf[17] [9]),
    .ZN(_08313_)
  );
  INV_X1 _15939_ (
    .A(\rf[17] [10]),
    .ZN(_08314_)
  );
  INV_X1 _15940_ (
    .A(\rf[17] [11]),
    .ZN(_08315_)
  );
  INV_X1 _15941_ (
    .A(\rf[17] [12]),
    .ZN(_08316_)
  );
  INV_X1 _15942_ (
    .A(\rf[17] [13]),
    .ZN(_08317_)
  );
  INV_X1 _15943_ (
    .A(\rf[17] [14]),
    .ZN(_08318_)
  );
  INV_X1 _15944_ (
    .A(\rf[17] [15]),
    .ZN(_08319_)
  );
  INV_X1 _15945_ (
    .A(\rf[17] [16]),
    .ZN(_08320_)
  );
  INV_X1 _15946_ (
    .A(\rf[17] [17]),
    .ZN(_08321_)
  );
  INV_X1 _15947_ (
    .A(\rf[17] [18]),
    .ZN(_08322_)
  );
  INV_X1 _15948_ (
    .A(\rf[17] [19]),
    .ZN(_08323_)
  );
  INV_X1 _15949_ (
    .A(\rf[17] [20]),
    .ZN(_08324_)
  );
  INV_X1 _15950_ (
    .A(\rf[17] [21]),
    .ZN(_08325_)
  );
  INV_X1 _15951_ (
    .A(\rf[17] [22]),
    .ZN(_08326_)
  );
  INV_X1 _15952_ (
    .A(\rf[17] [23]),
    .ZN(_08327_)
  );
  INV_X1 _15953_ (
    .A(\rf[17] [24]),
    .ZN(_08328_)
  );
  INV_X1 _15954_ (
    .A(\rf[17] [25]),
    .ZN(_08329_)
  );
  INV_X1 _15955_ (
    .A(\rf[17] [26]),
    .ZN(_08330_)
  );
  INV_X1 _15956_ (
    .A(\rf[17] [27]),
    .ZN(_08331_)
  );
  INV_X1 _15957_ (
    .A(\rf[17] [28]),
    .ZN(_08332_)
  );
  INV_X1 _15958_ (
    .A(\rf[17] [29]),
    .ZN(_08333_)
  );
  INV_X1 _15959_ (
    .A(\rf[17] [30]),
    .ZN(_08334_)
  );
  INV_X1 _15960_ (
    .A(\rf[10] [0]),
    .ZN(_08335_)
  );
  INV_X1 _15961_ (
    .A(\rf[10] [1]),
    .ZN(_08336_)
  );
  INV_X1 _15962_ (
    .A(\rf[10] [6]),
    .ZN(_08337_)
  );
  INV_X1 _15963_ (
    .A(\rf[10] [8]),
    .ZN(_08338_)
  );
  INV_X1 _15964_ (
    .A(\rf[10] [9]),
    .ZN(_08339_)
  );
  INV_X1 _15965_ (
    .A(\rf[10] [11]),
    .ZN(_08340_)
  );
  INV_X1 _15966_ (
    .A(\rf[10] [14]),
    .ZN(_08341_)
  );
  INV_X1 _15967_ (
    .A(\rf[10] [18]),
    .ZN(_08342_)
  );
  INV_X1 _15968_ (
    .A(\rf[10] [20]),
    .ZN(_08343_)
  );
  INV_X1 _15969_ (
    .A(\rf[10] [21]),
    .ZN(_08344_)
  );
  INV_X1 _15970_ (
    .A(\rf[10] [22]),
    .ZN(_08345_)
  );
  INV_X1 _15971_ (
    .A(\rf[10] [24]),
    .ZN(_08346_)
  );
  INV_X1 _15972_ (
    .A(\rf[10] [25]),
    .ZN(_08347_)
  );
  INV_X1 _15973_ (
    .A(\rf[10] [27]),
    .ZN(_08348_)
  );
  INV_X1 _15974_ (
    .A(\rf[10] [28]),
    .ZN(_08349_)
  );
  INV_X1 _15975_ (
    .A(\rf[10] [29]),
    .ZN(_08350_)
  );
  INV_X1 _15976_ (
    .A(\rf[10] [30]),
    .ZN(_08351_)
  );
  INV_X1 _15977_ (
    .A(\rf[18] [0]),
    .ZN(_08352_)
  );
  INV_X1 _15978_ (
    .A(\rf[18] [1]),
    .ZN(_08353_)
  );
  INV_X1 _15979_ (
    .A(\rf[18] [20]),
    .ZN(_08354_)
  );
  INV_X1 _15980_ (
    .A(\rf[18] [29]),
    .ZN(_08355_)
  );
  INV_X1 _15981_ (
    .A(\rf[12] [0]),
    .ZN(_08356_)
  );
  INV_X1 _15982_ (
    .A(\rf[12] [1]),
    .ZN(_08357_)
  );
  INV_X1 _15983_ (
    .A(\rf[12] [6]),
    .ZN(_08358_)
  );
  INV_X1 _15984_ (
    .A(\rf[12] [8]),
    .ZN(_08359_)
  );
  INV_X1 _15985_ (
    .A(\rf[12] [9]),
    .ZN(_08360_)
  );
  INV_X1 _15986_ (
    .A(\rf[12] [11]),
    .ZN(_08361_)
  );
  INV_X1 _15987_ (
    .A(\rf[12] [14]),
    .ZN(_08362_)
  );
  INV_X1 _15988_ (
    .A(\rf[12] [18]),
    .ZN(_08363_)
  );
  INV_X1 _15989_ (
    .A(\rf[12] [20]),
    .ZN(_08364_)
  );
  INV_X1 _15990_ (
    .A(\rf[12] [21]),
    .ZN(_08365_)
  );
  INV_X1 _15991_ (
    .A(\rf[12] [22]),
    .ZN(_08366_)
  );
  INV_X1 _15992_ (
    .A(\rf[12] [24]),
    .ZN(_08367_)
  );
  INV_X1 _15993_ (
    .A(\rf[12] [25]),
    .ZN(_08368_)
  );
  INV_X1 _15994_ (
    .A(\rf[12] [27]),
    .ZN(_08369_)
  );
  INV_X1 _15995_ (
    .A(\rf[12] [28]),
    .ZN(_08370_)
  );
  INV_X1 _15996_ (
    .A(\rf[12] [29]),
    .ZN(_08371_)
  );
  INV_X1 _15997_ (
    .A(\rf[12] [30]),
    .ZN(_08372_)
  );
  INV_X1 _15998_ (
    .A(\rf[20] [0]),
    .ZN(_08373_)
  );
  INV_X1 _15999_ (
    .A(\rf[20] [1]),
    .ZN(_08374_)
  );
  INV_X1 _16000_ (
    .A(\rf[20] [2]),
    .ZN(_08375_)
  );
  INV_X1 _16001_ (
    .A(\rf[20] [3]),
    .ZN(_08376_)
  );
  INV_X1 _16002_ (
    .A(\rf[20] [4]),
    .ZN(_08377_)
  );
  INV_X1 _16003_ (
    .A(\rf[20] [5]),
    .ZN(_08378_)
  );
  INV_X1 _16004_ (
    .A(\rf[20] [6]),
    .ZN(_08379_)
  );
  INV_X1 _16005_ (
    .A(\rf[20] [7]),
    .ZN(_08380_)
  );
  INV_X1 _16006_ (
    .A(\rf[20] [8]),
    .ZN(_08381_)
  );
  INV_X1 _16007_ (
    .A(\rf[20] [9]),
    .ZN(_08382_)
  );
  INV_X1 _16008_ (
    .A(\rf[20] [10]),
    .ZN(_08383_)
  );
  INV_X1 _16009_ (
    .A(\rf[20] [11]),
    .ZN(_08384_)
  );
  INV_X1 _16010_ (
    .A(\rf[20] [12]),
    .ZN(_08385_)
  );
  INV_X1 _16011_ (
    .A(\rf[20] [13]),
    .ZN(_08386_)
  );
  INV_X1 _16012_ (
    .A(\rf[20] [14]),
    .ZN(_08387_)
  );
  INV_X1 _16013_ (
    .A(\rf[20] [15]),
    .ZN(_08388_)
  );
  INV_X1 _16014_ (
    .A(\rf[20] [16]),
    .ZN(_08389_)
  );
  INV_X1 _16015_ (
    .A(\rf[20] [17]),
    .ZN(_08390_)
  );
  INV_X1 _16016_ (
    .A(\rf[20] [18]),
    .ZN(_08391_)
  );
  INV_X1 _16017_ (
    .A(\rf[20] [19]),
    .ZN(_08392_)
  );
  INV_X1 _16018_ (
    .A(\rf[20] [20]),
    .ZN(_08393_)
  );
  INV_X1 _16019_ (
    .A(\rf[20] [21]),
    .ZN(_08394_)
  );
  INV_X1 _16020_ (
    .A(\rf[20] [22]),
    .ZN(_08395_)
  );
  INV_X1 _16021_ (
    .A(\rf[20] [23]),
    .ZN(_08396_)
  );
  INV_X1 _16022_ (
    .A(\rf[20] [24]),
    .ZN(_08397_)
  );
  INV_X1 _16023_ (
    .A(\rf[20] [25]),
    .ZN(_08398_)
  );
  INV_X1 _16024_ (
    .A(\rf[20] [26]),
    .ZN(_08399_)
  );
  INV_X1 _16025_ (
    .A(\rf[20] [27]),
    .ZN(_08400_)
  );
  INV_X1 _16026_ (
    .A(\rf[20] [28]),
    .ZN(_08401_)
  );
  INV_X1 _16027_ (
    .A(\rf[20] [29]),
    .ZN(_08402_)
  );
  INV_X1 _16028_ (
    .A(\rf[20] [30]),
    .ZN(_08403_)
  );
  INV_X1 _16029_ (
    .A(\rf[21] [0]),
    .ZN(_08404_)
  );
  INV_X1 _16030_ (
    .A(\rf[21] [2]),
    .ZN(_08405_)
  );
  INV_X1 _16031_ (
    .A(\rf[21] [3]),
    .ZN(_08406_)
  );
  INV_X1 _16032_ (
    .A(\rf[21] [4]),
    .ZN(_08407_)
  );
  INV_X1 _16033_ (
    .A(\rf[21] [5]),
    .ZN(_08408_)
  );
  INV_X1 _16034_ (
    .A(\rf[21] [6]),
    .ZN(_08409_)
  );
  INV_X1 _16035_ (
    .A(\rf[21] [7]),
    .ZN(_08410_)
  );
  INV_X1 _16036_ (
    .A(\rf[21] [8]),
    .ZN(_08411_)
  );
  INV_X1 _16037_ (
    .A(\rf[21] [9]),
    .ZN(_08412_)
  );
  INV_X1 _16038_ (
    .A(\rf[21] [10]),
    .ZN(_08413_)
  );
  INV_X1 _16039_ (
    .A(\rf[21] [11]),
    .ZN(_08414_)
  );
  INV_X1 _16040_ (
    .A(\rf[21] [12]),
    .ZN(_08415_)
  );
  INV_X1 _16041_ (
    .A(\rf[21] [13]),
    .ZN(_08416_)
  );
  INV_X1 _16042_ (
    .A(\rf[21] [14]),
    .ZN(_08417_)
  );
  INV_X1 _16043_ (
    .A(\rf[21] [15]),
    .ZN(_08418_)
  );
  INV_X1 _16044_ (
    .A(\rf[21] [16]),
    .ZN(_08419_)
  );
  INV_X1 _16045_ (
    .A(\rf[21] [17]),
    .ZN(_08420_)
  );
  INV_X1 _16046_ (
    .A(\rf[21] [18]),
    .ZN(_08421_)
  );
  INV_X1 _16047_ (
    .A(\rf[21] [19]),
    .ZN(_08422_)
  );
  INV_X1 _16048_ (
    .A(\rf[21] [20]),
    .ZN(_08423_)
  );
  INV_X1 _16049_ (
    .A(\rf[21] [21]),
    .ZN(_08424_)
  );
  INV_X1 _16050_ (
    .A(\rf[21] [22]),
    .ZN(_08425_)
  );
  INV_X1 _16051_ (
    .A(\rf[21] [23]),
    .ZN(_08426_)
  );
  INV_X1 _16052_ (
    .A(\rf[21] [24]),
    .ZN(_08427_)
  );
  INV_X1 _16053_ (
    .A(\rf[21] [25]),
    .ZN(_08428_)
  );
  INV_X1 _16054_ (
    .A(\rf[21] [26]),
    .ZN(_08429_)
  );
  INV_X1 _16055_ (
    .A(\rf[21] [27]),
    .ZN(_08430_)
  );
  INV_X1 _16056_ (
    .A(\rf[21] [28]),
    .ZN(_08431_)
  );
  INV_X1 _16057_ (
    .A(\rf[21] [29]),
    .ZN(_08432_)
  );
  INV_X1 _16058_ (
    .A(\rf[21] [30]),
    .ZN(_08433_)
  );
  INV_X1 _16059_ (
    .A(\rf[28] [0]),
    .ZN(_08434_)
  );
  INV_X1 _16060_ (
    .A(\rf[28] [1]),
    .ZN(_08435_)
  );
  INV_X1 _16061_ (
    .A(\rf[28] [3]),
    .ZN(_08436_)
  );
  INV_X1 _16062_ (
    .A(\rf[28] [4]),
    .ZN(_08437_)
  );
  INV_X1 _16063_ (
    .A(\rf[28] [6]),
    .ZN(_08438_)
  );
  INV_X1 _16064_ (
    .A(\rf[28] [7]),
    .ZN(_08439_)
  );
  INV_X1 _16065_ (
    .A(\rf[28] [8]),
    .ZN(_08440_)
  );
  INV_X1 _16066_ (
    .A(\rf[28] [9]),
    .ZN(_08441_)
  );
  INV_X1 _16067_ (
    .A(\rf[28] [11]),
    .ZN(_08442_)
  );
  INV_X1 _16068_ (
    .A(\rf[28] [12]),
    .ZN(_08443_)
  );
  INV_X1 _16069_ (
    .A(\rf[28] [13]),
    .ZN(_08444_)
  );
  INV_X1 _16070_ (
    .A(\rf[28] [14]),
    .ZN(_08445_)
  );
  INV_X1 _16071_ (
    .A(\rf[28] [16]),
    .ZN(_08446_)
  );
  INV_X1 _16072_ (
    .A(\rf[28] [17]),
    .ZN(_08447_)
  );
  INV_X1 _16073_ (
    .A(\rf[28] [18]),
    .ZN(_08448_)
  );
  INV_X1 _16074_ (
    .A(\rf[28] [20]),
    .ZN(_08449_)
  );
  INV_X1 _16075_ (
    .A(\rf[28] [21]),
    .ZN(_08450_)
  );
  INV_X1 _16076_ (
    .A(\rf[28] [22]),
    .ZN(_08451_)
  );
  INV_X1 _16077_ (
    .A(\rf[28] [24]),
    .ZN(_08452_)
  );
  INV_X1 _16078_ (
    .A(\rf[28] [25]),
    .ZN(_08453_)
  );
  INV_X1 _16079_ (
    .A(\rf[28] [26]),
    .ZN(_08454_)
  );
  INV_X1 _16080_ (
    .A(\rf[28] [27]),
    .ZN(_08455_)
  );
  INV_X1 _16081_ (
    .A(\rf[28] [28]),
    .ZN(_08456_)
  );
  INV_X1 _16082_ (
    .A(\rf[28] [29]),
    .ZN(_08457_)
  );
  INV_X1 _16083_ (
    .A(\rf[28] [30]),
    .ZN(_08458_)
  );
  INV_X1 _16084_ (
    .A(\rf[29] [4]),
    .ZN(_08459_)
  );
  INV_X1 _16085_ (
    .A(\rf[29] [6]),
    .ZN(_08460_)
  );
  INV_X1 _16086_ (
    .A(\rf[29] [7]),
    .ZN(_08461_)
  );
  INV_X1 _16087_ (
    .A(\rf[29] [8]),
    .ZN(_08462_)
  );
  INV_X1 _16088_ (
    .A(\rf[29] [9]),
    .ZN(_08463_)
  );
  INV_X1 _16089_ (
    .A(\rf[29] [11]),
    .ZN(_08464_)
  );
  INV_X1 _16090_ (
    .A(\rf[29] [12]),
    .ZN(_08465_)
  );
  INV_X1 _16091_ (
    .A(\rf[29] [13]),
    .ZN(_08466_)
  );
  INV_X1 _16092_ (
    .A(\rf[30] [0]),
    .ZN(_08467_)
  );
  INV_X1 _16093_ (
    .A(\rf[30] [1]),
    .ZN(_08468_)
  );
  INV_X1 _16094_ (
    .A(\rf[30] [2]),
    .ZN(_08469_)
  );
  INV_X1 _16095_ (
    .A(\rf[30] [3]),
    .ZN(_08470_)
  );
  INV_X1 _16096_ (
    .A(\rf[30] [10]),
    .ZN(_08471_)
  );
  INV_X1 _16097_ (
    .A(\rf[30] [15]),
    .ZN(_08472_)
  );
  INV_X1 _16098_ (
    .A(\rf[14] [0]),
    .ZN(_08473_)
  );
  INV_X1 _16099_ (
    .A(\rf[14] [1]),
    .ZN(_08474_)
  );
  INV_X1 _16100_ (
    .A(\rf[14] [6]),
    .ZN(_08475_)
  );
  INV_X1 _16101_ (
    .A(\rf[14] [8]),
    .ZN(_08476_)
  );
  INV_X1 _16102_ (
    .A(\rf[14] [9]),
    .ZN(_08477_)
  );
  INV_X1 _16103_ (
    .A(\rf[14] [11]),
    .ZN(_08478_)
  );
  INV_X1 _16104_ (
    .A(\rf[14] [14]),
    .ZN(_08479_)
  );
  INV_X1 _16105_ (
    .A(\rf[14] [18]),
    .ZN(_08480_)
  );
  INV_X1 _16106_ (
    .A(\rf[14] [20]),
    .ZN(_08481_)
  );
  INV_X1 _16107_ (
    .A(\rf[14] [21]),
    .ZN(_08482_)
  );
  INV_X1 _16108_ (
    .A(\rf[14] [22]),
    .ZN(_08483_)
  );
  INV_X1 _16109_ (
    .A(\rf[14] [24]),
    .ZN(_08484_)
  );
  INV_X1 _16110_ (
    .A(\rf[14] [25]),
    .ZN(_08485_)
  );
  INV_X1 _16111_ (
    .A(\rf[14] [27]),
    .ZN(_08486_)
  );
  INV_X1 _16112_ (
    .A(\rf[14] [28]),
    .ZN(_08487_)
  );
  INV_X1 _16113_ (
    .A(\rf[14] [29]),
    .ZN(_08488_)
  );
  INV_X1 _16114_ (
    .A(\rf[14] [30]),
    .ZN(_08489_)
  );
  INV_X1 _16115_ (
    .A(\rf[22] [0]),
    .ZN(_08490_)
  );
  INV_X1 _16116_ (
    .A(\rf[22] [1]),
    .ZN(_08491_)
  );
  INV_X1 _16117_ (
    .A(\rf[22] [20]),
    .ZN(_08492_)
  );
  INV_X1 _16118_ (
    .A(\rf[22] [29]),
    .ZN(_08493_)
  );
  INV_X1 _16119_ (
    .A(\rf[26] [0]),
    .ZN(_08494_)
  );
  INV_X1 _16120_ (
    .A(\rf[26] [1]),
    .ZN(_08495_)
  );
  INV_X1 _16121_ (
    .A(\rf[26] [2]),
    .ZN(_08496_)
  );
  INV_X1 _16122_ (
    .A(\rf[26] [3]),
    .ZN(_08497_)
  );
  INV_X1 _16123_ (
    .A(\rf[26] [10]),
    .ZN(_08498_)
  );
  INV_X1 _16124_ (
    .A(\rf[26] [15]),
    .ZN(_08499_)
  );
  INV_X1 _16125_ (
    .A(\rf[2] [0]),
    .ZN(_08500_)
  );
  INV_X1 _16126_ (
    .A(\rf[2] [1]),
    .ZN(_08501_)
  );
  INV_X1 _16127_ (
    .A(\rf[2] [20]),
    .ZN(_08502_)
  );
  INV_X1 _16128_ (
    .A(\rf[2] [29]),
    .ZN(_08503_)
  );
  INV_X1 _16129_ (
    .A(\rf[24] [0]),
    .ZN(_08504_)
  );
  INV_X1 _16130_ (
    .A(\rf[24] [1]),
    .ZN(_08505_)
  );
  INV_X1 _16131_ (
    .A(\rf[24] [3]),
    .ZN(_08506_)
  );
  INV_X1 _16132_ (
    .A(\rf[24] [4]),
    .ZN(_08507_)
  );
  INV_X1 _16133_ (
    .A(\rf[24] [6]),
    .ZN(_08508_)
  );
  INV_X1 _16134_ (
    .A(\rf[24] [7]),
    .ZN(_08509_)
  );
  INV_X1 _16135_ (
    .A(\rf[24] [8]),
    .ZN(_08510_)
  );
  INV_X1 _16136_ (
    .A(\rf[24] [9]),
    .ZN(_08511_)
  );
  INV_X1 _16137_ (
    .A(\rf[24] [11]),
    .ZN(_08512_)
  );
  INV_X1 _16138_ (
    .A(\rf[24] [12]),
    .ZN(_08513_)
  );
  INV_X1 _16139_ (
    .A(\rf[24] [13]),
    .ZN(_08514_)
  );
  INV_X1 _16140_ (
    .A(\rf[24] [14]),
    .ZN(_08515_)
  );
  INV_X1 _16141_ (
    .A(\rf[24] [16]),
    .ZN(_08516_)
  );
  INV_X1 _16142_ (
    .A(\rf[24] [17]),
    .ZN(_08517_)
  );
  INV_X1 _16143_ (
    .A(\rf[24] [18]),
    .ZN(_08518_)
  );
  INV_X1 _16144_ (
    .A(\rf[24] [20]),
    .ZN(_08519_)
  );
  INV_X1 _16145_ (
    .A(\rf[24] [21]),
    .ZN(_08520_)
  );
  INV_X1 _16146_ (
    .A(\rf[24] [22]),
    .ZN(_08521_)
  );
  INV_X1 _16147_ (
    .A(\rf[24] [24]),
    .ZN(_08522_)
  );
  INV_X1 _16148_ (
    .A(\rf[24] [25]),
    .ZN(_08523_)
  );
  INV_X1 _16149_ (
    .A(\rf[24] [26]),
    .ZN(_08524_)
  );
  INV_X1 _16150_ (
    .A(\rf[24] [27]),
    .ZN(_08525_)
  );
  INV_X1 _16151_ (
    .A(\rf[24] [28]),
    .ZN(_08526_)
  );
  INV_X1 _16152_ (
    .A(\rf[24] [29]),
    .ZN(_08527_)
  );
  INV_X1 _16153_ (
    .A(\rf[24] [30]),
    .ZN(_08528_)
  );
  INV_X1 _16154_ (
    .A(csr_io_decode_0_inst[6]),
    .ZN(_08529_)
  );
  INV_X1 _16155_ (
    .A(csr_io_decode_0_inst[2]),
    .ZN(_08530_)
  );
  INV_X1 _16156_ (
    .A(csr_io_decode_0_inst[5]),
    .ZN(_08531_)
  );
  INV_X1 _16157_ (
    .A(csr_io_decode_0_inst[4]),
    .ZN(_08532_)
  );
  INV_X1 _16158_ (
    .A(csr_io_decode_0_inst[3]),
    .ZN(_08533_)
  );
  INV_X1 _16159_ (
    .A(_00023_),
    .ZN(_08534_)
  );
  INV_X1 _16160_ (
    .A(_00022_),
    .ZN(_08535_)
  );
  INV_X1 _16161_ (
    .A(_00021_),
    .ZN(_08536_)
  );
  INV_X1 _16162_ (
    .A(_00020_),
    .ZN(_08537_)
  );
  INV_X1 _16163_ (
    .A(_00012_),
    .ZN(_08538_)
  );
  INV_X1 _16164_ (
    .A(_00018_),
    .ZN(_08539_)
  );
  INV_X1 _16165_ (
    .A(ibuf_io_inst_0_bits_inst_rs1[0]),
    .ZN(_08540_)
  );
  INV_X1 _16166_ (
    .A(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_08541_)
  );
  INV_X1 _16167_ (
    .A(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_08542_)
  );
  INV_X1 _16168_ (
    .A(ibuf_io_inst_0_bits_inst_rs1[3]),
    .ZN(_08543_)
  );
  INV_X1 _16169_ (
    .A(ibuf_io_inst_0_bits_inst_rs2[0]),
    .ZN(_08544_)
  );
  INV_X1 _16170_ (
    .A(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_08545_)
  );
  INV_X1 _16171_ (
    .A(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08546_)
  );
  INV_X1 _16172_ (
    .A(ibuf_io_inst_0_bits_inst_rs2[3]),
    .ZN(_08547_)
  );
  INV_X1 _16173_ (
    .A(ibuf_io_inst_0_bits_inst_rd[0]),
    .ZN(_08548_)
  );
  INV_X1 _16174_ (
    .A(ibuf_io_inst_0_bits_inst_rd[1]),
    .ZN(_08549_)
  );
  INV_X1 _16175_ (
    .A(ibuf_io_inst_0_bits_inst_rd[2]),
    .ZN(_08550_)
  );
  INV_X1 _16176_ (
    .A(ibuf_io_inst_0_bits_inst_rd[3]),
    .ZN(_08551_)
  );
  INV_X1 _16177_ (
    .A(ibuf_io_inst_0_bits_inst_rd[4]),
    .ZN(_08552_)
  );
  INV_X1 _16178_ (
    .A(_00027_),
    .ZN(_08553_)
  );
  INV_X1 _16179_ (
    .A(_00026_),
    .ZN(_08554_)
  );
  INV_X1 _16180_ (
    .A(_00025_),
    .ZN(_08555_)
  );
  INV_X1 _16181_ (
    .A(_00024_),
    .ZN(_08556_)
  );
  INV_X1 _16182_ (
    .A(_15563_[0]),
    .ZN(_08557_)
  );
  INV_X1 _16183_ (
    .A(_00016_),
    .ZN(_08558_)
  );
  INV_X1 _16184_ (
    .A(_00015_),
    .ZN(_08559_)
  );
  INV_X1 _16185_ (
    .A(_00014_),
    .ZN(_08560_)
  );
  INV_X1 _16186_ (
    .A(_00013_),
    .ZN(_08561_)
  );
  INV_X1 _16187_ (
    .A(_00030_),
    .ZN(_08562_)
  );
  INV_X1 _16188_ (
    .A(_00019_),
    .ZN(_08563_)
  );
  INV_X1 _16189_ (
    .A(ibuf_io_inst_0_bits_xcpt1_ae_inst),
    .ZN(_08564_)
  );
  INV_X1 _16190_ (
    .A(ibuf_io_inst_0_bits_xcpt1_gf_inst),
    .ZN(_08565_)
  );
  INV_X1 _16191_ (
    .A(ibuf_io_inst_0_bits_xcpt1_pf_inst),
    .ZN(_08566_)
  );
  INV_X1 _16192_ (
    .A(_00032_),
    .ZN(_08567_)
  );
  INV_X1 _16193_ (
    .A(_00031_),
    .ZN(_08568_)
  );
  INV_X1 _16194_ (
    .A(_00017_),
    .ZN(_08569_)
  );
  INV_X1 _16195_ (
    .A(_00035_),
    .ZN(_08570_)
  );
  INV_X1 _16196_ (
    .A(ibuf_io_inst_0_bits_inst_rs1[4]),
    .ZN(_08571_)
  );
  INV_X1 _16197_ (
    .A(ibuf_io_inst_0_bits_inst_rs2[4]),
    .ZN(_08572_)
  );
  INV_X1 _16198_ (
    .A(csr_io_time[0]),
    .ZN(_08573_)
  );
  INV_X1 _16199_ (
    .A(csr_io_time[1]),
    .ZN(_08574_)
  );
  INV_X1 _16200_ (
    .A(csr_io_time[2]),
    .ZN(_08575_)
  );
  INV_X1 _16201_ (
    .A(csr_io_time[3]),
    .ZN(_08576_)
  );
  INV_X1 _16202_ (
    .A(csr_io_time[4]),
    .ZN(_08577_)
  );
  INV_X1 _16203_ (
    .A(ibuf_io_inst_0_bits_rvc),
    .ZN(_08578_)
  );
  INV_X1 _16204_ (
    .A(csr_io_interrupt_cause[1]),
    .ZN(_08579_)
  );
  INV_X1 _16205_ (
    .A(csr_io_interrupt_cause[2]),
    .ZN(_08580_)
  );
  INV_X1 _16206_ (
    .A(ibuf_io_inst_0_bits_xcpt0_ae_inst),
    .ZN(_08581_)
  );
  INV_X1 _16207_ (
    .A(bpu_io_xcpt_if),
    .ZN(_08582_)
  );
  INV_X1 _16208_ (
    .A(bpu_io_debug_if),
    .ZN(_08583_)
  );
  INV_X1 _16209_ (
    .A(div_io_resp_bits_tag[0]),
    .ZN(_08584_)
  );
  INV_X1 _16210_ (
    .A(io_dmem_resp_bits_tag[1]),
    .ZN(_08585_)
  );
  INV_X1 _16211_ (
    .A(div_io_resp_bits_tag[1]),
    .ZN(_08586_)
  );
  INV_X1 _16212_ (
    .A(io_dmem_resp_bits_tag[2]),
    .ZN(_08587_)
  );
  INV_X1 _16213_ (
    .A(div_io_resp_bits_tag[2]),
    .ZN(_08588_)
  );
  INV_X1 _16214_ (
    .A(io_dmem_resp_bits_tag[3]),
    .ZN(_08589_)
  );
  INV_X1 _16215_ (
    .A(div_io_resp_bits_tag[3]),
    .ZN(_08590_)
  );
  INV_X1 _16216_ (
    .A(io_dmem_resp_bits_tag[4]),
    .ZN(_08591_)
  );
  INV_X1 _16217_ (
    .A(div_io_resp_bits_tag[4]),
    .ZN(_08592_)
  );
  INV_X1 _16218_ (
    .A(io_dmem_resp_bits_tag[5]),
    .ZN(_08593_)
  );
  INV_X1 _16219_ (
    .A(csr_io_evec[1]),
    .ZN(_08594_)
  );
  INV_X1 _16220_ (
    .A(wb_reg_xcpt),
    .ZN(_08595_)
  );
  INV_X1 _16221_ (
    .A(mem_reg_xcpt),
    .ZN(_08596_)
  );
  INV_X1 _16222_ (
    .A(csr_io_status_isa[12]),
    .ZN(_08597_)
  );
  INV_X1 _16223_ (
    .A(csr_io_status_isa[0]),
    .ZN(_08598_)
  );
  INV_X1 _16224_ (
    .A(csr_io_status_isa[2]),
    .ZN(_08599_)
  );
  INV_X1 _16225_ (
    .A(io_dmem_resp_valid),
    .ZN(_08600_)
  );
  INV_X1 _16226_ (
    .A(io_dmem_resp_bits_tag[0]),
    .ZN(_08601_)
  );
  INV_X1 _16227_ (
    .A(io_dmem_perf_grant),
    .ZN(_08602_)
  );
  INV_X1 _16228_ (
    .A(ibuf_io_inst_0_valid),
    .ZN(_08603_)
  );
  INV_X1 _16229_ (
    .A(div_io_req_ready),
    .ZN(_08604_)
  );
  INV_X1 _16230_ (
    .A(io_dmem_req_ready),
    .ZN(_08605_)
  );
  INV_X1 _16231_ (
    .A(ex_reg_valid),
    .ZN(_08606_)
  );
  INV_X1 _16232_ (
    .A(mem_reg_valid),
    .ZN(_08607_)
  );
  INV_X1 _16233_ (
    .A(io_dmem_s2_nack),
    .ZN(_08608_)
  );
  INV_X1 _16234_ (
    .A(wb_reg_replay),
    .ZN(_08609_)
  );
  INV_X1 _16235_ (
    .A(wb_reg_valid),
    .ZN(_08610_)
  );
  INV_X1 _16236_ (
    .A(io_dmem_s2_xcpt_ae_ld),
    .ZN(_08611_)
  );
  INV_X1 _16237_ (
    .A(csr_io_eret),
    .ZN(_08612_)
  );
  INV_X1 _16238_ (
    .A(wb_reg_flush_pipe),
    .ZN(_08613_)
  );
  INV_X1 _16239_ (
    .A(csr_io_decode_0_read_illegal),
    .ZN(_08614_)
  );
  INV_X1 _16240_ (
    .A(blocked),
    .ZN(_08615_)
  );
  INV_X1 _16241_ (
    .A(csr_io_csr_stall),
    .ZN(_08616_)
  );
  INV_X1 _16242_ (
    .A(ibuf_io_inst_0_bits_replay),
    .ZN(_08617_)
  );
  INV_X1 _16243_ (
    .A(ex_reg_replay),
    .ZN(_08618_)
  );
  INV_X1 _16244_ (
    .A(ex_reg_xcpt_interrupt),
    .ZN(_08619_)
  );
  INV_X1 _16245_ (
    .A(_00034_),
    .ZN(_08620_)
  );
  INV_X1 _16246_ (
    .A(_15564_[1]),
    .ZN(_08621_)
  );
  INV_X1 _16247_ (
    .A(ex_reg_xcpt),
    .ZN(_08622_)
  );
  INV_X1 _16248_ (
    .A(mem_reg_replay),
    .ZN(_08623_)
  );
  INV_X1 _16249_ (
    .A(mem_reg_xcpt_interrupt),
    .ZN(_08624_)
  );
  INV_X1 _16250_ (
    .A(io_imem_resp_valid),
    .ZN(_08625_)
  );
  INV_X1 _16251_ (
    .A(_00033_),
    .ZN(_08626_)
  );
  INV_X1 _16252_ (
    .A(tval_dmem_addr),
    .ZN(_08627_)
  );
  INV_X1 _16253_ (
    .A(csr_io_inhibit_cycle),
    .ZN(_08628_)
  );
  INV_X1 _16254_ (
    .A(io_ptw_customCSRs_csrs_0_value[1]),
    .ZN(_08629_)
  );
  AND2_X1 _16255_ (
    .A1(io_dmem_resp_valid),
    .A2(io_dmem_resp_bits_has_data),
    .ZN(_08630_)
  );
  AND2_X1 _16256_ (
    .A1(_08601_),
    .A2(_08630_),
    .ZN(_08631_)
  );
  AND2_X1 _16257_ (
    .A1(io_dmem_resp_bits_replay),
    .A2(_08631_),
    .ZN(_08632_)
  );
  INV_X1 _16258_ (
    .A(_08632_),
    .ZN(_08633_)
  );
  MUX2_X1 _16259_ (
    .A(_08584_),
    .B(_08585_),
    .S(_08632_),
    .Z(_08634_)
  );
  MUX2_X1 _16260_ (
    .A(div_io_resp_bits_tag[0]),
    .B(io_dmem_resp_bits_tag[1]),
    .S(_08632_),
    .Z(_08635_)
  );
  MUX2_X1 _16261_ (
    .A(_08586_),
    .B(_08587_),
    .S(_08632_),
    .Z(_08636_)
  );
  MUX2_X1 _16262_ (
    .A(div_io_resp_bits_tag[1]),
    .B(io_dmem_resp_bits_tag[2]),
    .S(_08632_),
    .Z(_08637_)
  );
  AND2_X1 _16263_ (
    .A1(_08635_),
    .A2(_08636_),
    .ZN(_08638_)
  );
  MUX2_X1 _16264_ (
    .A(_08588_),
    .B(_08589_),
    .S(_08632_),
    .Z(_08639_)
  );
  MUX2_X1 _16265_ (
    .A(div_io_resp_bits_tag[2]),
    .B(io_dmem_resp_bits_tag[3]),
    .S(_08632_),
    .Z(_08640_)
  );
  AND2_X1 _16266_ (
    .A1(_08638_),
    .A2(_08639_),
    .ZN(_08641_)
  );
  MUX2_X1 _16267_ (
    .A(_08590_),
    .B(_08591_),
    .S(_08632_),
    .Z(_08642_)
  );
  MUX2_X1 _16268_ (
    .A(div_io_resp_bits_tag[3]),
    .B(io_dmem_resp_bits_tag[4]),
    .S(_08632_),
    .Z(_08643_)
  );
  MUX2_X1 _16269_ (
    .A(_08592_),
    .B(_08593_),
    .S(_08632_),
    .Z(_08644_)
  );
  MUX2_X1 _16270_ (
    .A(div_io_resp_bits_tag[4]),
    .B(io_dmem_resp_bits_tag[5]),
    .S(_08632_),
    .Z(_08645_)
  );
  AND2_X1 _16271_ (
    .A1(wb_ctrl_wxd),
    .A2(wb_reg_valid),
    .ZN(_08646_)
  );
  INV_X1 _16272_ (
    .A(_08646_),
    .ZN(_08647_)
  );
  AND2_X1 _16273_ (
    .A1(div_io_resp_valid),
    .A2(_08647_),
    .ZN(_08648_)
  );
  INV_X1 _16274_ (
    .A(_08648_),
    .ZN(_08649_)
  );
  AND2_X1 _16275_ (
    .A1(_08633_),
    .A2(_08649_),
    .ZN(_08650_)
  );
  INV_X1 _16276_ (
    .A(_08650_),
    .ZN(_08651_)
  );
  AND2_X1 _16277_ (
    .A1(_08644_),
    .A2(_08651_),
    .ZN(_08652_)
  );
  AND2_X1 _16278_ (
    .A1(_08642_),
    .A2(_08652_),
    .ZN(_08653_)
  );
  AND2_X1 _16279_ (
    .A1(_08641_),
    .A2(_08653_),
    .ZN(_08654_)
  );
  INV_X1 _16280_ (
    .A(_08654_),
    .ZN(_08655_)
  );
  AND2_X1 _16281_ (
    .A1(_r[1]),
    .A2(_08655_),
    .ZN(_08656_)
  );
  INV_X1 _16282_ (
    .A(_08656_),
    .ZN(_08657_)
  );
  AND2_X1 _16283_ (
    .A1(wb_reg_inst[7]),
    .A2(_08197_),
    .ZN(_08658_)
  );
  AND2_X1 _16284_ (
    .A1(_08198_),
    .A2(_08658_),
    .ZN(_08659_)
  );
  AND2_X1 _16285_ (
    .A1(_08199_),
    .A2(_08659_),
    .ZN(_08660_)
  );
  AND2_X1 _16286_ (
    .A1(wb_ctrl_mem),
    .A2(_08600_),
    .ZN(_08661_)
  );
  INV_X1 _16287_ (
    .A(_08661_),
    .ZN(_08662_)
  );
  AND2_X1 _16288_ (
    .A1(_08194_),
    .A2(_08662_),
    .ZN(_08663_)
  );
  INV_X1 _16289_ (
    .A(_08663_),
    .ZN(_08664_)
  );
  AND2_X1 _16290_ (
    .A1(wb_ctrl_mem),
    .A2(wb_reg_valid),
    .ZN(_08665_)
  );
  AND2_X1 _16291_ (
    .A1(io_dmem_s2_xcpt_pf_st),
    .A2(_08665_),
    .ZN(_08666_)
  );
  INV_X1 _16292_ (
    .A(_08666_),
    .ZN(_08667_)
  );
  AND2_X1 _16293_ (
    .A1(io_dmem_s2_xcpt_pf_ld),
    .A2(_08665_),
    .ZN(_08668_)
  );
  INV_X1 _16294_ (
    .A(_08668_),
    .ZN(_08669_)
  );
  AND2_X1 _16295_ (
    .A1(_08595_),
    .A2(_08669_),
    .ZN(_08670_)
  );
  AND2_X1 _16296_ (
    .A1(_08667_),
    .A2(_08670_),
    .ZN(_08671_)
  );
  INV_X1 _16297_ (
    .A(_08671_),
    .ZN(_08672_)
  );
  AND2_X1 _16298_ (
    .A1(io_dmem_s2_xcpt_ae_ld),
    .A2(_08665_),
    .ZN(_08673_)
  );
  INV_X1 _16299_ (
    .A(_08673_),
    .ZN(_08674_)
  );
  AND2_X1 _16300_ (
    .A1(io_dmem_s2_xcpt_ae_st),
    .A2(_08665_),
    .ZN(_08675_)
  );
  INV_X1 _16301_ (
    .A(_08675_),
    .ZN(_08676_)
  );
  AND2_X1 _16302_ (
    .A1(_08674_),
    .A2(_08676_),
    .ZN(_08677_)
  );
  AND2_X1 _16303_ (
    .A1(_08671_),
    .A2(_08677_),
    .ZN(_08678_)
  );
  INV_X1 _16304_ (
    .A(_08678_),
    .ZN(_08679_)
  );
  AND2_X1 _16305_ (
    .A1(io_dmem_s2_xcpt_ma_ld),
    .A2(_08665_),
    .ZN(_08680_)
  );
  INV_X1 _16306_ (
    .A(_08680_),
    .ZN(_08681_)
  );
  AND2_X1 _16307_ (
    .A1(io_dmem_s2_xcpt_ma_st),
    .A2(_08665_),
    .ZN(_08682_)
  );
  INV_X1 _16308_ (
    .A(_08682_),
    .ZN(_08683_)
  );
  AND2_X1 _16309_ (
    .A1(_08681_),
    .A2(_08683_),
    .ZN(_08684_)
  );
  AND2_X1 _16310_ (
    .A1(_08678_),
    .A2(_08684_),
    .ZN(_08685_)
  );
  INV_X1 _16311_ (
    .A(_08685_),
    .ZN(csr_io_exception)
  );
  AND2_X1 _16312_ (
    .A1(_08608_),
    .A2(_08609_),
    .ZN(_08686_)
  );
  INV_X1 _16313_ (
    .A(_08686_),
    .ZN(_08687_)
  );
  AND2_X1 _16314_ (
    .A1(wb_reg_valid),
    .A2(_08686_),
    .ZN(_08688_)
  );
  AND2_X1 _16315_ (
    .A1(_08685_),
    .A2(_08688_),
    .ZN(csr_io_retire)
  );
  AND2_X1 _16316_ (
    .A1(wb_ctrl_wxd),
    .A2(csr_io_retire),
    .ZN(_08689_)
  );
  INV_X1 _16317_ (
    .A(_08689_),
    .ZN(_08690_)
  );
  AND2_X1 _16318_ (
    .A1(_08664_),
    .A2(_08689_),
    .ZN(_08691_)
  );
  AND2_X1 _16319_ (
    .A1(_08200_),
    .A2(_08691_),
    .ZN(_08692_)
  );
  AND2_X1 _16320_ (
    .A1(_08660_),
    .A2(_08692_),
    .ZN(_08693_)
  );
  INV_X1 _16321_ (
    .A(_08693_),
    .ZN(_08694_)
  );
  AND2_X1 _16322_ (
    .A1(_08657_),
    .A2(_08694_),
    .ZN(_08695_)
  );
  INV_X1 _16323_ (
    .A(_08695_),
    .ZN(_08696_)
  );
  AND2_X1 _16324_ (
    .A1(_07954_),
    .A2(_08696_),
    .ZN(_00036_)
  );
  AND2_X1 _16325_ (
    .A1(_08634_),
    .A2(_08637_),
    .ZN(_08697_)
  );
  AND2_X1 _16326_ (
    .A1(_08639_),
    .A2(_08697_),
    .ZN(_08698_)
  );
  AND2_X1 _16327_ (
    .A1(_08653_),
    .A2(_08698_),
    .ZN(_08699_)
  );
  INV_X1 _16328_ (
    .A(_08699_),
    .ZN(_08700_)
  );
  AND2_X1 _16329_ (
    .A1(_r[2]),
    .A2(_08700_),
    .ZN(_08701_)
  );
  INV_X1 _16330_ (
    .A(_08701_),
    .ZN(_08702_)
  );
  AND2_X1 _16331_ (
    .A1(wb_reg_inst[8]),
    .A2(_00029_),
    .ZN(_08703_)
  );
  AND2_X1 _16332_ (
    .A1(_08198_),
    .A2(_08703_),
    .ZN(_08704_)
  );
  AND2_X1 _16333_ (
    .A1(_08199_),
    .A2(_08704_),
    .ZN(_08705_)
  );
  AND2_X1 _16334_ (
    .A1(_08692_),
    .A2(_08705_),
    .ZN(_08706_)
  );
  INV_X1 _16335_ (
    .A(_08706_),
    .ZN(_08707_)
  );
  AND2_X1 _16336_ (
    .A1(_08702_),
    .A2(_08707_),
    .ZN(_08708_)
  );
  INV_X1 _16337_ (
    .A(_08708_),
    .ZN(_08709_)
  );
  AND2_X1 _16338_ (
    .A1(_07954_),
    .A2(_08709_),
    .ZN(_00037_)
  );
  AND2_X1 _16339_ (
    .A1(_08635_),
    .A2(_08637_),
    .ZN(_08710_)
  );
  AND2_X1 _16340_ (
    .A1(_08639_),
    .A2(_08710_),
    .ZN(_08711_)
  );
  AND2_X1 _16341_ (
    .A1(_08653_),
    .A2(_08711_),
    .ZN(_08712_)
  );
  INV_X1 _16342_ (
    .A(_08712_),
    .ZN(_08713_)
  );
  AND2_X1 _16343_ (
    .A1(_r[3]),
    .A2(_08713_),
    .ZN(_08714_)
  );
  INV_X1 _16344_ (
    .A(_08714_),
    .ZN(_08715_)
  );
  AND2_X1 _16345_ (
    .A1(wb_reg_inst[7]),
    .A2(wb_reg_inst[8]),
    .ZN(_08716_)
  );
  AND2_X1 _16346_ (
    .A1(_08198_),
    .A2(_08716_),
    .ZN(_08717_)
  );
  AND2_X1 _16347_ (
    .A1(_08199_),
    .A2(_08717_),
    .ZN(_08718_)
  );
  AND2_X1 _16348_ (
    .A1(_08692_),
    .A2(_08718_),
    .ZN(_08719_)
  );
  INV_X1 _16349_ (
    .A(_08719_),
    .ZN(_08720_)
  );
  AND2_X1 _16350_ (
    .A1(_08715_),
    .A2(_08720_),
    .ZN(_08721_)
  );
  INV_X1 _16351_ (
    .A(_08721_),
    .ZN(_08722_)
  );
  AND2_X1 _16352_ (
    .A1(_07954_),
    .A2(_08722_),
    .ZN(_00038_)
  );
  AND2_X1 _16353_ (
    .A1(_08634_),
    .A2(_08636_),
    .ZN(_08723_)
  );
  AND2_X1 _16354_ (
    .A1(_08640_),
    .A2(_08723_),
    .ZN(_08724_)
  );
  AND2_X1 _16355_ (
    .A1(_08653_),
    .A2(_08724_),
    .ZN(_08725_)
  );
  INV_X1 _16356_ (
    .A(_08725_),
    .ZN(_08726_)
  );
  AND2_X1 _16357_ (
    .A1(_r[4]),
    .A2(_08726_),
    .ZN(_08727_)
  );
  INV_X1 _16358_ (
    .A(_08727_),
    .ZN(_08728_)
  );
  AND2_X1 _16359_ (
    .A1(_08197_),
    .A2(_00029_),
    .ZN(_08729_)
  );
  AND2_X1 _16360_ (
    .A1(wb_reg_inst[9]),
    .A2(_08729_),
    .ZN(_08730_)
  );
  AND2_X1 _16361_ (
    .A1(_08199_),
    .A2(_08730_),
    .ZN(_08731_)
  );
  AND2_X1 _16362_ (
    .A1(_08692_),
    .A2(_08731_),
    .ZN(_08732_)
  );
  INV_X1 _16363_ (
    .A(_08732_),
    .ZN(_08733_)
  );
  AND2_X1 _16364_ (
    .A1(_08728_),
    .A2(_08733_),
    .ZN(_08734_)
  );
  INV_X1 _16365_ (
    .A(_08734_),
    .ZN(_08735_)
  );
  AND2_X1 _16366_ (
    .A1(_07954_),
    .A2(_08735_),
    .ZN(_00039_)
  );
  AND2_X1 _16367_ (
    .A1(_08638_),
    .A2(_08640_),
    .ZN(_08736_)
  );
  AND2_X1 _16368_ (
    .A1(_08653_),
    .A2(_08736_),
    .ZN(_08737_)
  );
  INV_X1 _16369_ (
    .A(_08737_),
    .ZN(_08738_)
  );
  AND2_X1 _16370_ (
    .A1(_r[5]),
    .A2(_08738_),
    .ZN(_08739_)
  );
  INV_X1 _16371_ (
    .A(_08739_),
    .ZN(_08740_)
  );
  AND2_X1 _16372_ (
    .A1(wb_reg_inst[9]),
    .A2(_08658_),
    .ZN(_08741_)
  );
  AND2_X1 _16373_ (
    .A1(_08199_),
    .A2(_08741_),
    .ZN(_08742_)
  );
  AND2_X1 _16374_ (
    .A1(_08692_),
    .A2(_08742_),
    .ZN(_08743_)
  );
  INV_X1 _16375_ (
    .A(_08743_),
    .ZN(_08744_)
  );
  AND2_X1 _16376_ (
    .A1(_08740_),
    .A2(_08744_),
    .ZN(_08745_)
  );
  INV_X1 _16377_ (
    .A(_08745_),
    .ZN(_08746_)
  );
  AND2_X1 _16378_ (
    .A1(_07954_),
    .A2(_08746_),
    .ZN(_00040_)
  );
  AND2_X1 _16379_ (
    .A1(_08640_),
    .A2(_08697_),
    .ZN(_08747_)
  );
  AND2_X1 _16380_ (
    .A1(_08653_),
    .A2(_08747_),
    .ZN(_08748_)
  );
  INV_X1 _16381_ (
    .A(_08748_),
    .ZN(_08749_)
  );
  AND2_X1 _16382_ (
    .A1(_r[6]),
    .A2(_08749_),
    .ZN(_08750_)
  );
  INV_X1 _16383_ (
    .A(_08750_),
    .ZN(_08751_)
  );
  AND2_X1 _16384_ (
    .A1(wb_reg_inst[9]),
    .A2(_08703_),
    .ZN(_08752_)
  );
  AND2_X1 _16385_ (
    .A1(_08199_),
    .A2(_08752_),
    .ZN(_08753_)
  );
  AND2_X1 _16386_ (
    .A1(_08692_),
    .A2(_08753_),
    .ZN(_08754_)
  );
  INV_X1 _16387_ (
    .A(_08754_),
    .ZN(_08755_)
  );
  AND2_X1 _16388_ (
    .A1(_08751_),
    .A2(_08755_),
    .ZN(_08756_)
  );
  INV_X1 _16389_ (
    .A(_08756_),
    .ZN(_08757_)
  );
  AND2_X1 _16390_ (
    .A1(_07954_),
    .A2(_08757_),
    .ZN(_00041_)
  );
  AND2_X1 _16391_ (
    .A1(_08640_),
    .A2(_08710_),
    .ZN(_08758_)
  );
  AND2_X1 _16392_ (
    .A1(_08653_),
    .A2(_08758_),
    .ZN(_08759_)
  );
  INV_X1 _16393_ (
    .A(_08759_),
    .ZN(_08760_)
  );
  AND2_X1 _16394_ (
    .A1(_r[7]),
    .A2(_08760_),
    .ZN(_08761_)
  );
  INV_X1 _16395_ (
    .A(_08761_),
    .ZN(_08762_)
  );
  AND2_X1 _16396_ (
    .A1(wb_reg_inst[9]),
    .A2(_08716_),
    .ZN(_08763_)
  );
  AND2_X1 _16397_ (
    .A1(_08199_),
    .A2(_08763_),
    .ZN(_08764_)
  );
  AND2_X1 _16398_ (
    .A1(_08692_),
    .A2(_08764_),
    .ZN(_08765_)
  );
  INV_X1 _16399_ (
    .A(_08765_),
    .ZN(_08766_)
  );
  AND2_X1 _16400_ (
    .A1(_08762_),
    .A2(_08766_),
    .ZN(_08767_)
  );
  INV_X1 _16401_ (
    .A(_08767_),
    .ZN(_08768_)
  );
  AND2_X1 _16402_ (
    .A1(_07954_),
    .A2(_08768_),
    .ZN(_00042_)
  );
  AND2_X1 _16403_ (
    .A1(_08639_),
    .A2(_08723_),
    .ZN(_08769_)
  );
  AND2_X1 _16404_ (
    .A1(_08643_),
    .A2(_08769_),
    .ZN(_08770_)
  );
  AND2_X1 _16405_ (
    .A1(_08652_),
    .A2(_08770_),
    .ZN(_08771_)
  );
  INV_X1 _16406_ (
    .A(_08771_),
    .ZN(_08772_)
  );
  AND2_X1 _16407_ (
    .A1(_r[8]),
    .A2(_08772_),
    .ZN(_08773_)
  );
  INV_X1 _16408_ (
    .A(_08773_),
    .ZN(_08774_)
  );
  AND2_X1 _16409_ (
    .A1(_08198_),
    .A2(_08729_),
    .ZN(_08775_)
  );
  AND2_X1 _16410_ (
    .A1(wb_reg_inst[10]),
    .A2(_08691_),
    .ZN(_08776_)
  );
  AND2_X1 _16411_ (
    .A1(_08775_),
    .A2(_08776_),
    .ZN(_08777_)
  );
  AND2_X1 _16412_ (
    .A1(_08200_),
    .A2(_08777_),
    .ZN(_08778_)
  );
  INV_X1 _16413_ (
    .A(_08778_),
    .ZN(_08779_)
  );
  AND2_X1 _16414_ (
    .A1(_08774_),
    .A2(_08779_),
    .ZN(_08780_)
  );
  INV_X1 _16415_ (
    .A(_08780_),
    .ZN(_08781_)
  );
  AND2_X1 _16416_ (
    .A1(_07954_),
    .A2(_08781_),
    .ZN(_00043_)
  );
  AND2_X1 _16417_ (
    .A1(_08641_),
    .A2(_08643_),
    .ZN(_08782_)
  );
  AND2_X1 _16418_ (
    .A1(_08652_),
    .A2(_08782_),
    .ZN(_08783_)
  );
  INV_X1 _16419_ (
    .A(_08783_),
    .ZN(_08784_)
  );
  AND2_X1 _16420_ (
    .A1(_r[9]),
    .A2(_08784_),
    .ZN(_08785_)
  );
  INV_X1 _16421_ (
    .A(_08785_),
    .ZN(_08786_)
  );
  AND2_X1 _16422_ (
    .A1(_08659_),
    .A2(_08776_),
    .ZN(_08787_)
  );
  AND2_X1 _16423_ (
    .A1(_08200_),
    .A2(_08787_),
    .ZN(_08788_)
  );
  INV_X1 _16424_ (
    .A(_08788_),
    .ZN(_08789_)
  );
  AND2_X1 _16425_ (
    .A1(_08786_),
    .A2(_08789_),
    .ZN(_08790_)
  );
  INV_X1 _16426_ (
    .A(_08790_),
    .ZN(_08791_)
  );
  AND2_X1 _16427_ (
    .A1(_07954_),
    .A2(_08791_),
    .ZN(_00044_)
  );
  AND2_X1 _16428_ (
    .A1(_08643_),
    .A2(_08698_),
    .ZN(_08792_)
  );
  AND2_X1 _16429_ (
    .A1(_08652_),
    .A2(_08792_),
    .ZN(_08793_)
  );
  INV_X1 _16430_ (
    .A(_08793_),
    .ZN(_08794_)
  );
  AND2_X1 _16431_ (
    .A1(_r[10]),
    .A2(_08794_),
    .ZN(_08795_)
  );
  INV_X1 _16432_ (
    .A(_08795_),
    .ZN(_08796_)
  );
  AND2_X1 _16433_ (
    .A1(_08704_),
    .A2(_08776_),
    .ZN(_08797_)
  );
  AND2_X1 _16434_ (
    .A1(_08200_),
    .A2(_08797_),
    .ZN(_08798_)
  );
  INV_X1 _16435_ (
    .A(_08798_),
    .ZN(_08799_)
  );
  AND2_X1 _16436_ (
    .A1(_08796_),
    .A2(_08799_),
    .ZN(_08800_)
  );
  INV_X1 _16437_ (
    .A(_08800_),
    .ZN(_08801_)
  );
  AND2_X1 _16438_ (
    .A1(_07954_),
    .A2(_08801_),
    .ZN(_00045_)
  );
  AND2_X1 _16439_ (
    .A1(_08643_),
    .A2(_08711_),
    .ZN(_08802_)
  );
  AND2_X1 _16440_ (
    .A1(_08652_),
    .A2(_08802_),
    .ZN(_08803_)
  );
  INV_X1 _16441_ (
    .A(_08803_),
    .ZN(_08804_)
  );
  AND2_X1 _16442_ (
    .A1(_r[11]),
    .A2(_08804_),
    .ZN(_08805_)
  );
  INV_X1 _16443_ (
    .A(_08805_),
    .ZN(_08806_)
  );
  AND2_X1 _16444_ (
    .A1(_08717_),
    .A2(_08776_),
    .ZN(_08807_)
  );
  AND2_X1 _16445_ (
    .A1(_08200_),
    .A2(_08807_),
    .ZN(_08808_)
  );
  INV_X1 _16446_ (
    .A(_08808_),
    .ZN(_08809_)
  );
  AND2_X1 _16447_ (
    .A1(_08806_),
    .A2(_08809_),
    .ZN(_08810_)
  );
  INV_X1 _16448_ (
    .A(_08810_),
    .ZN(_08811_)
  );
  AND2_X1 _16449_ (
    .A1(_07954_),
    .A2(_08811_),
    .ZN(_00046_)
  );
  AND2_X1 _16450_ (
    .A1(_08643_),
    .A2(_08724_),
    .ZN(_08812_)
  );
  AND2_X1 _16451_ (
    .A1(_08652_),
    .A2(_08812_),
    .ZN(_08813_)
  );
  INV_X1 _16452_ (
    .A(_08813_),
    .ZN(_08814_)
  );
  AND2_X1 _16453_ (
    .A1(_r[12]),
    .A2(_08814_),
    .ZN(_08815_)
  );
  INV_X1 _16454_ (
    .A(_08815_),
    .ZN(_08816_)
  );
  AND2_X1 _16455_ (
    .A1(_08730_),
    .A2(_08776_),
    .ZN(_08817_)
  );
  AND2_X1 _16456_ (
    .A1(_08200_),
    .A2(_08817_),
    .ZN(_08818_)
  );
  INV_X1 _16457_ (
    .A(_08818_),
    .ZN(_08819_)
  );
  AND2_X1 _16458_ (
    .A1(_08816_),
    .A2(_08819_),
    .ZN(_08820_)
  );
  INV_X1 _16459_ (
    .A(_08820_),
    .ZN(_08821_)
  );
  AND2_X1 _16460_ (
    .A1(_07954_),
    .A2(_08821_),
    .ZN(_00047_)
  );
  AND2_X1 _16461_ (
    .A1(_08643_),
    .A2(_08736_),
    .ZN(_08822_)
  );
  AND2_X1 _16462_ (
    .A1(_08652_),
    .A2(_08822_),
    .ZN(_08823_)
  );
  INV_X1 _16463_ (
    .A(_08823_),
    .ZN(_08824_)
  );
  AND2_X1 _16464_ (
    .A1(_r[13]),
    .A2(_08824_),
    .ZN(_08825_)
  );
  INV_X1 _16465_ (
    .A(_08825_),
    .ZN(_08826_)
  );
  AND2_X1 _16466_ (
    .A1(_08741_),
    .A2(_08776_),
    .ZN(_08827_)
  );
  AND2_X1 _16467_ (
    .A1(_08200_),
    .A2(_08827_),
    .ZN(_08828_)
  );
  INV_X1 _16468_ (
    .A(_08828_),
    .ZN(_08829_)
  );
  AND2_X1 _16469_ (
    .A1(_08826_),
    .A2(_08829_),
    .ZN(_08830_)
  );
  INV_X1 _16470_ (
    .A(_08830_),
    .ZN(_08831_)
  );
  AND2_X1 _16471_ (
    .A1(_07954_),
    .A2(_08831_),
    .ZN(_00048_)
  );
  AND2_X1 _16472_ (
    .A1(_08643_),
    .A2(_08747_),
    .ZN(_08832_)
  );
  AND2_X1 _16473_ (
    .A1(_08652_),
    .A2(_08832_),
    .ZN(_08833_)
  );
  INV_X1 _16474_ (
    .A(_08833_),
    .ZN(_08834_)
  );
  AND2_X1 _16475_ (
    .A1(_r[14]),
    .A2(_08834_),
    .ZN(_08835_)
  );
  INV_X1 _16476_ (
    .A(_08835_),
    .ZN(_08836_)
  );
  AND2_X1 _16477_ (
    .A1(_08752_),
    .A2(_08776_),
    .ZN(_08837_)
  );
  AND2_X1 _16478_ (
    .A1(_08200_),
    .A2(_08837_),
    .ZN(_08838_)
  );
  INV_X1 _16479_ (
    .A(_08838_),
    .ZN(_08839_)
  );
  AND2_X1 _16480_ (
    .A1(_08836_),
    .A2(_08839_),
    .ZN(_08840_)
  );
  INV_X1 _16481_ (
    .A(_08840_),
    .ZN(_08841_)
  );
  AND2_X1 _16482_ (
    .A1(_07954_),
    .A2(_08841_),
    .ZN(_00049_)
  );
  AND2_X1 _16483_ (
    .A1(_08643_),
    .A2(_08758_),
    .ZN(_08842_)
  );
  AND2_X1 _16484_ (
    .A1(_08652_),
    .A2(_08842_),
    .ZN(_08843_)
  );
  INV_X1 _16485_ (
    .A(_08843_),
    .ZN(_08844_)
  );
  AND2_X1 _16486_ (
    .A1(_r[15]),
    .A2(_08844_),
    .ZN(_08845_)
  );
  INV_X1 _16487_ (
    .A(_08845_),
    .ZN(_08846_)
  );
  AND2_X1 _16488_ (
    .A1(_08763_),
    .A2(_08776_),
    .ZN(_08847_)
  );
  AND2_X1 _16489_ (
    .A1(_08200_),
    .A2(_08847_),
    .ZN(_08848_)
  );
  INV_X1 _16490_ (
    .A(_08848_),
    .ZN(_08849_)
  );
  AND2_X1 _16491_ (
    .A1(_08846_),
    .A2(_08849_),
    .ZN(_08850_)
  );
  INV_X1 _16492_ (
    .A(_08850_),
    .ZN(_08851_)
  );
  AND2_X1 _16493_ (
    .A1(_07954_),
    .A2(_08851_),
    .ZN(_00050_)
  );
  AND2_X1 _16494_ (
    .A1(_08645_),
    .A2(_08651_),
    .ZN(_08852_)
  );
  AND2_X1 _16495_ (
    .A1(_08642_),
    .A2(_08852_),
    .ZN(_08853_)
  );
  AND2_X1 _16496_ (
    .A1(_08769_),
    .A2(_08853_),
    .ZN(_08854_)
  );
  INV_X1 _16497_ (
    .A(_08854_),
    .ZN(_08855_)
  );
  AND2_X1 _16498_ (
    .A1(_r[16]),
    .A2(_08855_),
    .ZN(_08856_)
  );
  INV_X1 _16499_ (
    .A(_08856_),
    .ZN(_08857_)
  );
  AND2_X1 _16500_ (
    .A1(wb_reg_inst[11]),
    .A2(_08691_),
    .ZN(_08858_)
  );
  AND2_X1 _16501_ (
    .A1(_08775_),
    .A2(_08858_),
    .ZN(_08859_)
  );
  AND2_X1 _16502_ (
    .A1(_08199_),
    .A2(_08859_),
    .ZN(_08860_)
  );
  INV_X1 _16503_ (
    .A(_08860_),
    .ZN(_08861_)
  );
  AND2_X1 _16504_ (
    .A1(_08857_),
    .A2(_08861_),
    .ZN(_08862_)
  );
  INV_X1 _16505_ (
    .A(_08862_),
    .ZN(_08863_)
  );
  AND2_X1 _16506_ (
    .A1(_07954_),
    .A2(_08863_),
    .ZN(_00051_)
  );
  AND2_X1 _16507_ (
    .A1(_08641_),
    .A2(_08853_),
    .ZN(_08864_)
  );
  INV_X1 _16508_ (
    .A(_08864_),
    .ZN(_08865_)
  );
  AND2_X1 _16509_ (
    .A1(_r[17]),
    .A2(_08865_),
    .ZN(_08866_)
  );
  INV_X1 _16510_ (
    .A(_08866_),
    .ZN(_08867_)
  );
  AND2_X1 _16511_ (
    .A1(_08660_),
    .A2(_08858_),
    .ZN(_08868_)
  );
  INV_X1 _16512_ (
    .A(_08868_),
    .ZN(_08869_)
  );
  AND2_X1 _16513_ (
    .A1(_08867_),
    .A2(_08869_),
    .ZN(_08870_)
  );
  INV_X1 _16514_ (
    .A(_08870_),
    .ZN(_08871_)
  );
  AND2_X1 _16515_ (
    .A1(_07954_),
    .A2(_08871_),
    .ZN(_00052_)
  );
  AND2_X1 _16516_ (
    .A1(_08698_),
    .A2(_08853_),
    .ZN(_08872_)
  );
  INV_X1 _16517_ (
    .A(_08872_),
    .ZN(_08873_)
  );
  AND2_X1 _16518_ (
    .A1(_r[18]),
    .A2(_08873_),
    .ZN(_08874_)
  );
  INV_X1 _16519_ (
    .A(_08874_),
    .ZN(_08875_)
  );
  AND2_X1 _16520_ (
    .A1(_08705_),
    .A2(_08858_),
    .ZN(_08876_)
  );
  INV_X1 _16521_ (
    .A(_08876_),
    .ZN(_08877_)
  );
  AND2_X1 _16522_ (
    .A1(_08875_),
    .A2(_08877_),
    .ZN(_08878_)
  );
  INV_X1 _16523_ (
    .A(_08878_),
    .ZN(_08879_)
  );
  AND2_X1 _16524_ (
    .A1(_07954_),
    .A2(_08879_),
    .ZN(_00053_)
  );
  AND2_X1 _16525_ (
    .A1(_08711_),
    .A2(_08853_),
    .ZN(_08880_)
  );
  INV_X1 _16526_ (
    .A(_08880_),
    .ZN(_08881_)
  );
  AND2_X1 _16527_ (
    .A1(_r[19]),
    .A2(_08881_),
    .ZN(_08882_)
  );
  INV_X1 _16528_ (
    .A(_08882_),
    .ZN(_08883_)
  );
  AND2_X1 _16529_ (
    .A1(_08718_),
    .A2(_08858_),
    .ZN(_08884_)
  );
  INV_X1 _16530_ (
    .A(_08884_),
    .ZN(_08885_)
  );
  AND2_X1 _16531_ (
    .A1(_08883_),
    .A2(_08885_),
    .ZN(_08886_)
  );
  INV_X1 _16532_ (
    .A(_08886_),
    .ZN(_08887_)
  );
  AND2_X1 _16533_ (
    .A1(_07954_),
    .A2(_08887_),
    .ZN(_00054_)
  );
  AND2_X1 _16534_ (
    .A1(_08724_),
    .A2(_08853_),
    .ZN(_08888_)
  );
  INV_X1 _16535_ (
    .A(_08888_),
    .ZN(_08889_)
  );
  AND2_X1 _16536_ (
    .A1(_r[20]),
    .A2(_08889_),
    .ZN(_08890_)
  );
  INV_X1 _16537_ (
    .A(_08890_),
    .ZN(_08891_)
  );
  AND2_X1 _16538_ (
    .A1(_08731_),
    .A2(_08858_),
    .ZN(_08892_)
  );
  INV_X1 _16539_ (
    .A(_08892_),
    .ZN(_08893_)
  );
  AND2_X1 _16540_ (
    .A1(_08891_),
    .A2(_08893_),
    .ZN(_08894_)
  );
  INV_X1 _16541_ (
    .A(_08894_),
    .ZN(_08895_)
  );
  AND2_X1 _16542_ (
    .A1(_07954_),
    .A2(_08895_),
    .ZN(_00055_)
  );
  AND2_X1 _16543_ (
    .A1(_08736_),
    .A2(_08853_),
    .ZN(_08896_)
  );
  INV_X1 _16544_ (
    .A(_08896_),
    .ZN(_08897_)
  );
  AND2_X1 _16545_ (
    .A1(_r[21]),
    .A2(_08897_),
    .ZN(_08898_)
  );
  INV_X1 _16546_ (
    .A(_08898_),
    .ZN(_08899_)
  );
  AND2_X1 _16547_ (
    .A1(_08742_),
    .A2(_08858_),
    .ZN(_08900_)
  );
  INV_X1 _16548_ (
    .A(_08900_),
    .ZN(_08901_)
  );
  AND2_X1 _16549_ (
    .A1(_08899_),
    .A2(_08901_),
    .ZN(_08902_)
  );
  INV_X1 _16550_ (
    .A(_08902_),
    .ZN(_08903_)
  );
  AND2_X1 _16551_ (
    .A1(_07954_),
    .A2(_08903_),
    .ZN(_00056_)
  );
  AND2_X1 _16552_ (
    .A1(_08747_),
    .A2(_08853_),
    .ZN(_08904_)
  );
  INV_X1 _16553_ (
    .A(_08904_),
    .ZN(_08905_)
  );
  AND2_X1 _16554_ (
    .A1(_r[22]),
    .A2(_08905_),
    .ZN(_08906_)
  );
  INV_X1 _16555_ (
    .A(_08906_),
    .ZN(_08907_)
  );
  AND2_X1 _16556_ (
    .A1(_08753_),
    .A2(_08858_),
    .ZN(_08908_)
  );
  INV_X1 _16557_ (
    .A(_08908_),
    .ZN(_08909_)
  );
  AND2_X1 _16558_ (
    .A1(_08907_),
    .A2(_08909_),
    .ZN(_08910_)
  );
  INV_X1 _16559_ (
    .A(_08910_),
    .ZN(_08911_)
  );
  AND2_X1 _16560_ (
    .A1(_07954_),
    .A2(_08911_),
    .ZN(_00057_)
  );
  AND2_X1 _16561_ (
    .A1(_08758_),
    .A2(_08853_),
    .ZN(_08912_)
  );
  INV_X1 _16562_ (
    .A(_08912_),
    .ZN(_08913_)
  );
  AND2_X1 _16563_ (
    .A1(_r[23]),
    .A2(_08913_),
    .ZN(_08914_)
  );
  INV_X1 _16564_ (
    .A(_08914_),
    .ZN(_08915_)
  );
  AND2_X1 _16565_ (
    .A1(_08764_),
    .A2(_08858_),
    .ZN(_08916_)
  );
  INV_X1 _16566_ (
    .A(_08916_),
    .ZN(_08917_)
  );
  AND2_X1 _16567_ (
    .A1(_08915_),
    .A2(_08917_),
    .ZN(_08918_)
  );
  INV_X1 _16568_ (
    .A(_08918_),
    .ZN(_08919_)
  );
  AND2_X1 _16569_ (
    .A1(_07954_),
    .A2(_08919_),
    .ZN(_00058_)
  );
  AND2_X1 _16570_ (
    .A1(_08770_),
    .A2(_08852_),
    .ZN(_08920_)
  );
  INV_X1 _16571_ (
    .A(_08920_),
    .ZN(_08921_)
  );
  AND2_X1 _16572_ (
    .A1(_r[24]),
    .A2(_08921_),
    .ZN(_08922_)
  );
  INV_X1 _16573_ (
    .A(_08922_),
    .ZN(_08923_)
  );
  AND2_X1 _16574_ (
    .A1(wb_reg_inst[10]),
    .A2(_08859_),
    .ZN(_08924_)
  );
  INV_X1 _16575_ (
    .A(_08924_),
    .ZN(_08925_)
  );
  AND2_X1 _16576_ (
    .A1(_08923_),
    .A2(_08925_),
    .ZN(_08926_)
  );
  INV_X1 _16577_ (
    .A(_08926_),
    .ZN(_08927_)
  );
  AND2_X1 _16578_ (
    .A1(_07954_),
    .A2(_08927_),
    .ZN(_00059_)
  );
  AND2_X1 _16579_ (
    .A1(_08782_),
    .A2(_08852_),
    .ZN(_08928_)
  );
  INV_X1 _16580_ (
    .A(_08928_),
    .ZN(_08929_)
  );
  AND2_X1 _16581_ (
    .A1(_r[25]),
    .A2(_08929_),
    .ZN(_08930_)
  );
  INV_X1 _16582_ (
    .A(_08930_),
    .ZN(_08931_)
  );
  AND2_X1 _16583_ (
    .A1(wb_reg_inst[11]),
    .A2(_08787_),
    .ZN(_08932_)
  );
  INV_X1 _16584_ (
    .A(_08932_),
    .ZN(_08933_)
  );
  AND2_X1 _16585_ (
    .A1(_08931_),
    .A2(_08933_),
    .ZN(_08934_)
  );
  INV_X1 _16586_ (
    .A(_08934_),
    .ZN(_08935_)
  );
  AND2_X1 _16587_ (
    .A1(_07954_),
    .A2(_08935_),
    .ZN(_00060_)
  );
  AND2_X1 _16588_ (
    .A1(_08792_),
    .A2(_08852_),
    .ZN(_08936_)
  );
  INV_X1 _16589_ (
    .A(_08936_),
    .ZN(_08937_)
  );
  AND2_X1 _16590_ (
    .A1(_r[26]),
    .A2(_08937_),
    .ZN(_08938_)
  );
  INV_X1 _16591_ (
    .A(_08938_),
    .ZN(_08939_)
  );
  AND2_X1 _16592_ (
    .A1(wb_reg_inst[11]),
    .A2(_08797_),
    .ZN(_08940_)
  );
  INV_X1 _16593_ (
    .A(_08940_),
    .ZN(_08941_)
  );
  AND2_X1 _16594_ (
    .A1(_08939_),
    .A2(_08941_),
    .ZN(_08942_)
  );
  INV_X1 _16595_ (
    .A(_08942_),
    .ZN(_08943_)
  );
  AND2_X1 _16596_ (
    .A1(_07954_),
    .A2(_08943_),
    .ZN(_00061_)
  );
  AND2_X1 _16597_ (
    .A1(_08802_),
    .A2(_08852_),
    .ZN(_08944_)
  );
  INV_X1 _16598_ (
    .A(_08944_),
    .ZN(_08945_)
  );
  AND2_X1 _16599_ (
    .A1(_r[27]),
    .A2(_08945_),
    .ZN(_08946_)
  );
  INV_X1 _16600_ (
    .A(_08946_),
    .ZN(_08947_)
  );
  AND2_X1 _16601_ (
    .A1(wb_reg_inst[11]),
    .A2(_08807_),
    .ZN(_08948_)
  );
  INV_X1 _16602_ (
    .A(_08948_),
    .ZN(_08949_)
  );
  AND2_X1 _16603_ (
    .A1(_08947_),
    .A2(_08949_),
    .ZN(_08950_)
  );
  INV_X1 _16604_ (
    .A(_08950_),
    .ZN(_08951_)
  );
  AND2_X1 _16605_ (
    .A1(_07954_),
    .A2(_08951_),
    .ZN(_00062_)
  );
  AND2_X1 _16606_ (
    .A1(_08812_),
    .A2(_08852_),
    .ZN(_08952_)
  );
  INV_X1 _16607_ (
    .A(_08952_),
    .ZN(_08953_)
  );
  AND2_X1 _16608_ (
    .A1(_r[28]),
    .A2(_08953_),
    .ZN(_08954_)
  );
  INV_X1 _16609_ (
    .A(_08954_),
    .ZN(_08955_)
  );
  AND2_X1 _16610_ (
    .A1(wb_reg_inst[11]),
    .A2(_08817_),
    .ZN(_08956_)
  );
  INV_X1 _16611_ (
    .A(_08956_),
    .ZN(_08957_)
  );
  AND2_X1 _16612_ (
    .A1(_08955_),
    .A2(_08957_),
    .ZN(_08958_)
  );
  INV_X1 _16613_ (
    .A(_08958_),
    .ZN(_08959_)
  );
  AND2_X1 _16614_ (
    .A1(_07954_),
    .A2(_08959_),
    .ZN(_00063_)
  );
  AND2_X1 _16615_ (
    .A1(_08822_),
    .A2(_08852_),
    .ZN(_08960_)
  );
  INV_X1 _16616_ (
    .A(_08960_),
    .ZN(_08961_)
  );
  AND2_X1 _16617_ (
    .A1(_r[29]),
    .A2(_08961_),
    .ZN(_08962_)
  );
  INV_X1 _16618_ (
    .A(_08962_),
    .ZN(_08963_)
  );
  AND2_X1 _16619_ (
    .A1(wb_reg_inst[11]),
    .A2(_08827_),
    .ZN(_08964_)
  );
  INV_X1 _16620_ (
    .A(_08964_),
    .ZN(_08965_)
  );
  AND2_X1 _16621_ (
    .A1(_08963_),
    .A2(_08965_),
    .ZN(_08966_)
  );
  INV_X1 _16622_ (
    .A(_08966_),
    .ZN(_08967_)
  );
  AND2_X1 _16623_ (
    .A1(_07954_),
    .A2(_08967_),
    .ZN(_00064_)
  );
  AND2_X1 _16624_ (
    .A1(_08832_),
    .A2(_08852_),
    .ZN(_08968_)
  );
  INV_X1 _16625_ (
    .A(_08968_),
    .ZN(_08969_)
  );
  AND2_X1 _16626_ (
    .A1(_r[30]),
    .A2(_08969_),
    .ZN(_08970_)
  );
  INV_X1 _16627_ (
    .A(_08970_),
    .ZN(_08971_)
  );
  AND2_X1 _16628_ (
    .A1(wb_reg_inst[11]),
    .A2(_08837_),
    .ZN(_08972_)
  );
  INV_X1 _16629_ (
    .A(_08972_),
    .ZN(_08973_)
  );
  AND2_X1 _16630_ (
    .A1(_08971_),
    .A2(_08973_),
    .ZN(_08974_)
  );
  INV_X1 _16631_ (
    .A(_08974_),
    .ZN(_08975_)
  );
  AND2_X1 _16632_ (
    .A1(_07954_),
    .A2(_08975_),
    .ZN(_00065_)
  );
  AND2_X1 _16633_ (
    .A1(_08842_),
    .A2(_08852_),
    .ZN(_08976_)
  );
  INV_X1 _16634_ (
    .A(_08976_),
    .ZN(_08977_)
  );
  AND2_X1 _16635_ (
    .A1(_r[31]),
    .A2(_08977_),
    .ZN(_08978_)
  );
  INV_X1 _16636_ (
    .A(_08978_),
    .ZN(_08979_)
  );
  AND2_X1 _16637_ (
    .A1(wb_reg_inst[11]),
    .A2(_08847_),
    .ZN(_08980_)
  );
  INV_X1 _16638_ (
    .A(_08980_),
    .ZN(_08981_)
  );
  AND2_X1 _16639_ (
    .A1(_08979_),
    .A2(_08981_),
    .ZN(_08982_)
  );
  INV_X1 _16640_ (
    .A(_08982_),
    .ZN(_08983_)
  );
  AND2_X1 _16641_ (
    .A1(_07954_),
    .A2(_08983_),
    .ZN(_00066_)
  );
  AND2_X1 _16642_ (
    .A1(csr_io_decode_0_inst[1]),
    .A2(_08530_),
    .ZN(_08984_)
  );
  AND2_X1 _16643_ (
    .A1(_08533_),
    .A2(_08984_),
    .ZN(_08985_)
  );
  AND2_X1 _16644_ (
    .A1(csr_io_decode_0_inst[0]),
    .A2(csr_io_decode_0_inst[1]),
    .ZN(_08986_)
  );
  AND2_X1 _16645_ (
    .A1(csr_io_decode_0_inst[0]),
    .A2(_08985_),
    .ZN(_08987_)
  );
  AND2_X1 _16646_ (
    .A1(_08529_),
    .A2(_08987_),
    .ZN(_08988_)
  );
  AND2_X1 _16647_ (
    .A1(_08531_),
    .A2(_08988_),
    .ZN(_08989_)
  );
  AND2_X1 _16648_ (
    .A1(_08133_),
    .A2(_08134_),
    .ZN(_08990_)
  );
  INV_X1 _16649_ (
    .A(_08990_),
    .ZN(_08991_)
  );
  AND2_X1 _16650_ (
    .A1(_08989_),
    .A2(_08990_),
    .ZN(_08992_)
  );
  INV_X1 _16651_ (
    .A(_08992_),
    .ZN(_08993_)
  );
  AND2_X1 _16652_ (
    .A1(_08134_),
    .A2(_08532_),
    .ZN(_08994_)
  );
  INV_X1 _16653_ (
    .A(_08994_),
    .ZN(_08995_)
  );
  AND2_X1 _16654_ (
    .A1(_08134_),
    .A2(_08135_),
    .ZN(_08996_)
  );
  INV_X1 _16655_ (
    .A(_08996_),
    .ZN(_08997_)
  );
  AND2_X1 _16656_ (
    .A1(_08532_),
    .A2(_08996_),
    .ZN(_08998_)
  );
  INV_X1 _16657_ (
    .A(_08998_),
    .ZN(_08999_)
  );
  AND2_X1 _16658_ (
    .A1(_08133_),
    .A2(_08135_),
    .ZN(_09000_)
  );
  INV_X1 _16659_ (
    .A(_09000_),
    .ZN(_09001_)
  );
  AND2_X1 _16660_ (
    .A1(_08532_),
    .A2(_09000_),
    .ZN(_09002_)
  );
  INV_X1 _16661_ (
    .A(_09002_),
    .ZN(_09003_)
  );
  AND2_X1 _16662_ (
    .A1(_08531_),
    .A2(_08994_),
    .ZN(_09004_)
  );
  INV_X1 _16663_ (
    .A(_09004_),
    .ZN(_09005_)
  );
  AND2_X1 _16664_ (
    .A1(_09003_),
    .A2(_09005_),
    .ZN(_09006_)
  );
  AND2_X1 _16665_ (
    .A1(_08999_),
    .A2(_09006_),
    .ZN(_09007_)
  );
  INV_X1 _16666_ (
    .A(_09007_),
    .ZN(_09008_)
  );
  AND2_X1 _16667_ (
    .A1(_08988_),
    .A2(_09008_),
    .ZN(_09009_)
  );
  INV_X1 _16668_ (
    .A(_09009_),
    .ZN(_09010_)
  );
  AND2_X1 _16669_ (
    .A1(_08993_),
    .A2(_09010_),
    .ZN(_09011_)
  );
  AND2_X1 _16670_ (
    .A1(_08533_),
    .A2(_08986_),
    .ZN(_09012_)
  );
  AND2_X1 _16671_ (
    .A1(csr_io_decode_0_inst[6]),
    .A2(csr_io_decode_0_inst[5]),
    .ZN(_09013_)
  );
  AND2_X1 _16672_ (
    .A1(_08994_),
    .A2(_09013_),
    .ZN(_09014_)
  );
  AND2_X1 _16673_ (
    .A1(_09000_),
    .A2(_09014_),
    .ZN(_09015_)
  );
  AND2_X1 _16674_ (
    .A1(_09012_),
    .A2(_09015_),
    .ZN(_09016_)
  );
  INV_X1 _16675_ (
    .A(_09016_),
    .ZN(_09017_)
  );
  AND2_X1 _16676_ (
    .A1(csr_io_decode_0_inst[0]),
    .A2(csr_io_decode_0_inst[4]),
    .ZN(_09018_)
  );
  AND2_X1 _16677_ (
    .A1(_08985_),
    .A2(_09018_),
    .ZN(_09019_)
  );
  AND2_X1 _16678_ (
    .A1(csr_io_decode_0_inst[12]),
    .A2(_08529_),
    .ZN(_09020_)
  );
  AND2_X1 _16679_ (
    .A1(_09019_),
    .A2(_09020_),
    .ZN(_09021_)
  );
  AND2_X1 _16680_ (
    .A1(_08146_),
    .A2(_08147_),
    .ZN(_09022_)
  );
  AND2_X1 _16681_ (
    .A1(_08147_),
    .A2(_08148_),
    .ZN(_09023_)
  );
  AND2_X1 _16682_ (
    .A1(_08134_),
    .A2(_08146_),
    .ZN(_09024_)
  );
  AND2_X1 _16683_ (
    .A1(_09023_),
    .A2(_09024_),
    .ZN(_09025_)
  );
  AND2_X1 _16684_ (
    .A1(_08151_),
    .A2(_08152_),
    .ZN(_09026_)
  );
  AND2_X1 _16685_ (
    .A1(_08150_),
    .A2(_08152_),
    .ZN(_09027_)
  );
  AND2_X1 _16686_ (
    .A1(_08150_),
    .A2(_09026_),
    .ZN(_09028_)
  );
  AND2_X1 _16687_ (
    .A1(_08149_),
    .A2(_09027_),
    .ZN(_09029_)
  );
  AND2_X1 _16688_ (
    .A1(_08151_),
    .A2(_09029_),
    .ZN(_09030_)
  );
  AND2_X1 _16689_ (
    .A1(_09025_),
    .A2(_09030_),
    .ZN(_09031_)
  );
  AND2_X1 _16690_ (
    .A1(_09021_),
    .A2(_09031_),
    .ZN(_09032_)
  );
  INV_X1 _16691_ (
    .A(_09032_),
    .ZN(_09033_)
  );
  AND2_X1 _16692_ (
    .A1(_09017_),
    .A2(_09033_),
    .ZN(_09034_)
  );
  AND2_X1 _16693_ (
    .A1(_09011_),
    .A2(_09034_),
    .ZN(_09035_)
  );
  AND2_X1 _16694_ (
    .A1(_08532_),
    .A2(_08987_),
    .ZN(_09036_)
  );
  AND2_X1 _16695_ (
    .A1(_09013_),
    .A2(_09036_),
    .ZN(_09037_)
  );
  AND2_X1 _16696_ (
    .A1(csr_io_decode_0_inst[14]),
    .A2(_09013_),
    .ZN(_09038_)
  );
  AND2_X1 _16697_ (
    .A1(_09036_),
    .A2(_09038_),
    .ZN(_09039_)
  );
  INV_X1 _16698_ (
    .A(_09039_),
    .ZN(_09040_)
  );
  AND2_X1 _16699_ (
    .A1(csr_io_decode_0_inst[14]),
    .A2(_09025_),
    .ZN(_09041_)
  );
  AND2_X1 _16700_ (
    .A1(_09021_),
    .A2(_09041_),
    .ZN(_09042_)
  );
  INV_X1 _16701_ (
    .A(_09042_),
    .ZN(_09043_)
  );
  AND2_X1 _16702_ (
    .A1(_09029_),
    .A2(_09042_),
    .ZN(_09044_)
  );
  INV_X1 _16703_ (
    .A(_09044_),
    .ZN(_09045_)
  );
  AND2_X1 _16704_ (
    .A1(_09040_),
    .A2(_09045_),
    .ZN(_09046_)
  );
  AND2_X1 _16705_ (
    .A1(csr_io_decode_0_inst[13]),
    .A2(_08529_),
    .ZN(_09047_)
  );
  AND2_X1 _16706_ (
    .A1(_08531_),
    .A2(_09019_),
    .ZN(_09048_)
  );
  AND2_X1 _16707_ (
    .A1(_09047_),
    .A2(_09048_),
    .ZN(_09049_)
  );
  INV_X1 _16708_ (
    .A(_09049_),
    .ZN(_09050_)
  );
  AND2_X1 _16709_ (
    .A1(_08148_),
    .A2(_08149_),
    .ZN(_09051_)
  );
  AND2_X1 _16710_ (
    .A1(csr_io_decode_0_inst[5]),
    .A2(_09002_),
    .ZN(_09052_)
  );
  AND2_X1 _16711_ (
    .A1(csr_io_decode_0_inst[2]),
    .A2(csr_io_decode_0_inst[3]),
    .ZN(_09053_)
  );
  AND2_X1 _16712_ (
    .A1(_08986_),
    .A2(_09053_),
    .ZN(_09054_)
  );
  AND2_X1 _16713_ (
    .A1(_09047_),
    .A2(_09054_),
    .ZN(_09055_)
  );
  AND2_X1 _16714_ (
    .A1(_09052_),
    .A2(_09055_),
    .ZN(_09056_)
  );
  AND2_X1 _16715_ (
    .A1(_09051_),
    .A2(_09056_),
    .ZN(_09057_)
  );
  INV_X1 _16716_ (
    .A(_09057_),
    .ZN(_09058_)
  );
  AND2_X1 _16717_ (
    .A1(_09050_),
    .A2(_09058_),
    .ZN(_09059_)
  );
  AND2_X1 _16718_ (
    .A1(csr_io_decode_0_inst[13]),
    .A2(_08135_),
    .ZN(_09060_)
  );
  INV_X1 _16719_ (
    .A(_09060_),
    .ZN(_09061_)
  );
  AND2_X1 _16720_ (
    .A1(csr_io_decode_0_inst[5]),
    .A2(csr_io_decode_0_inst[4]),
    .ZN(_09062_)
  );
  AND2_X1 _16721_ (
    .A1(_09013_),
    .A2(_09018_),
    .ZN(_09063_)
  );
  AND2_X1 _16722_ (
    .A1(_08985_),
    .A2(_09063_),
    .ZN(_09064_)
  );
  AND2_X1 _16723_ (
    .A1(_09060_),
    .A2(_09064_),
    .ZN(_09065_)
  );
  INV_X1 _16724_ (
    .A(_09065_),
    .ZN(_09066_)
  );
  AND2_X1 _16725_ (
    .A1(csr_io_decode_0_inst[12]),
    .A2(_09013_),
    .ZN(_09067_)
  );
  AND2_X1 _16726_ (
    .A1(_08987_),
    .A2(_08996_),
    .ZN(_09068_)
  );
  AND2_X1 _16727_ (
    .A1(_09067_),
    .A2(_09068_),
    .ZN(_09069_)
  );
  INV_X1 _16728_ (
    .A(_09069_),
    .ZN(_09070_)
  );
  AND2_X1 _16729_ (
    .A1(_09066_),
    .A2(_09070_),
    .ZN(_09071_)
  );
  AND2_X1 _16730_ (
    .A1(_09059_),
    .A2(_09071_),
    .ZN(_09072_)
  );
  AND2_X1 _16731_ (
    .A1(csr_io_decode_0_inst[5]),
    .A2(_08532_),
    .ZN(_09073_)
  );
  AND2_X1 _16732_ (
    .A1(_09054_),
    .A2(_09073_),
    .ZN(_09074_)
  );
  AND2_X1 _16733_ (
    .A1(_08133_),
    .A2(_08529_),
    .ZN(_09075_)
  );
  AND2_X1 _16734_ (
    .A1(_09046_),
    .A2(_09072_),
    .ZN(_09076_)
  );
  AND2_X1 _16735_ (
    .A1(_08529_),
    .A2(_08531_),
    .ZN(_09077_)
  );
  AND2_X1 _16736_ (
    .A1(_09035_),
    .A2(_09076_),
    .ZN(_09078_)
  );
  AND2_X1 _16737_ (
    .A1(csr_io_decode_0_inst[28]),
    .A2(_09028_),
    .ZN(_09079_)
  );
  AND2_X1 _16738_ (
    .A1(_08145_),
    .A2(_08148_),
    .ZN(_09080_)
  );
  AND2_X1 _16739_ (
    .A1(_08142_),
    .A2(_08144_),
    .ZN(_09081_)
  );
  AND2_X1 _16740_ (
    .A1(_08141_),
    .A2(_08143_),
    .ZN(_09082_)
  );
  AND2_X1 _16741_ (
    .A1(_09081_),
    .A2(_09082_),
    .ZN(_09083_)
  );
  AND2_X1 _16742_ (
    .A1(_09080_),
    .A2(_09083_),
    .ZN(_09084_)
  );
  AND2_X1 _16743_ (
    .A1(_09079_),
    .A2(_09084_),
    .ZN(_09085_)
  );
  AND2_X1 _16744_ (
    .A1(_08529_),
    .A2(_09074_),
    .ZN(_09086_)
  );
  AND2_X1 _16745_ (
    .A1(_09085_),
    .A2(_09086_),
    .ZN(_09087_)
  );
  INV_X1 _16746_ (
    .A(_09087_),
    .ZN(_09088_)
  );
  AND2_X1 _16747_ (
    .A1(csr_io_decode_0_inst[27]),
    .A2(_09056_),
    .ZN(_09089_)
  );
  AND2_X1 _16748_ (
    .A1(_09028_),
    .A2(_09089_),
    .ZN(_09090_)
  );
  INV_X1 _16749_ (
    .A(_09090_),
    .ZN(_09091_)
  );
  AND2_X1 _16750_ (
    .A1(_09088_),
    .A2(_09091_),
    .ZN(_09092_)
  );
  AND2_X1 _16751_ (
    .A1(_09023_),
    .A2(_09030_),
    .ZN(_09093_)
  );
  AND2_X1 _16752_ (
    .A1(csr_io_decode_0_inst[5]),
    .A2(_09019_),
    .ZN(_09094_)
  );
  AND2_X1 _16753_ (
    .A1(_08529_),
    .A2(_09094_),
    .ZN(_09095_)
  );
  AND2_X1 _16754_ (
    .A1(_09093_),
    .A2(_09095_),
    .ZN(_09096_)
  );
  INV_X1 _16755_ (
    .A(_09096_),
    .ZN(_09097_)
  );
  AND2_X1 _16756_ (
    .A1(_08148_),
    .A2(_09075_),
    .ZN(_09098_)
  );
  AND2_X1 _16757_ (
    .A1(_08996_),
    .A2(_09022_),
    .ZN(_09099_)
  );
  AND2_X1 _16758_ (
    .A1(_09098_),
    .A2(_09099_),
    .ZN(_09100_)
  );
  AND2_X1 _16759_ (
    .A1(_09029_),
    .A2(_09100_),
    .ZN(_09101_)
  );
  AND2_X1 _16760_ (
    .A1(_09094_),
    .A2(_09101_),
    .ZN(_09102_)
  );
  INV_X1 _16761_ (
    .A(_09102_),
    .ZN(_09103_)
  );
  AND2_X1 _16762_ (
    .A1(_09097_),
    .A2(_09103_),
    .ZN(_09104_)
  );
  AND2_X1 _16763_ (
    .A1(_09092_),
    .A2(_09104_),
    .ZN(_09105_)
  );
  AND2_X1 _16764_ (
    .A1(_09035_),
    .A2(_09046_),
    .ZN(_09106_)
  );
  AND2_X1 _16765_ (
    .A1(_08532_),
    .A2(_09054_),
    .ZN(_09107_)
  );
  AND2_X1 _16766_ (
    .A1(_09078_),
    .A2(_09105_),
    .ZN(_09108_)
  );
  INV_X1 _16767_ (
    .A(_09108_),
    .ZN(_09109_)
  );
  AND2_X1 _16768_ (
    .A1(_08540_),
    .A2(_08543_),
    .ZN(_09110_)
  );
  AND2_X1 _16769_ (
    .A1(_08541_),
    .A2(_08542_),
    .ZN(_09111_)
  );
  AND2_X1 _16770_ (
    .A1(_08571_),
    .A2(_09111_),
    .ZN(_09112_)
  );
  AND2_X1 _16771_ (
    .A1(_09110_),
    .A2(_09112_),
    .ZN(_09113_)
  );
  INV_X1 _16772_ (
    .A(_09113_),
    .ZN(_09114_)
  );
  AND2_X1 _16773_ (
    .A1(ex_ctrl_wxd),
    .A2(ex_reg_valid),
    .ZN(_09115_)
  );
  AND2_X1 _16774_ (
    .A1(ex_reg_inst[7]),
    .A2(_08540_),
    .ZN(_09116_)
  );
  INV_X1 _16775_ (
    .A(_09116_),
    .ZN(_09117_)
  );
  AND2_X1 _16776_ (
    .A1(ex_reg_inst[8]),
    .A2(_08541_),
    .ZN(_09118_)
  );
  INV_X1 _16777_ (
    .A(_09118_),
    .ZN(_09119_)
  );
  AND2_X1 _16778_ (
    .A1(_08087_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_09120_)
  );
  INV_X1 _16779_ (
    .A(_09120_),
    .ZN(_09121_)
  );
  AND2_X1 _16780_ (
    .A1(_08085_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[0]),
    .ZN(_09122_)
  );
  INV_X1 _16781_ (
    .A(_09122_),
    .ZN(_09123_)
  );
  AND2_X1 _16782_ (
    .A1(ex_reg_inst[9]),
    .A2(_08542_),
    .ZN(_09124_)
  );
  INV_X1 _16783_ (
    .A(_09124_),
    .ZN(_09125_)
  );
  AND2_X1 _16784_ (
    .A1(_08089_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_09126_)
  );
  INV_X1 _16785_ (
    .A(_09126_),
    .ZN(_09127_)
  );
  AND2_X1 _16786_ (
    .A1(_09125_),
    .A2(_09127_),
    .ZN(_09128_)
  );
  AND2_X1 _16787_ (
    .A1(ex_reg_inst[11]),
    .A2(_08571_),
    .ZN(_09129_)
  );
  INV_X1 _16788_ (
    .A(_09129_),
    .ZN(_09130_)
  );
  AND2_X1 _16789_ (
    .A1(_08093_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[4]),
    .ZN(_09131_)
  );
  INV_X1 _16790_ (
    .A(_09131_),
    .ZN(_09132_)
  );
  AND2_X1 _16791_ (
    .A1(ex_reg_inst[10]),
    .A2(_08543_),
    .ZN(_09133_)
  );
  INV_X1 _16792_ (
    .A(_09133_),
    .ZN(_09134_)
  );
  AND2_X1 _16793_ (
    .A1(_08091_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[3]),
    .ZN(_09135_)
  );
  INV_X1 _16794_ (
    .A(_09135_),
    .ZN(_09136_)
  );
  AND2_X1 _16795_ (
    .A1(_09130_),
    .A2(_09134_),
    .ZN(_09137_)
  );
  AND2_X1 _16796_ (
    .A1(_09128_),
    .A2(_09132_),
    .ZN(_09138_)
  );
  AND2_X1 _16797_ (
    .A1(_09137_),
    .A2(_09138_),
    .ZN(_09139_)
  );
  AND2_X1 _16798_ (
    .A1(_09117_),
    .A2(_09136_),
    .ZN(_09140_)
  );
  AND2_X1 _16799_ (
    .A1(_09119_),
    .A2(_09123_),
    .ZN(_09141_)
  );
  AND2_X1 _16800_ (
    .A1(_09121_),
    .A2(_09141_),
    .ZN(_09142_)
  );
  AND2_X1 _16801_ (
    .A1(_09140_),
    .A2(_09142_),
    .ZN(_09143_)
  );
  AND2_X1 _16802_ (
    .A1(_09139_),
    .A2(_09143_),
    .ZN(_09144_)
  );
  AND2_X1 _16803_ (
    .A1(_09115_),
    .A2(_09144_),
    .ZN(_09145_)
  );
  INV_X1 _16804_ (
    .A(_09145_),
    .ZN(_09146_)
  );
  AND2_X1 _16805_ (
    .A1(_09114_),
    .A2(_09146_),
    .ZN(_09147_)
  );
  AND2_X1 _16806_ (
    .A1(mem_ctrl_wxd),
    .A2(mem_reg_valid),
    .ZN(_09148_)
  );
  AND2_X1 _16807_ (
    .A1(mem_reg_inst[7]),
    .A2(_08540_),
    .ZN(_09149_)
  );
  INV_X1 _16808_ (
    .A(_09149_),
    .ZN(_09150_)
  );
  AND2_X1 _16809_ (
    .A1(mem_reg_inst[8]),
    .A2(_08541_),
    .ZN(_09151_)
  );
  INV_X1 _16810_ (
    .A(_09151_),
    .ZN(_09152_)
  );
  AND2_X1 _16811_ (
    .A1(_08086_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_09153_)
  );
  INV_X1 _16812_ (
    .A(_09153_),
    .ZN(_09154_)
  );
  AND2_X1 _16813_ (
    .A1(_08084_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[0]),
    .ZN(_09155_)
  );
  INV_X1 _16814_ (
    .A(_09155_),
    .ZN(_09156_)
  );
  AND2_X1 _16815_ (
    .A1(mem_reg_inst[9]),
    .A2(_08542_),
    .ZN(_09157_)
  );
  INV_X1 _16816_ (
    .A(_09157_),
    .ZN(_09158_)
  );
  AND2_X1 _16817_ (
    .A1(_08088_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_09159_)
  );
  INV_X1 _16818_ (
    .A(_09159_),
    .ZN(_09160_)
  );
  AND2_X1 _16819_ (
    .A1(_09158_),
    .A2(_09160_),
    .ZN(_09161_)
  );
  AND2_X1 _16820_ (
    .A1(mem_reg_inst[11]),
    .A2(_08571_),
    .ZN(_09162_)
  );
  INV_X1 _16821_ (
    .A(_09162_),
    .ZN(_09163_)
  );
  AND2_X1 _16822_ (
    .A1(_08092_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[4]),
    .ZN(_09164_)
  );
  INV_X1 _16823_ (
    .A(_09164_),
    .ZN(_09165_)
  );
  AND2_X1 _16824_ (
    .A1(mem_reg_inst[10]),
    .A2(_08543_),
    .ZN(_09166_)
  );
  INV_X1 _16825_ (
    .A(_09166_),
    .ZN(_09167_)
  );
  AND2_X1 _16826_ (
    .A1(_08090_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[3]),
    .ZN(_09168_)
  );
  INV_X1 _16827_ (
    .A(_09168_),
    .ZN(_09169_)
  );
  AND2_X1 _16828_ (
    .A1(_09163_),
    .A2(_09167_),
    .ZN(_09170_)
  );
  AND2_X1 _16829_ (
    .A1(_09161_),
    .A2(_09165_),
    .ZN(_09171_)
  );
  AND2_X1 _16830_ (
    .A1(_09170_),
    .A2(_09171_),
    .ZN(_09172_)
  );
  AND2_X1 _16831_ (
    .A1(_09150_),
    .A2(_09169_),
    .ZN(_09173_)
  );
  AND2_X1 _16832_ (
    .A1(_09152_),
    .A2(_09156_),
    .ZN(_09174_)
  );
  AND2_X1 _16833_ (
    .A1(_09154_),
    .A2(_09174_),
    .ZN(_09175_)
  );
  AND2_X1 _16834_ (
    .A1(_09173_),
    .A2(_09175_),
    .ZN(_09176_)
  );
  AND2_X1 _16835_ (
    .A1(_09172_),
    .A2(_09176_),
    .ZN(_09177_)
  );
  AND2_X1 _16836_ (
    .A1(_09148_),
    .A2(_09177_),
    .ZN(_09178_)
  );
  INV_X1 _16837_ (
    .A(_09178_),
    .ZN(_09179_)
  );
  AND2_X1 _16838_ (
    .A1(_09147_),
    .A2(_09179_),
    .ZN(_09180_)
  );
  INV_X1 _16839_ (
    .A(_09180_),
    .ZN(_09181_)
  );
  AND2_X1 _16840_ (
    .A1(_09109_),
    .A2(_09180_),
    .ZN(_09182_)
  );
  INV_X1 _16841_ (
    .A(_09182_),
    .ZN(_09183_)
  );
  AND2_X1 _16842_ (
    .A1(_08529_),
    .A2(csr_io_decode_0_inst[4]),
    .ZN(_09184_)
  );
  AND2_X1 _16843_ (
    .A1(csr_io_decode_0_inst[2]),
    .A2(_09184_),
    .ZN(_09185_)
  );
  AND2_X1 _16844_ (
    .A1(_09012_),
    .A2(_09185_),
    .ZN(_09186_)
  );
  INV_X1 _16845_ (
    .A(_09186_),
    .ZN(_09187_)
  );
  AND2_X1 _16846_ (
    .A1(_09104_),
    .A2(_09187_),
    .ZN(_09188_)
  );
  AND2_X1 _16847_ (
    .A1(_09022_),
    .A2(_09080_),
    .ZN(_09189_)
  );
  AND2_X1 _16848_ (
    .A1(_09026_),
    .A2(_09081_),
    .ZN(_09190_)
  );
  AND2_X1 _16849_ (
    .A1(_09063_),
    .A2(_09190_),
    .ZN(_09191_)
  );
  AND2_X1 _16850_ (
    .A1(_09189_),
    .A2(_09191_),
    .ZN(_09192_)
  );
  AND2_X1 _16851_ (
    .A1(_08137_),
    .A2(_08138_),
    .ZN(_09193_)
  );
  AND2_X1 _16852_ (
    .A1(_08136_),
    .A2(_08139_),
    .ZN(_09194_)
  );
  AND2_X1 _16853_ (
    .A1(_09193_),
    .A2(_09194_),
    .ZN(_09195_)
  );
  AND2_X1 _16854_ (
    .A1(_08131_),
    .A2(_08135_),
    .ZN(_09196_)
  );
  AND2_X1 _16855_ (
    .A1(_08130_),
    .A2(_09196_),
    .ZN(_09197_)
  );
  AND2_X1 _16856_ (
    .A1(_09195_),
    .A2(_09197_),
    .ZN(_09198_)
  );
  AND2_X1 _16857_ (
    .A1(_08128_),
    .A2(_08129_),
    .ZN(_09199_)
  );
  AND2_X1 _16858_ (
    .A1(_08132_),
    .A2(_08140_),
    .ZN(_09200_)
  );
  AND2_X1 _16859_ (
    .A1(_09199_),
    .A2(_09200_),
    .ZN(_09201_)
  );
  AND2_X1 _16860_ (
    .A1(_08990_),
    .A2(_09201_),
    .ZN(_09202_)
  );
  AND2_X1 _16861_ (
    .A1(_09198_),
    .A2(_09202_),
    .ZN(_09203_)
  );
  AND2_X1 _16862_ (
    .A1(_08143_),
    .A2(_08149_),
    .ZN(_09204_)
  );
  AND2_X1 _16863_ (
    .A1(_08150_),
    .A2(_09204_),
    .ZN(_09205_)
  );
  INV_X1 _16864_ (
    .A(_09205_),
    .ZN(_09206_)
  );
  AND2_X1 _16865_ (
    .A1(csr_io_decode_0_inst[20]),
    .A2(csr_io_decode_0_inst[22]),
    .ZN(_09207_)
  );
  AND2_X1 _16866_ (
    .A1(csr_io_decode_0_inst[28]),
    .A2(_09207_),
    .ZN(_09208_)
  );
  INV_X1 _16867_ (
    .A(_09208_),
    .ZN(_09209_)
  );
  AND2_X1 _16868_ (
    .A1(_09206_),
    .A2(_09209_),
    .ZN(_09210_)
  );
  INV_X1 _16869_ (
    .A(_09210_),
    .ZN(_09211_)
  );
  AND2_X1 _16870_ (
    .A1(_09203_),
    .A2(_09211_),
    .ZN(_09212_)
  );
  AND2_X1 _16871_ (
    .A1(_09192_),
    .A2(_09212_),
    .ZN(_09213_)
  );
  INV_X1 _16872_ (
    .A(_09213_),
    .ZN(_09214_)
  );
  AND2_X1 _16873_ (
    .A1(_08985_),
    .A2(_09213_),
    .ZN(_09215_)
  );
  INV_X1 _16874_ (
    .A(_09215_),
    .ZN(_09216_)
  );
  AND2_X1 _16875_ (
    .A1(_09188_),
    .A2(_09216_),
    .ZN(_09217_)
  );
  AND2_X1 _16876_ (
    .A1(_09106_),
    .A2(_09217_),
    .ZN(_09218_)
  );
  AND2_X1 _16877_ (
    .A1(_08134_),
    .A2(_09067_),
    .ZN(_09219_)
  );
  INV_X1 _16878_ (
    .A(_09219_),
    .ZN(_09220_)
  );
  AND2_X1 _16879_ (
    .A1(csr_io_decode_0_inst[28]),
    .A2(csr_io_decode_0_inst[29]),
    .ZN(_09221_)
  );
  AND2_X1 _16880_ (
    .A1(_08152_),
    .A2(csr_io_decode_0_inst[6]),
    .ZN(_09222_)
  );
  AND2_X1 _16881_ (
    .A1(_09221_),
    .A2(_09222_),
    .ZN(_09223_)
  );
  AND2_X1 _16882_ (
    .A1(csr_io_decode_0_inst[21]),
    .A2(_08144_),
    .ZN(_09224_)
  );
  AND2_X1 _16883_ (
    .A1(_09082_),
    .A2(_09224_),
    .ZN(_09225_)
  );
  AND2_X1 _16884_ (
    .A1(_09062_),
    .A2(_09225_),
    .ZN(_09226_)
  );
  AND2_X1 _16885_ (
    .A1(_09223_),
    .A2(_09226_),
    .ZN(_09227_)
  );
  AND2_X1 _16886_ (
    .A1(csr_io_decode_0_inst[25]),
    .A2(csr_io_decode_0_inst[27]),
    .ZN(_09228_)
  );
  AND2_X1 _16887_ (
    .A1(csr_io_decode_0_inst[24]),
    .A2(_09228_),
    .ZN(_09229_)
  );
  AND2_X1 _16888_ (
    .A1(_08147_),
    .A2(_09229_),
    .ZN(_09230_)
  );
  MUX2_X1 _16889_ (
    .A(_09189_),
    .B(_09230_),
    .S(csr_io_decode_0_inst[30]),
    .Z(_09231_)
  );
  AND2_X1 _16890_ (
    .A1(_09203_),
    .A2(_09231_),
    .ZN(_09232_)
  );
  AND2_X1 _16891_ (
    .A1(_09227_),
    .A2(_09232_),
    .ZN(_09233_)
  );
  INV_X1 _16892_ (
    .A(_09233_),
    .ZN(_09234_)
  );
  AND2_X1 _16893_ (
    .A1(_09220_),
    .A2(_09234_),
    .ZN(_09235_)
  );
  INV_X1 _16894_ (
    .A(_09235_),
    .ZN(_09236_)
  );
  AND2_X1 _16895_ (
    .A1(_08987_),
    .A2(_09236_),
    .ZN(_09237_)
  );
  INV_X1 _16896_ (
    .A(_09237_),
    .ZN(_09238_)
  );
  AND2_X1 _16897_ (
    .A1(_09056_),
    .A2(_09085_),
    .ZN(_09239_)
  );
  INV_X1 _16898_ (
    .A(_09239_),
    .ZN(_09240_)
  );
  AND2_X1 _16899_ (
    .A1(csr_io_decode_0_inst[13]),
    .A2(_09064_),
    .ZN(_09241_)
  );
  INV_X1 _16900_ (
    .A(_09241_),
    .ZN(_09242_)
  );
  AND2_X1 _16901_ (
    .A1(csr_io_decode_0_inst[6]),
    .A2(_09074_),
    .ZN(_09243_)
  );
  INV_X1 _16902_ (
    .A(_09243_),
    .ZN(_09244_)
  );
  AND2_X1 _16903_ (
    .A1(_09013_),
    .A2(_09107_),
    .ZN(_09245_)
  );
  INV_X1 _16904_ (
    .A(_09245_),
    .ZN(_09246_)
  );
  AND2_X1 _16905_ (
    .A1(_09242_),
    .A2(_09246_),
    .ZN(_09247_)
  );
  AND2_X1 _16906_ (
    .A1(_08135_),
    .A2(_08529_),
    .ZN(_09248_)
  );
  AND2_X1 _16907_ (
    .A1(_09054_),
    .A2(_09248_),
    .ZN(_09249_)
  );
  AND2_X1 _16908_ (
    .A1(_09004_),
    .A2(_09249_),
    .ZN(_09250_)
  );
  INV_X1 _16909_ (
    .A(_09250_),
    .ZN(_09251_)
  );
  AND2_X1 _16910_ (
    .A1(_09247_),
    .A2(_09251_),
    .ZN(_09252_)
  );
  AND2_X1 _16911_ (
    .A1(_09240_),
    .A2(_09252_),
    .ZN(_09253_)
  );
  AND2_X1 _16912_ (
    .A1(_09059_),
    .A2(_09091_),
    .ZN(_09254_)
  );
  AND2_X1 _16913_ (
    .A1(_09253_),
    .A2(_09254_),
    .ZN(_09255_)
  );
  AND2_X1 _16914_ (
    .A1(_09238_),
    .A2(_09255_),
    .ZN(_09256_)
  );
  AND2_X1 _16915_ (
    .A1(_08996_),
    .A2(_09107_),
    .ZN(_09257_)
  );
  AND2_X1 _16916_ (
    .A1(_09077_),
    .A2(_09257_),
    .ZN(_09258_)
  );
  AND2_X1 _16917_ (
    .A1(_09218_),
    .A2(_09256_),
    .ZN(_09259_)
  );
  INV_X1 _16918_ (
    .A(_09259_),
    .ZN(_09260_)
  );
  AND2_X1 _16919_ (
    .A1(csr_io_decode_0_inst[12]),
    .A2(_09064_),
    .ZN(_09261_)
  );
  INV_X1 _16920_ (
    .A(_09261_),
    .ZN(_09262_)
  );
  AND2_X1 _16921_ (
    .A1(_08991_),
    .A2(_09064_),
    .ZN(_09263_)
  );
  AND2_X1 _16922_ (
    .A1(_09242_),
    .A2(_09262_),
    .ZN(_09264_)
  );
  AND2_X1 _16923_ (
    .A1(_09214_),
    .A2(_09264_),
    .ZN(_09265_)
  );
  AND2_X1 _16924_ (
    .A1(_09234_),
    .A2(_09265_),
    .ZN(_09266_)
  );
  INV_X1 _16925_ (
    .A(_09266_),
    .ZN(_09267_)
  );
  AND2_X1 _16926_ (
    .A1(_09264_),
    .A2(_09267_),
    .ZN(_09268_)
  );
  INV_X1 _16927_ (
    .A(_09268_),
    .ZN(_09269_)
  );
  AND2_X1 _16928_ (
    .A1(_08578_),
    .A2(csr_io_decode_0_system_illegal),
    .ZN(_09270_)
  );
  AND2_X1 _16929_ (
    .A1(_09268_),
    .A2(_09270_),
    .ZN(_09271_)
  );
  INV_X1 _16930_ (
    .A(_09271_),
    .ZN(_09272_)
  );
  AND2_X1 _16931_ (
    .A1(_09113_),
    .A2(_09241_),
    .ZN(_09273_)
  );
  INV_X1 _16932_ (
    .A(_09273_),
    .ZN(_09274_)
  );
  AND2_X1 _16933_ (
    .A1(csr_io_decode_0_write_illegal),
    .A2(_09274_),
    .ZN(_09275_)
  );
  INV_X1 _16934_ (
    .A(_09275_),
    .ZN(_09276_)
  );
  AND2_X1 _16935_ (
    .A1(_08614_),
    .A2(_09276_),
    .ZN(_09277_)
  );
  INV_X1 _16936_ (
    .A(_09277_),
    .ZN(_09278_)
  );
  AND2_X1 _16937_ (
    .A1(_09263_),
    .A2(_09278_),
    .ZN(_09279_)
  );
  INV_X1 _16938_ (
    .A(_09279_),
    .ZN(_09280_)
  );
  AND2_X1 _16939_ (
    .A1(ibuf_io_inst_0_bits_rvc),
    .A2(_08599_),
    .ZN(_09281_)
  );
  INV_X1 _16940_ (
    .A(_09281_),
    .ZN(_09282_)
  );
  AND2_X1 _16941_ (
    .A1(csr_io_decode_0_inst[25]),
    .A2(_09096_),
    .ZN(_09283_)
  );
  AND2_X1 _16942_ (
    .A1(_08597_),
    .A2(_09283_),
    .ZN(_09284_)
  );
  INV_X1 _16943_ (
    .A(_09284_),
    .ZN(_09285_)
  );
  AND2_X1 _16944_ (
    .A1(_09282_),
    .A2(_09285_),
    .ZN(_09286_)
  );
  AND2_X1 _16945_ (
    .A1(_09280_),
    .A2(_09286_),
    .ZN(_09287_)
  );
  AND2_X1 _16946_ (
    .A1(_09058_),
    .A2(_09092_),
    .ZN(_09288_)
  );
  INV_X1 _16947_ (
    .A(_09288_),
    .ZN(_09289_)
  );
  AND2_X1 _16948_ (
    .A1(_08598_),
    .A2(_09289_),
    .ZN(_09290_)
  );
  INV_X1 _16949_ (
    .A(_09290_),
    .ZN(_09291_)
  );
  AND2_X1 _16950_ (
    .A1(_09287_),
    .A2(_09291_),
    .ZN(_09292_)
  );
  AND2_X1 _16951_ (
    .A1(_09272_),
    .A2(_09292_),
    .ZN(_09293_)
  );
  AND2_X1 _16952_ (
    .A1(_09260_),
    .A2(_09293_),
    .ZN(_09294_)
  );
  INV_X1 _16953_ (
    .A(_09294_),
    .ZN(_09295_)
  );
  AND2_X1 _16954_ (
    .A1(_09183_),
    .A2(_09294_),
    .ZN(_09296_)
  );
  INV_X1 _16955_ (
    .A(_09296_),
    .ZN(_09297_)
  );
  AND2_X1 _16956_ (
    .A1(_07941_),
    .A2(_08617_),
    .ZN(_09298_)
  );
  AND2_X1 _16957_ (
    .A1(_09033_),
    .A2(_09045_),
    .ZN(_09299_)
  );
  INV_X1 _16958_ (
    .A(_09299_),
    .ZN(_09300_)
  );
  AND2_X1 _16959_ (
    .A1(_09187_),
    .A2(_09262_),
    .ZN(_09301_)
  );
  AND2_X1 _16960_ (
    .A1(_09247_),
    .A2(_09301_),
    .ZN(_09302_)
  );
  AND2_X1 _16961_ (
    .A1(csr_io_decode_0_inst[2]),
    .A2(_09016_),
    .ZN(_09303_)
  );
  INV_X1 _16962_ (
    .A(_09303_),
    .ZN(_09304_)
  );
  AND2_X1 _16963_ (
    .A1(csr_io_decode_0_inst[13]),
    .A2(csr_io_decode_0_inst[14]),
    .ZN(_09305_)
  );
  INV_X1 _16964_ (
    .A(_09305_),
    .ZN(_09306_)
  );
  AND2_X1 _16965_ (
    .A1(_08991_),
    .A2(_09001_),
    .ZN(_09307_)
  );
  AND2_X1 _16966_ (
    .A1(_08995_),
    .A2(_09307_),
    .ZN(_09308_)
  );
  INV_X1 _16967_ (
    .A(_09308_),
    .ZN(_09309_)
  );
  AND2_X1 _16968_ (
    .A1(_08989_),
    .A2(_09309_),
    .ZN(_09310_)
  );
  INV_X1 _16969_ (
    .A(_09310_),
    .ZN(_09311_)
  );
  AND2_X1 _16970_ (
    .A1(_09304_),
    .A2(_09311_),
    .ZN(_09312_)
  );
  AND2_X1 _16971_ (
    .A1(_09302_),
    .A2(_09312_),
    .ZN(_09313_)
  );
  AND2_X1 _16972_ (
    .A1(_09059_),
    .A2(_09313_),
    .ZN(_09314_)
  );
  AND2_X1 _16973_ (
    .A1(_09299_),
    .A2(_09314_),
    .ZN(_09315_)
  );
  AND2_X1 _16974_ (
    .A1(_09105_),
    .A2(_09315_),
    .ZN(_09316_)
  );
  INV_X1 _16975_ (
    .A(_09316_),
    .ZN(_09317_)
  );
  AND2_X1 _16976_ (
    .A1(_08548_),
    .A2(_08549_),
    .ZN(_09318_)
  );
  AND2_X1 _16977_ (
    .A1(_08550_),
    .A2(_08552_),
    .ZN(_09319_)
  );
  AND2_X1 _16978_ (
    .A1(_09318_),
    .A2(_09319_),
    .ZN(_09320_)
  );
  AND2_X1 _16979_ (
    .A1(_08551_),
    .A2(_09320_),
    .ZN(_09321_)
  );
  INV_X1 _16980_ (
    .A(_09321_),
    .ZN(_09322_)
  );
  AND2_X1 _16981_ (
    .A1(_09317_),
    .A2(_09322_),
    .ZN(_09323_)
  );
  AND2_X1 _16982_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[0]),
    .A2(_08634_),
    .ZN(_09324_)
  );
  INV_X1 _16983_ (
    .A(_09324_),
    .ZN(_09325_)
  );
  AND2_X1 _16984_ (
    .A1(_08551_),
    .A2(_08643_),
    .ZN(_09326_)
  );
  INV_X1 _16985_ (
    .A(_09326_),
    .ZN(_09327_)
  );
  AND2_X1 _16986_ (
    .A1(_08548_),
    .A2(_08635_),
    .ZN(_09328_)
  );
  INV_X1 _16987_ (
    .A(_09328_),
    .ZN(_09329_)
  );
  AND2_X1 _16988_ (
    .A1(_08550_),
    .A2(_08640_),
    .ZN(_09330_)
  );
  INV_X1 _16989_ (
    .A(_09330_),
    .ZN(_09331_)
  );
  AND2_X1 _16990_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[4]),
    .A2(_08644_),
    .ZN(_09332_)
  );
  INV_X1 _16991_ (
    .A(_09332_),
    .ZN(_09333_)
  );
  AND2_X1 _16992_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[2]),
    .A2(_08639_),
    .ZN(_09334_)
  );
  INV_X1 _16993_ (
    .A(_09334_),
    .ZN(_09335_)
  );
  AND2_X1 _16994_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[3]),
    .A2(_08642_),
    .ZN(_09336_)
  );
  INV_X1 _16995_ (
    .A(_09336_),
    .ZN(_09337_)
  );
  AND2_X1 _16996_ (
    .A1(_08549_),
    .A2(_08637_),
    .ZN(_09338_)
  );
  INV_X1 _16997_ (
    .A(_09338_),
    .ZN(_09339_)
  );
  AND2_X1 _16998_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[1]),
    .A2(_08636_),
    .ZN(_09340_)
  );
  INV_X1 _16999_ (
    .A(_09340_),
    .ZN(_09341_)
  );
  AND2_X1 _17000_ (
    .A1(_08552_),
    .A2(_08645_),
    .ZN(_09342_)
  );
  INV_X1 _17001_ (
    .A(_09342_),
    .ZN(_09343_)
  );
  AND2_X1 _17002_ (
    .A1(_09331_),
    .A2(_09335_),
    .ZN(_09344_)
  );
  AND2_X1 _17003_ (
    .A1(_09327_),
    .A2(_09337_),
    .ZN(_09345_)
  );
  AND2_X1 _17004_ (
    .A1(_09333_),
    .A2(_09343_),
    .ZN(_09346_)
  );
  AND2_X1 _17005_ (
    .A1(_09341_),
    .A2(_09344_),
    .ZN(_09347_)
  );
  AND2_X1 _17006_ (
    .A1(_09345_),
    .A2(_09346_),
    .ZN(_09348_)
  );
  AND2_X1 _17007_ (
    .A1(_09347_),
    .A2(_09348_),
    .ZN(_09349_)
  );
  AND2_X1 _17008_ (
    .A1(_08651_),
    .A2(_09329_),
    .ZN(_09350_)
  );
  AND2_X1 _17009_ (
    .A1(_09325_),
    .A2(_09350_),
    .ZN(_09351_)
  );
  AND2_X1 _17010_ (
    .A1(_09339_),
    .A2(_09351_),
    .ZN(_09352_)
  );
  AND2_X1 _17011_ (
    .A1(_09349_),
    .A2(_09352_),
    .ZN(_09353_)
  );
  INV_X1 _17012_ (
    .A(_09353_),
    .ZN(_09354_)
  );
  MUX2_X1 _17013_ (
    .A(_r[24]),
    .B(_r[25]),
    .S(ibuf_io_inst_0_bits_inst_rd[0]),
    .Z(_09355_)
  );
  AND2_X1 _17014_ (
    .A1(_08550_),
    .A2(_09355_),
    .ZN(_09356_)
  );
  INV_X1 _17015_ (
    .A(_09356_),
    .ZN(_09357_)
  );
  MUX2_X1 _17016_ (
    .A(_r[28]),
    .B(_r[29]),
    .S(ibuf_io_inst_0_bits_inst_rd[0]),
    .Z(_09358_)
  );
  AND2_X1 _17017_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[2]),
    .A2(_09358_),
    .ZN(_09359_)
  );
  INV_X1 _17018_ (
    .A(_09359_),
    .ZN(_09360_)
  );
  AND2_X1 _17019_ (
    .A1(_08549_),
    .A2(_09360_),
    .ZN(_09361_)
  );
  AND2_X1 _17020_ (
    .A1(_09357_),
    .A2(_09361_),
    .ZN(_09362_)
  );
  INV_X1 _17021_ (
    .A(_09362_),
    .ZN(_09363_)
  );
  MUX2_X1 _17022_ (
    .A(_r[26]),
    .B(_r[27]),
    .S(ibuf_io_inst_0_bits_inst_rd[0]),
    .Z(_09364_)
  );
  AND2_X1 _17023_ (
    .A1(_08550_),
    .A2(_09364_),
    .ZN(_09365_)
  );
  INV_X1 _17024_ (
    .A(_09365_),
    .ZN(_09366_)
  );
  MUX2_X1 _17025_ (
    .A(_r[30]),
    .B(_r[31]),
    .S(ibuf_io_inst_0_bits_inst_rd[0]),
    .Z(_09367_)
  );
  AND2_X1 _17026_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[2]),
    .A2(_09367_),
    .ZN(_09368_)
  );
  INV_X1 _17027_ (
    .A(_09368_),
    .ZN(_09369_)
  );
  AND2_X1 _17028_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[1]),
    .A2(_09369_),
    .ZN(_09370_)
  );
  AND2_X1 _17029_ (
    .A1(_09366_),
    .A2(_09370_),
    .ZN(_09371_)
  );
  INV_X1 _17030_ (
    .A(_09371_),
    .ZN(_09372_)
  );
  AND2_X1 _17031_ (
    .A1(_09363_),
    .A2(_09372_),
    .ZN(_09373_)
  );
  AND2_X1 _17032_ (
    .A1(_r[17]),
    .A2(_08549_),
    .ZN(_09374_)
  );
  INV_X1 _17033_ (
    .A(_09374_),
    .ZN(_09375_)
  );
  AND2_X1 _17034_ (
    .A1(_r[19]),
    .A2(ibuf_io_inst_0_bits_inst_rd[1]),
    .ZN(_09376_)
  );
  INV_X1 _17035_ (
    .A(_09376_),
    .ZN(_09377_)
  );
  AND2_X1 _17036_ (
    .A1(_08550_),
    .A2(_09377_),
    .ZN(_09378_)
  );
  AND2_X1 _17037_ (
    .A1(_09375_),
    .A2(_09378_),
    .ZN(_09379_)
  );
  INV_X1 _17038_ (
    .A(_09379_),
    .ZN(_09380_)
  );
  AND2_X1 _17039_ (
    .A1(_r[21]),
    .A2(_08549_),
    .ZN(_09381_)
  );
  INV_X1 _17040_ (
    .A(_09381_),
    .ZN(_09382_)
  );
  AND2_X1 _17041_ (
    .A1(_r[23]),
    .A2(ibuf_io_inst_0_bits_inst_rd[1]),
    .ZN(_09383_)
  );
  INV_X1 _17042_ (
    .A(_09383_),
    .ZN(_09384_)
  );
  AND2_X1 _17043_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[2]),
    .A2(_09384_),
    .ZN(_09385_)
  );
  AND2_X1 _17044_ (
    .A1(_09382_),
    .A2(_09385_),
    .ZN(_09386_)
  );
  INV_X1 _17045_ (
    .A(_09386_),
    .ZN(_09387_)
  );
  AND2_X1 _17046_ (
    .A1(_09380_),
    .A2(_09387_),
    .ZN(_09388_)
  );
  AND2_X1 _17047_ (
    .A1(_r[16]),
    .A2(_08549_),
    .ZN(_09389_)
  );
  INV_X1 _17048_ (
    .A(_09389_),
    .ZN(_09390_)
  );
  AND2_X1 _17049_ (
    .A1(_r[18]),
    .A2(ibuf_io_inst_0_bits_inst_rd[1]),
    .ZN(_09391_)
  );
  INV_X1 _17050_ (
    .A(_09391_),
    .ZN(_09392_)
  );
  AND2_X1 _17051_ (
    .A1(_08550_),
    .A2(_09392_),
    .ZN(_09393_)
  );
  AND2_X1 _17052_ (
    .A1(_09390_),
    .A2(_09393_),
    .ZN(_09394_)
  );
  INV_X1 _17053_ (
    .A(_09394_),
    .ZN(_09395_)
  );
  AND2_X1 _17054_ (
    .A1(_r[20]),
    .A2(_08549_),
    .ZN(_09396_)
  );
  INV_X1 _17055_ (
    .A(_09396_),
    .ZN(_09397_)
  );
  AND2_X1 _17056_ (
    .A1(_r[22]),
    .A2(ibuf_io_inst_0_bits_inst_rd[1]),
    .ZN(_09398_)
  );
  INV_X1 _17057_ (
    .A(_09398_),
    .ZN(_09399_)
  );
  AND2_X1 _17058_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[2]),
    .A2(_09399_),
    .ZN(_09400_)
  );
  AND2_X1 _17059_ (
    .A1(_09397_),
    .A2(_09400_),
    .ZN(_09401_)
  );
  INV_X1 _17060_ (
    .A(_09401_),
    .ZN(_09402_)
  );
  AND2_X1 _17061_ (
    .A1(_09395_),
    .A2(_09402_),
    .ZN(_09403_)
  );
  MUX2_X1 _17062_ (
    .A(_09388_),
    .B(_09403_),
    .S(_08548_),
    .Z(_09404_)
  );
  MUX2_X1 _17063_ (
    .A(_09373_),
    .B(_09404_),
    .S(_08551_),
    .Z(_09405_)
  );
  AND2_X1 _17064_ (
    .A1(_r[4]),
    .A2(_08548_),
    .ZN(_09406_)
  );
  AND2_X1 _17065_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[2]),
    .A2(_09406_),
    .ZN(_09407_)
  );
  INV_X1 _17066_ (
    .A(_09407_),
    .ZN(_09408_)
  );
  MUX2_X1 _17067_ (
    .A(_r[1]),
    .B(_r[5]),
    .S(ibuf_io_inst_0_bits_inst_rd[2]),
    .Z(_09409_)
  );
  AND2_X1 _17068_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[0]),
    .A2(_09409_),
    .ZN(_09410_)
  );
  INV_X1 _17069_ (
    .A(_09410_),
    .ZN(_09411_)
  );
  AND2_X1 _17070_ (
    .A1(_09408_),
    .A2(_09411_),
    .ZN(_09412_)
  );
  INV_X1 _17071_ (
    .A(_09412_),
    .ZN(_09413_)
  );
  AND2_X1 _17072_ (
    .A1(_08549_),
    .A2(_09413_),
    .ZN(_09414_)
  );
  INV_X1 _17073_ (
    .A(_09414_),
    .ZN(_09415_)
  );
  MUX2_X1 _17074_ (
    .A(_r[3]),
    .B(_r[7]),
    .S(ibuf_io_inst_0_bits_inst_rd[2]),
    .Z(_09416_)
  );
  MUX2_X1 _17075_ (
    .A(_r[2]),
    .B(_r[6]),
    .S(ibuf_io_inst_0_bits_inst_rd[2]),
    .Z(_09417_)
  );
  MUX2_X1 _17076_ (
    .A(_09416_),
    .B(_09417_),
    .S(_08548_),
    .Z(_09418_)
  );
  AND2_X1 _17077_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[1]),
    .A2(_09418_),
    .ZN(_09419_)
  );
  INV_X1 _17078_ (
    .A(_09419_),
    .ZN(_09420_)
  );
  AND2_X1 _17079_ (
    .A1(_08551_),
    .A2(_09420_),
    .ZN(_09421_)
  );
  AND2_X1 _17080_ (
    .A1(_09415_),
    .A2(_09421_),
    .ZN(_09422_)
  );
  INV_X1 _17081_ (
    .A(_09422_),
    .ZN(_09423_)
  );
  AND2_X1 _17082_ (
    .A1(_r[14]),
    .A2(_08548_),
    .ZN(_09424_)
  );
  INV_X1 _17083_ (
    .A(_09424_),
    .ZN(_09425_)
  );
  AND2_X1 _17084_ (
    .A1(_r[15]),
    .A2(ibuf_io_inst_0_bits_inst_rd[0]),
    .ZN(_09426_)
  );
  INV_X1 _17085_ (
    .A(_09426_),
    .ZN(_09427_)
  );
  AND2_X1 _17086_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[2]),
    .A2(_09427_),
    .ZN(_09428_)
  );
  AND2_X1 _17087_ (
    .A1(_09425_),
    .A2(_09428_),
    .ZN(_09429_)
  );
  INV_X1 _17088_ (
    .A(_09429_),
    .ZN(_09430_)
  );
  AND2_X1 _17089_ (
    .A1(_r[10]),
    .A2(_08548_),
    .ZN(_09431_)
  );
  INV_X1 _17090_ (
    .A(_09431_),
    .ZN(_09432_)
  );
  AND2_X1 _17091_ (
    .A1(_r[11]),
    .A2(ibuf_io_inst_0_bits_inst_rd[0]),
    .ZN(_09433_)
  );
  INV_X1 _17092_ (
    .A(_09433_),
    .ZN(_09434_)
  );
  AND2_X1 _17093_ (
    .A1(_08550_),
    .A2(_09434_),
    .ZN(_09435_)
  );
  AND2_X1 _17094_ (
    .A1(_09432_),
    .A2(_09435_),
    .ZN(_09436_)
  );
  INV_X1 _17095_ (
    .A(_09436_),
    .ZN(_09437_)
  );
  AND2_X1 _17096_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[1]),
    .A2(_09437_),
    .ZN(_09438_)
  );
  AND2_X1 _17097_ (
    .A1(_09430_),
    .A2(_09438_),
    .ZN(_09439_)
  );
  INV_X1 _17098_ (
    .A(_09439_),
    .ZN(_09440_)
  );
  AND2_X1 _17099_ (
    .A1(_r[12]),
    .A2(_08548_),
    .ZN(_09441_)
  );
  INV_X1 _17100_ (
    .A(_09441_),
    .ZN(_09442_)
  );
  AND2_X1 _17101_ (
    .A1(_r[13]),
    .A2(ibuf_io_inst_0_bits_inst_rd[0]),
    .ZN(_09443_)
  );
  INV_X1 _17102_ (
    .A(_09443_),
    .ZN(_09444_)
  );
  AND2_X1 _17103_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[2]),
    .A2(_09444_),
    .ZN(_09445_)
  );
  AND2_X1 _17104_ (
    .A1(_09442_),
    .A2(_09445_),
    .ZN(_09446_)
  );
  INV_X1 _17105_ (
    .A(_09446_),
    .ZN(_09447_)
  );
  AND2_X1 _17106_ (
    .A1(_r[8]),
    .A2(_08548_),
    .ZN(_09448_)
  );
  INV_X1 _17107_ (
    .A(_09448_),
    .ZN(_09449_)
  );
  AND2_X1 _17108_ (
    .A1(_r[9]),
    .A2(ibuf_io_inst_0_bits_inst_rd[0]),
    .ZN(_09450_)
  );
  INV_X1 _17109_ (
    .A(_09450_),
    .ZN(_09451_)
  );
  AND2_X1 _17110_ (
    .A1(_08550_),
    .A2(_09451_),
    .ZN(_09452_)
  );
  AND2_X1 _17111_ (
    .A1(_09449_),
    .A2(_09452_),
    .ZN(_09453_)
  );
  INV_X1 _17112_ (
    .A(_09453_),
    .ZN(_09454_)
  );
  AND2_X1 _17113_ (
    .A1(_08549_),
    .A2(_09454_),
    .ZN(_09455_)
  );
  AND2_X1 _17114_ (
    .A1(_09447_),
    .A2(_09455_),
    .ZN(_09456_)
  );
  INV_X1 _17115_ (
    .A(_09456_),
    .ZN(_09457_)
  );
  AND2_X1 _17116_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[3]),
    .A2(_09457_),
    .ZN(_09458_)
  );
  AND2_X1 _17117_ (
    .A1(_09440_),
    .A2(_09458_),
    .ZN(_09459_)
  );
  INV_X1 _17118_ (
    .A(_09459_),
    .ZN(_09460_)
  );
  AND2_X1 _17119_ (
    .A1(_09423_),
    .A2(_09460_),
    .ZN(_09461_)
  );
  MUX2_X1 _17120_ (
    .A(_09405_),
    .B(_09461_),
    .S(_08552_),
    .Z(_09462_)
  );
  AND2_X1 _17121_ (
    .A1(_09354_),
    .A2(_09462_),
    .ZN(_09463_)
  );
  AND2_X1 _17122_ (
    .A1(_09323_),
    .A2(_09463_),
    .ZN(_09464_)
  );
  INV_X1 _17123_ (
    .A(_09464_),
    .ZN(_09465_)
  );
  AND2_X1 _17124_ (
    .A1(ex_ctrl_mem),
    .A2(ex_reg_valid),
    .ZN(io_dmem_req_valid)
  );
  INV_X1 _17125_ (
    .A(io_dmem_req_valid),
    .ZN(_09466_)
  );
  AND2_X1 _17126_ (
    .A1(io_dmem_ordered),
    .A2(_09466_),
    .ZN(_09467_)
  );
  INV_X1 _17127_ (
    .A(_09467_),
    .ZN(_09468_)
  );
  AND2_X1 _17128_ (
    .A1(csr_io_decode_0_inst[25]),
    .A2(_09289_),
    .ZN(_09469_)
  );
  INV_X1 _17129_ (
    .A(_09469_),
    .ZN(_09470_)
  );
  AND2_X1 _17130_ (
    .A1(csr_io_decode_0_inst[12]),
    .A2(_09250_),
    .ZN(_09471_)
  );
  INV_X1 _17131_ (
    .A(_09471_),
    .ZN(_09472_)
  );
  AND2_X1 _17132_ (
    .A1(_09470_),
    .A2(_09472_),
    .ZN(_09473_)
  );
  INV_X1 _17133_ (
    .A(_09473_),
    .ZN(_09474_)
  );
  AND2_X1 _17134_ (
    .A1(_09468_),
    .A2(_09474_),
    .ZN(_09475_)
  );
  INV_X1 _17135_ (
    .A(_09475_),
    .ZN(_09476_)
  );
  AND2_X1 _17136_ (
    .A1(_08604_),
    .A2(_08649_),
    .ZN(_09477_)
  );
  INV_X1 _17137_ (
    .A(_09477_),
    .ZN(_09478_)
  );
  AND2_X1 _17138_ (
    .A1(ex_ctrl_div),
    .A2(ex_reg_valid),
    .ZN(div_io_req_valid)
  );
  INV_X1 _17139_ (
    .A(div_io_req_valid),
    .ZN(_09479_)
  );
  AND2_X1 _17140_ (
    .A1(_09478_),
    .A2(_09479_),
    .ZN(_09480_)
  );
  INV_X1 _17141_ (
    .A(_09480_),
    .ZN(_09481_)
  );
  AND2_X1 _17142_ (
    .A1(_09283_),
    .A2(_09481_),
    .ZN(_09482_)
  );
  INV_X1 _17143_ (
    .A(_09482_),
    .ZN(_09483_)
  );
  AND2_X1 _17144_ (
    .A1(_08606_),
    .A2(_08607_),
    .ZN(_09484_)
  );
  AND2_X1 _17145_ (
    .A1(_08610_),
    .A2(_09484_),
    .ZN(_09485_)
  );
  INV_X1 _17146_ (
    .A(_09485_),
    .ZN(_09486_)
  );
  AND2_X1 _17147_ (
    .A1(csr_io_singleStep),
    .A2(_09486_),
    .ZN(_09487_)
  );
  INV_X1 _17148_ (
    .A(_09487_),
    .ZN(_09488_)
  );
  AND2_X1 _17149_ (
    .A1(_07940_),
    .A2(_08616_),
    .ZN(_09489_)
  );
  AND2_X1 _17150_ (
    .A1(_09488_),
    .A2(_09489_),
    .ZN(_09490_)
  );
  AND2_X1 _17151_ (
    .A1(_09483_),
    .A2(_09490_),
    .ZN(_09491_)
  );
  AND2_X1 _17152_ (
    .A1(_08602_),
    .A2(blocked),
    .ZN(_09492_)
  );
  INV_X1 _17153_ (
    .A(_09492_),
    .ZN(_09493_)
  );
  AND2_X1 _17154_ (
    .A1(id_reg_fence),
    .A2(_09468_),
    .ZN(_09494_)
  );
  INV_X1 _17155_ (
    .A(_09494_),
    .ZN(_09495_)
  );
  AND2_X1 _17156_ (
    .A1(_09493_),
    .A2(_09495_),
    .ZN(_09496_)
  );
  INV_X1 _17157_ (
    .A(_09496_),
    .ZN(_09497_)
  );
  AND2_X1 _17158_ (
    .A1(_09010_),
    .A2(_09058_),
    .ZN(_09498_)
  );
  AND2_X1 _17159_ (
    .A1(_09240_),
    .A2(_09498_),
    .ZN(_09499_)
  );
  AND2_X1 _17160_ (
    .A1(_09091_),
    .A2(_09499_),
    .ZN(_09500_)
  );
  INV_X1 _17161_ (
    .A(_09500_),
    .ZN(_09501_)
  );
  AND2_X1 _17162_ (
    .A1(_09497_),
    .A2(_09501_),
    .ZN(_09502_)
  );
  INV_X1 _17163_ (
    .A(_09502_),
    .ZN(_09503_)
  );
  AND2_X1 _17164_ (
    .A1(_09491_),
    .A2(_09503_),
    .ZN(_09504_)
  );
  AND2_X1 _17165_ (
    .A1(_09476_),
    .A2(_09504_),
    .ZN(_09505_)
  );
  AND2_X1 _17166_ (
    .A1(_09465_),
    .A2(_09505_),
    .ZN(_09506_)
  );
  AND2_X1 _17167_ (
    .A1(_09109_),
    .A2(_09114_),
    .ZN(_09507_)
  );
  AND2_X1 _17168_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_08634_),
    .ZN(_09508_)
  );
  INV_X1 _17169_ (
    .A(_09508_),
    .ZN(_09509_)
  );
  AND2_X1 _17170_ (
    .A1(_08540_),
    .A2(_08635_),
    .ZN(_09510_)
  );
  INV_X1 _17171_ (
    .A(_09510_),
    .ZN(_09511_)
  );
  AND2_X1 _17172_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_08642_),
    .ZN(_09512_)
  );
  INV_X1 _17173_ (
    .A(_09512_),
    .ZN(_09513_)
  );
  AND2_X1 _17174_ (
    .A1(_09511_),
    .A2(_09513_),
    .ZN(_09514_)
  );
  AND2_X1 _17175_ (
    .A1(_09509_),
    .A2(_09514_),
    .ZN(_09515_)
  );
  AND2_X1 _17176_ (
    .A1(_08542_),
    .A2(_08640_),
    .ZN(_09516_)
  );
  INV_X1 _17177_ (
    .A(_09516_),
    .ZN(_09517_)
  );
  AND2_X1 _17178_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_08636_),
    .ZN(_09518_)
  );
  INV_X1 _17179_ (
    .A(_09518_),
    .ZN(_09519_)
  );
  AND2_X1 _17180_ (
    .A1(_09517_),
    .A2(_09519_),
    .ZN(_09520_)
  );
  AND2_X1 _17181_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_08639_),
    .ZN(_09521_)
  );
  INV_X1 _17182_ (
    .A(_09521_),
    .ZN(_09522_)
  );
  AND2_X1 _17183_ (
    .A1(_08543_),
    .A2(_08643_),
    .ZN(_09523_)
  );
  INV_X1 _17184_ (
    .A(_09523_),
    .ZN(_09524_)
  );
  AND2_X1 _17185_ (
    .A1(_09522_),
    .A2(_09524_),
    .ZN(_09525_)
  );
  AND2_X1 _17186_ (
    .A1(_09520_),
    .A2(_09525_),
    .ZN(_09526_)
  );
  AND2_X1 _17187_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_08644_),
    .ZN(_09527_)
  );
  INV_X1 _17188_ (
    .A(_09527_),
    .ZN(_09528_)
  );
  AND2_X1 _17189_ (
    .A1(_08571_),
    .A2(_08645_),
    .ZN(_09529_)
  );
  INV_X1 _17190_ (
    .A(_09529_),
    .ZN(_09530_)
  );
  AND2_X1 _17191_ (
    .A1(_09528_),
    .A2(_09530_),
    .ZN(_09531_)
  );
  AND2_X1 _17192_ (
    .A1(_08541_),
    .A2(_08637_),
    .ZN(_09532_)
  );
  INV_X1 _17193_ (
    .A(_09532_),
    .ZN(_09533_)
  );
  AND2_X1 _17194_ (
    .A1(_08651_),
    .A2(_09533_),
    .ZN(_09534_)
  );
  AND2_X1 _17195_ (
    .A1(_09531_),
    .A2(_09534_),
    .ZN(_09535_)
  );
  AND2_X1 _17196_ (
    .A1(_09526_),
    .A2(_09535_),
    .ZN(_09536_)
  );
  AND2_X1 _17197_ (
    .A1(_09515_),
    .A2(_09536_),
    .ZN(_09537_)
  );
  INV_X1 _17198_ (
    .A(_09537_),
    .ZN(_09538_)
  );
  MUX2_X1 _17199_ (
    .A(_r[26]),
    .B(_r[30]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_09539_)
  );
  AND2_X1 _17200_ (
    .A1(_08540_),
    .A2(_09539_),
    .ZN(_09540_)
  );
  INV_X1 _17201_ (
    .A(_09540_),
    .ZN(_09541_)
  );
  AND2_X1 _17202_ (
    .A1(_07944_),
    .A2(_08542_),
    .ZN(_09542_)
  );
  INV_X1 _17203_ (
    .A(_09542_),
    .ZN(_09543_)
  );
  AND2_X1 _17204_ (
    .A1(_07942_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_09544_)
  );
  INV_X1 _17205_ (
    .A(_09544_),
    .ZN(_09545_)
  );
  AND2_X1 _17206_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_09545_),
    .ZN(_09546_)
  );
  AND2_X1 _17207_ (
    .A1(_09543_),
    .A2(_09546_),
    .ZN(_09547_)
  );
  INV_X1 _17208_ (
    .A(_09547_),
    .ZN(_09548_)
  );
  AND2_X1 _17209_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_09548_),
    .ZN(_09549_)
  );
  AND2_X1 _17210_ (
    .A1(_09541_),
    .A2(_09549_),
    .ZN(_09550_)
  );
  INV_X1 _17211_ (
    .A(_09550_),
    .ZN(_09551_)
  );
  AND2_X1 _17212_ (
    .A1(_07943_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_09552_)
  );
  INV_X1 _17213_ (
    .A(_09552_),
    .ZN(_09553_)
  );
  AND2_X1 _17214_ (
    .A1(_07945_),
    .A2(_08542_),
    .ZN(_09554_)
  );
  INV_X1 _17215_ (
    .A(_09554_),
    .ZN(_09555_)
  );
  AND2_X1 _17216_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_09555_),
    .ZN(_09556_)
  );
  AND2_X1 _17217_ (
    .A1(_09553_),
    .A2(_09556_),
    .ZN(_09557_)
  );
  INV_X1 _17218_ (
    .A(_09557_),
    .ZN(_09558_)
  );
  MUX2_X1 _17219_ (
    .A(_r[24]),
    .B(_r[28]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_09559_)
  );
  AND2_X1 _17220_ (
    .A1(_08540_),
    .A2(_09559_),
    .ZN(_09560_)
  );
  INV_X1 _17221_ (
    .A(_09560_),
    .ZN(_09561_)
  );
  AND2_X1 _17222_ (
    .A1(_08541_),
    .A2(_09561_),
    .ZN(_09562_)
  );
  AND2_X1 _17223_ (
    .A1(_09558_),
    .A2(_09562_),
    .ZN(_09563_)
  );
  INV_X1 _17224_ (
    .A(_09563_),
    .ZN(_09564_)
  );
  AND2_X1 _17225_ (
    .A1(_09551_),
    .A2(_09564_),
    .ZN(_09565_)
  );
  AND2_X1 _17226_ (
    .A1(_r[17]),
    .A2(_08541_),
    .ZN(_09566_)
  );
  INV_X1 _17227_ (
    .A(_09566_),
    .ZN(_09567_)
  );
  AND2_X1 _17228_ (
    .A1(_r[19]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_09568_)
  );
  INV_X1 _17229_ (
    .A(_09568_),
    .ZN(_09569_)
  );
  AND2_X1 _17230_ (
    .A1(_08542_),
    .A2(_09569_),
    .ZN(_09570_)
  );
  AND2_X1 _17231_ (
    .A1(_09567_),
    .A2(_09570_),
    .ZN(_09571_)
  );
  INV_X1 _17232_ (
    .A(_09571_),
    .ZN(_09572_)
  );
  AND2_X1 _17233_ (
    .A1(_r[21]),
    .A2(_08541_),
    .ZN(_09573_)
  );
  INV_X1 _17234_ (
    .A(_09573_),
    .ZN(_09574_)
  );
  AND2_X1 _17235_ (
    .A1(_r[23]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_09575_)
  );
  INV_X1 _17236_ (
    .A(_09575_),
    .ZN(_09576_)
  );
  AND2_X1 _17237_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_09576_),
    .ZN(_09577_)
  );
  AND2_X1 _17238_ (
    .A1(_09574_),
    .A2(_09577_),
    .ZN(_09578_)
  );
  INV_X1 _17239_ (
    .A(_09578_),
    .ZN(_09579_)
  );
  AND2_X1 _17240_ (
    .A1(_09572_),
    .A2(_09579_),
    .ZN(_09580_)
  );
  AND2_X1 _17241_ (
    .A1(_r[16]),
    .A2(_08541_),
    .ZN(_09581_)
  );
  INV_X1 _17242_ (
    .A(_09581_),
    .ZN(_09582_)
  );
  AND2_X1 _17243_ (
    .A1(_r[18]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_09583_)
  );
  INV_X1 _17244_ (
    .A(_09583_),
    .ZN(_09584_)
  );
  AND2_X1 _17245_ (
    .A1(_08542_),
    .A2(_09584_),
    .ZN(_09585_)
  );
  AND2_X1 _17246_ (
    .A1(_09582_),
    .A2(_09585_),
    .ZN(_09586_)
  );
  INV_X1 _17247_ (
    .A(_09586_),
    .ZN(_09587_)
  );
  AND2_X1 _17248_ (
    .A1(_r[20]),
    .A2(_08541_),
    .ZN(_09588_)
  );
  INV_X1 _17249_ (
    .A(_09588_),
    .ZN(_09589_)
  );
  AND2_X1 _17250_ (
    .A1(_r[22]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_09590_)
  );
  INV_X1 _17251_ (
    .A(_09590_),
    .ZN(_09591_)
  );
  AND2_X1 _17252_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_09591_),
    .ZN(_09592_)
  );
  AND2_X1 _17253_ (
    .A1(_09589_),
    .A2(_09592_),
    .ZN(_09593_)
  );
  INV_X1 _17254_ (
    .A(_09593_),
    .ZN(_09594_)
  );
  AND2_X1 _17255_ (
    .A1(_09587_),
    .A2(_09594_),
    .ZN(_09595_)
  );
  MUX2_X1 _17256_ (
    .A(_09580_),
    .B(_09595_),
    .S(_08540_),
    .Z(_09596_)
  );
  MUX2_X1 _17257_ (
    .A(_09565_),
    .B(_09596_),
    .S(_08543_),
    .Z(_09597_)
  );
  MUX2_X1 _17258_ (
    .A(_r[6]),
    .B(_r[7]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_09598_)
  );
  MUX2_X1 _17259_ (
    .A(_r[2]),
    .B(_r[3]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_09599_)
  );
  MUX2_X1 _17260_ (
    .A(_09598_),
    .B(_09599_),
    .S(_08542_),
    .Z(_09600_)
  );
  AND2_X1 _17261_ (
    .A1(_07951_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_09601_)
  );
  INV_X1 _17262_ (
    .A(_09601_),
    .ZN(_09602_)
  );
  AND2_X1 _17263_ (
    .A1(_07953_),
    .A2(_08542_),
    .ZN(_09603_)
  );
  INV_X1 _17264_ (
    .A(_09603_),
    .ZN(_09604_)
  );
  AND2_X1 _17265_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_09604_),
    .ZN(_09605_)
  );
  AND2_X1 _17266_ (
    .A1(_09602_),
    .A2(_09605_),
    .ZN(_09606_)
  );
  INV_X1 _17267_ (
    .A(_09606_),
    .ZN(_09607_)
  );
  AND2_X1 _17268_ (
    .A1(_08540_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_09608_)
  );
  AND2_X1 _17269_ (
    .A1(_r[4]),
    .A2(_09608_),
    .ZN(_09609_)
  );
  INV_X1 _17270_ (
    .A(_09609_),
    .ZN(_09610_)
  );
  AND2_X1 _17271_ (
    .A1(_09607_),
    .A2(_09610_),
    .ZN(_09611_)
  );
  INV_X1 _17272_ (
    .A(_09611_),
    .ZN(_09612_)
  );
  MUX2_X1 _17273_ (
    .A(_09600_),
    .B(_09612_),
    .S(_08541_),
    .Z(_09613_)
  );
  AND2_X1 _17274_ (
    .A1(_07946_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_09614_)
  );
  INV_X1 _17275_ (
    .A(_09614_),
    .ZN(_09615_)
  );
  AND2_X1 _17276_ (
    .A1(_07948_),
    .A2(_08542_),
    .ZN(_09616_)
  );
  INV_X1 _17277_ (
    .A(_09616_),
    .ZN(_09617_)
  );
  AND2_X1 _17278_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_09617_),
    .ZN(_09618_)
  );
  AND2_X1 _17279_ (
    .A1(_09615_),
    .A2(_09618_),
    .ZN(_09619_)
  );
  INV_X1 _17280_ (
    .A(_09619_),
    .ZN(_09620_)
  );
  MUX2_X1 _17281_ (
    .A(_r[10]),
    .B(_r[14]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_09621_)
  );
  AND2_X1 _17282_ (
    .A1(_08540_),
    .A2(_09621_),
    .ZN(_09622_)
  );
  INV_X1 _17283_ (
    .A(_09622_),
    .ZN(_09623_)
  );
  AND2_X1 _17284_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_09623_),
    .ZN(_09624_)
  );
  AND2_X1 _17285_ (
    .A1(_09620_),
    .A2(_09624_),
    .ZN(_09625_)
  );
  INV_X1 _17286_ (
    .A(_09625_),
    .ZN(_09626_)
  );
  AND2_X1 _17287_ (
    .A1(_07947_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_09627_)
  );
  INV_X1 _17288_ (
    .A(_09627_),
    .ZN(_09628_)
  );
  AND2_X1 _17289_ (
    .A1(_07949_),
    .A2(_08542_),
    .ZN(_09629_)
  );
  INV_X1 _17290_ (
    .A(_09629_),
    .ZN(_09630_)
  );
  AND2_X1 _17291_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_09630_),
    .ZN(_09631_)
  );
  AND2_X1 _17292_ (
    .A1(_09628_),
    .A2(_09631_),
    .ZN(_09632_)
  );
  INV_X1 _17293_ (
    .A(_09632_),
    .ZN(_09633_)
  );
  MUX2_X1 _17294_ (
    .A(_r[8]),
    .B(_r[12]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_09634_)
  );
  AND2_X1 _17295_ (
    .A1(_08540_),
    .A2(_09634_),
    .ZN(_09635_)
  );
  INV_X1 _17296_ (
    .A(_09635_),
    .ZN(_09636_)
  );
  AND2_X1 _17297_ (
    .A1(_08541_),
    .A2(_09636_),
    .ZN(_09637_)
  );
  AND2_X1 _17298_ (
    .A1(_09633_),
    .A2(_09637_),
    .ZN(_09638_)
  );
  INV_X1 _17299_ (
    .A(_09638_),
    .ZN(_09639_)
  );
  AND2_X1 _17300_ (
    .A1(_09626_),
    .A2(_09639_),
    .ZN(_09640_)
  );
  MUX2_X1 _17301_ (
    .A(_09613_),
    .B(_09640_),
    .S(ibuf_io_inst_0_bits_inst_rs1[3]),
    .Z(_09641_)
  );
  MUX2_X1 _17302_ (
    .A(_09597_),
    .B(_09641_),
    .S(_08571_),
    .Z(_09642_)
  );
  AND2_X1 _17303_ (
    .A1(_09538_),
    .A2(_09642_),
    .ZN(_09643_)
  );
  AND2_X1 _17304_ (
    .A1(_09507_),
    .A2(_09643_),
    .ZN(_09644_)
  );
  INV_X1 _17305_ (
    .A(_09644_),
    .ZN(_09645_)
  );
  AND2_X1 _17306_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[2]),
    .A2(_08639_),
    .ZN(_09646_)
  );
  INV_X1 _17307_ (
    .A(_09646_),
    .ZN(_09647_)
  );
  AND2_X1 _17308_ (
    .A1(_08546_),
    .A2(_08640_),
    .ZN(_09648_)
  );
  INV_X1 _17309_ (
    .A(_09648_),
    .ZN(_09649_)
  );
  AND2_X1 _17310_ (
    .A1(_08544_),
    .A2(_08635_),
    .ZN(_09650_)
  );
  INV_X1 _17311_ (
    .A(_09650_),
    .ZN(_09651_)
  );
  AND2_X1 _17312_ (
    .A1(_09647_),
    .A2(_09649_),
    .ZN(_09652_)
  );
  AND2_X1 _17313_ (
    .A1(_09651_),
    .A2(_09652_),
    .ZN(_09653_)
  );
  AND2_X1 _17314_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[4]),
    .A2(_08644_),
    .ZN(_09654_)
  );
  INV_X1 _17315_ (
    .A(_09654_),
    .ZN(_09655_)
  );
  AND2_X1 _17316_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_08642_),
    .ZN(_09656_)
  );
  INV_X1 _17317_ (
    .A(_09656_),
    .ZN(_09657_)
  );
  AND2_X1 _17318_ (
    .A1(_09655_),
    .A2(_09657_),
    .ZN(_09658_)
  );
  AND2_X1 _17319_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08634_),
    .ZN(_09659_)
  );
  INV_X1 _17320_ (
    .A(_09659_),
    .ZN(_09660_)
  );
  AND2_X1 _17321_ (
    .A1(_08547_),
    .A2(_08643_),
    .ZN(_09661_)
  );
  INV_X1 _17322_ (
    .A(_09661_),
    .ZN(_09662_)
  );
  AND2_X1 _17323_ (
    .A1(_09660_),
    .A2(_09662_),
    .ZN(_09663_)
  );
  AND2_X1 _17324_ (
    .A1(_09658_),
    .A2(_09663_),
    .ZN(_09664_)
  );
  AND2_X1 _17325_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08636_),
    .ZN(_09665_)
  );
  INV_X1 _17326_ (
    .A(_09665_),
    .ZN(_09666_)
  );
  AND2_X1 _17327_ (
    .A1(_08651_),
    .A2(_09666_),
    .ZN(_09667_)
  );
  AND2_X1 _17328_ (
    .A1(_08545_),
    .A2(_08637_),
    .ZN(_09668_)
  );
  INV_X1 _17329_ (
    .A(_09668_),
    .ZN(_09669_)
  );
  AND2_X1 _17330_ (
    .A1(_08572_),
    .A2(_08645_),
    .ZN(_09670_)
  );
  INV_X1 _17331_ (
    .A(_09670_),
    .ZN(_09671_)
  );
  AND2_X1 _17332_ (
    .A1(_09669_),
    .A2(_09671_),
    .ZN(_09672_)
  );
  AND2_X1 _17333_ (
    .A1(_09667_),
    .A2(_09672_),
    .ZN(_09673_)
  );
  AND2_X1 _17334_ (
    .A1(_09664_),
    .A2(_09673_),
    .ZN(_09674_)
  );
  AND2_X1 _17335_ (
    .A1(_09653_),
    .A2(_09674_),
    .ZN(_09675_)
  );
  INV_X1 _17336_ (
    .A(_09675_),
    .ZN(_09676_)
  );
  AND2_X1 _17337_ (
    .A1(_09040_),
    .A2(_09058_),
    .ZN(_09677_)
  );
  AND2_X1 _17338_ (
    .A1(_09068_),
    .A2(_09073_),
    .ZN(_09678_)
  );
  INV_X1 _17339_ (
    .A(_09678_),
    .ZN(_09679_)
  );
  AND2_X1 _17340_ (
    .A1(_08988_),
    .A2(_09052_),
    .ZN(_09680_)
  );
  INV_X1 _17341_ (
    .A(_09680_),
    .ZN(_09681_)
  );
  AND2_X1 _17342_ (
    .A1(_09679_),
    .A2(_09681_),
    .ZN(_09682_)
  );
  INV_X1 _17343_ (
    .A(_09682_),
    .ZN(_09683_)
  );
  AND2_X1 _17344_ (
    .A1(_09020_),
    .A2(_09029_),
    .ZN(_09684_)
  );
  AND2_X1 _17345_ (
    .A1(_09094_),
    .A2(_09684_),
    .ZN(_09685_)
  );
  AND2_X1 _17346_ (
    .A1(_09041_),
    .A2(_09685_),
    .ZN(_09686_)
  );
  INV_X1 _17347_ (
    .A(_09686_),
    .ZN(_09687_)
  );
  AND2_X1 _17348_ (
    .A1(_09682_),
    .A2(_09687_),
    .ZN(_09688_)
  );
  AND2_X1 _17349_ (
    .A1(_09677_),
    .A2(_09688_),
    .ZN(_09689_)
  );
  AND2_X1 _17350_ (
    .A1(_09105_),
    .A2(_09689_),
    .ZN(_09690_)
  );
  INV_X1 _17351_ (
    .A(_09690_),
    .ZN(_09691_)
  );
  AND2_X1 _17352_ (
    .A1(_08544_),
    .A2(_08547_),
    .ZN(_09692_)
  );
  AND2_X1 _17353_ (
    .A1(_08545_),
    .A2(_08546_),
    .ZN(_09693_)
  );
  AND2_X1 _17354_ (
    .A1(_08572_),
    .A2(_09693_),
    .ZN(_09694_)
  );
  AND2_X1 _17355_ (
    .A1(_09692_),
    .A2(_09694_),
    .ZN(_09695_)
  );
  INV_X1 _17356_ (
    .A(_09695_),
    .ZN(_09696_)
  );
  AND2_X1 _17357_ (
    .A1(_09691_),
    .A2(_09696_),
    .ZN(_09697_)
  );
  AND2_X1 _17358_ (
    .A1(_07951_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_09698_)
  );
  INV_X1 _17359_ (
    .A(_09698_),
    .ZN(_09699_)
  );
  AND2_X1 _17360_ (
    .A1(_07953_),
    .A2(_08546_),
    .ZN(_09700_)
  );
  INV_X1 _17361_ (
    .A(_09700_),
    .ZN(_09701_)
  );
  AND2_X1 _17362_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_09701_),
    .ZN(_09702_)
  );
  AND2_X1 _17363_ (
    .A1(_09699_),
    .A2(_09702_),
    .ZN(_09703_)
  );
  INV_X1 _17364_ (
    .A(_09703_),
    .ZN(_09704_)
  );
  AND2_X1 _17365_ (
    .A1(_08544_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_09705_)
  );
  AND2_X1 _17366_ (
    .A1(_r[4]),
    .A2(_09705_),
    .ZN(_09706_)
  );
  INV_X1 _17367_ (
    .A(_09706_),
    .ZN(_09707_)
  );
  AND2_X1 _17368_ (
    .A1(_08545_),
    .A2(_09707_),
    .ZN(_09708_)
  );
  AND2_X1 _17369_ (
    .A1(_09704_),
    .A2(_09708_),
    .ZN(_09709_)
  );
  INV_X1 _17370_ (
    .A(_09709_),
    .ZN(_09710_)
  );
  AND2_X1 _17371_ (
    .A1(_07952_),
    .A2(_08546_),
    .ZN(_09711_)
  );
  INV_X1 _17372_ (
    .A(_09711_),
    .ZN(_09712_)
  );
  AND2_X1 _17373_ (
    .A1(_07950_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_09713_)
  );
  INV_X1 _17374_ (
    .A(_09713_),
    .ZN(_09714_)
  );
  AND2_X1 _17375_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_09714_),
    .ZN(_09715_)
  );
  AND2_X1 _17376_ (
    .A1(_09712_),
    .A2(_09715_),
    .ZN(_09716_)
  );
  INV_X1 _17377_ (
    .A(_09716_),
    .ZN(_09717_)
  );
  MUX2_X1 _17378_ (
    .A(_r[2]),
    .B(_r[6]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_09718_)
  );
  AND2_X1 _17379_ (
    .A1(_08544_),
    .A2(_09718_),
    .ZN(_09719_)
  );
  INV_X1 _17380_ (
    .A(_09719_),
    .ZN(_09720_)
  );
  AND2_X1 _17381_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_09720_),
    .ZN(_09721_)
  );
  AND2_X1 _17382_ (
    .A1(_09717_),
    .A2(_09721_),
    .ZN(_09722_)
  );
  INV_X1 _17383_ (
    .A(_09722_),
    .ZN(_09723_)
  );
  AND2_X1 _17384_ (
    .A1(_09710_),
    .A2(_09723_),
    .ZN(_09724_)
  );
  MUX2_X1 _17385_ (
    .A(_r[10]),
    .B(_r[14]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_09725_)
  );
  AND2_X1 _17386_ (
    .A1(_08544_),
    .A2(_09725_),
    .ZN(_09726_)
  );
  INV_X1 _17387_ (
    .A(_09726_),
    .ZN(_09727_)
  );
  AND2_X1 _17388_ (
    .A1(_07946_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_09728_)
  );
  INV_X1 _17389_ (
    .A(_09728_),
    .ZN(_09729_)
  );
  AND2_X1 _17390_ (
    .A1(_07948_),
    .A2(_08546_),
    .ZN(_09730_)
  );
  INV_X1 _17391_ (
    .A(_09730_),
    .ZN(_09731_)
  );
  AND2_X1 _17392_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_09731_),
    .ZN(_09732_)
  );
  AND2_X1 _17393_ (
    .A1(_09729_),
    .A2(_09732_),
    .ZN(_09733_)
  );
  INV_X1 _17394_ (
    .A(_09733_),
    .ZN(_09734_)
  );
  AND2_X1 _17395_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_09734_),
    .ZN(_09735_)
  );
  AND2_X1 _17396_ (
    .A1(_09727_),
    .A2(_09735_),
    .ZN(_09736_)
  );
  INV_X1 _17397_ (
    .A(_09736_),
    .ZN(_09737_)
  );
  MUX2_X1 _17398_ (
    .A(_r[8]),
    .B(_r[12]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_09738_)
  );
  AND2_X1 _17399_ (
    .A1(_08544_),
    .A2(_09738_),
    .ZN(_09739_)
  );
  INV_X1 _17400_ (
    .A(_09739_),
    .ZN(_09740_)
  );
  AND2_X1 _17401_ (
    .A1(_07947_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_09741_)
  );
  INV_X1 _17402_ (
    .A(_09741_),
    .ZN(_09742_)
  );
  AND2_X1 _17403_ (
    .A1(_07949_),
    .A2(_08546_),
    .ZN(_09743_)
  );
  INV_X1 _17404_ (
    .A(_09743_),
    .ZN(_09744_)
  );
  AND2_X1 _17405_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_09744_),
    .ZN(_09745_)
  );
  AND2_X1 _17406_ (
    .A1(_09742_),
    .A2(_09745_),
    .ZN(_09746_)
  );
  INV_X1 _17407_ (
    .A(_09746_),
    .ZN(_09747_)
  );
  AND2_X1 _17408_ (
    .A1(_09740_),
    .A2(_09747_),
    .ZN(_09748_)
  );
  AND2_X1 _17409_ (
    .A1(_08545_),
    .A2(_09748_),
    .ZN(_09749_)
  );
  INV_X1 _17410_ (
    .A(_09749_),
    .ZN(_09750_)
  );
  AND2_X1 _17411_ (
    .A1(_09737_),
    .A2(_09750_),
    .ZN(_09751_)
  );
  MUX2_X1 _17412_ (
    .A(_09724_),
    .B(_09751_),
    .S(ibuf_io_inst_0_bits_inst_rs2[3]),
    .Z(_09752_)
  );
  AND2_X1 _17413_ (
    .A1(_08572_),
    .A2(_09752_),
    .ZN(_09753_)
  );
  INV_X1 _17414_ (
    .A(_09753_),
    .ZN(_09754_)
  );
  MUX2_X1 _17415_ (
    .A(_r[17]),
    .B(_r[21]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_09755_)
  );
  MUX2_X1 _17416_ (
    .A(_r[16]),
    .B(_r[20]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_09756_)
  );
  MUX2_X1 _17417_ (
    .A(_r[19]),
    .B(_r[23]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_09757_)
  );
  MUX2_X1 _17418_ (
    .A(_r[18]),
    .B(_r[22]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_09758_)
  );
  MUX2_X1 _17419_ (
    .A(_09755_),
    .B(_09756_),
    .S(_08544_),
    .Z(_09759_)
  );
  MUX2_X1 _17420_ (
    .A(_09757_),
    .B(_09758_),
    .S(_08544_),
    .Z(_09760_)
  );
  MUX2_X1 _17421_ (
    .A(_09759_),
    .B(_09760_),
    .S(ibuf_io_inst_0_bits_inst_rs2[1]),
    .Z(_09761_)
  );
  INV_X1 _17422_ (
    .A(_09761_),
    .ZN(_09762_)
  );
  AND2_X1 _17423_ (
    .A1(_08547_),
    .A2(_09762_),
    .ZN(_09763_)
  );
  INV_X1 _17424_ (
    .A(_09763_),
    .ZN(_09764_)
  );
  AND2_X1 _17425_ (
    .A1(_07943_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_09765_)
  );
  INV_X1 _17426_ (
    .A(_09765_),
    .ZN(_09766_)
  );
  AND2_X1 _17427_ (
    .A1(_07945_),
    .A2(_08546_),
    .ZN(_09767_)
  );
  INV_X1 _17428_ (
    .A(_09767_),
    .ZN(_09768_)
  );
  AND2_X1 _17429_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_09768_),
    .ZN(_09769_)
  );
  AND2_X1 _17430_ (
    .A1(_09766_),
    .A2(_09769_),
    .ZN(_09770_)
  );
  INV_X1 _17431_ (
    .A(_09770_),
    .ZN(_09771_)
  );
  MUX2_X1 _17432_ (
    .A(_r[24]),
    .B(_r[28]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_09772_)
  );
  AND2_X1 _17433_ (
    .A1(_08544_),
    .A2(_09772_),
    .ZN(_09773_)
  );
  INV_X1 _17434_ (
    .A(_09773_),
    .ZN(_09774_)
  );
  AND2_X1 _17435_ (
    .A1(_08545_),
    .A2(_09774_),
    .ZN(_09775_)
  );
  AND2_X1 _17436_ (
    .A1(_09771_),
    .A2(_09775_),
    .ZN(_09776_)
  );
  INV_X1 _17437_ (
    .A(_09776_),
    .ZN(_09777_)
  );
  AND2_X1 _17438_ (
    .A1(_07944_),
    .A2(_08546_),
    .ZN(_09778_)
  );
  INV_X1 _17439_ (
    .A(_09778_),
    .ZN(_09779_)
  );
  AND2_X1 _17440_ (
    .A1(_07942_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_09780_)
  );
  INV_X1 _17441_ (
    .A(_09780_),
    .ZN(_09781_)
  );
  AND2_X1 _17442_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_09781_),
    .ZN(_09782_)
  );
  AND2_X1 _17443_ (
    .A1(_09779_),
    .A2(_09782_),
    .ZN(_09783_)
  );
  INV_X1 _17444_ (
    .A(_09783_),
    .ZN(_09784_)
  );
  MUX2_X1 _17445_ (
    .A(_r[26]),
    .B(_r[30]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_09785_)
  );
  AND2_X1 _17446_ (
    .A1(_08544_),
    .A2(_09785_),
    .ZN(_09786_)
  );
  INV_X1 _17447_ (
    .A(_09786_),
    .ZN(_09787_)
  );
  AND2_X1 _17448_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_09787_),
    .ZN(_09788_)
  );
  AND2_X1 _17449_ (
    .A1(_09784_),
    .A2(_09788_),
    .ZN(_09789_)
  );
  INV_X1 _17450_ (
    .A(_09789_),
    .ZN(_09790_)
  );
  AND2_X1 _17451_ (
    .A1(_09777_),
    .A2(_09790_),
    .ZN(_09791_)
  );
  INV_X1 _17452_ (
    .A(_09791_),
    .ZN(_09792_)
  );
  AND2_X1 _17453_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_09792_),
    .ZN(_09793_)
  );
  INV_X1 _17454_ (
    .A(_09793_),
    .ZN(_09794_)
  );
  AND2_X1 _17455_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[4]),
    .A2(_09764_),
    .ZN(_09795_)
  );
  AND2_X1 _17456_ (
    .A1(_09794_),
    .A2(_09795_),
    .ZN(_09796_)
  );
  INV_X1 _17457_ (
    .A(_09796_),
    .ZN(_09797_)
  );
  AND2_X1 _17458_ (
    .A1(_09754_),
    .A2(_09797_),
    .ZN(_09798_)
  );
  INV_X1 _17459_ (
    .A(_09798_),
    .ZN(_09799_)
  );
  AND2_X1 _17460_ (
    .A1(_09697_),
    .A2(_09799_),
    .ZN(_09800_)
  );
  AND2_X1 _17461_ (
    .A1(_09676_),
    .A2(_09800_),
    .ZN(_09801_)
  );
  INV_X1 _17462_ (
    .A(_09801_),
    .ZN(_09802_)
  );
  AND2_X1 _17463_ (
    .A1(_09645_),
    .A2(_09802_),
    .ZN(_09803_)
  );
  AND2_X1 _17464_ (
    .A1(_09506_),
    .A2(_09803_),
    .ZN(_09804_)
  );
  AND2_X1 _17465_ (
    .A1(mem_reg_slow_bypass),
    .A2(mem_ctrl_mem),
    .ZN(_09805_)
  );
  INV_X1 _17466_ (
    .A(_09805_),
    .ZN(_09806_)
  );
  AND2_X1 _17467_ (
    .A1(_08189_),
    .A2(_08191_),
    .ZN(_09807_)
  );
  AND2_X1 _17468_ (
    .A1(_08193_),
    .A2(_08195_),
    .ZN(_09808_)
  );
  AND2_X1 _17469_ (
    .A1(_09807_),
    .A2(_09808_),
    .ZN(_09809_)
  );
  AND2_X1 _17470_ (
    .A1(_09806_),
    .A2(_09809_),
    .ZN(_09810_)
  );
  INV_X1 _17471_ (
    .A(_09810_),
    .ZN(_09811_)
  );
  AND2_X1 _17472_ (
    .A1(mem_reg_inst[8]),
    .A2(_08545_),
    .ZN(_09812_)
  );
  INV_X1 _17473_ (
    .A(_09812_),
    .ZN(_09813_)
  );
  AND2_X1 _17474_ (
    .A1(mem_reg_inst[11]),
    .A2(_08572_),
    .ZN(_09814_)
  );
  INV_X1 _17475_ (
    .A(_09814_),
    .ZN(_09815_)
  );
  AND2_X1 _17476_ (
    .A1(_08086_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_09816_)
  );
  INV_X1 _17477_ (
    .A(_09816_),
    .ZN(_09817_)
  );
  AND2_X1 _17478_ (
    .A1(_08092_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[4]),
    .ZN(_09818_)
  );
  INV_X1 _17479_ (
    .A(_09818_),
    .ZN(_09819_)
  );
  AND2_X1 _17480_ (
    .A1(mem_reg_inst[7]),
    .A2(_08544_),
    .ZN(_09820_)
  );
  INV_X1 _17481_ (
    .A(_09820_),
    .ZN(_09821_)
  );
  AND2_X1 _17482_ (
    .A1(_08084_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[0]),
    .ZN(_09822_)
  );
  INV_X1 _17483_ (
    .A(_09822_),
    .ZN(_09823_)
  );
  AND2_X1 _17484_ (
    .A1(_09821_),
    .A2(_09823_),
    .ZN(_09824_)
  );
  AND2_X1 _17485_ (
    .A1(mem_reg_inst[9]),
    .A2(_08546_),
    .ZN(_09825_)
  );
  INV_X1 _17486_ (
    .A(_09825_),
    .ZN(_09826_)
  );
  AND2_X1 _17487_ (
    .A1(_08088_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_09827_)
  );
  INV_X1 _17488_ (
    .A(_09827_),
    .ZN(_09828_)
  );
  AND2_X1 _17489_ (
    .A1(_09826_),
    .A2(_09828_),
    .ZN(_09829_)
  );
  AND2_X1 _17490_ (
    .A1(_08090_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[3]),
    .ZN(_09830_)
  );
  INV_X1 _17491_ (
    .A(_09830_),
    .ZN(_09831_)
  );
  AND2_X1 _17492_ (
    .A1(mem_reg_inst[10]),
    .A2(_08547_),
    .ZN(_09832_)
  );
  INV_X1 _17493_ (
    .A(_09832_),
    .ZN(_09833_)
  );
  AND2_X1 _17494_ (
    .A1(_09813_),
    .A2(_09831_),
    .ZN(_09834_)
  );
  AND2_X1 _17495_ (
    .A1(_09824_),
    .A2(_09834_),
    .ZN(_09835_)
  );
  AND2_X1 _17496_ (
    .A1(_09819_),
    .A2(_09829_),
    .ZN(_09836_)
  );
  AND2_X1 _17497_ (
    .A1(_09817_),
    .A2(_09836_),
    .ZN(_09837_)
  );
  AND2_X1 _17498_ (
    .A1(_09815_),
    .A2(_09833_),
    .ZN(_09838_)
  );
  AND2_X1 _17499_ (
    .A1(_09835_),
    .A2(_09838_),
    .ZN(_09839_)
  );
  AND2_X1 _17500_ (
    .A1(_09837_),
    .A2(_09839_),
    .ZN(_09840_)
  );
  AND2_X1 _17501_ (
    .A1(_09148_),
    .A2(_09840_),
    .ZN(_09841_)
  );
  INV_X1 _17502_ (
    .A(_09841_),
    .ZN(_09842_)
  );
  AND2_X1 _17503_ (
    .A1(_09697_),
    .A2(_09841_),
    .ZN(_09843_)
  );
  INV_X1 _17504_ (
    .A(_09843_),
    .ZN(_09844_)
  );
  AND2_X1 _17505_ (
    .A1(_09178_),
    .A2(_09507_),
    .ZN(_09845_)
  );
  INV_X1 _17506_ (
    .A(_09845_),
    .ZN(_09846_)
  );
  AND2_X1 _17507_ (
    .A1(_09844_),
    .A2(_09846_),
    .ZN(_09847_)
  );
  AND2_X1 _17508_ (
    .A1(_08090_),
    .A2(ibuf_io_inst_0_bits_inst_rd[3]),
    .ZN(_09848_)
  );
  INV_X1 _17509_ (
    .A(_09848_),
    .ZN(_09849_)
  );
  AND2_X1 _17510_ (
    .A1(mem_reg_inst[9]),
    .A2(_08550_),
    .ZN(_09850_)
  );
  INV_X1 _17511_ (
    .A(_09850_),
    .ZN(_09851_)
  );
  AND2_X1 _17512_ (
    .A1(mem_reg_inst[10]),
    .A2(_08551_),
    .ZN(_09852_)
  );
  INV_X1 _17513_ (
    .A(_09852_),
    .ZN(_09853_)
  );
  AND2_X1 _17514_ (
    .A1(_09851_),
    .A2(_09853_),
    .ZN(_09854_)
  );
  AND2_X1 _17515_ (
    .A1(_09849_),
    .A2(_09854_),
    .ZN(_09855_)
  );
  AND2_X1 _17516_ (
    .A1(_08084_),
    .A2(ibuf_io_inst_0_bits_inst_rd[0]),
    .ZN(_09856_)
  );
  INV_X1 _17517_ (
    .A(_09856_),
    .ZN(_09857_)
  );
  AND2_X1 _17518_ (
    .A1(mem_reg_inst[8]),
    .A2(_08549_),
    .ZN(_09858_)
  );
  INV_X1 _17519_ (
    .A(_09858_),
    .ZN(_09859_)
  );
  AND2_X1 _17520_ (
    .A1(_09857_),
    .A2(_09859_),
    .ZN(_09860_)
  );
  AND2_X1 _17521_ (
    .A1(_08088_),
    .A2(ibuf_io_inst_0_bits_inst_rd[2]),
    .ZN(_09861_)
  );
  INV_X1 _17522_ (
    .A(_09861_),
    .ZN(_09862_)
  );
  AND2_X1 _17523_ (
    .A1(_08086_),
    .A2(ibuf_io_inst_0_bits_inst_rd[1]),
    .ZN(_09863_)
  );
  INV_X1 _17524_ (
    .A(_09863_),
    .ZN(_09864_)
  );
  AND2_X1 _17525_ (
    .A1(_09862_),
    .A2(_09864_),
    .ZN(_09865_)
  );
  AND2_X1 _17526_ (
    .A1(_09860_),
    .A2(_09865_),
    .ZN(_09866_)
  );
  AND2_X1 _17527_ (
    .A1(mem_reg_inst[11]),
    .A2(_08552_),
    .ZN(_09867_)
  );
  INV_X1 _17528_ (
    .A(_09867_),
    .ZN(_09868_)
  );
  AND2_X1 _17529_ (
    .A1(_08092_),
    .A2(ibuf_io_inst_0_bits_inst_rd[4]),
    .ZN(_09869_)
  );
  INV_X1 _17530_ (
    .A(_09869_),
    .ZN(_09870_)
  );
  AND2_X1 _17531_ (
    .A1(_09868_),
    .A2(_09870_),
    .ZN(_09871_)
  );
  AND2_X1 _17532_ (
    .A1(mem_reg_inst[7]),
    .A2(_08548_),
    .ZN(_09872_)
  );
  INV_X1 _17533_ (
    .A(_09872_),
    .ZN(_09873_)
  );
  AND2_X1 _17534_ (
    .A1(_09148_),
    .A2(_09873_),
    .ZN(_09874_)
  );
  AND2_X1 _17535_ (
    .A1(_09871_),
    .A2(_09874_),
    .ZN(_09875_)
  );
  AND2_X1 _17536_ (
    .A1(_09866_),
    .A2(_09875_),
    .ZN(_09876_)
  );
  AND2_X1 _17537_ (
    .A1(_09855_),
    .A2(_09876_),
    .ZN(_09877_)
  );
  AND2_X1 _17538_ (
    .A1(_09323_),
    .A2(_09877_),
    .ZN(_09878_)
  );
  INV_X1 _17539_ (
    .A(_09878_),
    .ZN(_09879_)
  );
  AND2_X1 _17540_ (
    .A1(_09847_),
    .A2(_09879_),
    .ZN(_09880_)
  );
  INV_X1 _17541_ (
    .A(_09880_),
    .ZN(_09881_)
  );
  AND2_X1 _17542_ (
    .A1(_09811_),
    .A2(_09881_),
    .ZN(_09882_)
  );
  INV_X1 _17543_ (
    .A(_09882_),
    .ZN(_09883_)
  );
  AND2_X1 _17544_ (
    .A1(_09804_),
    .A2(_09883_),
    .ZN(_09884_)
  );
  AND2_X1 _17545_ (
    .A1(_08646_),
    .A2(_08664_),
    .ZN(_09885_)
  );
  AND2_X1 _17546_ (
    .A1(_08198_),
    .A2(_08546_),
    .ZN(_09886_)
  );
  INV_X1 _17547_ (
    .A(_09886_),
    .ZN(_09887_)
  );
  AND2_X1 _17548_ (
    .A1(wb_reg_inst[9]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_09888_)
  );
  INV_X1 _17549_ (
    .A(_09888_),
    .ZN(_09889_)
  );
  AND2_X1 _17550_ (
    .A1(_09887_),
    .A2(_09889_),
    .ZN(_09890_)
  );
  INV_X1 _17551_ (
    .A(_09890_),
    .ZN(_09891_)
  );
  AND2_X1 _17552_ (
    .A1(_08197_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_09892_)
  );
  INV_X1 _17553_ (
    .A(_09892_),
    .ZN(_09893_)
  );
  AND2_X1 _17554_ (
    .A1(wb_reg_inst[7]),
    .A2(_08544_),
    .ZN(_09894_)
  );
  INV_X1 _17555_ (
    .A(_09894_),
    .ZN(_09895_)
  );
  AND2_X1 _17556_ (
    .A1(wb_reg_inst[8]),
    .A2(_08545_),
    .ZN(_09896_)
  );
  INV_X1 _17557_ (
    .A(_09896_),
    .ZN(_09897_)
  );
  AND2_X1 _17558_ (
    .A1(_09895_),
    .A2(_09897_),
    .ZN(_09898_)
  );
  AND2_X1 _17559_ (
    .A1(_09893_),
    .A2(_09898_),
    .ZN(_09899_)
  );
  AND2_X1 _17560_ (
    .A1(_08199_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[3]),
    .ZN(_09900_)
  );
  INV_X1 _17561_ (
    .A(_09900_),
    .ZN(_09901_)
  );
  AND2_X1 _17562_ (
    .A1(_08196_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[0]),
    .ZN(_09902_)
  );
  INV_X1 _17563_ (
    .A(_09902_),
    .ZN(_09903_)
  );
  AND2_X1 _17564_ (
    .A1(_08200_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[4]),
    .ZN(_09904_)
  );
  INV_X1 _17565_ (
    .A(_09904_),
    .ZN(_09905_)
  );
  AND2_X1 _17566_ (
    .A1(_09901_),
    .A2(_09905_),
    .ZN(_09906_)
  );
  AND2_X1 _17567_ (
    .A1(wb_reg_inst[11]),
    .A2(_08572_),
    .ZN(_09907_)
  );
  INV_X1 _17568_ (
    .A(_09907_),
    .ZN(_09908_)
  );
  AND2_X1 _17569_ (
    .A1(_09903_),
    .A2(_09908_),
    .ZN(_09909_)
  );
  AND2_X1 _17570_ (
    .A1(_09906_),
    .A2(_09909_),
    .ZN(_09910_)
  );
  AND2_X1 _17571_ (
    .A1(wb_reg_inst[10]),
    .A2(_08547_),
    .ZN(_09911_)
  );
  INV_X1 _17572_ (
    .A(_09911_),
    .ZN(_09912_)
  );
  AND2_X1 _17573_ (
    .A1(_09891_),
    .A2(_09912_),
    .ZN(_09913_)
  );
  AND2_X1 _17574_ (
    .A1(_09910_),
    .A2(_09913_),
    .ZN(_09914_)
  );
  AND2_X1 _17575_ (
    .A1(_09899_),
    .A2(_09914_),
    .ZN(_09915_)
  );
  AND2_X1 _17576_ (
    .A1(_09697_),
    .A2(_09915_),
    .ZN(_09916_)
  );
  INV_X1 _17577_ (
    .A(_09916_),
    .ZN(_09917_)
  );
  AND2_X1 _17578_ (
    .A1(_08197_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_09918_)
  );
  INV_X1 _17579_ (
    .A(_09918_),
    .ZN(_09919_)
  );
  AND2_X1 _17580_ (
    .A1(_08199_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[3]),
    .ZN(_09920_)
  );
  INV_X1 _17581_ (
    .A(_09920_),
    .ZN(_09921_)
  );
  AND2_X1 _17582_ (
    .A1(wb_reg_inst[9]),
    .A2(_08542_),
    .ZN(_09922_)
  );
  INV_X1 _17583_ (
    .A(_09922_),
    .ZN(_09923_)
  );
  AND2_X1 _17584_ (
    .A1(_08198_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_09924_)
  );
  INV_X1 _17585_ (
    .A(_09924_),
    .ZN(_09925_)
  );
  AND2_X1 _17586_ (
    .A1(wb_reg_inst[11]),
    .A2(_08571_),
    .ZN(_09926_)
  );
  INV_X1 _17587_ (
    .A(_09926_),
    .ZN(_09927_)
  );
  AND2_X1 _17588_ (
    .A1(_08200_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[4]),
    .ZN(_09928_)
  );
  INV_X1 _17589_ (
    .A(_09928_),
    .ZN(_09929_)
  );
  AND2_X1 _17590_ (
    .A1(_08196_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[0]),
    .ZN(_09930_)
  );
  INV_X1 _17591_ (
    .A(_09930_),
    .ZN(_09931_)
  );
  AND2_X1 _17592_ (
    .A1(wb_reg_inst[7]),
    .A2(_08540_),
    .ZN(_09932_)
  );
  INV_X1 _17593_ (
    .A(_09932_),
    .ZN(_09933_)
  );
  AND2_X1 _17594_ (
    .A1(_09931_),
    .A2(_09933_),
    .ZN(_09934_)
  );
  AND2_X1 _17595_ (
    .A1(wb_reg_inst[8]),
    .A2(_08541_),
    .ZN(_09935_)
  );
  INV_X1 _17596_ (
    .A(_09935_),
    .ZN(_09936_)
  );
  AND2_X1 _17597_ (
    .A1(wb_reg_inst[10]),
    .A2(_08543_),
    .ZN(_09937_)
  );
  INV_X1 _17598_ (
    .A(_09937_),
    .ZN(_09938_)
  );
  AND2_X1 _17599_ (
    .A1(_09923_),
    .A2(_09938_),
    .ZN(_09939_)
  );
  AND2_X1 _17600_ (
    .A1(_09934_),
    .A2(_09939_),
    .ZN(_09940_)
  );
  AND2_X1 _17601_ (
    .A1(_09919_),
    .A2(_09936_),
    .ZN(_09941_)
  );
  AND2_X1 _17602_ (
    .A1(_09925_),
    .A2(_09927_),
    .ZN(_09942_)
  );
  AND2_X1 _17603_ (
    .A1(_09921_),
    .A2(_09929_),
    .ZN(_09943_)
  );
  AND2_X1 _17604_ (
    .A1(_09942_),
    .A2(_09943_),
    .ZN(_09944_)
  );
  AND2_X1 _17605_ (
    .A1(_09940_),
    .A2(_09944_),
    .ZN(_09945_)
  );
  AND2_X1 _17606_ (
    .A1(_09941_),
    .A2(_09945_),
    .ZN(_09946_)
  );
  AND2_X1 _17607_ (
    .A1(_09507_),
    .A2(_09946_),
    .ZN(_09947_)
  );
  INV_X1 _17608_ (
    .A(_09947_),
    .ZN(_09948_)
  );
  AND2_X1 _17609_ (
    .A1(_09917_),
    .A2(_09948_),
    .ZN(_09949_)
  );
  AND2_X1 _17610_ (
    .A1(_08199_),
    .A2(ibuf_io_inst_0_bits_inst_rd[3]),
    .ZN(_09950_)
  );
  INV_X1 _17611_ (
    .A(_09950_),
    .ZN(_09951_)
  );
  AND2_X1 _17612_ (
    .A1(_08197_),
    .A2(ibuf_io_inst_0_bits_inst_rd[1]),
    .ZN(_09952_)
  );
  INV_X1 _17613_ (
    .A(_09952_),
    .ZN(_09953_)
  );
  AND2_X1 _17614_ (
    .A1(_08200_),
    .A2(ibuf_io_inst_0_bits_inst_rd[4]),
    .ZN(_09954_)
  );
  INV_X1 _17615_ (
    .A(_09954_),
    .ZN(_09955_)
  );
  AND2_X1 _17616_ (
    .A1(wb_reg_inst[11]),
    .A2(_08552_),
    .ZN(_09956_)
  );
  INV_X1 _17617_ (
    .A(_09956_),
    .ZN(_09957_)
  );
  AND2_X1 _17618_ (
    .A1(wb_reg_inst[9]),
    .A2(_08550_),
    .ZN(_09958_)
  );
  INV_X1 _17619_ (
    .A(_09958_),
    .ZN(_09959_)
  );
  AND2_X1 _17620_ (
    .A1(_08198_),
    .A2(ibuf_io_inst_0_bits_inst_rd[2]),
    .ZN(_09960_)
  );
  INV_X1 _17621_ (
    .A(_09960_),
    .ZN(_09961_)
  );
  AND2_X1 _17622_ (
    .A1(_09959_),
    .A2(_09961_),
    .ZN(_09962_)
  );
  AND2_X1 _17623_ (
    .A1(wb_reg_inst[7]),
    .A2(_08548_),
    .ZN(_09963_)
  );
  INV_X1 _17624_ (
    .A(_09963_),
    .ZN(_09964_)
  );
  AND2_X1 _17625_ (
    .A1(_08196_),
    .A2(ibuf_io_inst_0_bits_inst_rd[0]),
    .ZN(_09965_)
  );
  INV_X1 _17626_ (
    .A(_09965_),
    .ZN(_09966_)
  );
  AND2_X1 _17627_ (
    .A1(_09964_),
    .A2(_09966_),
    .ZN(_09967_)
  );
  AND2_X1 _17628_ (
    .A1(wb_reg_inst[8]),
    .A2(_08549_),
    .ZN(_09968_)
  );
  INV_X1 _17629_ (
    .A(_09968_),
    .ZN(_09969_)
  );
  AND2_X1 _17630_ (
    .A1(wb_reg_inst[10]),
    .A2(_08551_),
    .ZN(_09970_)
  );
  INV_X1 _17631_ (
    .A(_09970_),
    .ZN(_09971_)
  );
  AND2_X1 _17632_ (
    .A1(_09957_),
    .A2(_09971_),
    .ZN(_09972_)
  );
  AND2_X1 _17633_ (
    .A1(_09967_),
    .A2(_09972_),
    .ZN(_09973_)
  );
  AND2_X1 _17634_ (
    .A1(_09953_),
    .A2(_09969_),
    .ZN(_09974_)
  );
  AND2_X1 _17635_ (
    .A1(_09951_),
    .A2(_09955_),
    .ZN(_09975_)
  );
  AND2_X1 _17636_ (
    .A1(_09962_),
    .A2(_09975_),
    .ZN(_09976_)
  );
  AND2_X1 _17637_ (
    .A1(_09974_),
    .A2(_09976_),
    .ZN(_09977_)
  );
  AND2_X1 _17638_ (
    .A1(_09973_),
    .A2(_09977_),
    .ZN(_09978_)
  );
  AND2_X1 _17639_ (
    .A1(_09323_),
    .A2(_09978_),
    .ZN(_09979_)
  );
  INV_X1 _17640_ (
    .A(_09979_),
    .ZN(_09980_)
  );
  AND2_X1 _17641_ (
    .A1(_09949_),
    .A2(_09980_),
    .ZN(_09981_)
  );
  INV_X1 _17642_ (
    .A(_09981_),
    .ZN(_09982_)
  );
  AND2_X1 _17643_ (
    .A1(_09885_),
    .A2(_09982_),
    .ZN(_09983_)
  );
  INV_X1 _17644_ (
    .A(_09983_),
    .ZN(_09984_)
  );
  AND2_X1 _17645_ (
    .A1(_08201_),
    .A2(_08202_),
    .ZN(_09985_)
  );
  AND2_X1 _17646_ (
    .A1(_08203_),
    .A2(_08207_),
    .ZN(_09986_)
  );
  AND2_X1 _17647_ (
    .A1(_08204_),
    .A2(_08205_),
    .ZN(_09987_)
  );
  AND2_X1 _17648_ (
    .A1(_09985_),
    .A2(_09987_),
    .ZN(_09988_)
  );
  AND2_X1 _17649_ (
    .A1(_09986_),
    .A2(_09988_),
    .ZN(_09989_)
  );
  INV_X1 _17650_ (
    .A(_09989_),
    .ZN(_09990_)
  );
  AND2_X1 _17651_ (
    .A1(_09115_),
    .A2(_09990_),
    .ZN(_09991_)
  );
  AND2_X1 _17652_ (
    .A1(_09144_),
    .A2(_09507_),
    .ZN(_09992_)
  );
  INV_X1 _17653_ (
    .A(_09992_),
    .ZN(_09993_)
  );
  AND2_X1 _17654_ (
    .A1(ex_reg_inst[8]),
    .A2(_08545_),
    .ZN(_09994_)
  );
  INV_X1 _17655_ (
    .A(_09994_),
    .ZN(_09995_)
  );
  AND2_X1 _17656_ (
    .A1(ex_reg_inst[11]),
    .A2(_08572_),
    .ZN(_09996_)
  );
  INV_X1 _17657_ (
    .A(_09996_),
    .ZN(_09997_)
  );
  AND2_X1 _17658_ (
    .A1(_08087_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_09998_)
  );
  INV_X1 _17659_ (
    .A(_09998_),
    .ZN(_09999_)
  );
  AND2_X1 _17660_ (
    .A1(_08093_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[4]),
    .ZN(_10000_)
  );
  INV_X1 _17661_ (
    .A(_10000_),
    .ZN(_10001_)
  );
  AND2_X1 _17662_ (
    .A1(ex_reg_inst[7]),
    .A2(_08544_),
    .ZN(_10002_)
  );
  INV_X1 _17663_ (
    .A(_10002_),
    .ZN(_10003_)
  );
  AND2_X1 _17664_ (
    .A1(_08085_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[0]),
    .ZN(_10004_)
  );
  INV_X1 _17665_ (
    .A(_10004_),
    .ZN(_10005_)
  );
  AND2_X1 _17666_ (
    .A1(_10003_),
    .A2(_10005_),
    .ZN(_10006_)
  );
  AND2_X1 _17667_ (
    .A1(ex_reg_inst[9]),
    .A2(_08546_),
    .ZN(_10007_)
  );
  INV_X1 _17668_ (
    .A(_10007_),
    .ZN(_10008_)
  );
  AND2_X1 _17669_ (
    .A1(_08089_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_10009_)
  );
  INV_X1 _17670_ (
    .A(_10009_),
    .ZN(_10010_)
  );
  AND2_X1 _17671_ (
    .A1(_10008_),
    .A2(_10010_),
    .ZN(_10011_)
  );
  AND2_X1 _17672_ (
    .A1(_08091_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[3]),
    .ZN(_10012_)
  );
  INV_X1 _17673_ (
    .A(_10012_),
    .ZN(_10013_)
  );
  AND2_X1 _17674_ (
    .A1(ex_reg_inst[10]),
    .A2(_08547_),
    .ZN(_10014_)
  );
  INV_X1 _17675_ (
    .A(_10014_),
    .ZN(_10015_)
  );
  AND2_X1 _17676_ (
    .A1(_09995_),
    .A2(_10013_),
    .ZN(_10016_)
  );
  AND2_X1 _17677_ (
    .A1(_10006_),
    .A2(_10016_),
    .ZN(_10017_)
  );
  AND2_X1 _17678_ (
    .A1(_10001_),
    .A2(_10011_),
    .ZN(_10018_)
  );
  AND2_X1 _17679_ (
    .A1(_09999_),
    .A2(_10018_),
    .ZN(_10019_)
  );
  AND2_X1 _17680_ (
    .A1(_09997_),
    .A2(_10015_),
    .ZN(_10020_)
  );
  AND2_X1 _17681_ (
    .A1(_10017_),
    .A2(_10020_),
    .ZN(_10021_)
  );
  AND2_X1 _17682_ (
    .A1(_10019_),
    .A2(_10021_),
    .ZN(_10022_)
  );
  AND2_X1 _17683_ (
    .A1(_09697_),
    .A2(_10022_),
    .ZN(_10023_)
  );
  INV_X1 _17684_ (
    .A(_10023_),
    .ZN(_10024_)
  );
  AND2_X1 _17685_ (
    .A1(_08093_),
    .A2(ibuf_io_inst_0_bits_inst_rd[4]),
    .ZN(_10025_)
  );
  INV_X1 _17686_ (
    .A(_10025_),
    .ZN(_10026_)
  );
  AND2_X1 _17687_ (
    .A1(ex_reg_inst[11]),
    .A2(_08552_),
    .ZN(_10027_)
  );
  INV_X1 _17688_ (
    .A(_10027_),
    .ZN(_10028_)
  );
  AND2_X1 _17689_ (
    .A1(_10026_),
    .A2(_10028_),
    .ZN(_10029_)
  );
  AND2_X1 _17690_ (
    .A1(_08091_),
    .A2(ibuf_io_inst_0_bits_inst_rd[3]),
    .ZN(_10030_)
  );
  INV_X1 _17691_ (
    .A(_10030_),
    .ZN(_10031_)
  );
  AND2_X1 _17692_ (
    .A1(_08085_),
    .A2(ibuf_io_inst_0_bits_inst_rd[0]),
    .ZN(_10032_)
  );
  INV_X1 _17693_ (
    .A(_10032_),
    .ZN(_10033_)
  );
  AND2_X1 _17694_ (
    .A1(_10031_),
    .A2(_10033_),
    .ZN(_10034_)
  );
  AND2_X1 _17695_ (
    .A1(_10029_),
    .A2(_10034_),
    .ZN(_10035_)
  );
  AND2_X1 _17696_ (
    .A1(_08089_),
    .A2(_08550_),
    .ZN(_10036_)
  );
  INV_X1 _17697_ (
    .A(_10036_),
    .ZN(_10037_)
  );
  AND2_X1 _17698_ (
    .A1(ex_reg_inst[9]),
    .A2(ibuf_io_inst_0_bits_inst_rd[2]),
    .ZN(_10038_)
  );
  INV_X1 _17699_ (
    .A(_10038_),
    .ZN(_10039_)
  );
  AND2_X1 _17700_ (
    .A1(_10037_),
    .A2(_10039_),
    .ZN(_10040_)
  );
  INV_X1 _17701_ (
    .A(_10040_),
    .ZN(_10041_)
  );
  AND2_X1 _17702_ (
    .A1(ex_reg_inst[8]),
    .A2(_08549_),
    .ZN(_10042_)
  );
  INV_X1 _17703_ (
    .A(_10042_),
    .ZN(_10043_)
  );
  AND2_X1 _17704_ (
    .A1(_08087_),
    .A2(ibuf_io_inst_0_bits_inst_rd[1]),
    .ZN(_10044_)
  );
  INV_X1 _17705_ (
    .A(_10044_),
    .ZN(_10045_)
  );
  AND2_X1 _17706_ (
    .A1(_10043_),
    .A2(_10045_),
    .ZN(_10046_)
  );
  AND2_X1 _17707_ (
    .A1(ex_reg_inst[10]),
    .A2(_08551_),
    .ZN(_10047_)
  );
  INV_X1 _17708_ (
    .A(_10047_),
    .ZN(_10048_)
  );
  AND2_X1 _17709_ (
    .A1(ex_reg_inst[7]),
    .A2(_08548_),
    .ZN(_10049_)
  );
  INV_X1 _17710_ (
    .A(_10049_),
    .ZN(_10050_)
  );
  AND2_X1 _17711_ (
    .A1(_10048_),
    .A2(_10050_),
    .ZN(_10051_)
  );
  AND2_X1 _17712_ (
    .A1(_10046_),
    .A2(_10051_),
    .ZN(_10052_)
  );
  AND2_X1 _17713_ (
    .A1(_10041_),
    .A2(_10052_),
    .ZN(_10053_)
  );
  AND2_X1 _17714_ (
    .A1(_10035_),
    .A2(_10053_),
    .ZN(_10054_)
  );
  AND2_X1 _17715_ (
    .A1(_09323_),
    .A2(_10054_),
    .ZN(_10055_)
  );
  INV_X1 _17716_ (
    .A(_10055_),
    .ZN(_10056_)
  );
  AND2_X1 _17717_ (
    .A1(_10024_),
    .A2(_10056_),
    .ZN(_10057_)
  );
  AND2_X1 _17718_ (
    .A1(_09993_),
    .A2(_10057_),
    .ZN(_10058_)
  );
  INV_X1 _17719_ (
    .A(_10058_),
    .ZN(_10059_)
  );
  AND2_X1 _17720_ (
    .A1(_09991_),
    .A2(_10059_),
    .ZN(_10060_)
  );
  INV_X1 _17721_ (
    .A(_10060_),
    .ZN(_10061_)
  );
  AND2_X1 _17722_ (
    .A1(_09984_),
    .A2(_10061_),
    .ZN(_10062_)
  );
  AND2_X1 _17723_ (
    .A1(_09884_),
    .A2(_10062_),
    .ZN(ibuf_io_inst_0_ready)
  );
  AND2_X1 _17724_ (
    .A1(_08612_),
    .A2(_08685_),
    .ZN(_10063_)
  );
  INV_X1 _17725_ (
    .A(_10063_),
    .ZN(_10064_)
  );
  AND2_X1 _17726_ (
    .A1(_08613_),
    .A2(_08686_),
    .ZN(_10065_)
  );
  AND2_X1 _17727_ (
    .A1(_10063_),
    .A2(_10065_),
    .ZN(io_imem_req_bits_speculative)
  );
  AND2_X1 _17728_ (
    .A1(mem_br_taken),
    .A2(mem_ctrl_branch),
    .ZN(_10066_)
  );
  INV_X1 _17729_ (
    .A(_10066_),
    .ZN(_10067_)
  );
  AND2_X1 _17730_ (
    .A1(_08208_),
    .A2(_10067_),
    .ZN(_10068_)
  );
  INV_X1 _17731_ (
    .A(_10068_),
    .ZN(_10069_)
  );
  AND2_X1 _17732_ (
    .A1(_08206_),
    .A2(_10068_),
    .ZN(_10070_)
  );
  INV_X1 _17733_ (
    .A(_10070_),
    .ZN(_10071_)
  );
  AND2_X1 _17734_ (
    .A1(mem_reg_valid),
    .A2(_take_pc_mem_T),
    .ZN(_10072_)
  );
  AND2_X1 _17735_ (
    .A1(_10071_),
    .A2(_10072_),
    .ZN(_10073_)
  );
  INV_X1 _17736_ (
    .A(_10073_),
    .ZN(_10074_)
  );
  AND2_X1 _17737_ (
    .A1(io_imem_req_bits_speculative),
    .A2(_10074_),
    .ZN(_10075_)
  );
  INV_X1 _17738_ (
    .A(_10075_),
    .ZN(ibuf_io_kill)
  );
  AND2_X1 _17739_ (
    .A1(ibuf_io_inst_0_valid),
    .A2(_10075_),
    .ZN(_10076_)
  );
  AND2_X1 _17740_ (
    .A1(ibuf_io_inst_0_ready),
    .A2(_10076_),
    .ZN(_10077_)
  );
  AND2_X1 _17741_ (
    .A1(_09298_),
    .A2(_10077_),
    .ZN(_ex_reg_valid_T)
  );
  INV_X1 _17742_ (
    .A(_ex_reg_valid_T),
    .ZN(_10078_)
  );
  AND2_X1 _17743_ (
    .A1(_09297_),
    .A2(_ex_reg_valid_T),
    .ZN(_10079_)
  );
  AND2_X1 _17744_ (
    .A1(ibuf_io_inst_0_bits_raw[2]),
    .A2(_09295_),
    .ZN(_10080_)
  );
  INV_X1 _17745_ (
    .A(_10080_),
    .ZN(_10081_)
  );
  AND2_X1 _17746_ (
    .A1(_09182_),
    .A2(_09294_),
    .ZN(_10082_)
  );
  AND2_X1 _17747_ (
    .A1(_08650_),
    .A2(_08690_),
    .ZN(_10083_)
  );
  INV_X1 _17748_ (
    .A(_10083_),
    .ZN(_10084_)
  );
  MUX2_X1 _17749_ (
    .A(_08636_),
    .B(_08197_),
    .S(_08650_),
    .Z(_10085_)
  );
  MUX2_X1 _17750_ (
    .A(_08637_),
    .B(wb_reg_inst[8]),
    .S(_08650_),
    .Z(_10086_)
  );
  MUX2_X1 _17751_ (
    .A(_08635_),
    .B(wb_reg_inst[7]),
    .S(_08650_),
    .Z(_10087_)
  );
  MUX2_X1 _17752_ (
    .A(_08634_),
    .B(_08196_),
    .S(_08650_),
    .Z(_10088_)
  );
  AND2_X1 _17753_ (
    .A1(_10085_),
    .A2(_10088_),
    .ZN(_10089_)
  );
  MUX2_X1 _17754_ (
    .A(_08639_),
    .B(_08198_),
    .S(_08650_),
    .Z(_10090_)
  );
  MUX2_X1 _17755_ (
    .A(_08640_),
    .B(wb_reg_inst[9]),
    .S(_08650_),
    .Z(_10091_)
  );
  MUX2_X1 _17756_ (
    .A(_08644_),
    .B(_08200_),
    .S(_08650_),
    .Z(_10092_)
  );
  MUX2_X1 _17757_ (
    .A(_08645_),
    .B(wb_reg_inst[11]),
    .S(_08650_),
    .Z(_10093_)
  );
  MUX2_X1 _17758_ (
    .A(_08643_),
    .B(wb_reg_inst[10]),
    .S(_08650_),
    .Z(_10094_)
  );
  MUX2_X1 _17759_ (
    .A(_08642_),
    .B(_08199_),
    .S(_08650_),
    .Z(_10095_)
  );
  AND2_X1 _17760_ (
    .A1(_10092_),
    .A2(_10095_),
    .ZN(_10096_)
  );
  AND2_X1 _17761_ (
    .A1(_10090_),
    .A2(_10096_),
    .ZN(_10097_)
  );
  AND2_X1 _17762_ (
    .A1(_10089_),
    .A2(_10097_),
    .ZN(_10098_)
  );
  INV_X1 _17763_ (
    .A(_10098_),
    .ZN(_10099_)
  );
  AND2_X1 _17764_ (
    .A1(_10084_),
    .A2(_10099_),
    .ZN(_10100_)
  );
  AND2_X1 _17765_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_10092_),
    .ZN(_10101_)
  );
  INV_X1 _17766_ (
    .A(_10101_),
    .ZN(_10102_)
  );
  AND2_X1 _17767_ (
    .A1(_08571_),
    .A2(_10093_),
    .ZN(_10103_)
  );
  INV_X1 _17768_ (
    .A(_10103_),
    .ZN(_10104_)
  );
  AND2_X1 _17769_ (
    .A1(_10102_),
    .A2(_10104_),
    .ZN(_10105_)
  );
  AND2_X1 _17770_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_10090_),
    .ZN(_10106_)
  );
  INV_X1 _17771_ (
    .A(_10106_),
    .ZN(_10107_)
  );
  AND2_X1 _17772_ (
    .A1(_08542_),
    .A2(_10091_),
    .ZN(_10108_)
  );
  INV_X1 _17773_ (
    .A(_10108_),
    .ZN(_10109_)
  );
  AND2_X1 _17774_ (
    .A1(_10107_),
    .A2(_10109_),
    .ZN(_10110_)
  );
  AND2_X1 _17775_ (
    .A1(_10105_),
    .A2(_10110_),
    .ZN(_10111_)
  );
  AND2_X1 _17776_ (
    .A1(_08541_),
    .A2(_10086_),
    .ZN(_10112_)
  );
  INV_X1 _17777_ (
    .A(_10112_),
    .ZN(_10113_)
  );
  AND2_X1 _17778_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10085_),
    .ZN(_10114_)
  );
  INV_X1 _17779_ (
    .A(_10114_),
    .ZN(_10115_)
  );
  AND2_X1 _17780_ (
    .A1(_10113_),
    .A2(_10115_),
    .ZN(_10116_)
  );
  AND2_X1 _17781_ (
    .A1(_08543_),
    .A2(_10095_),
    .ZN(_10117_)
  );
  INV_X1 _17782_ (
    .A(_10117_),
    .ZN(_10118_)
  );
  AND2_X1 _17783_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_10094_),
    .ZN(_10119_)
  );
  INV_X1 _17784_ (
    .A(_10119_),
    .ZN(_10120_)
  );
  AND2_X1 _17785_ (
    .A1(_10118_),
    .A2(_10120_),
    .ZN(_10121_)
  );
  INV_X1 _17786_ (
    .A(_10121_),
    .ZN(_10122_)
  );
  AND2_X1 _17787_ (
    .A1(_08540_),
    .A2(_10087_),
    .ZN(_10123_)
  );
  INV_X1 _17788_ (
    .A(_10123_),
    .ZN(_10124_)
  );
  AND2_X1 _17789_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_10088_),
    .ZN(_10125_)
  );
  INV_X1 _17790_ (
    .A(_10125_),
    .ZN(_10126_)
  );
  AND2_X1 _17791_ (
    .A1(_10124_),
    .A2(_10126_),
    .ZN(_10127_)
  );
  AND2_X1 _17792_ (
    .A1(_10122_),
    .A2(_10127_),
    .ZN(_10128_)
  );
  AND2_X1 _17793_ (
    .A1(_10116_),
    .A2(_10128_),
    .ZN(_10129_)
  );
  AND2_X1 _17794_ (
    .A1(_10111_),
    .A2(_10129_),
    .ZN(_10130_)
  );
  AND2_X1 _17795_ (
    .A1(_10100_),
    .A2(_10130_),
    .ZN(_10131_)
  );
  INV_X1 _17796_ (
    .A(_10131_),
    .ZN(_10132_)
  );
  AND2_X1 _17797_ (
    .A1(_08188_),
    .A2(_08190_),
    .ZN(_10133_)
  );
  AND2_X1 _17798_ (
    .A1(_08192_),
    .A2(_10133_),
    .ZN(_10134_)
  );
  MUX2_X1 _17799_ (
    .A(csr_io_rw_rdata[2]),
    .B(wb_reg_wdata[2]),
    .S(_10134_),
    .Z(_10135_)
  );
  MUX2_X1 _17800_ (
    .A(div_io_resp_bits_data[2]),
    .B(_10135_),
    .S(_08649_),
    .Z(_10136_)
  );
  MUX2_X1 _17801_ (
    .A(_10136_),
    .B(io_dmem_resp_bits_data[2]),
    .S(_08631_),
    .Z(_10137_)
  );
  MUX2_X1 _17802_ (
    .A(\rf[23] [2]),
    .B(\rf[22] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_10138_)
  );
  INV_X1 _17803_ (
    .A(_10138_),
    .ZN(_10139_)
  );
  AND2_X1 _17804_ (
    .A1(_08542_),
    .A2(_10139_),
    .ZN(_10140_)
  );
  INV_X1 _17805_ (
    .A(_10140_),
    .ZN(_10141_)
  );
  MUX2_X1 _17806_ (
    .A(\rf[19] [2]),
    .B(\rf[18] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_10142_)
  );
  INV_X1 _17807_ (
    .A(_10142_),
    .ZN(_10143_)
  );
  AND2_X1 _17808_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_10143_),
    .ZN(_10144_)
  );
  INV_X1 _17809_ (
    .A(_10144_),
    .ZN(_10145_)
  );
  AND2_X1 _17810_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_10145_),
    .ZN(_10146_)
  );
  AND2_X1 _17811_ (
    .A1(_10141_),
    .A2(_10146_),
    .ZN(_10147_)
  );
  INV_X1 _17812_ (
    .A(_10147_),
    .ZN(_10148_)
  );
  AND2_X1 _17813_ (
    .A1(_08496_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10149_)
  );
  INV_X1 _17814_ (
    .A(_10149_),
    .ZN(_10150_)
  );
  AND2_X1 _17815_ (
    .A1(_08469_),
    .A2(_08542_),
    .ZN(_10151_)
  );
  INV_X1 _17816_ (
    .A(_10151_),
    .ZN(_10152_)
  );
  AND2_X1 _17817_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_10152_),
    .ZN(_10153_)
  );
  AND2_X1 _17818_ (
    .A1(_10150_),
    .A2(_10153_),
    .ZN(_10154_)
  );
  INV_X1 _17819_ (
    .A(_10154_),
    .ZN(_10155_)
  );
  AND2_X1 _17820_ (
    .A1(\rf[27] [2]),
    .A2(_09608_),
    .ZN(_10156_)
  );
  INV_X1 _17821_ (
    .A(_10156_),
    .ZN(_10157_)
  );
  AND2_X1 _17822_ (
    .A1(_10155_),
    .A2(_10157_),
    .ZN(_10158_)
  );
  INV_X1 _17823_ (
    .A(_10158_),
    .ZN(_10159_)
  );
  AND2_X1 _17824_ (
    .A1(_08543_),
    .A2(_10159_),
    .ZN(_10160_)
  );
  INV_X1 _17825_ (
    .A(_10160_),
    .ZN(_10161_)
  );
  AND2_X1 _17826_ (
    .A1(_08541_),
    .A2(_10161_),
    .ZN(_10162_)
  );
  AND2_X1 _17827_ (
    .A1(_10148_),
    .A2(_10162_),
    .ZN(_10163_)
  );
  INV_X1 _17828_ (
    .A(_10163_),
    .ZN(_10164_)
  );
  AND2_X1 _17829_ (
    .A1(\rf[20] [2]),
    .A2(_08542_),
    .ZN(_10165_)
  );
  INV_X1 _17830_ (
    .A(_10165_),
    .ZN(_10166_)
  );
  AND2_X1 _17831_ (
    .A1(\rf[16] [2]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10167_)
  );
  INV_X1 _17832_ (
    .A(_10167_),
    .ZN(_10168_)
  );
  AND2_X1 _17833_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_10168_),
    .ZN(_10169_)
  );
  AND2_X1 _17834_ (
    .A1(_10166_),
    .A2(_10169_),
    .ZN(_10170_)
  );
  INV_X1 _17835_ (
    .A(_10170_),
    .ZN(_10171_)
  );
  AND2_X1 _17836_ (
    .A1(\rf[21] [2]),
    .A2(_08542_),
    .ZN(_10172_)
  );
  INV_X1 _17837_ (
    .A(_10172_),
    .ZN(_10173_)
  );
  AND2_X1 _17838_ (
    .A1(\rf[17] [2]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10174_)
  );
  INV_X1 _17839_ (
    .A(_10174_),
    .ZN(_10175_)
  );
  AND2_X1 _17840_ (
    .A1(_08540_),
    .A2(_10175_),
    .ZN(_10176_)
  );
  AND2_X1 _17841_ (
    .A1(_10173_),
    .A2(_10176_),
    .ZN(_10177_)
  );
  INV_X1 _17842_ (
    .A(_10177_),
    .ZN(_10178_)
  );
  AND2_X1 _17843_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_10178_),
    .ZN(_10179_)
  );
  AND2_X1 _17844_ (
    .A1(_10171_),
    .A2(_10179_),
    .ZN(_10180_)
  );
  INV_X1 _17845_ (
    .A(_10180_),
    .ZN(_10181_)
  );
  AND2_X1 _17846_ (
    .A1(\rf[28] [2]),
    .A2(_08542_),
    .ZN(_10182_)
  );
  INV_X1 _17847_ (
    .A(_10182_),
    .ZN(_10183_)
  );
  AND2_X1 _17848_ (
    .A1(\rf[24] [2]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10184_)
  );
  INV_X1 _17849_ (
    .A(_10184_),
    .ZN(_10185_)
  );
  AND2_X1 _17850_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_10185_),
    .ZN(_10186_)
  );
  AND2_X1 _17851_ (
    .A1(_10183_),
    .A2(_10186_),
    .ZN(_10187_)
  );
  INV_X1 _17852_ (
    .A(_10187_),
    .ZN(_10188_)
  );
  AND2_X1 _17853_ (
    .A1(\rf[29] [2]),
    .A2(_08542_),
    .ZN(_10189_)
  );
  INV_X1 _17854_ (
    .A(_10189_),
    .ZN(_10190_)
  );
  AND2_X1 _17855_ (
    .A1(\rf[25] [2]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10191_)
  );
  INV_X1 _17856_ (
    .A(_10191_),
    .ZN(_10192_)
  );
  AND2_X1 _17857_ (
    .A1(_08540_),
    .A2(_10192_),
    .ZN(_10193_)
  );
  AND2_X1 _17858_ (
    .A1(_10190_),
    .A2(_10193_),
    .ZN(_10194_)
  );
  INV_X1 _17859_ (
    .A(_10194_),
    .ZN(_10195_)
  );
  AND2_X1 _17860_ (
    .A1(_08543_),
    .A2(_10195_),
    .ZN(_10196_)
  );
  AND2_X1 _17861_ (
    .A1(_10188_),
    .A2(_10196_),
    .ZN(_10197_)
  );
  INV_X1 _17862_ (
    .A(_10197_),
    .ZN(_10198_)
  );
  AND2_X1 _17863_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10198_),
    .ZN(_10199_)
  );
  AND2_X1 _17864_ (
    .A1(_10181_),
    .A2(_10199_),
    .ZN(_10200_)
  );
  INV_X1 _17865_ (
    .A(_10200_),
    .ZN(_10201_)
  );
  AND2_X1 _17866_ (
    .A1(_10164_),
    .A2(_10201_),
    .ZN(_10202_)
  );
  MUX2_X1 _17867_ (
    .A(\rf[1] [2]),
    .B(\rf[0] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_10203_)
  );
  MUX2_X1 _17868_ (
    .A(\rf[5] [2]),
    .B(\rf[4] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_10204_)
  );
  MUX2_X1 _17869_ (
    .A(_10203_),
    .B(_10204_),
    .S(_08542_),
    .Z(_10205_)
  );
  INV_X1 _17870_ (
    .A(_10205_),
    .ZN(_10206_)
  );
  AND2_X1 _17871_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_10206_),
    .ZN(_10207_)
  );
  INV_X1 _17872_ (
    .A(_10207_),
    .ZN(_10208_)
  );
  MUX2_X1 _17873_ (
    .A(\rf[13] [2]),
    .B(\rf[9] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10209_)
  );
  INV_X1 _17874_ (
    .A(_10209_),
    .ZN(_10210_)
  );
  AND2_X1 _17875_ (
    .A1(_09110_),
    .A2(_10210_),
    .ZN(_10211_)
  );
  INV_X1 _17876_ (
    .A(_10211_),
    .ZN(_10212_)
  );
  AND2_X1 _17877_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_08543_),
    .ZN(_10213_)
  );
  MUX2_X1 _17878_ (
    .A(\rf[12] [2]),
    .B(\rf[8] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10214_)
  );
  INV_X1 _17879_ (
    .A(_10214_),
    .ZN(_10215_)
  );
  AND2_X1 _17880_ (
    .A1(_10213_),
    .A2(_10215_),
    .ZN(_10216_)
  );
  INV_X1 _17881_ (
    .A(_10216_),
    .ZN(_10217_)
  );
  AND2_X1 _17882_ (
    .A1(_10212_),
    .A2(_10217_),
    .ZN(_10218_)
  );
  AND2_X1 _17883_ (
    .A1(_10208_),
    .A2(_10218_),
    .ZN(_10219_)
  );
  MUX2_X1 _17884_ (
    .A(\rf[3] [2]),
    .B(\rf[2] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_10220_)
  );
  MUX2_X1 _17885_ (
    .A(\rf[7] [2]),
    .B(\rf[6] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_10221_)
  );
  MUX2_X1 _17886_ (
    .A(_10220_),
    .B(_10221_),
    .S(_08542_),
    .Z(_10222_)
  );
  INV_X1 _17887_ (
    .A(_10222_),
    .ZN(_10223_)
  );
  AND2_X1 _17888_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_10223_),
    .ZN(_10224_)
  );
  INV_X1 _17889_ (
    .A(_10224_),
    .ZN(_10225_)
  );
  MUX2_X1 _17890_ (
    .A(\rf[14] [2]),
    .B(\rf[10] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10226_)
  );
  INV_X1 _17891_ (
    .A(_10226_),
    .ZN(_10227_)
  );
  AND2_X1 _17892_ (
    .A1(_10213_),
    .A2(_10227_),
    .ZN(_10228_)
  );
  INV_X1 _17893_ (
    .A(_10228_),
    .ZN(_10229_)
  );
  MUX2_X1 _17894_ (
    .A(\rf[15] [2]),
    .B(\rf[11] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10230_)
  );
  INV_X1 _17895_ (
    .A(_10230_),
    .ZN(_10231_)
  );
  AND2_X1 _17896_ (
    .A1(_09110_),
    .A2(_10231_),
    .ZN(_10232_)
  );
  INV_X1 _17897_ (
    .A(_10232_),
    .ZN(_10233_)
  );
  AND2_X1 _17898_ (
    .A1(_10229_),
    .A2(_10233_),
    .ZN(_10234_)
  );
  AND2_X1 _17899_ (
    .A1(_10225_),
    .A2(_10234_),
    .ZN(_10235_)
  );
  MUX2_X1 _17900_ (
    .A(_10219_),
    .B(_10235_),
    .S(_08541_),
    .Z(_10236_)
  );
  MUX2_X1 _17901_ (
    .A(_10202_),
    .B(_10236_),
    .S(ibuf_io_inst_0_bits_inst_rs1[4]),
    .Z(_10237_)
  );
  MUX2_X1 _17902_ (
    .A(_10137_),
    .B(_10237_),
    .S(_10132_),
    .Z(_10238_)
  );
  AND2_X1 _17903_ (
    .A1(_10082_),
    .A2(_10238_),
    .ZN(_10239_)
  );
  INV_X1 _17904_ (
    .A(_10239_),
    .ZN(_10240_)
  );
  AND2_X1 _17905_ (
    .A1(_10081_),
    .A2(_10240_),
    .ZN(_10241_)
  );
  INV_X1 _17906_ (
    .A(_10241_),
    .ZN(_10242_)
  );
  AND2_X1 _17907_ (
    .A1(_09298_),
    .A2(_10076_),
    .ZN(_10243_)
  );
  AND2_X1 _17908_ (
    .A1(ibuf_io_inst_0_ready),
    .A2(_10243_),
    .ZN(_10244_)
  );
  INV_X1 _17909_ (
    .A(_10244_),
    .ZN(_10245_)
  );
  MUX2_X1 _17910_ (
    .A(ex_reg_rs_msb_0[0]),
    .B(_10242_),
    .S(_10079_),
    .Z(_00067_)
  );
  AND2_X1 _17911_ (
    .A1(ibuf_io_inst_0_bits_raw[3]),
    .A2(_09295_),
    .ZN(_10246_)
  );
  INV_X1 _17912_ (
    .A(_10246_),
    .ZN(_10247_)
  );
  MUX2_X1 _17913_ (
    .A(csr_io_rw_rdata[3]),
    .B(wb_reg_wdata[3]),
    .S(_10134_),
    .Z(_10248_)
  );
  MUX2_X1 _17914_ (
    .A(div_io_resp_bits_data[3]),
    .B(_10248_),
    .S(_08649_),
    .Z(_10249_)
  );
  MUX2_X1 _17915_ (
    .A(_10249_),
    .B(io_dmem_resp_bits_data[3]),
    .S(_08631_),
    .Z(_10250_)
  );
  AND2_X1 _17916_ (
    .A1(\rf[2] [3]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10251_)
  );
  INV_X1 _17917_ (
    .A(_10251_),
    .ZN(_10252_)
  );
  AND2_X1 _17918_ (
    .A1(\rf[6] [3]),
    .A2(_08542_),
    .ZN(_10253_)
  );
  INV_X1 _17919_ (
    .A(_10253_),
    .ZN(_10254_)
  );
  AND2_X1 _17920_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_10254_),
    .ZN(_10255_)
  );
  AND2_X1 _17921_ (
    .A1(_10252_),
    .A2(_10255_),
    .ZN(_10256_)
  );
  INV_X1 _17922_ (
    .A(_10256_),
    .ZN(_10257_)
  );
  AND2_X1 _17923_ (
    .A1(\rf[3] [3]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10258_)
  );
  INV_X1 _17924_ (
    .A(_10258_),
    .ZN(_10259_)
  );
  AND2_X1 _17925_ (
    .A1(\rf[7] [3]),
    .A2(_08542_),
    .ZN(_10260_)
  );
  INV_X1 _17926_ (
    .A(_10260_),
    .ZN(_10261_)
  );
  AND2_X1 _17927_ (
    .A1(_08540_),
    .A2(_10261_),
    .ZN(_10262_)
  );
  AND2_X1 _17928_ (
    .A1(_10259_),
    .A2(_10262_),
    .ZN(_10263_)
  );
  INV_X1 _17929_ (
    .A(_10263_),
    .ZN(_10264_)
  );
  AND2_X1 _17930_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_10264_),
    .ZN(_10265_)
  );
  AND2_X1 _17931_ (
    .A1(_10257_),
    .A2(_10265_),
    .ZN(_10266_)
  );
  INV_X1 _17932_ (
    .A(_10266_),
    .ZN(_10267_)
  );
  MUX2_X1 _17933_ (
    .A(\rf[15] [3]),
    .B(\rf[11] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10268_)
  );
  INV_X1 _17934_ (
    .A(_10268_),
    .ZN(_10269_)
  );
  AND2_X1 _17935_ (
    .A1(_08540_),
    .A2(_10269_),
    .ZN(_10270_)
  );
  INV_X1 _17936_ (
    .A(_10270_),
    .ZN(_10271_)
  );
  MUX2_X1 _17937_ (
    .A(\rf[14] [3]),
    .B(\rf[10] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10272_)
  );
  INV_X1 _17938_ (
    .A(_10272_),
    .ZN(_10273_)
  );
  AND2_X1 _17939_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_10273_),
    .ZN(_10274_)
  );
  INV_X1 _17940_ (
    .A(_10274_),
    .ZN(_10275_)
  );
  AND2_X1 _17941_ (
    .A1(_08543_),
    .A2(_10275_),
    .ZN(_10276_)
  );
  AND2_X1 _17942_ (
    .A1(_10271_),
    .A2(_10276_),
    .ZN(_10277_)
  );
  INV_X1 _17943_ (
    .A(_10277_),
    .ZN(_10278_)
  );
  AND2_X1 _17944_ (
    .A1(_08541_),
    .A2(_10278_),
    .ZN(_10279_)
  );
  AND2_X1 _17945_ (
    .A1(_10267_),
    .A2(_10279_),
    .ZN(_10280_)
  );
  INV_X1 _17946_ (
    .A(_10280_),
    .ZN(_10281_)
  );
  AND2_X1 _17947_ (
    .A1(\rf[4] [3]),
    .A2(_08542_),
    .ZN(_10282_)
  );
  INV_X1 _17948_ (
    .A(_10282_),
    .ZN(_10283_)
  );
  AND2_X1 _17949_ (
    .A1(\rf[0] [3]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10284_)
  );
  INV_X1 _17950_ (
    .A(_10284_),
    .ZN(_10285_)
  );
  AND2_X1 _17951_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_10285_),
    .ZN(_10286_)
  );
  AND2_X1 _17952_ (
    .A1(_10283_),
    .A2(_10286_),
    .ZN(_10287_)
  );
  INV_X1 _17953_ (
    .A(_10287_),
    .ZN(_10288_)
  );
  AND2_X1 _17954_ (
    .A1(\rf[5] [3]),
    .A2(_08542_),
    .ZN(_10289_)
  );
  INV_X1 _17955_ (
    .A(_10289_),
    .ZN(_10290_)
  );
  AND2_X1 _17956_ (
    .A1(\rf[1] [3]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10291_)
  );
  INV_X1 _17957_ (
    .A(_10291_),
    .ZN(_10292_)
  );
  AND2_X1 _17958_ (
    .A1(_08540_),
    .A2(_10292_),
    .ZN(_10293_)
  );
  AND2_X1 _17959_ (
    .A1(_10290_),
    .A2(_10293_),
    .ZN(_10294_)
  );
  INV_X1 _17960_ (
    .A(_10294_),
    .ZN(_10295_)
  );
  AND2_X1 _17961_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_10295_),
    .ZN(_10296_)
  );
  AND2_X1 _17962_ (
    .A1(_10288_),
    .A2(_10296_),
    .ZN(_10297_)
  );
  INV_X1 _17963_ (
    .A(_10297_),
    .ZN(_10298_)
  );
  MUX2_X1 _17964_ (
    .A(\rf[13] [3]),
    .B(\rf[9] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10299_)
  );
  INV_X1 _17965_ (
    .A(_10299_),
    .ZN(_10300_)
  );
  AND2_X1 _17966_ (
    .A1(_08540_),
    .A2(_10300_),
    .ZN(_10301_)
  );
  INV_X1 _17967_ (
    .A(_10301_),
    .ZN(_10302_)
  );
  MUX2_X1 _17968_ (
    .A(\rf[12] [3]),
    .B(\rf[8] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10303_)
  );
  INV_X1 _17969_ (
    .A(_10303_),
    .ZN(_10304_)
  );
  AND2_X1 _17970_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_10304_),
    .ZN(_10305_)
  );
  INV_X1 _17971_ (
    .A(_10305_),
    .ZN(_10306_)
  );
  AND2_X1 _17972_ (
    .A1(_08543_),
    .A2(_10306_),
    .ZN(_10307_)
  );
  AND2_X1 _17973_ (
    .A1(_10302_),
    .A2(_10307_),
    .ZN(_10308_)
  );
  INV_X1 _17974_ (
    .A(_10308_),
    .ZN(_10309_)
  );
  AND2_X1 _17975_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10309_),
    .ZN(_10310_)
  );
  AND2_X1 _17976_ (
    .A1(_10298_),
    .A2(_10310_),
    .ZN(_10311_)
  );
  INV_X1 _17977_ (
    .A(_10311_),
    .ZN(_10312_)
  );
  AND2_X1 _17978_ (
    .A1(_10281_),
    .A2(_10312_),
    .ZN(_10313_)
  );
  AND2_X1 _17979_ (
    .A1(\rf[22] [3]),
    .A2(_08542_),
    .ZN(_10314_)
  );
  INV_X1 _17980_ (
    .A(_10314_),
    .ZN(_10315_)
  );
  AND2_X1 _17981_ (
    .A1(\rf[18] [3]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10316_)
  );
  INV_X1 _17982_ (
    .A(_10316_),
    .ZN(_10317_)
  );
  AND2_X1 _17983_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_10317_),
    .ZN(_10318_)
  );
  AND2_X1 _17984_ (
    .A1(_10315_),
    .A2(_10318_),
    .ZN(_10319_)
  );
  INV_X1 _17985_ (
    .A(_10319_),
    .ZN(_10320_)
  );
  AND2_X1 _17986_ (
    .A1(\rf[23] [3]),
    .A2(_08542_),
    .ZN(_10321_)
  );
  INV_X1 _17987_ (
    .A(_10321_),
    .ZN(_10322_)
  );
  AND2_X1 _17988_ (
    .A1(\rf[19] [3]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10323_)
  );
  INV_X1 _17989_ (
    .A(_10323_),
    .ZN(_10324_)
  );
  AND2_X1 _17990_ (
    .A1(_08540_),
    .A2(_10324_),
    .ZN(_10325_)
  );
  AND2_X1 _17991_ (
    .A1(_10322_),
    .A2(_10325_),
    .ZN(_10326_)
  );
  INV_X1 _17992_ (
    .A(_10326_),
    .ZN(_10327_)
  );
  AND2_X1 _17993_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_10327_),
    .ZN(_10328_)
  );
  AND2_X1 _17994_ (
    .A1(_10320_),
    .A2(_10328_),
    .ZN(_10329_)
  );
  INV_X1 _17995_ (
    .A(_10329_),
    .ZN(_10330_)
  );
  AND2_X1 _17996_ (
    .A1(_08497_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10331_)
  );
  INV_X1 _17997_ (
    .A(_10331_),
    .ZN(_10332_)
  );
  AND2_X1 _17998_ (
    .A1(_08470_),
    .A2(_08542_),
    .ZN(_10333_)
  );
  INV_X1 _17999_ (
    .A(_10333_),
    .ZN(_10334_)
  );
  AND2_X1 _18000_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_10334_),
    .ZN(_10335_)
  );
  AND2_X1 _18001_ (
    .A1(_10332_),
    .A2(_10335_),
    .ZN(_10336_)
  );
  INV_X1 _18002_ (
    .A(_10336_),
    .ZN(_10337_)
  );
  AND2_X1 _18003_ (
    .A1(\rf[27] [3]),
    .A2(_09608_),
    .ZN(_10338_)
  );
  INV_X1 _18004_ (
    .A(_10338_),
    .ZN(_10339_)
  );
  AND2_X1 _18005_ (
    .A1(_10337_),
    .A2(_10339_),
    .ZN(_10340_)
  );
  INV_X1 _18006_ (
    .A(_10340_),
    .ZN(_10341_)
  );
  AND2_X1 _18007_ (
    .A1(_08543_),
    .A2(_10341_),
    .ZN(_10342_)
  );
  INV_X1 _18008_ (
    .A(_10342_),
    .ZN(_10343_)
  );
  AND2_X1 _18009_ (
    .A1(_08541_),
    .A2(_10343_),
    .ZN(_10344_)
  );
  AND2_X1 _18010_ (
    .A1(_10330_),
    .A2(_10344_),
    .ZN(_10345_)
  );
  INV_X1 _18011_ (
    .A(_10345_),
    .ZN(_10346_)
  );
  MUX2_X1 _18012_ (
    .A(\rf[29] [3]),
    .B(\rf[28] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_10347_)
  );
  INV_X1 _18013_ (
    .A(_10347_),
    .ZN(_10348_)
  );
  AND2_X1 _18014_ (
    .A1(_08542_),
    .A2(_10348_),
    .ZN(_10349_)
  );
  INV_X1 _18015_ (
    .A(_10349_),
    .ZN(_10350_)
  );
  MUX2_X1 _18016_ (
    .A(\rf[25] [3]),
    .B(\rf[24] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_10351_)
  );
  INV_X1 _18017_ (
    .A(_10351_),
    .ZN(_10352_)
  );
  AND2_X1 _18018_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_10352_),
    .ZN(_10353_)
  );
  INV_X1 _18019_ (
    .A(_10353_),
    .ZN(_10354_)
  );
  AND2_X1 _18020_ (
    .A1(_08543_),
    .A2(_10354_),
    .ZN(_10355_)
  );
  AND2_X1 _18021_ (
    .A1(_10350_),
    .A2(_10355_),
    .ZN(_10356_)
  );
  INV_X1 _18022_ (
    .A(_10356_),
    .ZN(_10357_)
  );
  AND2_X1 _18023_ (
    .A1(\rf[20] [3]),
    .A2(_08542_),
    .ZN(_10358_)
  );
  INV_X1 _18024_ (
    .A(_10358_),
    .ZN(_10359_)
  );
  AND2_X1 _18025_ (
    .A1(\rf[16] [3]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10360_)
  );
  INV_X1 _18026_ (
    .A(_10360_),
    .ZN(_10361_)
  );
  AND2_X1 _18027_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_10361_),
    .ZN(_10362_)
  );
  AND2_X1 _18028_ (
    .A1(_10359_),
    .A2(_10362_),
    .ZN(_10363_)
  );
  INV_X1 _18029_ (
    .A(_10363_),
    .ZN(_10364_)
  );
  AND2_X1 _18030_ (
    .A1(\rf[21] [3]),
    .A2(_08542_),
    .ZN(_10365_)
  );
  INV_X1 _18031_ (
    .A(_10365_),
    .ZN(_10366_)
  );
  AND2_X1 _18032_ (
    .A1(\rf[17] [3]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10367_)
  );
  INV_X1 _18033_ (
    .A(_10367_),
    .ZN(_10368_)
  );
  AND2_X1 _18034_ (
    .A1(_08540_),
    .A2(_10368_),
    .ZN(_10369_)
  );
  AND2_X1 _18035_ (
    .A1(_10366_),
    .A2(_10369_),
    .ZN(_10370_)
  );
  INV_X1 _18036_ (
    .A(_10370_),
    .ZN(_10371_)
  );
  AND2_X1 _18037_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_10371_),
    .ZN(_10372_)
  );
  AND2_X1 _18038_ (
    .A1(_10364_),
    .A2(_10372_),
    .ZN(_10373_)
  );
  INV_X1 _18039_ (
    .A(_10373_),
    .ZN(_10374_)
  );
  AND2_X1 _18040_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10374_),
    .ZN(_10375_)
  );
  AND2_X1 _18041_ (
    .A1(_10357_),
    .A2(_10375_),
    .ZN(_10376_)
  );
  INV_X1 _18042_ (
    .A(_10376_),
    .ZN(_10377_)
  );
  AND2_X1 _18043_ (
    .A1(_10346_),
    .A2(_10377_),
    .ZN(_10378_)
  );
  MUX2_X1 _18044_ (
    .A(_10313_),
    .B(_10378_),
    .S(_08571_),
    .Z(_10379_)
  );
  MUX2_X1 _18045_ (
    .A(_10250_),
    .B(_10379_),
    .S(_10132_),
    .Z(_10380_)
  );
  AND2_X1 _18046_ (
    .A1(_10082_),
    .A2(_10380_),
    .ZN(_10381_)
  );
  INV_X1 _18047_ (
    .A(_10381_),
    .ZN(_10382_)
  );
  AND2_X1 _18048_ (
    .A1(_10247_),
    .A2(_10382_),
    .ZN(_10383_)
  );
  INV_X1 _18049_ (
    .A(_10383_),
    .ZN(_10384_)
  );
  MUX2_X1 _18050_ (
    .A(ex_reg_rs_msb_0[1]),
    .B(_10384_),
    .S(_10079_),
    .Z(_00068_)
  );
  AND2_X1 _18051_ (
    .A1(ibuf_io_inst_0_bits_raw[4]),
    .A2(_09295_),
    .ZN(_10385_)
  );
  INV_X1 _18052_ (
    .A(_10385_),
    .ZN(_10386_)
  );
  MUX2_X1 _18053_ (
    .A(csr_io_rw_rdata[4]),
    .B(wb_reg_wdata[4]),
    .S(_10134_),
    .Z(_10387_)
  );
  MUX2_X1 _18054_ (
    .A(div_io_resp_bits_data[4]),
    .B(_10387_),
    .S(_08649_),
    .Z(_10388_)
  );
  MUX2_X1 _18055_ (
    .A(_10388_),
    .B(io_dmem_resp_bits_data[4]),
    .S(_08631_),
    .Z(_10389_)
  );
  MUX2_X1 _18056_ (
    .A(\rf[3] [4]),
    .B(\rf[1] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_10390_)
  );
  MUX2_X1 _18057_ (
    .A(\rf[7] [4]),
    .B(\rf[5] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_10391_)
  );
  MUX2_X1 _18058_ (
    .A(_10390_),
    .B(_10391_),
    .S(_08542_),
    .Z(_10392_)
  );
  AND2_X1 _18059_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_10392_),
    .ZN(_10393_)
  );
  INV_X1 _18060_ (
    .A(_10393_),
    .ZN(_10394_)
  );
  MUX2_X1 _18061_ (
    .A(\rf[13] [4]),
    .B(\rf[9] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10395_)
  );
  INV_X1 _18062_ (
    .A(_10395_),
    .ZN(_10396_)
  );
  AND2_X1 _18063_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10396_),
    .ZN(_10397_)
  );
  INV_X1 _18064_ (
    .A(_10397_),
    .ZN(_10398_)
  );
  MUX2_X1 _18065_ (
    .A(\rf[15] [4]),
    .B(\rf[11] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10399_)
  );
  INV_X1 _18066_ (
    .A(_10399_),
    .ZN(_10400_)
  );
  AND2_X1 _18067_ (
    .A1(_08541_),
    .A2(_10400_),
    .ZN(_10401_)
  );
  INV_X1 _18068_ (
    .A(_10401_),
    .ZN(_10402_)
  );
  AND2_X1 _18069_ (
    .A1(_08543_),
    .A2(_10402_),
    .ZN(_10403_)
  );
  AND2_X1 _18070_ (
    .A1(_10398_),
    .A2(_10403_),
    .ZN(_10404_)
  );
  INV_X1 _18071_ (
    .A(_10404_),
    .ZN(_10405_)
  );
  AND2_X1 _18072_ (
    .A1(_08540_),
    .A2(_10405_),
    .ZN(_10406_)
  );
  AND2_X1 _18073_ (
    .A1(_10394_),
    .A2(_10406_),
    .ZN(_10407_)
  );
  INV_X1 _18074_ (
    .A(_10407_),
    .ZN(_10408_)
  );
  MUX2_X1 _18075_ (
    .A(\rf[2] [4]),
    .B(\rf[0] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_10409_)
  );
  MUX2_X1 _18076_ (
    .A(\rf[6] [4]),
    .B(\rf[4] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_10410_)
  );
  MUX2_X1 _18077_ (
    .A(_10409_),
    .B(_10410_),
    .S(_08542_),
    .Z(_10411_)
  );
  AND2_X1 _18078_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_10411_),
    .ZN(_10412_)
  );
  INV_X1 _18079_ (
    .A(_10412_),
    .ZN(_10413_)
  );
  MUX2_X1 _18080_ (
    .A(\rf[12] [4]),
    .B(\rf[8] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10414_)
  );
  INV_X1 _18081_ (
    .A(_10414_),
    .ZN(_10415_)
  );
  AND2_X1 _18082_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10415_),
    .ZN(_10416_)
  );
  INV_X1 _18083_ (
    .A(_10416_),
    .ZN(_10417_)
  );
  MUX2_X1 _18084_ (
    .A(\rf[14] [4]),
    .B(\rf[10] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10418_)
  );
  INV_X1 _18085_ (
    .A(_10418_),
    .ZN(_10419_)
  );
  AND2_X1 _18086_ (
    .A1(_08541_),
    .A2(_10419_),
    .ZN(_10420_)
  );
  INV_X1 _18087_ (
    .A(_10420_),
    .ZN(_10421_)
  );
  AND2_X1 _18088_ (
    .A1(_08543_),
    .A2(_10421_),
    .ZN(_10422_)
  );
  AND2_X1 _18089_ (
    .A1(_10417_),
    .A2(_10422_),
    .ZN(_10423_)
  );
  INV_X1 _18090_ (
    .A(_10423_),
    .ZN(_10424_)
  );
  AND2_X1 _18091_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_10424_),
    .ZN(_10425_)
  );
  AND2_X1 _18092_ (
    .A1(_10413_),
    .A2(_10425_),
    .ZN(_10426_)
  );
  INV_X1 _18093_ (
    .A(_10426_),
    .ZN(_10427_)
  );
  AND2_X1 _18094_ (
    .A1(_10408_),
    .A2(_10427_),
    .ZN(_10428_)
  );
  AND2_X1 _18095_ (
    .A1(\rf[21] [4]),
    .A2(_08542_),
    .ZN(_10429_)
  );
  INV_X1 _18096_ (
    .A(_10429_),
    .ZN(_10430_)
  );
  AND2_X1 _18097_ (
    .A1(\rf[17] [4]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10431_)
  );
  INV_X1 _18098_ (
    .A(_10431_),
    .ZN(_10432_)
  );
  AND2_X1 _18099_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10432_),
    .ZN(_10433_)
  );
  AND2_X1 _18100_ (
    .A1(_10430_),
    .A2(_10433_),
    .ZN(_10434_)
  );
  INV_X1 _18101_ (
    .A(_10434_),
    .ZN(_10435_)
  );
  AND2_X1 _18102_ (
    .A1(\rf[19] [4]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10436_)
  );
  INV_X1 _18103_ (
    .A(_10436_),
    .ZN(_10437_)
  );
  AND2_X1 _18104_ (
    .A1(\rf[23] [4]),
    .A2(_08542_),
    .ZN(_10438_)
  );
  INV_X1 _18105_ (
    .A(_10438_),
    .ZN(_10439_)
  );
  AND2_X1 _18106_ (
    .A1(_08541_),
    .A2(_10439_),
    .ZN(_10440_)
  );
  AND2_X1 _18107_ (
    .A1(_10437_),
    .A2(_10440_),
    .ZN(_10441_)
  );
  INV_X1 _18108_ (
    .A(_10441_),
    .ZN(_10442_)
  );
  AND2_X1 _18109_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_10442_),
    .ZN(_10443_)
  );
  AND2_X1 _18110_ (
    .A1(_10435_),
    .A2(_10443_),
    .ZN(_10444_)
  );
  INV_X1 _18111_ (
    .A(_10444_),
    .ZN(_10445_)
  );
  AND2_X1 _18112_ (
    .A1(_08236_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10446_)
  );
  INV_X1 _18113_ (
    .A(_10446_),
    .ZN(_10447_)
  );
  AND2_X1 _18114_ (
    .A1(_08459_),
    .A2(_08542_),
    .ZN(_10448_)
  );
  INV_X1 _18115_ (
    .A(_10448_),
    .ZN(_10449_)
  );
  AND2_X1 _18116_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10449_),
    .ZN(_10450_)
  );
  AND2_X1 _18117_ (
    .A1(_10447_),
    .A2(_10450_),
    .ZN(_10451_)
  );
  INV_X1 _18118_ (
    .A(_10451_),
    .ZN(_10452_)
  );
  AND2_X1 _18119_ (
    .A1(_08541_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10453_)
  );
  AND2_X1 _18120_ (
    .A1(\rf[27] [4]),
    .A2(_10453_),
    .ZN(_10454_)
  );
  INV_X1 _18121_ (
    .A(_10454_),
    .ZN(_10455_)
  );
  AND2_X1 _18122_ (
    .A1(_10452_),
    .A2(_10455_),
    .ZN(_10456_)
  );
  INV_X1 _18123_ (
    .A(_10456_),
    .ZN(_10457_)
  );
  AND2_X1 _18124_ (
    .A1(_08543_),
    .A2(_10457_),
    .ZN(_10458_)
  );
  INV_X1 _18125_ (
    .A(_10458_),
    .ZN(_10459_)
  );
  AND2_X1 _18126_ (
    .A1(_08540_),
    .A2(_10459_),
    .ZN(_10460_)
  );
  AND2_X1 _18127_ (
    .A1(_10445_),
    .A2(_10460_),
    .ZN(_10461_)
  );
  INV_X1 _18128_ (
    .A(_10461_),
    .ZN(_10462_)
  );
  MUX2_X1 _18129_ (
    .A(\rf[30] [4]),
    .B(\rf[26] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10463_)
  );
  INV_X1 _18130_ (
    .A(_10463_),
    .ZN(_10464_)
  );
  AND2_X1 _18131_ (
    .A1(_08541_),
    .A2(_10464_),
    .ZN(_10465_)
  );
  INV_X1 _18132_ (
    .A(_10465_),
    .ZN(_10466_)
  );
  MUX2_X1 _18133_ (
    .A(\rf[28] [4]),
    .B(\rf[24] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10467_)
  );
  INV_X1 _18134_ (
    .A(_10467_),
    .ZN(_10468_)
  );
  AND2_X1 _18135_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10468_),
    .ZN(_10469_)
  );
  INV_X1 _18136_ (
    .A(_10469_),
    .ZN(_10470_)
  );
  AND2_X1 _18137_ (
    .A1(_08543_),
    .A2(_10470_),
    .ZN(_10471_)
  );
  AND2_X1 _18138_ (
    .A1(_10466_),
    .A2(_10471_),
    .ZN(_10472_)
  );
  INV_X1 _18139_ (
    .A(_10472_),
    .ZN(_10473_)
  );
  AND2_X1 _18140_ (
    .A1(\rf[16] [4]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10474_)
  );
  INV_X1 _18141_ (
    .A(_10474_),
    .ZN(_10475_)
  );
  AND2_X1 _18142_ (
    .A1(\rf[20] [4]),
    .A2(_08542_),
    .ZN(_10476_)
  );
  INV_X1 _18143_ (
    .A(_10476_),
    .ZN(_10477_)
  );
  AND2_X1 _18144_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10477_),
    .ZN(_10478_)
  );
  AND2_X1 _18145_ (
    .A1(_10475_),
    .A2(_10478_),
    .ZN(_10479_)
  );
  INV_X1 _18146_ (
    .A(_10479_),
    .ZN(_10480_)
  );
  AND2_X1 _18147_ (
    .A1(\rf[18] [4]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10481_)
  );
  INV_X1 _18148_ (
    .A(_10481_),
    .ZN(_10482_)
  );
  AND2_X1 _18149_ (
    .A1(\rf[22] [4]),
    .A2(_08542_),
    .ZN(_10483_)
  );
  INV_X1 _18150_ (
    .A(_10483_),
    .ZN(_10484_)
  );
  AND2_X1 _18151_ (
    .A1(_08541_),
    .A2(_10484_),
    .ZN(_10485_)
  );
  AND2_X1 _18152_ (
    .A1(_10482_),
    .A2(_10485_),
    .ZN(_10486_)
  );
  INV_X1 _18153_ (
    .A(_10486_),
    .ZN(_10487_)
  );
  AND2_X1 _18154_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_10487_),
    .ZN(_10488_)
  );
  AND2_X1 _18155_ (
    .A1(_10480_),
    .A2(_10488_),
    .ZN(_10489_)
  );
  INV_X1 _18156_ (
    .A(_10489_),
    .ZN(_10490_)
  );
  AND2_X1 _18157_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_10490_),
    .ZN(_10491_)
  );
  AND2_X1 _18158_ (
    .A1(_10473_),
    .A2(_10491_),
    .ZN(_10492_)
  );
  INV_X1 _18159_ (
    .A(_10492_),
    .ZN(_10493_)
  );
  AND2_X1 _18160_ (
    .A1(_10462_),
    .A2(_10493_),
    .ZN(_10494_)
  );
  MUX2_X1 _18161_ (
    .A(_10428_),
    .B(_10494_),
    .S(_08571_),
    .Z(_10495_)
  );
  MUX2_X1 _18162_ (
    .A(_10389_),
    .B(_10495_),
    .S(_10132_),
    .Z(_10496_)
  );
  AND2_X1 _18163_ (
    .A1(_10082_),
    .A2(_10496_),
    .ZN(_10497_)
  );
  INV_X1 _18164_ (
    .A(_10497_),
    .ZN(_10498_)
  );
  AND2_X1 _18165_ (
    .A1(_10386_),
    .A2(_10498_),
    .ZN(_10499_)
  );
  INV_X1 _18166_ (
    .A(_10499_),
    .ZN(_10500_)
  );
  MUX2_X1 _18167_ (
    .A(ex_reg_rs_msb_0[2]),
    .B(_10500_),
    .S(_10079_),
    .Z(_00069_)
  );
  AND2_X1 _18168_ (
    .A1(ibuf_io_inst_0_bits_raw[5]),
    .A2(_09295_),
    .ZN(_10501_)
  );
  INV_X1 _18169_ (
    .A(_10501_),
    .ZN(_10502_)
  );
  MUX2_X1 _18170_ (
    .A(csr_io_rw_rdata[5]),
    .B(wb_reg_wdata[5]),
    .S(_10134_),
    .Z(_10503_)
  );
  MUX2_X1 _18171_ (
    .A(div_io_resp_bits_data[5]),
    .B(_10503_),
    .S(_08649_),
    .Z(_10504_)
  );
  MUX2_X1 _18172_ (
    .A(_10504_),
    .B(io_dmem_resp_bits_data[5]),
    .S(_08631_),
    .Z(_10505_)
  );
  MUX2_X1 _18173_ (
    .A(\rf[5] [5]),
    .B(\rf[1] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10506_)
  );
  MUX2_X1 _18174_ (
    .A(\rf[7] [5]),
    .B(\rf[3] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10507_)
  );
  MUX2_X1 _18175_ (
    .A(_10506_),
    .B(_10507_),
    .S(_08541_),
    .Z(_10508_)
  );
  AND2_X1 _18176_ (
    .A1(_08540_),
    .A2(_10508_),
    .ZN(_10509_)
  );
  INV_X1 _18177_ (
    .A(_10509_),
    .ZN(_10510_)
  );
  MUX2_X1 _18178_ (
    .A(\rf[4] [5]),
    .B(\rf[0] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10511_)
  );
  MUX2_X1 _18179_ (
    .A(\rf[6] [5]),
    .B(\rf[2] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10512_)
  );
  MUX2_X1 _18180_ (
    .A(_10511_),
    .B(_10512_),
    .S(_08541_),
    .Z(_10513_)
  );
  AND2_X1 _18181_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_10513_),
    .ZN(_10514_)
  );
  INV_X1 _18182_ (
    .A(_10514_),
    .ZN(_10515_)
  );
  AND2_X1 _18183_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_10515_),
    .ZN(_10516_)
  );
  AND2_X1 _18184_ (
    .A1(_10510_),
    .A2(_10516_),
    .ZN(_10517_)
  );
  INV_X1 _18185_ (
    .A(_10517_),
    .ZN(_10518_)
  );
  AND2_X1 _18186_ (
    .A1(_08378_),
    .A2(_08542_),
    .ZN(_10519_)
  );
  INV_X1 _18187_ (
    .A(_10519_),
    .ZN(_10520_)
  );
  AND2_X1 _18188_ (
    .A1(_08279_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10521_)
  );
  INV_X1 _18189_ (
    .A(_10521_),
    .ZN(_10522_)
  );
  AND2_X1 _18190_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10522_),
    .ZN(_10523_)
  );
  AND2_X1 _18191_ (
    .A1(_10520_),
    .A2(_10523_),
    .ZN(_10524_)
  );
  INV_X1 _18192_ (
    .A(_10524_),
    .ZN(_10525_)
  );
  MUX2_X1 _18193_ (
    .A(\rf[22] [5]),
    .B(\rf[18] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10526_)
  );
  AND2_X1 _18194_ (
    .A1(_08541_),
    .A2(_10526_),
    .ZN(_10527_)
  );
  INV_X1 _18195_ (
    .A(_10527_),
    .ZN(_10528_)
  );
  AND2_X1 _18196_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_10528_),
    .ZN(_10529_)
  );
  AND2_X1 _18197_ (
    .A1(_10525_),
    .A2(_10529_),
    .ZN(_10530_)
  );
  INV_X1 _18198_ (
    .A(_10530_),
    .ZN(_10531_)
  );
  AND2_X1 _18199_ (
    .A1(_08309_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10532_)
  );
  INV_X1 _18200_ (
    .A(_10532_),
    .ZN(_10533_)
  );
  AND2_X1 _18201_ (
    .A1(_08408_),
    .A2(_08542_),
    .ZN(_10534_)
  );
  INV_X1 _18202_ (
    .A(_10534_),
    .ZN(_10535_)
  );
  AND2_X1 _18203_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10535_),
    .ZN(_10536_)
  );
  AND2_X1 _18204_ (
    .A1(_10533_),
    .A2(_10536_),
    .ZN(_10537_)
  );
  INV_X1 _18205_ (
    .A(_10537_),
    .ZN(_10538_)
  );
  MUX2_X1 _18206_ (
    .A(\rf[23] [5]),
    .B(\rf[19] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10539_)
  );
  AND2_X1 _18207_ (
    .A1(_08541_),
    .A2(_10539_),
    .ZN(_10540_)
  );
  INV_X1 _18208_ (
    .A(_10540_),
    .ZN(_10541_)
  );
  AND2_X1 _18209_ (
    .A1(_08540_),
    .A2(_10541_),
    .ZN(_10542_)
  );
  AND2_X1 _18210_ (
    .A1(_10538_),
    .A2(_10542_),
    .ZN(_10543_)
  );
  INV_X1 _18211_ (
    .A(_10543_),
    .ZN(_10544_)
  );
  AND2_X1 _18212_ (
    .A1(_10531_),
    .A2(_10544_),
    .ZN(_10545_)
  );
  INV_X1 _18213_ (
    .A(_10545_),
    .ZN(_10546_)
  );
  AND2_X1 _18214_ (
    .A1(_08571_),
    .A2(_10546_),
    .ZN(_10547_)
  );
  INV_X1 _18215_ (
    .A(_10547_),
    .ZN(_10548_)
  );
  AND2_X1 _18216_ (
    .A1(_10518_),
    .A2(_10548_),
    .ZN(_10549_)
  );
  AND2_X1 _18217_ (
    .A1(\rf[10] [5]),
    .A2(_08541_),
    .ZN(_10550_)
  );
  INV_X1 _18218_ (
    .A(_10550_),
    .ZN(_10551_)
  );
  AND2_X1 _18219_ (
    .A1(\rf[8] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_10552_)
  );
  INV_X1 _18220_ (
    .A(_10552_),
    .ZN(_10553_)
  );
  AND2_X1 _18221_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_10553_),
    .ZN(_10554_)
  );
  AND2_X1 _18222_ (
    .A1(_10551_),
    .A2(_10554_),
    .ZN(_10555_)
  );
  INV_X1 _18223_ (
    .A(_10555_),
    .ZN(_10556_)
  );
  AND2_X1 _18224_ (
    .A1(\rf[14] [5]),
    .A2(_08541_),
    .ZN(_10557_)
  );
  INV_X1 _18225_ (
    .A(_10557_),
    .ZN(_10558_)
  );
  AND2_X1 _18226_ (
    .A1(\rf[12] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_10559_)
  );
  INV_X1 _18227_ (
    .A(_10559_),
    .ZN(_10560_)
  );
  AND2_X1 _18228_ (
    .A1(_08542_),
    .A2(_10560_),
    .ZN(_10561_)
  );
  AND2_X1 _18229_ (
    .A1(_10558_),
    .A2(_10561_),
    .ZN(_10562_)
  );
  INV_X1 _18230_ (
    .A(_10562_),
    .ZN(_10563_)
  );
  AND2_X1 _18231_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_10563_),
    .ZN(_10564_)
  );
  AND2_X1 _18232_ (
    .A1(_10556_),
    .A2(_10564_),
    .ZN(_10565_)
  );
  INV_X1 _18233_ (
    .A(_10565_),
    .ZN(_10566_)
  );
  AND2_X1 _18234_ (
    .A1(\rf[11] [5]),
    .A2(_08541_),
    .ZN(_10567_)
  );
  INV_X1 _18235_ (
    .A(_10567_),
    .ZN(_10568_)
  );
  AND2_X1 _18236_ (
    .A1(\rf[9] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_10569_)
  );
  INV_X1 _18237_ (
    .A(_10569_),
    .ZN(_10570_)
  );
  AND2_X1 _18238_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_10570_),
    .ZN(_10571_)
  );
  AND2_X1 _18239_ (
    .A1(_10568_),
    .A2(_10571_),
    .ZN(_10572_)
  );
  INV_X1 _18240_ (
    .A(_10572_),
    .ZN(_10573_)
  );
  AND2_X1 _18241_ (
    .A1(\rf[15] [5]),
    .A2(_08541_),
    .ZN(_10574_)
  );
  INV_X1 _18242_ (
    .A(_10574_),
    .ZN(_10575_)
  );
  AND2_X1 _18243_ (
    .A1(\rf[13] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_10576_)
  );
  INV_X1 _18244_ (
    .A(_10576_),
    .ZN(_10577_)
  );
  AND2_X1 _18245_ (
    .A1(_08542_),
    .A2(_10577_),
    .ZN(_10578_)
  );
  AND2_X1 _18246_ (
    .A1(_10575_),
    .A2(_10578_),
    .ZN(_10579_)
  );
  INV_X1 _18247_ (
    .A(_10579_),
    .ZN(_10580_)
  );
  AND2_X1 _18248_ (
    .A1(_08540_),
    .A2(_10580_),
    .ZN(_10581_)
  );
  AND2_X1 _18249_ (
    .A1(_10573_),
    .A2(_10581_),
    .ZN(_10582_)
  );
  INV_X1 _18250_ (
    .A(_10582_),
    .ZN(_10583_)
  );
  AND2_X1 _18251_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_10583_),
    .ZN(_10584_)
  );
  AND2_X1 _18252_ (
    .A1(_10566_),
    .A2(_10584_),
    .ZN(_10585_)
  );
  INV_X1 _18253_ (
    .A(_10585_),
    .ZN(_10586_)
  );
  AND2_X1 _18254_ (
    .A1(\rf[30] [5]),
    .A2(_08542_),
    .ZN(_10587_)
  );
  INV_X1 _18255_ (
    .A(_10587_),
    .ZN(_10588_)
  );
  AND2_X1 _18256_ (
    .A1(\rf[26] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10589_)
  );
  INV_X1 _18257_ (
    .A(_10589_),
    .ZN(_10590_)
  );
  AND2_X1 _18258_ (
    .A1(_08541_),
    .A2(_10590_),
    .ZN(_10591_)
  );
  AND2_X1 _18259_ (
    .A1(_10588_),
    .A2(_10591_),
    .ZN(_10592_)
  );
  INV_X1 _18260_ (
    .A(_10592_),
    .ZN(_10593_)
  );
  AND2_X1 _18261_ (
    .A1(\rf[24] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10594_)
  );
  INV_X1 _18262_ (
    .A(_10594_),
    .ZN(_10595_)
  );
  AND2_X1 _18263_ (
    .A1(\rf[28] [5]),
    .A2(_08542_),
    .ZN(_10596_)
  );
  INV_X1 _18264_ (
    .A(_10596_),
    .ZN(_10597_)
  );
  AND2_X1 _18265_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10597_),
    .ZN(_10598_)
  );
  AND2_X1 _18266_ (
    .A1(_10595_),
    .A2(_10598_),
    .ZN(_10599_)
  );
  INV_X1 _18267_ (
    .A(_10599_),
    .ZN(_10600_)
  );
  AND2_X1 _18268_ (
    .A1(_10593_),
    .A2(_10600_),
    .ZN(_10601_)
  );
  MUX2_X1 _18269_ (
    .A(\rf[29] [5]),
    .B(\rf[25] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10602_)
  );
  AND2_X1 _18270_ (
    .A1(\rf[27] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10603_)
  );
  MUX2_X1 _18271_ (
    .A(_10602_),
    .B(_10603_),
    .S(_08541_),
    .Z(_10604_)
  );
  MUX2_X1 _18272_ (
    .A(_10601_),
    .B(_10604_),
    .S(_08540_),
    .Z(_10605_)
  );
  INV_X1 _18273_ (
    .A(_10605_),
    .ZN(_10606_)
  );
  AND2_X1 _18274_ (
    .A1(_08571_),
    .A2(_10606_),
    .ZN(_10607_)
  );
  INV_X1 _18275_ (
    .A(_10607_),
    .ZN(_10608_)
  );
  AND2_X1 _18276_ (
    .A1(_10586_),
    .A2(_10608_),
    .ZN(_10609_)
  );
  MUX2_X1 _18277_ (
    .A(_10549_),
    .B(_10609_),
    .S(_08543_),
    .Z(_10610_)
  );
  MUX2_X1 _18278_ (
    .A(_10610_),
    .B(_10505_),
    .S(_10131_),
    .Z(_10611_)
  );
  AND2_X1 _18279_ (
    .A1(_10082_),
    .A2(_10611_),
    .ZN(_10612_)
  );
  INV_X1 _18280_ (
    .A(_10612_),
    .ZN(_10613_)
  );
  AND2_X1 _18281_ (
    .A1(_10502_),
    .A2(_10613_),
    .ZN(_10614_)
  );
  INV_X1 _18282_ (
    .A(_10614_),
    .ZN(_10615_)
  );
  MUX2_X1 _18283_ (
    .A(ex_reg_rs_msb_0[3]),
    .B(_10615_),
    .S(_10079_),
    .Z(_00070_)
  );
  AND2_X1 _18284_ (
    .A1(ibuf_io_inst_0_bits_raw[6]),
    .A2(_09295_),
    .ZN(_10616_)
  );
  INV_X1 _18285_ (
    .A(_10616_),
    .ZN(_10617_)
  );
  MUX2_X1 _18286_ (
    .A(csr_io_rw_rdata[6]),
    .B(wb_reg_wdata[6]),
    .S(_10134_),
    .Z(_10618_)
  );
  MUX2_X1 _18287_ (
    .A(div_io_resp_bits_data[6]),
    .B(_10618_),
    .S(_08649_),
    .Z(_10619_)
  );
  MUX2_X1 _18288_ (
    .A(_10619_),
    .B(io_dmem_resp_bits_data[6]),
    .S(_08631_),
    .Z(_10620_)
  );
  MUX2_X1 _18289_ (
    .A(\rf[3] [6]),
    .B(\rf[1] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_10621_)
  );
  MUX2_X1 _18290_ (
    .A(\rf[7] [6]),
    .B(\rf[5] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_10622_)
  );
  MUX2_X1 _18291_ (
    .A(_10621_),
    .B(_10622_),
    .S(_08542_),
    .Z(_10623_)
  );
  AND2_X1 _18292_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_10623_),
    .ZN(_10624_)
  );
  INV_X1 _18293_ (
    .A(_10624_),
    .ZN(_10625_)
  );
  MUX2_X1 _18294_ (
    .A(\rf[13] [6]),
    .B(\rf[9] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10626_)
  );
  INV_X1 _18295_ (
    .A(_10626_),
    .ZN(_10627_)
  );
  AND2_X1 _18296_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10627_),
    .ZN(_10628_)
  );
  INV_X1 _18297_ (
    .A(_10628_),
    .ZN(_10629_)
  );
  MUX2_X1 _18298_ (
    .A(\rf[15] [6]),
    .B(\rf[11] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10630_)
  );
  INV_X1 _18299_ (
    .A(_10630_),
    .ZN(_10631_)
  );
  AND2_X1 _18300_ (
    .A1(_08541_),
    .A2(_10631_),
    .ZN(_10632_)
  );
  INV_X1 _18301_ (
    .A(_10632_),
    .ZN(_10633_)
  );
  AND2_X1 _18302_ (
    .A1(_08543_),
    .A2(_10633_),
    .ZN(_10634_)
  );
  AND2_X1 _18303_ (
    .A1(_10629_),
    .A2(_10634_),
    .ZN(_10635_)
  );
  INV_X1 _18304_ (
    .A(_10635_),
    .ZN(_10636_)
  );
  AND2_X1 _18305_ (
    .A1(_08540_),
    .A2(_10636_),
    .ZN(_10637_)
  );
  AND2_X1 _18306_ (
    .A1(_10625_),
    .A2(_10637_),
    .ZN(_10638_)
  );
  INV_X1 _18307_ (
    .A(_10638_),
    .ZN(_10639_)
  );
  MUX2_X1 _18308_ (
    .A(\rf[2] [6]),
    .B(\rf[0] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_10640_)
  );
  MUX2_X1 _18309_ (
    .A(\rf[6] [6]),
    .B(\rf[4] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_10641_)
  );
  MUX2_X1 _18310_ (
    .A(_10640_),
    .B(_10641_),
    .S(_08542_),
    .Z(_10642_)
  );
  AND2_X1 _18311_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_10642_),
    .ZN(_10643_)
  );
  INV_X1 _18312_ (
    .A(_10643_),
    .ZN(_10644_)
  );
  MUX2_X1 _18313_ (
    .A(\rf[12] [6]),
    .B(\rf[8] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10645_)
  );
  INV_X1 _18314_ (
    .A(_10645_),
    .ZN(_10646_)
  );
  AND2_X1 _18315_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10646_),
    .ZN(_10647_)
  );
  INV_X1 _18316_ (
    .A(_10647_),
    .ZN(_10648_)
  );
  MUX2_X1 _18317_ (
    .A(\rf[14] [6]),
    .B(\rf[10] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10649_)
  );
  INV_X1 _18318_ (
    .A(_10649_),
    .ZN(_10650_)
  );
  AND2_X1 _18319_ (
    .A1(_08541_),
    .A2(_10650_),
    .ZN(_10651_)
  );
  INV_X1 _18320_ (
    .A(_10651_),
    .ZN(_10652_)
  );
  AND2_X1 _18321_ (
    .A1(_08543_),
    .A2(_10652_),
    .ZN(_10653_)
  );
  AND2_X1 _18322_ (
    .A1(_10648_),
    .A2(_10653_),
    .ZN(_10654_)
  );
  INV_X1 _18323_ (
    .A(_10654_),
    .ZN(_10655_)
  );
  AND2_X1 _18324_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_10655_),
    .ZN(_10656_)
  );
  AND2_X1 _18325_ (
    .A1(_10644_),
    .A2(_10656_),
    .ZN(_10657_)
  );
  INV_X1 _18326_ (
    .A(_10657_),
    .ZN(_10658_)
  );
  AND2_X1 _18327_ (
    .A1(_10639_),
    .A2(_10658_),
    .ZN(_10659_)
  );
  INV_X1 _18328_ (
    .A(_10659_),
    .ZN(_10660_)
  );
  AND2_X1 _18329_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_10660_),
    .ZN(_10661_)
  );
  INV_X1 _18330_ (
    .A(_10661_),
    .ZN(_10662_)
  );
  AND2_X1 _18331_ (
    .A1(_08237_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10663_)
  );
  INV_X1 _18332_ (
    .A(_10663_),
    .ZN(_10664_)
  );
  AND2_X1 _18333_ (
    .A1(_08460_),
    .A2(_08542_),
    .ZN(_10665_)
  );
  INV_X1 _18334_ (
    .A(_10665_),
    .ZN(_10666_)
  );
  AND2_X1 _18335_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10666_),
    .ZN(_10667_)
  );
  AND2_X1 _18336_ (
    .A1(_10664_),
    .A2(_10667_),
    .ZN(_10668_)
  );
  INV_X1 _18337_ (
    .A(_10668_),
    .ZN(_10669_)
  );
  AND2_X1 _18338_ (
    .A1(\rf[27] [6]),
    .A2(_10453_),
    .ZN(_10670_)
  );
  INV_X1 _18339_ (
    .A(_10670_),
    .ZN(_10671_)
  );
  MUX2_X1 _18340_ (
    .A(\rf[30] [6]),
    .B(\rf[26] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10672_)
  );
  AND2_X1 _18341_ (
    .A1(_08508_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10673_)
  );
  INV_X1 _18342_ (
    .A(_10673_),
    .ZN(_10674_)
  );
  AND2_X1 _18343_ (
    .A1(_08438_),
    .A2(_08542_),
    .ZN(_10675_)
  );
  INV_X1 _18344_ (
    .A(_10675_),
    .ZN(_10676_)
  );
  AND2_X1 _18345_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10674_),
    .ZN(_10677_)
  );
  AND2_X1 _18346_ (
    .A1(_10676_),
    .A2(_10677_),
    .ZN(_10678_)
  );
  INV_X1 _18347_ (
    .A(_10678_),
    .ZN(_10679_)
  );
  AND2_X1 _18348_ (
    .A1(_08541_),
    .A2(_10672_),
    .ZN(_10680_)
  );
  INV_X1 _18349_ (
    .A(_10680_),
    .ZN(_10681_)
  );
  AND2_X1 _18350_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_10681_),
    .ZN(_10682_)
  );
  AND2_X1 _18351_ (
    .A1(_10679_),
    .A2(_10682_),
    .ZN(_10683_)
  );
  INV_X1 _18352_ (
    .A(_10683_),
    .ZN(_10684_)
  );
  AND2_X1 _18353_ (
    .A1(_08540_),
    .A2(_10671_),
    .ZN(_10685_)
  );
  AND2_X1 _18354_ (
    .A1(_10669_),
    .A2(_10685_),
    .ZN(_10686_)
  );
  INV_X1 _18355_ (
    .A(_10686_),
    .ZN(_10687_)
  );
  AND2_X1 _18356_ (
    .A1(_10684_),
    .A2(_10687_),
    .ZN(_10688_)
  );
  AND2_X1 _18357_ (
    .A1(_08543_),
    .A2(_10688_),
    .ZN(_10689_)
  );
  INV_X1 _18358_ (
    .A(_10689_),
    .ZN(_10690_)
  );
  AND2_X1 _18359_ (
    .A1(_08379_),
    .A2(_08542_),
    .ZN(_10691_)
  );
  INV_X1 _18360_ (
    .A(_10691_),
    .ZN(_10692_)
  );
  AND2_X1 _18361_ (
    .A1(_08280_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10693_)
  );
  INV_X1 _18362_ (
    .A(_10693_),
    .ZN(_10694_)
  );
  AND2_X1 _18363_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10694_),
    .ZN(_10695_)
  );
  AND2_X1 _18364_ (
    .A1(_10692_),
    .A2(_10695_),
    .ZN(_10696_)
  );
  INV_X1 _18365_ (
    .A(_10696_),
    .ZN(_10697_)
  );
  MUX2_X1 _18366_ (
    .A(\rf[22] [6]),
    .B(\rf[18] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10698_)
  );
  AND2_X1 _18367_ (
    .A1(_08541_),
    .A2(_10698_),
    .ZN(_10699_)
  );
  INV_X1 _18368_ (
    .A(_10699_),
    .ZN(_10700_)
  );
  AND2_X1 _18369_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_10700_),
    .ZN(_10701_)
  );
  AND2_X1 _18370_ (
    .A1(_10697_),
    .A2(_10701_),
    .ZN(_10702_)
  );
  INV_X1 _18371_ (
    .A(_10702_),
    .ZN(_10703_)
  );
  AND2_X1 _18372_ (
    .A1(_08310_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10704_)
  );
  INV_X1 _18373_ (
    .A(_10704_),
    .ZN(_10705_)
  );
  AND2_X1 _18374_ (
    .A1(_08409_),
    .A2(_08542_),
    .ZN(_10706_)
  );
  INV_X1 _18375_ (
    .A(_10706_),
    .ZN(_10707_)
  );
  AND2_X1 _18376_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10707_),
    .ZN(_10708_)
  );
  AND2_X1 _18377_ (
    .A1(_10705_),
    .A2(_10708_),
    .ZN(_10709_)
  );
  INV_X1 _18378_ (
    .A(_10709_),
    .ZN(_10710_)
  );
  MUX2_X1 _18379_ (
    .A(\rf[23] [6]),
    .B(\rf[19] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10711_)
  );
  AND2_X1 _18380_ (
    .A1(_08541_),
    .A2(_10711_),
    .ZN(_10712_)
  );
  INV_X1 _18381_ (
    .A(_10712_),
    .ZN(_10713_)
  );
  AND2_X1 _18382_ (
    .A1(_08540_),
    .A2(_10713_),
    .ZN(_10714_)
  );
  AND2_X1 _18383_ (
    .A1(_10710_),
    .A2(_10714_),
    .ZN(_10715_)
  );
  INV_X1 _18384_ (
    .A(_10715_),
    .ZN(_10716_)
  );
  AND2_X1 _18385_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_10716_),
    .ZN(_10717_)
  );
  AND2_X1 _18386_ (
    .A1(_10703_),
    .A2(_10717_),
    .ZN(_10718_)
  );
  INV_X1 _18387_ (
    .A(_10718_),
    .ZN(_10719_)
  );
  AND2_X1 _18388_ (
    .A1(_08571_),
    .A2(_10719_),
    .ZN(_10720_)
  );
  AND2_X1 _18389_ (
    .A1(_10690_),
    .A2(_10720_),
    .ZN(_10721_)
  );
  INV_X1 _18390_ (
    .A(_10721_),
    .ZN(_10722_)
  );
  AND2_X1 _18391_ (
    .A1(_10662_),
    .A2(_10722_),
    .ZN(_10723_)
  );
  MUX2_X1 _18392_ (
    .A(_10620_),
    .B(_10723_),
    .S(_10132_),
    .Z(_10724_)
  );
  AND2_X1 _18393_ (
    .A1(_10082_),
    .A2(_10724_),
    .ZN(_10725_)
  );
  INV_X1 _18394_ (
    .A(_10725_),
    .ZN(_10726_)
  );
  AND2_X1 _18395_ (
    .A1(_10617_),
    .A2(_10726_),
    .ZN(_10727_)
  );
  INV_X1 _18396_ (
    .A(_10727_),
    .ZN(_10728_)
  );
  MUX2_X1 _18397_ (
    .A(ex_reg_rs_msb_0[4]),
    .B(_10728_),
    .S(_10079_),
    .Z(_00071_)
  );
  AND2_X1 _18398_ (
    .A1(ibuf_io_inst_0_bits_raw[7]),
    .A2(_09295_),
    .ZN(_10729_)
  );
  INV_X1 _18399_ (
    .A(_10729_),
    .ZN(_10730_)
  );
  MUX2_X1 _18400_ (
    .A(csr_io_rw_rdata[7]),
    .B(wb_reg_wdata[7]),
    .S(_10134_),
    .Z(_10731_)
  );
  MUX2_X1 _18401_ (
    .A(div_io_resp_bits_data[7]),
    .B(_10731_),
    .S(_08649_),
    .Z(_10732_)
  );
  MUX2_X1 _18402_ (
    .A(_10732_),
    .B(io_dmem_resp_bits_data[7]),
    .S(_08631_),
    .Z(_10733_)
  );
  MUX2_X1 _18403_ (
    .A(\rf[3] [7]),
    .B(\rf[1] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_10734_)
  );
  MUX2_X1 _18404_ (
    .A(\rf[7] [7]),
    .B(\rf[5] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_10735_)
  );
  MUX2_X1 _18405_ (
    .A(_10734_),
    .B(_10735_),
    .S(_08542_),
    .Z(_10736_)
  );
  AND2_X1 _18406_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_10736_),
    .ZN(_10737_)
  );
  INV_X1 _18407_ (
    .A(_10737_),
    .ZN(_10738_)
  );
  MUX2_X1 _18408_ (
    .A(\rf[13] [7]),
    .B(\rf[9] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10739_)
  );
  INV_X1 _18409_ (
    .A(_10739_),
    .ZN(_10740_)
  );
  AND2_X1 _18410_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10740_),
    .ZN(_10741_)
  );
  INV_X1 _18411_ (
    .A(_10741_),
    .ZN(_10742_)
  );
  MUX2_X1 _18412_ (
    .A(\rf[15] [7]),
    .B(\rf[11] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10743_)
  );
  INV_X1 _18413_ (
    .A(_10743_),
    .ZN(_10744_)
  );
  AND2_X1 _18414_ (
    .A1(_08541_),
    .A2(_10744_),
    .ZN(_10745_)
  );
  INV_X1 _18415_ (
    .A(_10745_),
    .ZN(_10746_)
  );
  AND2_X1 _18416_ (
    .A1(_08543_),
    .A2(_10746_),
    .ZN(_10747_)
  );
  AND2_X1 _18417_ (
    .A1(_10742_),
    .A2(_10747_),
    .ZN(_10748_)
  );
  INV_X1 _18418_ (
    .A(_10748_),
    .ZN(_10749_)
  );
  AND2_X1 _18419_ (
    .A1(_08540_),
    .A2(_10749_),
    .ZN(_10750_)
  );
  AND2_X1 _18420_ (
    .A1(_10738_),
    .A2(_10750_),
    .ZN(_10751_)
  );
  INV_X1 _18421_ (
    .A(_10751_),
    .ZN(_10752_)
  );
  MUX2_X1 _18422_ (
    .A(\rf[2] [7]),
    .B(\rf[0] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_10753_)
  );
  MUX2_X1 _18423_ (
    .A(\rf[6] [7]),
    .B(\rf[4] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_10754_)
  );
  MUX2_X1 _18424_ (
    .A(_10753_),
    .B(_10754_),
    .S(_08542_),
    .Z(_10755_)
  );
  AND2_X1 _18425_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_10755_),
    .ZN(_10756_)
  );
  INV_X1 _18426_ (
    .A(_10756_),
    .ZN(_10757_)
  );
  MUX2_X1 _18427_ (
    .A(\rf[12] [7]),
    .B(\rf[8] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10758_)
  );
  INV_X1 _18428_ (
    .A(_10758_),
    .ZN(_10759_)
  );
  AND2_X1 _18429_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10759_),
    .ZN(_10760_)
  );
  INV_X1 _18430_ (
    .A(_10760_),
    .ZN(_10761_)
  );
  MUX2_X1 _18431_ (
    .A(\rf[14] [7]),
    .B(\rf[10] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10762_)
  );
  INV_X1 _18432_ (
    .A(_10762_),
    .ZN(_10763_)
  );
  AND2_X1 _18433_ (
    .A1(_08541_),
    .A2(_10763_),
    .ZN(_10764_)
  );
  INV_X1 _18434_ (
    .A(_10764_),
    .ZN(_10765_)
  );
  AND2_X1 _18435_ (
    .A1(_08543_),
    .A2(_10765_),
    .ZN(_10766_)
  );
  AND2_X1 _18436_ (
    .A1(_10761_),
    .A2(_10766_),
    .ZN(_10767_)
  );
  INV_X1 _18437_ (
    .A(_10767_),
    .ZN(_10768_)
  );
  AND2_X1 _18438_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_10768_),
    .ZN(_10769_)
  );
  AND2_X1 _18439_ (
    .A1(_10757_),
    .A2(_10769_),
    .ZN(_10770_)
  );
  INV_X1 _18440_ (
    .A(_10770_),
    .ZN(_10771_)
  );
  AND2_X1 _18441_ (
    .A1(_10752_),
    .A2(_10771_),
    .ZN(_10772_)
  );
  INV_X1 _18442_ (
    .A(_10772_),
    .ZN(_10773_)
  );
  AND2_X1 _18443_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_10773_),
    .ZN(_10774_)
  );
  INV_X1 _18444_ (
    .A(_10774_),
    .ZN(_10775_)
  );
  AND2_X1 _18445_ (
    .A1(_08238_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10776_)
  );
  INV_X1 _18446_ (
    .A(_10776_),
    .ZN(_10777_)
  );
  AND2_X1 _18447_ (
    .A1(_08461_),
    .A2(_08542_),
    .ZN(_10778_)
  );
  INV_X1 _18448_ (
    .A(_10778_),
    .ZN(_10779_)
  );
  AND2_X1 _18449_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10779_),
    .ZN(_10780_)
  );
  AND2_X1 _18450_ (
    .A1(_10777_),
    .A2(_10780_),
    .ZN(_10781_)
  );
  INV_X1 _18451_ (
    .A(_10781_),
    .ZN(_10782_)
  );
  AND2_X1 _18452_ (
    .A1(\rf[27] [7]),
    .A2(_10453_),
    .ZN(_10783_)
  );
  INV_X1 _18453_ (
    .A(_10783_),
    .ZN(_10784_)
  );
  MUX2_X1 _18454_ (
    .A(\rf[30] [7]),
    .B(\rf[26] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10785_)
  );
  AND2_X1 _18455_ (
    .A1(_08509_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10786_)
  );
  INV_X1 _18456_ (
    .A(_10786_),
    .ZN(_10787_)
  );
  AND2_X1 _18457_ (
    .A1(_08439_),
    .A2(_08542_),
    .ZN(_10788_)
  );
  INV_X1 _18458_ (
    .A(_10788_),
    .ZN(_10789_)
  );
  AND2_X1 _18459_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10787_),
    .ZN(_10790_)
  );
  AND2_X1 _18460_ (
    .A1(_10789_),
    .A2(_10790_),
    .ZN(_10791_)
  );
  INV_X1 _18461_ (
    .A(_10791_),
    .ZN(_10792_)
  );
  AND2_X1 _18462_ (
    .A1(_08541_),
    .A2(_10785_),
    .ZN(_10793_)
  );
  INV_X1 _18463_ (
    .A(_10793_),
    .ZN(_10794_)
  );
  AND2_X1 _18464_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_10794_),
    .ZN(_10795_)
  );
  AND2_X1 _18465_ (
    .A1(_10792_),
    .A2(_10795_),
    .ZN(_10796_)
  );
  INV_X1 _18466_ (
    .A(_10796_),
    .ZN(_10797_)
  );
  AND2_X1 _18467_ (
    .A1(_08540_),
    .A2(_10784_),
    .ZN(_10798_)
  );
  AND2_X1 _18468_ (
    .A1(_10782_),
    .A2(_10798_),
    .ZN(_10799_)
  );
  INV_X1 _18469_ (
    .A(_10799_),
    .ZN(_10800_)
  );
  AND2_X1 _18470_ (
    .A1(_10797_),
    .A2(_10800_),
    .ZN(_10801_)
  );
  AND2_X1 _18471_ (
    .A1(_08543_),
    .A2(_10801_),
    .ZN(_10802_)
  );
  INV_X1 _18472_ (
    .A(_10802_),
    .ZN(_10803_)
  );
  AND2_X1 _18473_ (
    .A1(_08380_),
    .A2(_08542_),
    .ZN(_10804_)
  );
  INV_X1 _18474_ (
    .A(_10804_),
    .ZN(_10805_)
  );
  AND2_X1 _18475_ (
    .A1(_08281_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10806_)
  );
  INV_X1 _18476_ (
    .A(_10806_),
    .ZN(_10807_)
  );
  AND2_X1 _18477_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10807_),
    .ZN(_10808_)
  );
  AND2_X1 _18478_ (
    .A1(_10805_),
    .A2(_10808_),
    .ZN(_10809_)
  );
  INV_X1 _18479_ (
    .A(_10809_),
    .ZN(_10810_)
  );
  MUX2_X1 _18480_ (
    .A(\rf[22] [7]),
    .B(\rf[18] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10811_)
  );
  AND2_X1 _18481_ (
    .A1(_08541_),
    .A2(_10811_),
    .ZN(_10812_)
  );
  INV_X1 _18482_ (
    .A(_10812_),
    .ZN(_10813_)
  );
  AND2_X1 _18483_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_10813_),
    .ZN(_10814_)
  );
  AND2_X1 _18484_ (
    .A1(_10810_),
    .A2(_10814_),
    .ZN(_10815_)
  );
  INV_X1 _18485_ (
    .A(_10815_),
    .ZN(_10816_)
  );
  AND2_X1 _18486_ (
    .A1(_08311_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10817_)
  );
  INV_X1 _18487_ (
    .A(_10817_),
    .ZN(_10818_)
  );
  AND2_X1 _18488_ (
    .A1(_08410_),
    .A2(_08542_),
    .ZN(_10819_)
  );
  INV_X1 _18489_ (
    .A(_10819_),
    .ZN(_10820_)
  );
  AND2_X1 _18490_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10820_),
    .ZN(_10821_)
  );
  AND2_X1 _18491_ (
    .A1(_10818_),
    .A2(_10821_),
    .ZN(_10822_)
  );
  INV_X1 _18492_ (
    .A(_10822_),
    .ZN(_10823_)
  );
  MUX2_X1 _18493_ (
    .A(\rf[23] [7]),
    .B(\rf[19] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10824_)
  );
  AND2_X1 _18494_ (
    .A1(_08541_),
    .A2(_10824_),
    .ZN(_10825_)
  );
  INV_X1 _18495_ (
    .A(_10825_),
    .ZN(_10826_)
  );
  AND2_X1 _18496_ (
    .A1(_08540_),
    .A2(_10826_),
    .ZN(_10827_)
  );
  AND2_X1 _18497_ (
    .A1(_10823_),
    .A2(_10827_),
    .ZN(_10828_)
  );
  INV_X1 _18498_ (
    .A(_10828_),
    .ZN(_10829_)
  );
  AND2_X1 _18499_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_10829_),
    .ZN(_10830_)
  );
  AND2_X1 _18500_ (
    .A1(_10816_),
    .A2(_10830_),
    .ZN(_10831_)
  );
  INV_X1 _18501_ (
    .A(_10831_),
    .ZN(_10832_)
  );
  AND2_X1 _18502_ (
    .A1(_08571_),
    .A2(_10832_),
    .ZN(_10833_)
  );
  AND2_X1 _18503_ (
    .A1(_10803_),
    .A2(_10833_),
    .ZN(_10834_)
  );
  INV_X1 _18504_ (
    .A(_10834_),
    .ZN(_10835_)
  );
  AND2_X1 _18505_ (
    .A1(_10775_),
    .A2(_10835_),
    .ZN(_10836_)
  );
  MUX2_X1 _18506_ (
    .A(_10733_),
    .B(_10836_),
    .S(_10132_),
    .Z(_10837_)
  );
  AND2_X1 _18507_ (
    .A1(_10082_),
    .A2(_10837_),
    .ZN(_10838_)
  );
  INV_X1 _18508_ (
    .A(_10838_),
    .ZN(_10839_)
  );
  AND2_X1 _18509_ (
    .A1(_10730_),
    .A2(_10839_),
    .ZN(_10840_)
  );
  INV_X1 _18510_ (
    .A(_10840_),
    .ZN(_10841_)
  );
  MUX2_X1 _18511_ (
    .A(ex_reg_rs_msb_0[5]),
    .B(_10841_),
    .S(_10079_),
    .Z(_00072_)
  );
  AND2_X1 _18512_ (
    .A1(ibuf_io_inst_0_bits_raw[8]),
    .A2(_09295_),
    .ZN(_10842_)
  );
  INV_X1 _18513_ (
    .A(_10842_),
    .ZN(_10843_)
  );
  MUX2_X1 _18514_ (
    .A(csr_io_rw_rdata[8]),
    .B(wb_reg_wdata[8]),
    .S(_10134_),
    .Z(_10844_)
  );
  MUX2_X1 _18515_ (
    .A(div_io_resp_bits_data[8]),
    .B(_10844_),
    .S(_08649_),
    .Z(_10845_)
  );
  MUX2_X1 _18516_ (
    .A(_10845_),
    .B(io_dmem_resp_bits_data[8]),
    .S(_08631_),
    .Z(_10846_)
  );
  AND2_X1 _18517_ (
    .A1(_08239_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10847_)
  );
  INV_X1 _18518_ (
    .A(_10847_),
    .ZN(_10848_)
  );
  AND2_X1 _18519_ (
    .A1(_08462_),
    .A2(_08542_),
    .ZN(_10849_)
  );
  INV_X1 _18520_ (
    .A(_10849_),
    .ZN(_10850_)
  );
  AND2_X1 _18521_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10850_),
    .ZN(_10851_)
  );
  AND2_X1 _18522_ (
    .A1(_10848_),
    .A2(_10851_),
    .ZN(_10852_)
  );
  INV_X1 _18523_ (
    .A(_10852_),
    .ZN(_10853_)
  );
  AND2_X1 _18524_ (
    .A1(\rf[27] [8]),
    .A2(_10453_),
    .ZN(_10854_)
  );
  INV_X1 _18525_ (
    .A(_10854_),
    .ZN(_10855_)
  );
  MUX2_X1 _18526_ (
    .A(\rf[30] [8]),
    .B(\rf[26] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10856_)
  );
  AND2_X1 _18527_ (
    .A1(_08510_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10857_)
  );
  INV_X1 _18528_ (
    .A(_10857_),
    .ZN(_10858_)
  );
  AND2_X1 _18529_ (
    .A1(_08440_),
    .A2(_08542_),
    .ZN(_10859_)
  );
  INV_X1 _18530_ (
    .A(_10859_),
    .ZN(_10860_)
  );
  AND2_X1 _18531_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10858_),
    .ZN(_10861_)
  );
  AND2_X1 _18532_ (
    .A1(_10860_),
    .A2(_10861_),
    .ZN(_10862_)
  );
  INV_X1 _18533_ (
    .A(_10862_),
    .ZN(_10863_)
  );
  AND2_X1 _18534_ (
    .A1(_08541_),
    .A2(_10856_),
    .ZN(_10864_)
  );
  INV_X1 _18535_ (
    .A(_10864_),
    .ZN(_10865_)
  );
  AND2_X1 _18536_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_10865_),
    .ZN(_10866_)
  );
  AND2_X1 _18537_ (
    .A1(_10863_),
    .A2(_10866_),
    .ZN(_10867_)
  );
  INV_X1 _18538_ (
    .A(_10867_),
    .ZN(_10868_)
  );
  AND2_X1 _18539_ (
    .A1(_08540_),
    .A2(_10855_),
    .ZN(_10869_)
  );
  AND2_X1 _18540_ (
    .A1(_10853_),
    .A2(_10869_),
    .ZN(_10870_)
  );
  INV_X1 _18541_ (
    .A(_10870_),
    .ZN(_10871_)
  );
  AND2_X1 _18542_ (
    .A1(_10868_),
    .A2(_10871_),
    .ZN(_10872_)
  );
  AND2_X1 _18543_ (
    .A1(_08543_),
    .A2(_10872_),
    .ZN(_10873_)
  );
  INV_X1 _18544_ (
    .A(_10873_),
    .ZN(_10874_)
  );
  AND2_X1 _18545_ (
    .A1(_08381_),
    .A2(_08542_),
    .ZN(_10875_)
  );
  INV_X1 _18546_ (
    .A(_10875_),
    .ZN(_10876_)
  );
  AND2_X1 _18547_ (
    .A1(_08282_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10877_)
  );
  INV_X1 _18548_ (
    .A(_10877_),
    .ZN(_10878_)
  );
  AND2_X1 _18549_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10878_),
    .ZN(_10879_)
  );
  AND2_X1 _18550_ (
    .A1(_10876_),
    .A2(_10879_),
    .ZN(_10880_)
  );
  INV_X1 _18551_ (
    .A(_10880_),
    .ZN(_10881_)
  );
  MUX2_X1 _18552_ (
    .A(\rf[22] [8]),
    .B(\rf[18] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10882_)
  );
  AND2_X1 _18553_ (
    .A1(_08541_),
    .A2(_10882_),
    .ZN(_10883_)
  );
  INV_X1 _18554_ (
    .A(_10883_),
    .ZN(_10884_)
  );
  AND2_X1 _18555_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_10884_),
    .ZN(_10885_)
  );
  AND2_X1 _18556_ (
    .A1(_10881_),
    .A2(_10885_),
    .ZN(_10886_)
  );
  INV_X1 _18557_ (
    .A(_10886_),
    .ZN(_10887_)
  );
  AND2_X1 _18558_ (
    .A1(_08312_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10888_)
  );
  INV_X1 _18559_ (
    .A(_10888_),
    .ZN(_10889_)
  );
  AND2_X1 _18560_ (
    .A1(_08411_),
    .A2(_08542_),
    .ZN(_10890_)
  );
  INV_X1 _18561_ (
    .A(_10890_),
    .ZN(_10891_)
  );
  AND2_X1 _18562_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10891_),
    .ZN(_10892_)
  );
  AND2_X1 _18563_ (
    .A1(_10889_),
    .A2(_10892_),
    .ZN(_10893_)
  );
  INV_X1 _18564_ (
    .A(_10893_),
    .ZN(_10894_)
  );
  MUX2_X1 _18565_ (
    .A(\rf[23] [8]),
    .B(\rf[19] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10895_)
  );
  AND2_X1 _18566_ (
    .A1(_08541_),
    .A2(_10895_),
    .ZN(_10896_)
  );
  INV_X1 _18567_ (
    .A(_10896_),
    .ZN(_10897_)
  );
  AND2_X1 _18568_ (
    .A1(_08540_),
    .A2(_10897_),
    .ZN(_10898_)
  );
  AND2_X1 _18569_ (
    .A1(_10894_),
    .A2(_10898_),
    .ZN(_10899_)
  );
  INV_X1 _18570_ (
    .A(_10899_),
    .ZN(_10900_)
  );
  AND2_X1 _18571_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_10900_),
    .ZN(_10901_)
  );
  AND2_X1 _18572_ (
    .A1(_10887_),
    .A2(_10901_),
    .ZN(_10902_)
  );
  INV_X1 _18573_ (
    .A(_10902_),
    .ZN(_10903_)
  );
  AND2_X1 _18574_ (
    .A1(_08571_),
    .A2(_10903_),
    .ZN(_10904_)
  );
  AND2_X1 _18575_ (
    .A1(_10874_),
    .A2(_10904_),
    .ZN(_10905_)
  );
  INV_X1 _18576_ (
    .A(_10905_),
    .ZN(_10906_)
  );
  MUX2_X1 _18577_ (
    .A(\rf[1] [8]),
    .B(\rf[0] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_10907_)
  );
  MUX2_X1 _18578_ (
    .A(\rf[5] [8]),
    .B(\rf[4] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_10908_)
  );
  MUX2_X1 _18579_ (
    .A(_10907_),
    .B(_10908_),
    .S(_08542_),
    .Z(_10909_)
  );
  INV_X1 _18580_ (
    .A(_10909_),
    .ZN(_10910_)
  );
  AND2_X1 _18581_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_10910_),
    .ZN(_10911_)
  );
  INV_X1 _18582_ (
    .A(_10911_),
    .ZN(_10912_)
  );
  MUX2_X1 _18583_ (
    .A(\rf[12] [8]),
    .B(\rf[8] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10913_)
  );
  INV_X1 _18584_ (
    .A(_10913_),
    .ZN(_10914_)
  );
  AND2_X1 _18585_ (
    .A1(_10213_),
    .A2(_10914_),
    .ZN(_10915_)
  );
  INV_X1 _18586_ (
    .A(_10915_),
    .ZN(_10916_)
  );
  MUX2_X1 _18587_ (
    .A(\rf[13] [8]),
    .B(\rf[9] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10917_)
  );
  INV_X1 _18588_ (
    .A(_10917_),
    .ZN(_10918_)
  );
  AND2_X1 _18589_ (
    .A1(_09110_),
    .A2(_10918_),
    .ZN(_10919_)
  );
  INV_X1 _18590_ (
    .A(_10919_),
    .ZN(_10920_)
  );
  AND2_X1 _18591_ (
    .A1(_10916_),
    .A2(_10920_),
    .ZN(_10921_)
  );
  AND2_X1 _18592_ (
    .A1(_10912_),
    .A2(_10921_),
    .ZN(_10922_)
  );
  AND2_X1 _18593_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10922_),
    .ZN(_10923_)
  );
  INV_X1 _18594_ (
    .A(_10923_),
    .ZN(_10924_)
  );
  MUX2_X1 _18595_ (
    .A(\rf[3] [8]),
    .B(\rf[2] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_10925_)
  );
  MUX2_X1 _18596_ (
    .A(\rf[7] [8]),
    .B(\rf[6] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_10926_)
  );
  MUX2_X1 _18597_ (
    .A(_10925_),
    .B(_10926_),
    .S(_08542_),
    .Z(_10927_)
  );
  INV_X1 _18598_ (
    .A(_10927_),
    .ZN(_10928_)
  );
  AND2_X1 _18599_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_10928_),
    .ZN(_10929_)
  );
  INV_X1 _18600_ (
    .A(_10929_),
    .ZN(_10930_)
  );
  MUX2_X1 _18601_ (
    .A(\rf[15] [8]),
    .B(\rf[11] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10931_)
  );
  INV_X1 _18602_ (
    .A(_10931_),
    .ZN(_10932_)
  );
  AND2_X1 _18603_ (
    .A1(_09110_),
    .A2(_10932_),
    .ZN(_10933_)
  );
  INV_X1 _18604_ (
    .A(_10933_),
    .ZN(_10934_)
  );
  MUX2_X1 _18605_ (
    .A(\rf[14] [8]),
    .B(\rf[10] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10935_)
  );
  INV_X1 _18606_ (
    .A(_10935_),
    .ZN(_10936_)
  );
  AND2_X1 _18607_ (
    .A1(_10213_),
    .A2(_10936_),
    .ZN(_10937_)
  );
  INV_X1 _18608_ (
    .A(_10937_),
    .ZN(_10938_)
  );
  AND2_X1 _18609_ (
    .A1(_10934_),
    .A2(_10938_),
    .ZN(_10939_)
  );
  AND2_X1 _18610_ (
    .A1(_10930_),
    .A2(_10939_),
    .ZN(_10940_)
  );
  AND2_X1 _18611_ (
    .A1(_08541_),
    .A2(_10940_),
    .ZN(_10941_)
  );
  INV_X1 _18612_ (
    .A(_10941_),
    .ZN(_10942_)
  );
  AND2_X1 _18613_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_10924_),
    .ZN(_10943_)
  );
  AND2_X1 _18614_ (
    .A1(_10942_),
    .A2(_10943_),
    .ZN(_10944_)
  );
  INV_X1 _18615_ (
    .A(_10944_),
    .ZN(_10945_)
  );
  AND2_X1 _18616_ (
    .A1(_10906_),
    .A2(_10945_),
    .ZN(_10946_)
  );
  MUX2_X1 _18617_ (
    .A(_10846_),
    .B(_10946_),
    .S(_10132_),
    .Z(_10947_)
  );
  AND2_X1 _18618_ (
    .A1(_10082_),
    .A2(_10947_),
    .ZN(_10948_)
  );
  INV_X1 _18619_ (
    .A(_10948_),
    .ZN(_10949_)
  );
  AND2_X1 _18620_ (
    .A1(_10843_),
    .A2(_10949_),
    .ZN(_10950_)
  );
  INV_X1 _18621_ (
    .A(_10950_),
    .ZN(_10951_)
  );
  MUX2_X1 _18622_ (
    .A(ex_reg_rs_msb_0[6]),
    .B(_10951_),
    .S(_10079_),
    .Z(_00073_)
  );
  AND2_X1 _18623_ (
    .A1(ibuf_io_inst_0_bits_raw[9]),
    .A2(_09295_),
    .ZN(_10952_)
  );
  INV_X1 _18624_ (
    .A(_10952_),
    .ZN(_10953_)
  );
  MUX2_X1 _18625_ (
    .A(csr_io_rw_rdata[9]),
    .B(wb_reg_wdata[9]),
    .S(_10134_),
    .Z(_10954_)
  );
  MUX2_X1 _18626_ (
    .A(div_io_resp_bits_data[9]),
    .B(_10954_),
    .S(_08649_),
    .Z(_10955_)
  );
  MUX2_X1 _18627_ (
    .A(_10955_),
    .B(io_dmem_resp_bits_data[9]),
    .S(_08631_),
    .Z(_10956_)
  );
  AND2_X1 _18628_ (
    .A1(_08240_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10957_)
  );
  INV_X1 _18629_ (
    .A(_10957_),
    .ZN(_10958_)
  );
  AND2_X1 _18630_ (
    .A1(_08463_),
    .A2(_08542_),
    .ZN(_10959_)
  );
  INV_X1 _18631_ (
    .A(_10959_),
    .ZN(_10960_)
  );
  AND2_X1 _18632_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10960_),
    .ZN(_10961_)
  );
  AND2_X1 _18633_ (
    .A1(_10958_),
    .A2(_10961_),
    .ZN(_10962_)
  );
  INV_X1 _18634_ (
    .A(_10962_),
    .ZN(_10963_)
  );
  AND2_X1 _18635_ (
    .A1(\rf[27] [9]),
    .A2(_10453_),
    .ZN(_10964_)
  );
  INV_X1 _18636_ (
    .A(_10964_),
    .ZN(_10965_)
  );
  MUX2_X1 _18637_ (
    .A(\rf[30] [9]),
    .B(\rf[26] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10966_)
  );
  AND2_X1 _18638_ (
    .A1(_08511_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10967_)
  );
  INV_X1 _18639_ (
    .A(_10967_),
    .ZN(_10968_)
  );
  AND2_X1 _18640_ (
    .A1(_08441_),
    .A2(_08542_),
    .ZN(_10969_)
  );
  INV_X1 _18641_ (
    .A(_10969_),
    .ZN(_10970_)
  );
  AND2_X1 _18642_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10968_),
    .ZN(_10971_)
  );
  AND2_X1 _18643_ (
    .A1(_10970_),
    .A2(_10971_),
    .ZN(_10972_)
  );
  INV_X1 _18644_ (
    .A(_10972_),
    .ZN(_10973_)
  );
  AND2_X1 _18645_ (
    .A1(_08541_),
    .A2(_10966_),
    .ZN(_10974_)
  );
  INV_X1 _18646_ (
    .A(_10974_),
    .ZN(_10975_)
  );
  AND2_X1 _18647_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_10975_),
    .ZN(_10976_)
  );
  AND2_X1 _18648_ (
    .A1(_10973_),
    .A2(_10976_),
    .ZN(_10977_)
  );
  INV_X1 _18649_ (
    .A(_10977_),
    .ZN(_10978_)
  );
  AND2_X1 _18650_ (
    .A1(_08540_),
    .A2(_10965_),
    .ZN(_10979_)
  );
  AND2_X1 _18651_ (
    .A1(_10963_),
    .A2(_10979_),
    .ZN(_10980_)
  );
  INV_X1 _18652_ (
    .A(_10980_),
    .ZN(_10981_)
  );
  AND2_X1 _18653_ (
    .A1(_10978_),
    .A2(_10981_),
    .ZN(_10982_)
  );
  AND2_X1 _18654_ (
    .A1(_08543_),
    .A2(_10982_),
    .ZN(_10983_)
  );
  INV_X1 _18655_ (
    .A(_10983_),
    .ZN(_10984_)
  );
  AND2_X1 _18656_ (
    .A1(_08382_),
    .A2(_08542_),
    .ZN(_10985_)
  );
  INV_X1 _18657_ (
    .A(_10985_),
    .ZN(_10986_)
  );
  AND2_X1 _18658_ (
    .A1(_08283_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10987_)
  );
  INV_X1 _18659_ (
    .A(_10987_),
    .ZN(_10988_)
  );
  AND2_X1 _18660_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_10988_),
    .ZN(_10989_)
  );
  AND2_X1 _18661_ (
    .A1(_10986_),
    .A2(_10989_),
    .ZN(_10990_)
  );
  INV_X1 _18662_ (
    .A(_10990_),
    .ZN(_10991_)
  );
  MUX2_X1 _18663_ (
    .A(\rf[22] [9]),
    .B(\rf[18] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_10992_)
  );
  AND2_X1 _18664_ (
    .A1(_08541_),
    .A2(_10992_),
    .ZN(_10993_)
  );
  INV_X1 _18665_ (
    .A(_10993_),
    .ZN(_10994_)
  );
  AND2_X1 _18666_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_10994_),
    .ZN(_10995_)
  );
  AND2_X1 _18667_ (
    .A1(_10991_),
    .A2(_10995_),
    .ZN(_10996_)
  );
  INV_X1 _18668_ (
    .A(_10996_),
    .ZN(_10997_)
  );
  AND2_X1 _18669_ (
    .A1(_08313_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_10998_)
  );
  INV_X1 _18670_ (
    .A(_10998_),
    .ZN(_10999_)
  );
  AND2_X1 _18671_ (
    .A1(_08412_),
    .A2(_08542_),
    .ZN(_11000_)
  );
  INV_X1 _18672_ (
    .A(_11000_),
    .ZN(_11001_)
  );
  AND2_X1 _18673_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11001_),
    .ZN(_11002_)
  );
  AND2_X1 _18674_ (
    .A1(_10999_),
    .A2(_11002_),
    .ZN(_11003_)
  );
  INV_X1 _18675_ (
    .A(_11003_),
    .ZN(_11004_)
  );
  MUX2_X1 _18676_ (
    .A(\rf[23] [9]),
    .B(\rf[19] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11005_)
  );
  AND2_X1 _18677_ (
    .A1(_08541_),
    .A2(_11005_),
    .ZN(_11006_)
  );
  INV_X1 _18678_ (
    .A(_11006_),
    .ZN(_11007_)
  );
  AND2_X1 _18679_ (
    .A1(_08540_),
    .A2(_11007_),
    .ZN(_11008_)
  );
  AND2_X1 _18680_ (
    .A1(_11004_),
    .A2(_11008_),
    .ZN(_11009_)
  );
  INV_X1 _18681_ (
    .A(_11009_),
    .ZN(_11010_)
  );
  AND2_X1 _18682_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_11010_),
    .ZN(_11011_)
  );
  AND2_X1 _18683_ (
    .A1(_10997_),
    .A2(_11011_),
    .ZN(_11012_)
  );
  INV_X1 _18684_ (
    .A(_11012_),
    .ZN(_11013_)
  );
  AND2_X1 _18685_ (
    .A1(_08571_),
    .A2(_11013_),
    .ZN(_11014_)
  );
  AND2_X1 _18686_ (
    .A1(_10984_),
    .A2(_11014_),
    .ZN(_11015_)
  );
  INV_X1 _18687_ (
    .A(_11015_),
    .ZN(_11016_)
  );
  MUX2_X1 _18688_ (
    .A(\rf[1] [9]),
    .B(\rf[0] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_11017_)
  );
  MUX2_X1 _18689_ (
    .A(\rf[5] [9]),
    .B(\rf[4] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_11018_)
  );
  MUX2_X1 _18690_ (
    .A(_11017_),
    .B(_11018_),
    .S(_08542_),
    .Z(_11019_)
  );
  INV_X1 _18691_ (
    .A(_11019_),
    .ZN(_11020_)
  );
  AND2_X1 _18692_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_11020_),
    .ZN(_11021_)
  );
  INV_X1 _18693_ (
    .A(_11021_),
    .ZN(_11022_)
  );
  MUX2_X1 _18694_ (
    .A(\rf[12] [9]),
    .B(\rf[8] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11023_)
  );
  INV_X1 _18695_ (
    .A(_11023_),
    .ZN(_11024_)
  );
  AND2_X1 _18696_ (
    .A1(_10213_),
    .A2(_11024_),
    .ZN(_11025_)
  );
  INV_X1 _18697_ (
    .A(_11025_),
    .ZN(_11026_)
  );
  MUX2_X1 _18698_ (
    .A(\rf[13] [9]),
    .B(\rf[9] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11027_)
  );
  INV_X1 _18699_ (
    .A(_11027_),
    .ZN(_11028_)
  );
  AND2_X1 _18700_ (
    .A1(_09110_),
    .A2(_11028_),
    .ZN(_11029_)
  );
  INV_X1 _18701_ (
    .A(_11029_),
    .ZN(_11030_)
  );
  AND2_X1 _18702_ (
    .A1(_11026_),
    .A2(_11030_),
    .ZN(_11031_)
  );
  AND2_X1 _18703_ (
    .A1(_11022_),
    .A2(_11031_),
    .ZN(_11032_)
  );
  AND2_X1 _18704_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11032_),
    .ZN(_11033_)
  );
  INV_X1 _18705_ (
    .A(_11033_),
    .ZN(_11034_)
  );
  MUX2_X1 _18706_ (
    .A(\rf[3] [9]),
    .B(\rf[2] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_11035_)
  );
  MUX2_X1 _18707_ (
    .A(\rf[7] [9]),
    .B(\rf[6] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_11036_)
  );
  MUX2_X1 _18708_ (
    .A(_11035_),
    .B(_11036_),
    .S(_08542_),
    .Z(_11037_)
  );
  INV_X1 _18709_ (
    .A(_11037_),
    .ZN(_11038_)
  );
  AND2_X1 _18710_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_11038_),
    .ZN(_11039_)
  );
  INV_X1 _18711_ (
    .A(_11039_),
    .ZN(_11040_)
  );
  MUX2_X1 _18712_ (
    .A(\rf[14] [9]),
    .B(\rf[10] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11041_)
  );
  INV_X1 _18713_ (
    .A(_11041_),
    .ZN(_11042_)
  );
  AND2_X1 _18714_ (
    .A1(_10213_),
    .A2(_11042_),
    .ZN(_11043_)
  );
  INV_X1 _18715_ (
    .A(_11043_),
    .ZN(_11044_)
  );
  MUX2_X1 _18716_ (
    .A(\rf[15] [9]),
    .B(\rf[11] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11045_)
  );
  INV_X1 _18717_ (
    .A(_11045_),
    .ZN(_11046_)
  );
  AND2_X1 _18718_ (
    .A1(_09110_),
    .A2(_11046_),
    .ZN(_11047_)
  );
  INV_X1 _18719_ (
    .A(_11047_),
    .ZN(_11048_)
  );
  AND2_X1 _18720_ (
    .A1(_11044_),
    .A2(_11048_),
    .ZN(_11049_)
  );
  AND2_X1 _18721_ (
    .A1(_11040_),
    .A2(_11049_),
    .ZN(_11050_)
  );
  AND2_X1 _18722_ (
    .A1(_08541_),
    .A2(_11050_),
    .ZN(_11051_)
  );
  INV_X1 _18723_ (
    .A(_11051_),
    .ZN(_11052_)
  );
  AND2_X1 _18724_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_11034_),
    .ZN(_11053_)
  );
  AND2_X1 _18725_ (
    .A1(_11052_),
    .A2(_11053_),
    .ZN(_11054_)
  );
  INV_X1 _18726_ (
    .A(_11054_),
    .ZN(_11055_)
  );
  AND2_X1 _18727_ (
    .A1(_11016_),
    .A2(_11055_),
    .ZN(_11056_)
  );
  MUX2_X1 _18728_ (
    .A(_10956_),
    .B(_11056_),
    .S(_10132_),
    .Z(_11057_)
  );
  AND2_X1 _18729_ (
    .A1(_10082_),
    .A2(_11057_),
    .ZN(_11058_)
  );
  INV_X1 _18730_ (
    .A(_11058_),
    .ZN(_11059_)
  );
  AND2_X1 _18731_ (
    .A1(_10953_),
    .A2(_11059_),
    .ZN(_11060_)
  );
  INV_X1 _18732_ (
    .A(_11060_),
    .ZN(_11061_)
  );
  MUX2_X1 _18733_ (
    .A(ex_reg_rs_msb_0[7]),
    .B(_11061_),
    .S(_10079_),
    .Z(_00074_)
  );
  AND2_X1 _18734_ (
    .A1(ibuf_io_inst_0_bits_raw[10]),
    .A2(_09295_),
    .ZN(_11062_)
  );
  INV_X1 _18735_ (
    .A(_11062_),
    .ZN(_11063_)
  );
  MUX2_X1 _18736_ (
    .A(csr_io_rw_rdata[10]),
    .B(wb_reg_wdata[10]),
    .S(_10134_),
    .Z(_11064_)
  );
  MUX2_X1 _18737_ (
    .A(div_io_resp_bits_data[10]),
    .B(_11064_),
    .S(_08649_),
    .Z(_11065_)
  );
  MUX2_X1 _18738_ (
    .A(_11065_),
    .B(io_dmem_resp_bits_data[10]),
    .S(_08631_),
    .Z(_11066_)
  );
  AND2_X1 _18739_ (
    .A1(\rf[2] [10]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11067_)
  );
  INV_X1 _18740_ (
    .A(_11067_),
    .ZN(_11068_)
  );
  AND2_X1 _18741_ (
    .A1(\rf[6] [10]),
    .A2(_08542_),
    .ZN(_11069_)
  );
  INV_X1 _18742_ (
    .A(_11069_),
    .ZN(_11070_)
  );
  AND2_X1 _18743_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_11070_),
    .ZN(_11071_)
  );
  AND2_X1 _18744_ (
    .A1(_11068_),
    .A2(_11071_),
    .ZN(_11072_)
  );
  INV_X1 _18745_ (
    .A(_11072_),
    .ZN(_11073_)
  );
  AND2_X1 _18746_ (
    .A1(\rf[3] [10]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11074_)
  );
  INV_X1 _18747_ (
    .A(_11074_),
    .ZN(_11075_)
  );
  AND2_X1 _18748_ (
    .A1(\rf[7] [10]),
    .A2(_08542_),
    .ZN(_11076_)
  );
  INV_X1 _18749_ (
    .A(_11076_),
    .ZN(_11077_)
  );
  AND2_X1 _18750_ (
    .A1(_08540_),
    .A2(_11077_),
    .ZN(_11078_)
  );
  AND2_X1 _18751_ (
    .A1(_11075_),
    .A2(_11078_),
    .ZN(_11079_)
  );
  INV_X1 _18752_ (
    .A(_11079_),
    .ZN(_11080_)
  );
  AND2_X1 _18753_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_11080_),
    .ZN(_11081_)
  );
  AND2_X1 _18754_ (
    .A1(_11073_),
    .A2(_11081_),
    .ZN(_11082_)
  );
  INV_X1 _18755_ (
    .A(_11082_),
    .ZN(_11083_)
  );
  MUX2_X1 _18756_ (
    .A(\rf[15] [10]),
    .B(\rf[11] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11084_)
  );
  INV_X1 _18757_ (
    .A(_11084_),
    .ZN(_11085_)
  );
  AND2_X1 _18758_ (
    .A1(_08540_),
    .A2(_11085_),
    .ZN(_11086_)
  );
  INV_X1 _18759_ (
    .A(_11086_),
    .ZN(_11087_)
  );
  MUX2_X1 _18760_ (
    .A(\rf[14] [10]),
    .B(\rf[10] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11088_)
  );
  INV_X1 _18761_ (
    .A(_11088_),
    .ZN(_11089_)
  );
  AND2_X1 _18762_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_11089_),
    .ZN(_11090_)
  );
  INV_X1 _18763_ (
    .A(_11090_),
    .ZN(_11091_)
  );
  AND2_X1 _18764_ (
    .A1(_08543_),
    .A2(_11091_),
    .ZN(_11092_)
  );
  AND2_X1 _18765_ (
    .A1(_11087_),
    .A2(_11092_),
    .ZN(_11093_)
  );
  INV_X1 _18766_ (
    .A(_11093_),
    .ZN(_11094_)
  );
  AND2_X1 _18767_ (
    .A1(_08541_),
    .A2(_11094_),
    .ZN(_11095_)
  );
  AND2_X1 _18768_ (
    .A1(_11083_),
    .A2(_11095_),
    .ZN(_11096_)
  );
  INV_X1 _18769_ (
    .A(_11096_),
    .ZN(_11097_)
  );
  AND2_X1 _18770_ (
    .A1(\rf[4] [10]),
    .A2(_08542_),
    .ZN(_11098_)
  );
  INV_X1 _18771_ (
    .A(_11098_),
    .ZN(_11099_)
  );
  AND2_X1 _18772_ (
    .A1(\rf[0] [10]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11100_)
  );
  INV_X1 _18773_ (
    .A(_11100_),
    .ZN(_11101_)
  );
  AND2_X1 _18774_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_11101_),
    .ZN(_11102_)
  );
  AND2_X1 _18775_ (
    .A1(_11099_),
    .A2(_11102_),
    .ZN(_11103_)
  );
  INV_X1 _18776_ (
    .A(_11103_),
    .ZN(_11104_)
  );
  AND2_X1 _18777_ (
    .A1(\rf[5] [10]),
    .A2(_08542_),
    .ZN(_11105_)
  );
  INV_X1 _18778_ (
    .A(_11105_),
    .ZN(_11106_)
  );
  AND2_X1 _18779_ (
    .A1(\rf[1] [10]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11107_)
  );
  INV_X1 _18780_ (
    .A(_11107_),
    .ZN(_11108_)
  );
  AND2_X1 _18781_ (
    .A1(_08540_),
    .A2(_11108_),
    .ZN(_11109_)
  );
  AND2_X1 _18782_ (
    .A1(_11106_),
    .A2(_11109_),
    .ZN(_11110_)
  );
  INV_X1 _18783_ (
    .A(_11110_),
    .ZN(_11111_)
  );
  AND2_X1 _18784_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_11111_),
    .ZN(_11112_)
  );
  AND2_X1 _18785_ (
    .A1(_11104_),
    .A2(_11112_),
    .ZN(_11113_)
  );
  INV_X1 _18786_ (
    .A(_11113_),
    .ZN(_11114_)
  );
  MUX2_X1 _18787_ (
    .A(\rf[13] [10]),
    .B(\rf[9] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11115_)
  );
  INV_X1 _18788_ (
    .A(_11115_),
    .ZN(_11116_)
  );
  AND2_X1 _18789_ (
    .A1(_08540_),
    .A2(_11116_),
    .ZN(_11117_)
  );
  INV_X1 _18790_ (
    .A(_11117_),
    .ZN(_11118_)
  );
  MUX2_X1 _18791_ (
    .A(\rf[12] [10]),
    .B(\rf[8] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11119_)
  );
  INV_X1 _18792_ (
    .A(_11119_),
    .ZN(_11120_)
  );
  AND2_X1 _18793_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_11120_),
    .ZN(_11121_)
  );
  INV_X1 _18794_ (
    .A(_11121_),
    .ZN(_11122_)
  );
  AND2_X1 _18795_ (
    .A1(_08543_),
    .A2(_11122_),
    .ZN(_11123_)
  );
  AND2_X1 _18796_ (
    .A1(_11118_),
    .A2(_11123_),
    .ZN(_11124_)
  );
  INV_X1 _18797_ (
    .A(_11124_),
    .ZN(_11125_)
  );
  AND2_X1 _18798_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11125_),
    .ZN(_11126_)
  );
  AND2_X1 _18799_ (
    .A1(_11114_),
    .A2(_11126_),
    .ZN(_11127_)
  );
  INV_X1 _18800_ (
    .A(_11127_),
    .ZN(_11128_)
  );
  AND2_X1 _18801_ (
    .A1(_11097_),
    .A2(_11128_),
    .ZN(_11129_)
  );
  AND2_X1 _18802_ (
    .A1(\rf[22] [10]),
    .A2(_08542_),
    .ZN(_11130_)
  );
  INV_X1 _18803_ (
    .A(_11130_),
    .ZN(_11131_)
  );
  AND2_X1 _18804_ (
    .A1(\rf[18] [10]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11132_)
  );
  INV_X1 _18805_ (
    .A(_11132_),
    .ZN(_11133_)
  );
  AND2_X1 _18806_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_11133_),
    .ZN(_11134_)
  );
  AND2_X1 _18807_ (
    .A1(_11131_),
    .A2(_11134_),
    .ZN(_11135_)
  );
  INV_X1 _18808_ (
    .A(_11135_),
    .ZN(_11136_)
  );
  AND2_X1 _18809_ (
    .A1(\rf[23] [10]),
    .A2(_08542_),
    .ZN(_11137_)
  );
  INV_X1 _18810_ (
    .A(_11137_),
    .ZN(_11138_)
  );
  AND2_X1 _18811_ (
    .A1(\rf[19] [10]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11139_)
  );
  INV_X1 _18812_ (
    .A(_11139_),
    .ZN(_11140_)
  );
  AND2_X1 _18813_ (
    .A1(_08540_),
    .A2(_11140_),
    .ZN(_11141_)
  );
  AND2_X1 _18814_ (
    .A1(_11138_),
    .A2(_11141_),
    .ZN(_11142_)
  );
  INV_X1 _18815_ (
    .A(_11142_),
    .ZN(_11143_)
  );
  AND2_X1 _18816_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_11143_),
    .ZN(_11144_)
  );
  AND2_X1 _18817_ (
    .A1(_11136_),
    .A2(_11144_),
    .ZN(_11145_)
  );
  INV_X1 _18818_ (
    .A(_11145_),
    .ZN(_11146_)
  );
  AND2_X1 _18819_ (
    .A1(_08498_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11147_)
  );
  INV_X1 _18820_ (
    .A(_11147_),
    .ZN(_11148_)
  );
  AND2_X1 _18821_ (
    .A1(_08471_),
    .A2(_08542_),
    .ZN(_11149_)
  );
  INV_X1 _18822_ (
    .A(_11149_),
    .ZN(_11150_)
  );
  AND2_X1 _18823_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_11150_),
    .ZN(_11151_)
  );
  AND2_X1 _18824_ (
    .A1(_11148_),
    .A2(_11151_),
    .ZN(_11152_)
  );
  INV_X1 _18825_ (
    .A(_11152_),
    .ZN(_11153_)
  );
  AND2_X1 _18826_ (
    .A1(\rf[27] [10]),
    .A2(_09608_),
    .ZN(_11154_)
  );
  INV_X1 _18827_ (
    .A(_11154_),
    .ZN(_11155_)
  );
  AND2_X1 _18828_ (
    .A1(_11153_),
    .A2(_11155_),
    .ZN(_11156_)
  );
  INV_X1 _18829_ (
    .A(_11156_),
    .ZN(_11157_)
  );
  AND2_X1 _18830_ (
    .A1(_08543_),
    .A2(_11157_),
    .ZN(_11158_)
  );
  INV_X1 _18831_ (
    .A(_11158_),
    .ZN(_11159_)
  );
  AND2_X1 _18832_ (
    .A1(_08541_),
    .A2(_11159_),
    .ZN(_11160_)
  );
  AND2_X1 _18833_ (
    .A1(_11146_),
    .A2(_11160_),
    .ZN(_11161_)
  );
  INV_X1 _18834_ (
    .A(_11161_),
    .ZN(_11162_)
  );
  MUX2_X1 _18835_ (
    .A(\rf[29] [10]),
    .B(\rf[28] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_11163_)
  );
  INV_X1 _18836_ (
    .A(_11163_),
    .ZN(_11164_)
  );
  AND2_X1 _18837_ (
    .A1(_08542_),
    .A2(_11164_),
    .ZN(_11165_)
  );
  INV_X1 _18838_ (
    .A(_11165_),
    .ZN(_11166_)
  );
  MUX2_X1 _18839_ (
    .A(\rf[25] [10]),
    .B(\rf[24] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_11167_)
  );
  INV_X1 _18840_ (
    .A(_11167_),
    .ZN(_11168_)
  );
  AND2_X1 _18841_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_11168_),
    .ZN(_11169_)
  );
  INV_X1 _18842_ (
    .A(_11169_),
    .ZN(_11170_)
  );
  AND2_X1 _18843_ (
    .A1(_08543_),
    .A2(_11170_),
    .ZN(_11171_)
  );
  AND2_X1 _18844_ (
    .A1(_11166_),
    .A2(_11171_),
    .ZN(_11172_)
  );
  INV_X1 _18845_ (
    .A(_11172_),
    .ZN(_11173_)
  );
  AND2_X1 _18846_ (
    .A1(\rf[20] [10]),
    .A2(_08542_),
    .ZN(_11174_)
  );
  INV_X1 _18847_ (
    .A(_11174_),
    .ZN(_11175_)
  );
  AND2_X1 _18848_ (
    .A1(\rf[16] [10]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11176_)
  );
  INV_X1 _18849_ (
    .A(_11176_),
    .ZN(_11177_)
  );
  AND2_X1 _18850_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_11177_),
    .ZN(_11178_)
  );
  AND2_X1 _18851_ (
    .A1(_11175_),
    .A2(_11178_),
    .ZN(_11179_)
  );
  INV_X1 _18852_ (
    .A(_11179_),
    .ZN(_11180_)
  );
  AND2_X1 _18853_ (
    .A1(\rf[21] [10]),
    .A2(_08542_),
    .ZN(_11181_)
  );
  INV_X1 _18854_ (
    .A(_11181_),
    .ZN(_11182_)
  );
  AND2_X1 _18855_ (
    .A1(\rf[17] [10]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11183_)
  );
  INV_X1 _18856_ (
    .A(_11183_),
    .ZN(_11184_)
  );
  AND2_X1 _18857_ (
    .A1(_08540_),
    .A2(_11184_),
    .ZN(_11185_)
  );
  AND2_X1 _18858_ (
    .A1(_11182_),
    .A2(_11185_),
    .ZN(_11186_)
  );
  INV_X1 _18859_ (
    .A(_11186_),
    .ZN(_11187_)
  );
  AND2_X1 _18860_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_11187_),
    .ZN(_11188_)
  );
  AND2_X1 _18861_ (
    .A1(_11180_),
    .A2(_11188_),
    .ZN(_11189_)
  );
  INV_X1 _18862_ (
    .A(_11189_),
    .ZN(_11190_)
  );
  AND2_X1 _18863_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11190_),
    .ZN(_11191_)
  );
  AND2_X1 _18864_ (
    .A1(_11173_),
    .A2(_11191_),
    .ZN(_11192_)
  );
  INV_X1 _18865_ (
    .A(_11192_),
    .ZN(_11193_)
  );
  AND2_X1 _18866_ (
    .A1(_11162_),
    .A2(_11193_),
    .ZN(_11194_)
  );
  MUX2_X1 _18867_ (
    .A(_11129_),
    .B(_11194_),
    .S(_08571_),
    .Z(_11195_)
  );
  MUX2_X1 _18868_ (
    .A(_11066_),
    .B(_11195_),
    .S(_10132_),
    .Z(_11196_)
  );
  AND2_X1 _18869_ (
    .A1(_10082_),
    .A2(_11196_),
    .ZN(_11197_)
  );
  INV_X1 _18870_ (
    .A(_11197_),
    .ZN(_11198_)
  );
  AND2_X1 _18871_ (
    .A1(_11063_),
    .A2(_11198_),
    .ZN(_11199_)
  );
  INV_X1 _18872_ (
    .A(_11199_),
    .ZN(_11200_)
  );
  MUX2_X1 _18873_ (
    .A(ex_reg_rs_msb_0[8]),
    .B(_11200_),
    .S(_10079_),
    .Z(_00075_)
  );
  AND2_X1 _18874_ (
    .A1(ibuf_io_inst_0_bits_raw[11]),
    .A2(_09295_),
    .ZN(_11201_)
  );
  INV_X1 _18875_ (
    .A(_11201_),
    .ZN(_11202_)
  );
  MUX2_X1 _18876_ (
    .A(csr_io_rw_rdata[11]),
    .B(wb_reg_wdata[11]),
    .S(_10134_),
    .Z(_11203_)
  );
  MUX2_X1 _18877_ (
    .A(div_io_resp_bits_data[11]),
    .B(_11203_),
    .S(_08649_),
    .Z(_11204_)
  );
  MUX2_X1 _18878_ (
    .A(_11204_),
    .B(io_dmem_resp_bits_data[11]),
    .S(_08631_),
    .Z(_11205_)
  );
  AND2_X1 _18879_ (
    .A1(_08241_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11206_)
  );
  INV_X1 _18880_ (
    .A(_11206_),
    .ZN(_11207_)
  );
  AND2_X1 _18881_ (
    .A1(_08464_),
    .A2(_08542_),
    .ZN(_11208_)
  );
  INV_X1 _18882_ (
    .A(_11208_),
    .ZN(_11209_)
  );
  AND2_X1 _18883_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11209_),
    .ZN(_11210_)
  );
  AND2_X1 _18884_ (
    .A1(_11207_),
    .A2(_11210_),
    .ZN(_11211_)
  );
  INV_X1 _18885_ (
    .A(_11211_),
    .ZN(_11212_)
  );
  AND2_X1 _18886_ (
    .A1(\rf[27] [11]),
    .A2(_10453_),
    .ZN(_11213_)
  );
  INV_X1 _18887_ (
    .A(_11213_),
    .ZN(_11214_)
  );
  MUX2_X1 _18888_ (
    .A(\rf[30] [11]),
    .B(\rf[26] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11215_)
  );
  AND2_X1 _18889_ (
    .A1(_08512_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11216_)
  );
  INV_X1 _18890_ (
    .A(_11216_),
    .ZN(_11217_)
  );
  AND2_X1 _18891_ (
    .A1(_08442_),
    .A2(_08542_),
    .ZN(_11218_)
  );
  INV_X1 _18892_ (
    .A(_11218_),
    .ZN(_11219_)
  );
  AND2_X1 _18893_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11217_),
    .ZN(_11220_)
  );
  AND2_X1 _18894_ (
    .A1(_11219_),
    .A2(_11220_),
    .ZN(_11221_)
  );
  INV_X1 _18895_ (
    .A(_11221_),
    .ZN(_11222_)
  );
  AND2_X1 _18896_ (
    .A1(_08541_),
    .A2(_11215_),
    .ZN(_11223_)
  );
  INV_X1 _18897_ (
    .A(_11223_),
    .ZN(_11224_)
  );
  AND2_X1 _18898_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_11224_),
    .ZN(_11225_)
  );
  AND2_X1 _18899_ (
    .A1(_11222_),
    .A2(_11225_),
    .ZN(_11226_)
  );
  INV_X1 _18900_ (
    .A(_11226_),
    .ZN(_11227_)
  );
  AND2_X1 _18901_ (
    .A1(_08540_),
    .A2(_11214_),
    .ZN(_11228_)
  );
  AND2_X1 _18902_ (
    .A1(_11212_),
    .A2(_11228_),
    .ZN(_11229_)
  );
  INV_X1 _18903_ (
    .A(_11229_),
    .ZN(_11230_)
  );
  AND2_X1 _18904_ (
    .A1(_11227_),
    .A2(_11230_),
    .ZN(_11231_)
  );
  AND2_X1 _18905_ (
    .A1(_08543_),
    .A2(_11231_),
    .ZN(_11232_)
  );
  INV_X1 _18906_ (
    .A(_11232_),
    .ZN(_11233_)
  );
  AND2_X1 _18907_ (
    .A1(_08384_),
    .A2(_08542_),
    .ZN(_11234_)
  );
  INV_X1 _18908_ (
    .A(_11234_),
    .ZN(_11235_)
  );
  AND2_X1 _18909_ (
    .A1(_08285_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11236_)
  );
  INV_X1 _18910_ (
    .A(_11236_),
    .ZN(_11237_)
  );
  AND2_X1 _18911_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11237_),
    .ZN(_11238_)
  );
  AND2_X1 _18912_ (
    .A1(_11235_),
    .A2(_11238_),
    .ZN(_11239_)
  );
  INV_X1 _18913_ (
    .A(_11239_),
    .ZN(_11240_)
  );
  MUX2_X1 _18914_ (
    .A(\rf[22] [11]),
    .B(\rf[18] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11241_)
  );
  AND2_X1 _18915_ (
    .A1(_08541_),
    .A2(_11241_),
    .ZN(_11242_)
  );
  INV_X1 _18916_ (
    .A(_11242_),
    .ZN(_11243_)
  );
  AND2_X1 _18917_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_11243_),
    .ZN(_11244_)
  );
  AND2_X1 _18918_ (
    .A1(_11240_),
    .A2(_11244_),
    .ZN(_11245_)
  );
  INV_X1 _18919_ (
    .A(_11245_),
    .ZN(_11246_)
  );
  AND2_X1 _18920_ (
    .A1(_08315_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11247_)
  );
  INV_X1 _18921_ (
    .A(_11247_),
    .ZN(_11248_)
  );
  AND2_X1 _18922_ (
    .A1(_08414_),
    .A2(_08542_),
    .ZN(_11249_)
  );
  INV_X1 _18923_ (
    .A(_11249_),
    .ZN(_11250_)
  );
  AND2_X1 _18924_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11250_),
    .ZN(_11251_)
  );
  AND2_X1 _18925_ (
    .A1(_11248_),
    .A2(_11251_),
    .ZN(_11252_)
  );
  INV_X1 _18926_ (
    .A(_11252_),
    .ZN(_11253_)
  );
  MUX2_X1 _18927_ (
    .A(\rf[23] [11]),
    .B(\rf[19] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11254_)
  );
  AND2_X1 _18928_ (
    .A1(_08541_),
    .A2(_11254_),
    .ZN(_11255_)
  );
  INV_X1 _18929_ (
    .A(_11255_),
    .ZN(_11256_)
  );
  AND2_X1 _18930_ (
    .A1(_08540_),
    .A2(_11256_),
    .ZN(_11257_)
  );
  AND2_X1 _18931_ (
    .A1(_11253_),
    .A2(_11257_),
    .ZN(_11258_)
  );
  INV_X1 _18932_ (
    .A(_11258_),
    .ZN(_11259_)
  );
  AND2_X1 _18933_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_11259_),
    .ZN(_11260_)
  );
  AND2_X1 _18934_ (
    .A1(_11246_),
    .A2(_11260_),
    .ZN(_11261_)
  );
  INV_X1 _18935_ (
    .A(_11261_),
    .ZN(_11262_)
  );
  AND2_X1 _18936_ (
    .A1(_08571_),
    .A2(_11262_),
    .ZN(_11263_)
  );
  AND2_X1 _18937_ (
    .A1(_11233_),
    .A2(_11263_),
    .ZN(_11264_)
  );
  INV_X1 _18938_ (
    .A(_11264_),
    .ZN(_11265_)
  );
  MUX2_X1 _18939_ (
    .A(\rf[1] [11]),
    .B(\rf[0] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_11266_)
  );
  MUX2_X1 _18940_ (
    .A(\rf[5] [11]),
    .B(\rf[4] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_11267_)
  );
  MUX2_X1 _18941_ (
    .A(_11266_),
    .B(_11267_),
    .S(_08542_),
    .Z(_11268_)
  );
  INV_X1 _18942_ (
    .A(_11268_),
    .ZN(_11269_)
  );
  AND2_X1 _18943_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_11269_),
    .ZN(_11270_)
  );
  INV_X1 _18944_ (
    .A(_11270_),
    .ZN(_11271_)
  );
  MUX2_X1 _18945_ (
    .A(\rf[12] [11]),
    .B(\rf[8] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11272_)
  );
  INV_X1 _18946_ (
    .A(_11272_),
    .ZN(_11273_)
  );
  AND2_X1 _18947_ (
    .A1(_10213_),
    .A2(_11273_),
    .ZN(_11274_)
  );
  INV_X1 _18948_ (
    .A(_11274_),
    .ZN(_11275_)
  );
  MUX2_X1 _18949_ (
    .A(\rf[13] [11]),
    .B(\rf[9] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11276_)
  );
  INV_X1 _18950_ (
    .A(_11276_),
    .ZN(_11277_)
  );
  AND2_X1 _18951_ (
    .A1(_09110_),
    .A2(_11277_),
    .ZN(_11278_)
  );
  INV_X1 _18952_ (
    .A(_11278_),
    .ZN(_11279_)
  );
  AND2_X1 _18953_ (
    .A1(_11275_),
    .A2(_11279_),
    .ZN(_11280_)
  );
  AND2_X1 _18954_ (
    .A1(_11271_),
    .A2(_11280_),
    .ZN(_11281_)
  );
  AND2_X1 _18955_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11281_),
    .ZN(_11282_)
  );
  INV_X1 _18956_ (
    .A(_11282_),
    .ZN(_11283_)
  );
  MUX2_X1 _18957_ (
    .A(\rf[3] [11]),
    .B(\rf[2] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_11284_)
  );
  MUX2_X1 _18958_ (
    .A(\rf[7] [11]),
    .B(\rf[6] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_11285_)
  );
  MUX2_X1 _18959_ (
    .A(_11284_),
    .B(_11285_),
    .S(_08542_),
    .Z(_11286_)
  );
  INV_X1 _18960_ (
    .A(_11286_),
    .ZN(_11287_)
  );
  AND2_X1 _18961_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_11287_),
    .ZN(_11288_)
  );
  INV_X1 _18962_ (
    .A(_11288_),
    .ZN(_11289_)
  );
  MUX2_X1 _18963_ (
    .A(\rf[14] [11]),
    .B(\rf[10] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11290_)
  );
  INV_X1 _18964_ (
    .A(_11290_),
    .ZN(_11291_)
  );
  AND2_X1 _18965_ (
    .A1(_10213_),
    .A2(_11291_),
    .ZN(_11292_)
  );
  INV_X1 _18966_ (
    .A(_11292_),
    .ZN(_11293_)
  );
  MUX2_X1 _18967_ (
    .A(\rf[15] [11]),
    .B(\rf[11] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11294_)
  );
  INV_X1 _18968_ (
    .A(_11294_),
    .ZN(_11295_)
  );
  AND2_X1 _18969_ (
    .A1(_09110_),
    .A2(_11295_),
    .ZN(_11296_)
  );
  INV_X1 _18970_ (
    .A(_11296_),
    .ZN(_11297_)
  );
  AND2_X1 _18971_ (
    .A1(_11293_),
    .A2(_11297_),
    .ZN(_11298_)
  );
  AND2_X1 _18972_ (
    .A1(_11289_),
    .A2(_11298_),
    .ZN(_11299_)
  );
  AND2_X1 _18973_ (
    .A1(_08541_),
    .A2(_11299_),
    .ZN(_11300_)
  );
  INV_X1 _18974_ (
    .A(_11300_),
    .ZN(_11301_)
  );
  AND2_X1 _18975_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_11283_),
    .ZN(_11302_)
  );
  AND2_X1 _18976_ (
    .A1(_11301_),
    .A2(_11302_),
    .ZN(_11303_)
  );
  INV_X1 _18977_ (
    .A(_11303_),
    .ZN(_11304_)
  );
  AND2_X1 _18978_ (
    .A1(_11265_),
    .A2(_11304_),
    .ZN(_11305_)
  );
  MUX2_X1 _18979_ (
    .A(_11205_),
    .B(_11305_),
    .S(_10132_),
    .Z(_11306_)
  );
  AND2_X1 _18980_ (
    .A1(_10082_),
    .A2(_11306_),
    .ZN(_11307_)
  );
  INV_X1 _18981_ (
    .A(_11307_),
    .ZN(_11308_)
  );
  AND2_X1 _18982_ (
    .A1(_11202_),
    .A2(_11308_),
    .ZN(_11309_)
  );
  INV_X1 _18983_ (
    .A(_11309_),
    .ZN(_11310_)
  );
  MUX2_X1 _18984_ (
    .A(ex_reg_rs_msb_0[9]),
    .B(_11310_),
    .S(_10079_),
    .Z(_00076_)
  );
  AND2_X1 _18985_ (
    .A1(ibuf_io_inst_0_bits_raw[12]),
    .A2(_09295_),
    .ZN(_11311_)
  );
  INV_X1 _18986_ (
    .A(_11311_),
    .ZN(_11312_)
  );
  MUX2_X1 _18987_ (
    .A(csr_io_rw_rdata[12]),
    .B(wb_reg_wdata[12]),
    .S(_10134_),
    .Z(_11313_)
  );
  MUX2_X1 _18988_ (
    .A(div_io_resp_bits_data[12]),
    .B(_11313_),
    .S(_08649_),
    .Z(_11314_)
  );
  MUX2_X1 _18989_ (
    .A(_11314_),
    .B(io_dmem_resp_bits_data[12]),
    .S(_08631_),
    .Z(_11315_)
  );
  MUX2_X1 _18990_ (
    .A(\rf[3] [12]),
    .B(\rf[1] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_11316_)
  );
  MUX2_X1 _18991_ (
    .A(\rf[7] [12]),
    .B(\rf[5] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_11317_)
  );
  MUX2_X1 _18992_ (
    .A(_11316_),
    .B(_11317_),
    .S(_08542_),
    .Z(_11318_)
  );
  AND2_X1 _18993_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_11318_),
    .ZN(_11319_)
  );
  INV_X1 _18994_ (
    .A(_11319_),
    .ZN(_11320_)
  );
  MUX2_X1 _18995_ (
    .A(\rf[13] [12]),
    .B(\rf[9] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11321_)
  );
  INV_X1 _18996_ (
    .A(_11321_),
    .ZN(_11322_)
  );
  AND2_X1 _18997_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11322_),
    .ZN(_11323_)
  );
  INV_X1 _18998_ (
    .A(_11323_),
    .ZN(_11324_)
  );
  MUX2_X1 _18999_ (
    .A(\rf[15] [12]),
    .B(\rf[11] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11325_)
  );
  INV_X1 _19000_ (
    .A(_11325_),
    .ZN(_11326_)
  );
  AND2_X1 _19001_ (
    .A1(_08541_),
    .A2(_11326_),
    .ZN(_11327_)
  );
  INV_X1 _19002_ (
    .A(_11327_),
    .ZN(_11328_)
  );
  AND2_X1 _19003_ (
    .A1(_08543_),
    .A2(_11328_),
    .ZN(_11329_)
  );
  AND2_X1 _19004_ (
    .A1(_11324_),
    .A2(_11329_),
    .ZN(_11330_)
  );
  INV_X1 _19005_ (
    .A(_11330_),
    .ZN(_11331_)
  );
  AND2_X1 _19006_ (
    .A1(_08540_),
    .A2(_11331_),
    .ZN(_11332_)
  );
  AND2_X1 _19007_ (
    .A1(_11320_),
    .A2(_11332_),
    .ZN(_11333_)
  );
  INV_X1 _19008_ (
    .A(_11333_),
    .ZN(_11334_)
  );
  MUX2_X1 _19009_ (
    .A(\rf[2] [12]),
    .B(\rf[0] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_11335_)
  );
  MUX2_X1 _19010_ (
    .A(\rf[6] [12]),
    .B(\rf[4] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_11336_)
  );
  MUX2_X1 _19011_ (
    .A(_11335_),
    .B(_11336_),
    .S(_08542_),
    .Z(_11337_)
  );
  AND2_X1 _19012_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_11337_),
    .ZN(_11338_)
  );
  INV_X1 _19013_ (
    .A(_11338_),
    .ZN(_11339_)
  );
  MUX2_X1 _19014_ (
    .A(\rf[12] [12]),
    .B(\rf[8] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11340_)
  );
  INV_X1 _19015_ (
    .A(_11340_),
    .ZN(_11341_)
  );
  AND2_X1 _19016_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11341_),
    .ZN(_11342_)
  );
  INV_X1 _19017_ (
    .A(_11342_),
    .ZN(_11343_)
  );
  MUX2_X1 _19018_ (
    .A(\rf[14] [12]),
    .B(\rf[10] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11344_)
  );
  INV_X1 _19019_ (
    .A(_11344_),
    .ZN(_11345_)
  );
  AND2_X1 _19020_ (
    .A1(_08541_),
    .A2(_11345_),
    .ZN(_11346_)
  );
  INV_X1 _19021_ (
    .A(_11346_),
    .ZN(_11347_)
  );
  AND2_X1 _19022_ (
    .A1(_08543_),
    .A2(_11347_),
    .ZN(_11348_)
  );
  AND2_X1 _19023_ (
    .A1(_11343_),
    .A2(_11348_),
    .ZN(_11349_)
  );
  INV_X1 _19024_ (
    .A(_11349_),
    .ZN(_11350_)
  );
  AND2_X1 _19025_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_11350_),
    .ZN(_11351_)
  );
  AND2_X1 _19026_ (
    .A1(_11339_),
    .A2(_11351_),
    .ZN(_11352_)
  );
  INV_X1 _19027_ (
    .A(_11352_),
    .ZN(_11353_)
  );
  AND2_X1 _19028_ (
    .A1(_11334_),
    .A2(_11353_),
    .ZN(_11354_)
  );
  INV_X1 _19029_ (
    .A(_11354_),
    .ZN(_11355_)
  );
  AND2_X1 _19030_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_11355_),
    .ZN(_11356_)
  );
  INV_X1 _19031_ (
    .A(_11356_),
    .ZN(_11357_)
  );
  AND2_X1 _19032_ (
    .A1(_08242_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11358_)
  );
  INV_X1 _19033_ (
    .A(_11358_),
    .ZN(_11359_)
  );
  AND2_X1 _19034_ (
    .A1(_08465_),
    .A2(_08542_),
    .ZN(_11360_)
  );
  INV_X1 _19035_ (
    .A(_11360_),
    .ZN(_11361_)
  );
  AND2_X1 _19036_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11361_),
    .ZN(_11362_)
  );
  AND2_X1 _19037_ (
    .A1(_11359_),
    .A2(_11362_),
    .ZN(_11363_)
  );
  INV_X1 _19038_ (
    .A(_11363_),
    .ZN(_11364_)
  );
  AND2_X1 _19039_ (
    .A1(\rf[27] [12]),
    .A2(_10453_),
    .ZN(_11365_)
  );
  INV_X1 _19040_ (
    .A(_11365_),
    .ZN(_11366_)
  );
  MUX2_X1 _19041_ (
    .A(\rf[30] [12]),
    .B(\rf[26] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11367_)
  );
  AND2_X1 _19042_ (
    .A1(_08513_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11368_)
  );
  INV_X1 _19043_ (
    .A(_11368_),
    .ZN(_11369_)
  );
  AND2_X1 _19044_ (
    .A1(_08443_),
    .A2(_08542_),
    .ZN(_11370_)
  );
  INV_X1 _19045_ (
    .A(_11370_),
    .ZN(_11371_)
  );
  AND2_X1 _19046_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11369_),
    .ZN(_11372_)
  );
  AND2_X1 _19047_ (
    .A1(_11371_),
    .A2(_11372_),
    .ZN(_11373_)
  );
  INV_X1 _19048_ (
    .A(_11373_),
    .ZN(_11374_)
  );
  AND2_X1 _19049_ (
    .A1(_08541_),
    .A2(_11367_),
    .ZN(_11375_)
  );
  INV_X1 _19050_ (
    .A(_11375_),
    .ZN(_11376_)
  );
  AND2_X1 _19051_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_11376_),
    .ZN(_11377_)
  );
  AND2_X1 _19052_ (
    .A1(_11374_),
    .A2(_11377_),
    .ZN(_11378_)
  );
  INV_X1 _19053_ (
    .A(_11378_),
    .ZN(_11379_)
  );
  AND2_X1 _19054_ (
    .A1(_08540_),
    .A2(_11366_),
    .ZN(_11380_)
  );
  AND2_X1 _19055_ (
    .A1(_11364_),
    .A2(_11380_),
    .ZN(_11381_)
  );
  INV_X1 _19056_ (
    .A(_11381_),
    .ZN(_11382_)
  );
  AND2_X1 _19057_ (
    .A1(_11379_),
    .A2(_11382_),
    .ZN(_11383_)
  );
  AND2_X1 _19058_ (
    .A1(_08543_),
    .A2(_11383_),
    .ZN(_11384_)
  );
  INV_X1 _19059_ (
    .A(_11384_),
    .ZN(_11385_)
  );
  AND2_X1 _19060_ (
    .A1(_08385_),
    .A2(_08542_),
    .ZN(_11386_)
  );
  INV_X1 _19061_ (
    .A(_11386_),
    .ZN(_11387_)
  );
  AND2_X1 _19062_ (
    .A1(_08286_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11388_)
  );
  INV_X1 _19063_ (
    .A(_11388_),
    .ZN(_11389_)
  );
  AND2_X1 _19064_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11389_),
    .ZN(_11390_)
  );
  AND2_X1 _19065_ (
    .A1(_11387_),
    .A2(_11390_),
    .ZN(_11391_)
  );
  INV_X1 _19066_ (
    .A(_11391_),
    .ZN(_11392_)
  );
  MUX2_X1 _19067_ (
    .A(\rf[22] [12]),
    .B(\rf[18] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11393_)
  );
  AND2_X1 _19068_ (
    .A1(_08541_),
    .A2(_11393_),
    .ZN(_11394_)
  );
  INV_X1 _19069_ (
    .A(_11394_),
    .ZN(_11395_)
  );
  AND2_X1 _19070_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_11395_),
    .ZN(_11396_)
  );
  AND2_X1 _19071_ (
    .A1(_11392_),
    .A2(_11396_),
    .ZN(_11397_)
  );
  INV_X1 _19072_ (
    .A(_11397_),
    .ZN(_11398_)
  );
  AND2_X1 _19073_ (
    .A1(_08316_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11399_)
  );
  INV_X1 _19074_ (
    .A(_11399_),
    .ZN(_11400_)
  );
  AND2_X1 _19075_ (
    .A1(_08415_),
    .A2(_08542_),
    .ZN(_11401_)
  );
  INV_X1 _19076_ (
    .A(_11401_),
    .ZN(_11402_)
  );
  AND2_X1 _19077_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11402_),
    .ZN(_11403_)
  );
  AND2_X1 _19078_ (
    .A1(_11400_),
    .A2(_11403_),
    .ZN(_11404_)
  );
  INV_X1 _19079_ (
    .A(_11404_),
    .ZN(_11405_)
  );
  MUX2_X1 _19080_ (
    .A(\rf[23] [12]),
    .B(\rf[19] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11406_)
  );
  AND2_X1 _19081_ (
    .A1(_08541_),
    .A2(_11406_),
    .ZN(_11407_)
  );
  INV_X1 _19082_ (
    .A(_11407_),
    .ZN(_11408_)
  );
  AND2_X1 _19083_ (
    .A1(_08540_),
    .A2(_11408_),
    .ZN(_11409_)
  );
  AND2_X1 _19084_ (
    .A1(_11405_),
    .A2(_11409_),
    .ZN(_11410_)
  );
  INV_X1 _19085_ (
    .A(_11410_),
    .ZN(_11411_)
  );
  AND2_X1 _19086_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_11411_),
    .ZN(_11412_)
  );
  AND2_X1 _19087_ (
    .A1(_11398_),
    .A2(_11412_),
    .ZN(_11413_)
  );
  INV_X1 _19088_ (
    .A(_11413_),
    .ZN(_11414_)
  );
  AND2_X1 _19089_ (
    .A1(_08571_),
    .A2(_11414_),
    .ZN(_11415_)
  );
  AND2_X1 _19090_ (
    .A1(_11385_),
    .A2(_11415_),
    .ZN(_11416_)
  );
  INV_X1 _19091_ (
    .A(_11416_),
    .ZN(_11417_)
  );
  AND2_X1 _19092_ (
    .A1(_11357_),
    .A2(_11417_),
    .ZN(_11418_)
  );
  MUX2_X1 _19093_ (
    .A(_11315_),
    .B(_11418_),
    .S(_10132_),
    .Z(_11419_)
  );
  AND2_X1 _19094_ (
    .A1(_10082_),
    .A2(_11419_),
    .ZN(_11420_)
  );
  INV_X1 _19095_ (
    .A(_11420_),
    .ZN(_11421_)
  );
  AND2_X1 _19096_ (
    .A1(_11312_),
    .A2(_11421_),
    .ZN(_11422_)
  );
  INV_X1 _19097_ (
    .A(_11422_),
    .ZN(_11423_)
  );
  MUX2_X1 _19098_ (
    .A(ex_reg_rs_msb_0[10]),
    .B(_11423_),
    .S(_10079_),
    .Z(_00077_)
  );
  AND2_X1 _19099_ (
    .A1(ibuf_io_inst_0_bits_raw[13]),
    .A2(_09295_),
    .ZN(_11424_)
  );
  INV_X1 _19100_ (
    .A(_11424_),
    .ZN(_11425_)
  );
  MUX2_X1 _19101_ (
    .A(csr_io_rw_rdata[13]),
    .B(wb_reg_wdata[13]),
    .S(_10134_),
    .Z(_11426_)
  );
  MUX2_X1 _19102_ (
    .A(div_io_resp_bits_data[13]),
    .B(_11426_),
    .S(_08649_),
    .Z(_11427_)
  );
  MUX2_X1 _19103_ (
    .A(_11427_),
    .B(io_dmem_resp_bits_data[13]),
    .S(_08631_),
    .Z(_11428_)
  );
  MUX2_X1 _19104_ (
    .A(\rf[3] [13]),
    .B(\rf[1] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_11429_)
  );
  MUX2_X1 _19105_ (
    .A(\rf[7] [13]),
    .B(\rf[5] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_11430_)
  );
  MUX2_X1 _19106_ (
    .A(_11429_),
    .B(_11430_),
    .S(_08542_),
    .Z(_11431_)
  );
  AND2_X1 _19107_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_11431_),
    .ZN(_11432_)
  );
  INV_X1 _19108_ (
    .A(_11432_),
    .ZN(_11433_)
  );
  MUX2_X1 _19109_ (
    .A(\rf[13] [13]),
    .B(\rf[9] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11434_)
  );
  INV_X1 _19110_ (
    .A(_11434_),
    .ZN(_11435_)
  );
  AND2_X1 _19111_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11435_),
    .ZN(_11436_)
  );
  INV_X1 _19112_ (
    .A(_11436_),
    .ZN(_11437_)
  );
  MUX2_X1 _19113_ (
    .A(\rf[15] [13]),
    .B(\rf[11] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11438_)
  );
  INV_X1 _19114_ (
    .A(_11438_),
    .ZN(_11439_)
  );
  AND2_X1 _19115_ (
    .A1(_08541_),
    .A2(_11439_),
    .ZN(_11440_)
  );
  INV_X1 _19116_ (
    .A(_11440_),
    .ZN(_11441_)
  );
  AND2_X1 _19117_ (
    .A1(_08543_),
    .A2(_11441_),
    .ZN(_11442_)
  );
  AND2_X1 _19118_ (
    .A1(_11437_),
    .A2(_11442_),
    .ZN(_11443_)
  );
  INV_X1 _19119_ (
    .A(_11443_),
    .ZN(_11444_)
  );
  AND2_X1 _19120_ (
    .A1(_08540_),
    .A2(_11444_),
    .ZN(_11445_)
  );
  AND2_X1 _19121_ (
    .A1(_11433_),
    .A2(_11445_),
    .ZN(_11446_)
  );
  INV_X1 _19122_ (
    .A(_11446_),
    .ZN(_11447_)
  );
  MUX2_X1 _19123_ (
    .A(\rf[2] [13]),
    .B(\rf[0] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_11448_)
  );
  MUX2_X1 _19124_ (
    .A(\rf[6] [13]),
    .B(\rf[4] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_11449_)
  );
  MUX2_X1 _19125_ (
    .A(_11448_),
    .B(_11449_),
    .S(_08542_),
    .Z(_11450_)
  );
  AND2_X1 _19126_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_11450_),
    .ZN(_11451_)
  );
  INV_X1 _19127_ (
    .A(_11451_),
    .ZN(_11452_)
  );
  MUX2_X1 _19128_ (
    .A(\rf[12] [13]),
    .B(\rf[8] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11453_)
  );
  INV_X1 _19129_ (
    .A(_11453_),
    .ZN(_11454_)
  );
  AND2_X1 _19130_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11454_),
    .ZN(_11455_)
  );
  INV_X1 _19131_ (
    .A(_11455_),
    .ZN(_11456_)
  );
  MUX2_X1 _19132_ (
    .A(\rf[14] [13]),
    .B(\rf[10] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11457_)
  );
  INV_X1 _19133_ (
    .A(_11457_),
    .ZN(_11458_)
  );
  AND2_X1 _19134_ (
    .A1(_08541_),
    .A2(_11458_),
    .ZN(_11459_)
  );
  INV_X1 _19135_ (
    .A(_11459_),
    .ZN(_11460_)
  );
  AND2_X1 _19136_ (
    .A1(_08543_),
    .A2(_11460_),
    .ZN(_11461_)
  );
  AND2_X1 _19137_ (
    .A1(_11456_),
    .A2(_11461_),
    .ZN(_11462_)
  );
  INV_X1 _19138_ (
    .A(_11462_),
    .ZN(_11463_)
  );
  AND2_X1 _19139_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_11463_),
    .ZN(_11464_)
  );
  AND2_X1 _19140_ (
    .A1(_11452_),
    .A2(_11464_),
    .ZN(_11465_)
  );
  INV_X1 _19141_ (
    .A(_11465_),
    .ZN(_11466_)
  );
  AND2_X1 _19142_ (
    .A1(_11447_),
    .A2(_11466_),
    .ZN(_11467_)
  );
  INV_X1 _19143_ (
    .A(_11467_),
    .ZN(_11468_)
  );
  AND2_X1 _19144_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_11468_),
    .ZN(_11469_)
  );
  INV_X1 _19145_ (
    .A(_11469_),
    .ZN(_11470_)
  );
  AND2_X1 _19146_ (
    .A1(_08243_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11471_)
  );
  INV_X1 _19147_ (
    .A(_11471_),
    .ZN(_11472_)
  );
  AND2_X1 _19148_ (
    .A1(_08466_),
    .A2(_08542_),
    .ZN(_11473_)
  );
  INV_X1 _19149_ (
    .A(_11473_),
    .ZN(_11474_)
  );
  AND2_X1 _19150_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11474_),
    .ZN(_11475_)
  );
  AND2_X1 _19151_ (
    .A1(_11472_),
    .A2(_11475_),
    .ZN(_11476_)
  );
  INV_X1 _19152_ (
    .A(_11476_),
    .ZN(_11477_)
  );
  AND2_X1 _19153_ (
    .A1(\rf[27] [13]),
    .A2(_10453_),
    .ZN(_11478_)
  );
  INV_X1 _19154_ (
    .A(_11478_),
    .ZN(_11479_)
  );
  MUX2_X1 _19155_ (
    .A(\rf[30] [13]),
    .B(\rf[26] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11480_)
  );
  AND2_X1 _19156_ (
    .A1(_08514_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11481_)
  );
  INV_X1 _19157_ (
    .A(_11481_),
    .ZN(_11482_)
  );
  AND2_X1 _19158_ (
    .A1(_08444_),
    .A2(_08542_),
    .ZN(_11483_)
  );
  INV_X1 _19159_ (
    .A(_11483_),
    .ZN(_11484_)
  );
  AND2_X1 _19160_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11482_),
    .ZN(_11485_)
  );
  AND2_X1 _19161_ (
    .A1(_11484_),
    .A2(_11485_),
    .ZN(_11486_)
  );
  INV_X1 _19162_ (
    .A(_11486_),
    .ZN(_11487_)
  );
  AND2_X1 _19163_ (
    .A1(_08541_),
    .A2(_11480_),
    .ZN(_11488_)
  );
  INV_X1 _19164_ (
    .A(_11488_),
    .ZN(_11489_)
  );
  AND2_X1 _19165_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_11489_),
    .ZN(_11490_)
  );
  AND2_X1 _19166_ (
    .A1(_11487_),
    .A2(_11490_),
    .ZN(_11491_)
  );
  INV_X1 _19167_ (
    .A(_11491_),
    .ZN(_11492_)
  );
  AND2_X1 _19168_ (
    .A1(_08540_),
    .A2(_11479_),
    .ZN(_11493_)
  );
  AND2_X1 _19169_ (
    .A1(_11477_),
    .A2(_11493_),
    .ZN(_11494_)
  );
  INV_X1 _19170_ (
    .A(_11494_),
    .ZN(_11495_)
  );
  AND2_X1 _19171_ (
    .A1(_11492_),
    .A2(_11495_),
    .ZN(_11496_)
  );
  AND2_X1 _19172_ (
    .A1(_08543_),
    .A2(_11496_),
    .ZN(_11497_)
  );
  INV_X1 _19173_ (
    .A(_11497_),
    .ZN(_11498_)
  );
  AND2_X1 _19174_ (
    .A1(_08386_),
    .A2(_08542_),
    .ZN(_11499_)
  );
  INV_X1 _19175_ (
    .A(_11499_),
    .ZN(_11500_)
  );
  AND2_X1 _19176_ (
    .A1(_08287_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11501_)
  );
  INV_X1 _19177_ (
    .A(_11501_),
    .ZN(_11502_)
  );
  AND2_X1 _19178_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11502_),
    .ZN(_11503_)
  );
  AND2_X1 _19179_ (
    .A1(_11500_),
    .A2(_11503_),
    .ZN(_11504_)
  );
  INV_X1 _19180_ (
    .A(_11504_),
    .ZN(_11505_)
  );
  MUX2_X1 _19181_ (
    .A(\rf[22] [13]),
    .B(\rf[18] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11506_)
  );
  AND2_X1 _19182_ (
    .A1(_08541_),
    .A2(_11506_),
    .ZN(_11507_)
  );
  INV_X1 _19183_ (
    .A(_11507_),
    .ZN(_11508_)
  );
  AND2_X1 _19184_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_11508_),
    .ZN(_11509_)
  );
  AND2_X1 _19185_ (
    .A1(_11505_),
    .A2(_11509_),
    .ZN(_11510_)
  );
  INV_X1 _19186_ (
    .A(_11510_),
    .ZN(_11511_)
  );
  AND2_X1 _19187_ (
    .A1(_08317_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11512_)
  );
  INV_X1 _19188_ (
    .A(_11512_),
    .ZN(_11513_)
  );
  AND2_X1 _19189_ (
    .A1(_08416_),
    .A2(_08542_),
    .ZN(_11514_)
  );
  INV_X1 _19190_ (
    .A(_11514_),
    .ZN(_11515_)
  );
  AND2_X1 _19191_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11515_),
    .ZN(_11516_)
  );
  AND2_X1 _19192_ (
    .A1(_11513_),
    .A2(_11516_),
    .ZN(_11517_)
  );
  INV_X1 _19193_ (
    .A(_11517_),
    .ZN(_11518_)
  );
  MUX2_X1 _19194_ (
    .A(\rf[23] [13]),
    .B(\rf[19] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11519_)
  );
  AND2_X1 _19195_ (
    .A1(_08541_),
    .A2(_11519_),
    .ZN(_11520_)
  );
  INV_X1 _19196_ (
    .A(_11520_),
    .ZN(_11521_)
  );
  AND2_X1 _19197_ (
    .A1(_08540_),
    .A2(_11521_),
    .ZN(_11522_)
  );
  AND2_X1 _19198_ (
    .A1(_11518_),
    .A2(_11522_),
    .ZN(_11523_)
  );
  INV_X1 _19199_ (
    .A(_11523_),
    .ZN(_11524_)
  );
  AND2_X1 _19200_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_11524_),
    .ZN(_11525_)
  );
  AND2_X1 _19201_ (
    .A1(_11511_),
    .A2(_11525_),
    .ZN(_11526_)
  );
  INV_X1 _19202_ (
    .A(_11526_),
    .ZN(_11527_)
  );
  AND2_X1 _19203_ (
    .A1(_08571_),
    .A2(_11527_),
    .ZN(_11528_)
  );
  AND2_X1 _19204_ (
    .A1(_11498_),
    .A2(_11528_),
    .ZN(_11529_)
  );
  INV_X1 _19205_ (
    .A(_11529_),
    .ZN(_11530_)
  );
  AND2_X1 _19206_ (
    .A1(_11470_),
    .A2(_11530_),
    .ZN(_11531_)
  );
  MUX2_X1 _19207_ (
    .A(_11428_),
    .B(_11531_),
    .S(_10132_),
    .Z(_11532_)
  );
  AND2_X1 _19208_ (
    .A1(_10082_),
    .A2(_11532_),
    .ZN(_11533_)
  );
  INV_X1 _19209_ (
    .A(_11533_),
    .ZN(_11534_)
  );
  AND2_X1 _19210_ (
    .A1(_11425_),
    .A2(_11534_),
    .ZN(_11535_)
  );
  INV_X1 _19211_ (
    .A(_11535_),
    .ZN(_11536_)
  );
  MUX2_X1 _19212_ (
    .A(ex_reg_rs_msb_0[11]),
    .B(_11536_),
    .S(_10079_),
    .Z(_00078_)
  );
  AND2_X1 _19213_ (
    .A1(ibuf_io_inst_0_bits_raw[14]),
    .A2(_09295_),
    .ZN(_11537_)
  );
  INV_X1 _19214_ (
    .A(_11537_),
    .ZN(_11538_)
  );
  MUX2_X1 _19215_ (
    .A(csr_io_rw_rdata[14]),
    .B(wb_reg_wdata[14]),
    .S(_10134_),
    .Z(_11539_)
  );
  MUX2_X1 _19216_ (
    .A(div_io_resp_bits_data[14]),
    .B(_11539_),
    .S(_08649_),
    .Z(_11540_)
  );
  MUX2_X1 _19217_ (
    .A(_11540_),
    .B(io_dmem_resp_bits_data[14]),
    .S(_08631_),
    .Z(_11541_)
  );
  MUX2_X1 _19218_ (
    .A(\rf[5] [14]),
    .B(\rf[1] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11542_)
  );
  MUX2_X1 _19219_ (
    .A(\rf[7] [14]),
    .B(\rf[3] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11543_)
  );
  MUX2_X1 _19220_ (
    .A(_11542_),
    .B(_11543_),
    .S(_08541_),
    .Z(_11544_)
  );
  AND2_X1 _19221_ (
    .A1(_08540_),
    .A2(_11544_),
    .ZN(_11545_)
  );
  INV_X1 _19222_ (
    .A(_11545_),
    .ZN(_11546_)
  );
  MUX2_X1 _19223_ (
    .A(\rf[4] [14]),
    .B(\rf[0] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11547_)
  );
  MUX2_X1 _19224_ (
    .A(\rf[6] [14]),
    .B(\rf[2] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11548_)
  );
  MUX2_X1 _19225_ (
    .A(_11547_),
    .B(_11548_),
    .S(_08541_),
    .Z(_11549_)
  );
  AND2_X1 _19226_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_11549_),
    .ZN(_11550_)
  );
  INV_X1 _19227_ (
    .A(_11550_),
    .ZN(_11551_)
  );
  AND2_X1 _19228_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_11551_),
    .ZN(_11552_)
  );
  AND2_X1 _19229_ (
    .A1(_11546_),
    .A2(_11552_),
    .ZN(_11553_)
  );
  INV_X1 _19230_ (
    .A(_11553_),
    .ZN(_11554_)
  );
  AND2_X1 _19231_ (
    .A1(_08387_),
    .A2(_08542_),
    .ZN(_11555_)
  );
  INV_X1 _19232_ (
    .A(_11555_),
    .ZN(_11556_)
  );
  AND2_X1 _19233_ (
    .A1(_08288_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11557_)
  );
  INV_X1 _19234_ (
    .A(_11557_),
    .ZN(_11558_)
  );
  AND2_X1 _19235_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11558_),
    .ZN(_11559_)
  );
  AND2_X1 _19236_ (
    .A1(_11556_),
    .A2(_11559_),
    .ZN(_11560_)
  );
  INV_X1 _19237_ (
    .A(_11560_),
    .ZN(_11561_)
  );
  MUX2_X1 _19238_ (
    .A(\rf[22] [14]),
    .B(\rf[18] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11562_)
  );
  AND2_X1 _19239_ (
    .A1(_08541_),
    .A2(_11562_),
    .ZN(_11563_)
  );
  INV_X1 _19240_ (
    .A(_11563_),
    .ZN(_11564_)
  );
  AND2_X1 _19241_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_11564_),
    .ZN(_11565_)
  );
  AND2_X1 _19242_ (
    .A1(_11561_),
    .A2(_11565_),
    .ZN(_11566_)
  );
  INV_X1 _19243_ (
    .A(_11566_),
    .ZN(_11567_)
  );
  AND2_X1 _19244_ (
    .A1(_08318_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11568_)
  );
  INV_X1 _19245_ (
    .A(_11568_),
    .ZN(_11569_)
  );
  AND2_X1 _19246_ (
    .A1(_08417_),
    .A2(_08542_),
    .ZN(_11570_)
  );
  INV_X1 _19247_ (
    .A(_11570_),
    .ZN(_11571_)
  );
  AND2_X1 _19248_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11571_),
    .ZN(_11572_)
  );
  AND2_X1 _19249_ (
    .A1(_11569_),
    .A2(_11572_),
    .ZN(_11573_)
  );
  INV_X1 _19250_ (
    .A(_11573_),
    .ZN(_11574_)
  );
  MUX2_X1 _19251_ (
    .A(\rf[23] [14]),
    .B(\rf[19] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11575_)
  );
  AND2_X1 _19252_ (
    .A1(_08541_),
    .A2(_11575_),
    .ZN(_11576_)
  );
  INV_X1 _19253_ (
    .A(_11576_),
    .ZN(_11577_)
  );
  AND2_X1 _19254_ (
    .A1(_08540_),
    .A2(_11577_),
    .ZN(_11578_)
  );
  AND2_X1 _19255_ (
    .A1(_11574_),
    .A2(_11578_),
    .ZN(_11579_)
  );
  INV_X1 _19256_ (
    .A(_11579_),
    .ZN(_11580_)
  );
  AND2_X1 _19257_ (
    .A1(_11567_),
    .A2(_11580_),
    .ZN(_11581_)
  );
  INV_X1 _19258_ (
    .A(_11581_),
    .ZN(_11582_)
  );
  AND2_X1 _19259_ (
    .A1(_08571_),
    .A2(_11582_),
    .ZN(_11583_)
  );
  INV_X1 _19260_ (
    .A(_11583_),
    .ZN(_11584_)
  );
  AND2_X1 _19261_ (
    .A1(_11554_),
    .A2(_11584_),
    .ZN(_11585_)
  );
  AND2_X1 _19262_ (
    .A1(\rf[10] [14]),
    .A2(_08541_),
    .ZN(_11586_)
  );
  INV_X1 _19263_ (
    .A(_11586_),
    .ZN(_11587_)
  );
  AND2_X1 _19264_ (
    .A1(\rf[8] [14]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_11588_)
  );
  INV_X1 _19265_ (
    .A(_11588_),
    .ZN(_11589_)
  );
  AND2_X1 _19266_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_11589_),
    .ZN(_11590_)
  );
  AND2_X1 _19267_ (
    .A1(_11587_),
    .A2(_11590_),
    .ZN(_11591_)
  );
  INV_X1 _19268_ (
    .A(_11591_),
    .ZN(_11592_)
  );
  AND2_X1 _19269_ (
    .A1(\rf[14] [14]),
    .A2(_08541_),
    .ZN(_11593_)
  );
  INV_X1 _19270_ (
    .A(_11593_),
    .ZN(_11594_)
  );
  AND2_X1 _19271_ (
    .A1(\rf[12] [14]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_11595_)
  );
  INV_X1 _19272_ (
    .A(_11595_),
    .ZN(_11596_)
  );
  AND2_X1 _19273_ (
    .A1(_08542_),
    .A2(_11596_),
    .ZN(_11597_)
  );
  AND2_X1 _19274_ (
    .A1(_11594_),
    .A2(_11597_),
    .ZN(_11598_)
  );
  INV_X1 _19275_ (
    .A(_11598_),
    .ZN(_11599_)
  );
  AND2_X1 _19276_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_11599_),
    .ZN(_11600_)
  );
  AND2_X1 _19277_ (
    .A1(_11592_),
    .A2(_11600_),
    .ZN(_11601_)
  );
  INV_X1 _19278_ (
    .A(_11601_),
    .ZN(_11602_)
  );
  AND2_X1 _19279_ (
    .A1(\rf[11] [14]),
    .A2(_08541_),
    .ZN(_11603_)
  );
  INV_X1 _19280_ (
    .A(_11603_),
    .ZN(_11604_)
  );
  AND2_X1 _19281_ (
    .A1(\rf[9] [14]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_11605_)
  );
  INV_X1 _19282_ (
    .A(_11605_),
    .ZN(_11606_)
  );
  AND2_X1 _19283_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_11606_),
    .ZN(_11607_)
  );
  AND2_X1 _19284_ (
    .A1(_11604_),
    .A2(_11607_),
    .ZN(_11608_)
  );
  INV_X1 _19285_ (
    .A(_11608_),
    .ZN(_11609_)
  );
  AND2_X1 _19286_ (
    .A1(\rf[15] [14]),
    .A2(_08541_),
    .ZN(_11610_)
  );
  INV_X1 _19287_ (
    .A(_11610_),
    .ZN(_11611_)
  );
  AND2_X1 _19288_ (
    .A1(\rf[13] [14]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_11612_)
  );
  INV_X1 _19289_ (
    .A(_11612_),
    .ZN(_11613_)
  );
  AND2_X1 _19290_ (
    .A1(_08542_),
    .A2(_11613_),
    .ZN(_11614_)
  );
  AND2_X1 _19291_ (
    .A1(_11611_),
    .A2(_11614_),
    .ZN(_11615_)
  );
  INV_X1 _19292_ (
    .A(_11615_),
    .ZN(_11616_)
  );
  AND2_X1 _19293_ (
    .A1(_08540_),
    .A2(_11616_),
    .ZN(_11617_)
  );
  AND2_X1 _19294_ (
    .A1(_11609_),
    .A2(_11617_),
    .ZN(_11618_)
  );
  INV_X1 _19295_ (
    .A(_11618_),
    .ZN(_11619_)
  );
  AND2_X1 _19296_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_11619_),
    .ZN(_11620_)
  );
  AND2_X1 _19297_ (
    .A1(_11602_),
    .A2(_11620_),
    .ZN(_11621_)
  );
  INV_X1 _19298_ (
    .A(_11621_),
    .ZN(_11622_)
  );
  AND2_X1 _19299_ (
    .A1(\rf[30] [14]),
    .A2(_08542_),
    .ZN(_11623_)
  );
  INV_X1 _19300_ (
    .A(_11623_),
    .ZN(_11624_)
  );
  AND2_X1 _19301_ (
    .A1(\rf[26] [14]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11625_)
  );
  INV_X1 _19302_ (
    .A(_11625_),
    .ZN(_11626_)
  );
  AND2_X1 _19303_ (
    .A1(_08541_),
    .A2(_11626_),
    .ZN(_11627_)
  );
  AND2_X1 _19304_ (
    .A1(_11624_),
    .A2(_11627_),
    .ZN(_11628_)
  );
  INV_X1 _19305_ (
    .A(_11628_),
    .ZN(_11629_)
  );
  AND2_X1 _19306_ (
    .A1(\rf[24] [14]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11630_)
  );
  INV_X1 _19307_ (
    .A(_11630_),
    .ZN(_11631_)
  );
  AND2_X1 _19308_ (
    .A1(\rf[28] [14]),
    .A2(_08542_),
    .ZN(_11632_)
  );
  INV_X1 _19309_ (
    .A(_11632_),
    .ZN(_11633_)
  );
  AND2_X1 _19310_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11633_),
    .ZN(_11634_)
  );
  AND2_X1 _19311_ (
    .A1(_11631_),
    .A2(_11634_),
    .ZN(_11635_)
  );
  INV_X1 _19312_ (
    .A(_11635_),
    .ZN(_11636_)
  );
  AND2_X1 _19313_ (
    .A1(_11629_),
    .A2(_11636_),
    .ZN(_11637_)
  );
  MUX2_X1 _19314_ (
    .A(\rf[29] [14]),
    .B(\rf[25] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11638_)
  );
  AND2_X1 _19315_ (
    .A1(\rf[27] [14]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11639_)
  );
  MUX2_X1 _19316_ (
    .A(_11638_),
    .B(_11639_),
    .S(_08541_),
    .Z(_11640_)
  );
  MUX2_X1 _19317_ (
    .A(_11637_),
    .B(_11640_),
    .S(_08540_),
    .Z(_11641_)
  );
  INV_X1 _19318_ (
    .A(_11641_),
    .ZN(_11642_)
  );
  AND2_X1 _19319_ (
    .A1(_08571_),
    .A2(_11642_),
    .ZN(_11643_)
  );
  INV_X1 _19320_ (
    .A(_11643_),
    .ZN(_11644_)
  );
  AND2_X1 _19321_ (
    .A1(_11622_),
    .A2(_11644_),
    .ZN(_11645_)
  );
  MUX2_X1 _19322_ (
    .A(_11585_),
    .B(_11645_),
    .S(_08543_),
    .Z(_11646_)
  );
  MUX2_X1 _19323_ (
    .A(_11646_),
    .B(_11541_),
    .S(_10131_),
    .Z(_11647_)
  );
  AND2_X1 _19324_ (
    .A1(_10082_),
    .A2(_11647_),
    .ZN(_11648_)
  );
  INV_X1 _19325_ (
    .A(_11648_),
    .ZN(_11649_)
  );
  AND2_X1 _19326_ (
    .A1(_11538_),
    .A2(_11649_),
    .ZN(_11650_)
  );
  INV_X1 _19327_ (
    .A(_11650_),
    .ZN(_11651_)
  );
  MUX2_X1 _19328_ (
    .A(ex_reg_rs_msb_0[12]),
    .B(_11651_),
    .S(_10079_),
    .Z(_00079_)
  );
  AND2_X1 _19329_ (
    .A1(ibuf_io_inst_0_bits_raw[15]),
    .A2(_09295_),
    .ZN(_11652_)
  );
  INV_X1 _19330_ (
    .A(_11652_),
    .ZN(_11653_)
  );
  MUX2_X1 _19331_ (
    .A(csr_io_rw_rdata[15]),
    .B(wb_reg_wdata[15]),
    .S(_10134_),
    .Z(_11654_)
  );
  MUX2_X1 _19332_ (
    .A(div_io_resp_bits_data[15]),
    .B(_11654_),
    .S(_08649_),
    .Z(_11655_)
  );
  MUX2_X1 _19333_ (
    .A(_11655_),
    .B(io_dmem_resp_bits_data[15]),
    .S(_08631_),
    .Z(_11656_)
  );
  MUX2_X1 _19334_ (
    .A(\rf[23] [15]),
    .B(\rf[22] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_11657_)
  );
  INV_X1 _19335_ (
    .A(_11657_),
    .ZN(_11658_)
  );
  AND2_X1 _19336_ (
    .A1(_08542_),
    .A2(_11658_),
    .ZN(_11659_)
  );
  INV_X1 _19337_ (
    .A(_11659_),
    .ZN(_11660_)
  );
  MUX2_X1 _19338_ (
    .A(\rf[19] [15]),
    .B(\rf[18] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_11661_)
  );
  INV_X1 _19339_ (
    .A(_11661_),
    .ZN(_11662_)
  );
  AND2_X1 _19340_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_11662_),
    .ZN(_11663_)
  );
  INV_X1 _19341_ (
    .A(_11663_),
    .ZN(_11664_)
  );
  AND2_X1 _19342_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_11664_),
    .ZN(_11665_)
  );
  AND2_X1 _19343_ (
    .A1(_11660_),
    .A2(_11665_),
    .ZN(_11666_)
  );
  INV_X1 _19344_ (
    .A(_11666_),
    .ZN(_11667_)
  );
  AND2_X1 _19345_ (
    .A1(_08499_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11668_)
  );
  INV_X1 _19346_ (
    .A(_11668_),
    .ZN(_11669_)
  );
  AND2_X1 _19347_ (
    .A1(_08472_),
    .A2(_08542_),
    .ZN(_11670_)
  );
  INV_X1 _19348_ (
    .A(_11670_),
    .ZN(_11671_)
  );
  AND2_X1 _19349_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_11671_),
    .ZN(_11672_)
  );
  AND2_X1 _19350_ (
    .A1(_11669_),
    .A2(_11672_),
    .ZN(_11673_)
  );
  INV_X1 _19351_ (
    .A(_11673_),
    .ZN(_11674_)
  );
  AND2_X1 _19352_ (
    .A1(\rf[27] [15]),
    .A2(_09608_),
    .ZN(_11675_)
  );
  INV_X1 _19353_ (
    .A(_11675_),
    .ZN(_11676_)
  );
  AND2_X1 _19354_ (
    .A1(_11674_),
    .A2(_11676_),
    .ZN(_11677_)
  );
  INV_X1 _19355_ (
    .A(_11677_),
    .ZN(_11678_)
  );
  AND2_X1 _19356_ (
    .A1(_08543_),
    .A2(_11678_),
    .ZN(_11679_)
  );
  INV_X1 _19357_ (
    .A(_11679_),
    .ZN(_11680_)
  );
  AND2_X1 _19358_ (
    .A1(_08541_),
    .A2(_11680_),
    .ZN(_11681_)
  );
  AND2_X1 _19359_ (
    .A1(_11667_),
    .A2(_11681_),
    .ZN(_11682_)
  );
  INV_X1 _19360_ (
    .A(_11682_),
    .ZN(_11683_)
  );
  AND2_X1 _19361_ (
    .A1(\rf[20] [15]),
    .A2(_08542_),
    .ZN(_11684_)
  );
  INV_X1 _19362_ (
    .A(_11684_),
    .ZN(_11685_)
  );
  AND2_X1 _19363_ (
    .A1(\rf[16] [15]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11686_)
  );
  INV_X1 _19364_ (
    .A(_11686_),
    .ZN(_11687_)
  );
  AND2_X1 _19365_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_11687_),
    .ZN(_11688_)
  );
  AND2_X1 _19366_ (
    .A1(_11685_),
    .A2(_11688_),
    .ZN(_11689_)
  );
  INV_X1 _19367_ (
    .A(_11689_),
    .ZN(_11690_)
  );
  AND2_X1 _19368_ (
    .A1(\rf[21] [15]),
    .A2(_08542_),
    .ZN(_11691_)
  );
  INV_X1 _19369_ (
    .A(_11691_),
    .ZN(_11692_)
  );
  AND2_X1 _19370_ (
    .A1(\rf[17] [15]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11693_)
  );
  INV_X1 _19371_ (
    .A(_11693_),
    .ZN(_11694_)
  );
  AND2_X1 _19372_ (
    .A1(_08540_),
    .A2(_11694_),
    .ZN(_11695_)
  );
  AND2_X1 _19373_ (
    .A1(_11692_),
    .A2(_11695_),
    .ZN(_11696_)
  );
  INV_X1 _19374_ (
    .A(_11696_),
    .ZN(_11697_)
  );
  AND2_X1 _19375_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_11697_),
    .ZN(_11698_)
  );
  AND2_X1 _19376_ (
    .A1(_11690_),
    .A2(_11698_),
    .ZN(_11699_)
  );
  INV_X1 _19377_ (
    .A(_11699_),
    .ZN(_11700_)
  );
  AND2_X1 _19378_ (
    .A1(\rf[28] [15]),
    .A2(_08542_),
    .ZN(_11701_)
  );
  INV_X1 _19379_ (
    .A(_11701_),
    .ZN(_11702_)
  );
  AND2_X1 _19380_ (
    .A1(\rf[24] [15]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11703_)
  );
  INV_X1 _19381_ (
    .A(_11703_),
    .ZN(_11704_)
  );
  AND2_X1 _19382_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_11704_),
    .ZN(_11705_)
  );
  AND2_X1 _19383_ (
    .A1(_11702_),
    .A2(_11705_),
    .ZN(_11706_)
  );
  INV_X1 _19384_ (
    .A(_11706_),
    .ZN(_11707_)
  );
  AND2_X1 _19385_ (
    .A1(\rf[29] [15]),
    .A2(_08542_),
    .ZN(_11708_)
  );
  INV_X1 _19386_ (
    .A(_11708_),
    .ZN(_11709_)
  );
  AND2_X1 _19387_ (
    .A1(\rf[25] [15]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11710_)
  );
  INV_X1 _19388_ (
    .A(_11710_),
    .ZN(_11711_)
  );
  AND2_X1 _19389_ (
    .A1(_08540_),
    .A2(_11711_),
    .ZN(_11712_)
  );
  AND2_X1 _19390_ (
    .A1(_11709_),
    .A2(_11712_),
    .ZN(_11713_)
  );
  INV_X1 _19391_ (
    .A(_11713_),
    .ZN(_11714_)
  );
  AND2_X1 _19392_ (
    .A1(_08543_),
    .A2(_11714_),
    .ZN(_11715_)
  );
  AND2_X1 _19393_ (
    .A1(_11707_),
    .A2(_11715_),
    .ZN(_11716_)
  );
  INV_X1 _19394_ (
    .A(_11716_),
    .ZN(_11717_)
  );
  AND2_X1 _19395_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11717_),
    .ZN(_11718_)
  );
  AND2_X1 _19396_ (
    .A1(_11700_),
    .A2(_11718_),
    .ZN(_11719_)
  );
  INV_X1 _19397_ (
    .A(_11719_),
    .ZN(_11720_)
  );
  AND2_X1 _19398_ (
    .A1(_11683_),
    .A2(_11720_),
    .ZN(_11721_)
  );
  MUX2_X1 _19399_ (
    .A(\rf[1] [15]),
    .B(\rf[0] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_11722_)
  );
  MUX2_X1 _19400_ (
    .A(\rf[5] [15]),
    .B(\rf[4] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_11723_)
  );
  MUX2_X1 _19401_ (
    .A(_11722_),
    .B(_11723_),
    .S(_08542_),
    .Z(_11724_)
  );
  INV_X1 _19402_ (
    .A(_11724_),
    .ZN(_11725_)
  );
  AND2_X1 _19403_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_11725_),
    .ZN(_11726_)
  );
  INV_X1 _19404_ (
    .A(_11726_),
    .ZN(_11727_)
  );
  MUX2_X1 _19405_ (
    .A(\rf[12] [15]),
    .B(\rf[8] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11728_)
  );
  INV_X1 _19406_ (
    .A(_11728_),
    .ZN(_11729_)
  );
  AND2_X1 _19407_ (
    .A1(_10213_),
    .A2(_11729_),
    .ZN(_11730_)
  );
  INV_X1 _19408_ (
    .A(_11730_),
    .ZN(_11731_)
  );
  MUX2_X1 _19409_ (
    .A(\rf[13] [15]),
    .B(\rf[9] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11732_)
  );
  INV_X1 _19410_ (
    .A(_11732_),
    .ZN(_11733_)
  );
  AND2_X1 _19411_ (
    .A1(_09110_),
    .A2(_11733_),
    .ZN(_11734_)
  );
  INV_X1 _19412_ (
    .A(_11734_),
    .ZN(_11735_)
  );
  AND2_X1 _19413_ (
    .A1(_11731_),
    .A2(_11735_),
    .ZN(_11736_)
  );
  AND2_X1 _19414_ (
    .A1(_11727_),
    .A2(_11736_),
    .ZN(_11737_)
  );
  MUX2_X1 _19415_ (
    .A(\rf[3] [15]),
    .B(\rf[2] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_11738_)
  );
  MUX2_X1 _19416_ (
    .A(\rf[7] [15]),
    .B(\rf[6] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_11739_)
  );
  MUX2_X1 _19417_ (
    .A(_11738_),
    .B(_11739_),
    .S(_08542_),
    .Z(_11740_)
  );
  INV_X1 _19418_ (
    .A(_11740_),
    .ZN(_11741_)
  );
  AND2_X1 _19419_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_11741_),
    .ZN(_11742_)
  );
  INV_X1 _19420_ (
    .A(_11742_),
    .ZN(_11743_)
  );
  MUX2_X1 _19421_ (
    .A(\rf[14] [15]),
    .B(\rf[10] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11744_)
  );
  INV_X1 _19422_ (
    .A(_11744_),
    .ZN(_11745_)
  );
  AND2_X1 _19423_ (
    .A1(_10213_),
    .A2(_11745_),
    .ZN(_11746_)
  );
  INV_X1 _19424_ (
    .A(_11746_),
    .ZN(_11747_)
  );
  MUX2_X1 _19425_ (
    .A(\rf[15] [15]),
    .B(\rf[11] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11748_)
  );
  INV_X1 _19426_ (
    .A(_11748_),
    .ZN(_11749_)
  );
  AND2_X1 _19427_ (
    .A1(_09110_),
    .A2(_11749_),
    .ZN(_11750_)
  );
  INV_X1 _19428_ (
    .A(_11750_),
    .ZN(_11751_)
  );
  AND2_X1 _19429_ (
    .A1(_11747_),
    .A2(_11751_),
    .ZN(_11752_)
  );
  AND2_X1 _19430_ (
    .A1(_11743_),
    .A2(_11752_),
    .ZN(_11753_)
  );
  MUX2_X1 _19431_ (
    .A(_11737_),
    .B(_11753_),
    .S(_08541_),
    .Z(_11754_)
  );
  MUX2_X1 _19432_ (
    .A(_11721_),
    .B(_11754_),
    .S(ibuf_io_inst_0_bits_inst_rs1[4]),
    .Z(_11755_)
  );
  MUX2_X1 _19433_ (
    .A(_11656_),
    .B(_11755_),
    .S(_10132_),
    .Z(_11756_)
  );
  AND2_X1 _19434_ (
    .A1(_10082_),
    .A2(_11756_),
    .ZN(_11757_)
  );
  INV_X1 _19435_ (
    .A(_11757_),
    .ZN(_11758_)
  );
  AND2_X1 _19436_ (
    .A1(_11653_),
    .A2(_11758_),
    .ZN(_11759_)
  );
  INV_X1 _19437_ (
    .A(_11759_),
    .ZN(_11760_)
  );
  MUX2_X1 _19438_ (
    .A(ex_reg_rs_msb_0[13]),
    .B(_11760_),
    .S(_10079_),
    .Z(_00080_)
  );
  AND2_X1 _19439_ (
    .A1(_08578_),
    .A2(ibuf_io_inst_0_bits_raw[16]),
    .ZN(_11761_)
  );
  AND2_X1 _19440_ (
    .A1(_09295_),
    .A2(_11761_),
    .ZN(_11762_)
  );
  INV_X1 _19441_ (
    .A(_11762_),
    .ZN(_11763_)
  );
  MUX2_X1 _19442_ (
    .A(csr_io_rw_rdata[16]),
    .B(wb_reg_wdata[16]),
    .S(_10134_),
    .Z(_11764_)
  );
  MUX2_X1 _19443_ (
    .A(div_io_resp_bits_data[16]),
    .B(_11764_),
    .S(_08649_),
    .Z(_11765_)
  );
  MUX2_X1 _19444_ (
    .A(_11765_),
    .B(io_dmem_resp_bits_data[16]),
    .S(_08631_),
    .Z(_11766_)
  );
  MUX2_X1 _19445_ (
    .A(\rf[5] [16]),
    .B(\rf[1] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11767_)
  );
  MUX2_X1 _19446_ (
    .A(\rf[7] [16]),
    .B(\rf[3] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11768_)
  );
  MUX2_X1 _19447_ (
    .A(_11767_),
    .B(_11768_),
    .S(_08541_),
    .Z(_11769_)
  );
  AND2_X1 _19448_ (
    .A1(_08540_),
    .A2(_11769_),
    .ZN(_11770_)
  );
  INV_X1 _19449_ (
    .A(_11770_),
    .ZN(_11771_)
  );
  MUX2_X1 _19450_ (
    .A(\rf[4] [16]),
    .B(\rf[0] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11772_)
  );
  MUX2_X1 _19451_ (
    .A(\rf[6] [16]),
    .B(\rf[2] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11773_)
  );
  MUX2_X1 _19452_ (
    .A(_11772_),
    .B(_11773_),
    .S(_08541_),
    .Z(_11774_)
  );
  AND2_X1 _19453_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_11774_),
    .ZN(_11775_)
  );
  INV_X1 _19454_ (
    .A(_11775_),
    .ZN(_11776_)
  );
  AND2_X1 _19455_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_11776_),
    .ZN(_11777_)
  );
  AND2_X1 _19456_ (
    .A1(_11771_),
    .A2(_11777_),
    .ZN(_11778_)
  );
  INV_X1 _19457_ (
    .A(_11778_),
    .ZN(_11779_)
  );
  AND2_X1 _19458_ (
    .A1(_08389_),
    .A2(_08542_),
    .ZN(_11780_)
  );
  INV_X1 _19459_ (
    .A(_11780_),
    .ZN(_11781_)
  );
  AND2_X1 _19460_ (
    .A1(_08290_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11782_)
  );
  INV_X1 _19461_ (
    .A(_11782_),
    .ZN(_11783_)
  );
  AND2_X1 _19462_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11783_),
    .ZN(_11784_)
  );
  AND2_X1 _19463_ (
    .A1(_11781_),
    .A2(_11784_),
    .ZN(_11785_)
  );
  INV_X1 _19464_ (
    .A(_11785_),
    .ZN(_11786_)
  );
  MUX2_X1 _19465_ (
    .A(\rf[22] [16]),
    .B(\rf[18] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11787_)
  );
  AND2_X1 _19466_ (
    .A1(_08541_),
    .A2(_11787_),
    .ZN(_11788_)
  );
  INV_X1 _19467_ (
    .A(_11788_),
    .ZN(_11789_)
  );
  AND2_X1 _19468_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_11789_),
    .ZN(_11790_)
  );
  AND2_X1 _19469_ (
    .A1(_11786_),
    .A2(_11790_),
    .ZN(_11791_)
  );
  INV_X1 _19470_ (
    .A(_11791_),
    .ZN(_11792_)
  );
  AND2_X1 _19471_ (
    .A1(_08320_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11793_)
  );
  INV_X1 _19472_ (
    .A(_11793_),
    .ZN(_11794_)
  );
  AND2_X1 _19473_ (
    .A1(_08419_),
    .A2(_08542_),
    .ZN(_11795_)
  );
  INV_X1 _19474_ (
    .A(_11795_),
    .ZN(_11796_)
  );
  AND2_X1 _19475_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11796_),
    .ZN(_11797_)
  );
  AND2_X1 _19476_ (
    .A1(_11794_),
    .A2(_11797_),
    .ZN(_11798_)
  );
  INV_X1 _19477_ (
    .A(_11798_),
    .ZN(_11799_)
  );
  MUX2_X1 _19478_ (
    .A(\rf[23] [16]),
    .B(\rf[19] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11800_)
  );
  AND2_X1 _19479_ (
    .A1(_08541_),
    .A2(_11800_),
    .ZN(_11801_)
  );
  INV_X1 _19480_ (
    .A(_11801_),
    .ZN(_11802_)
  );
  AND2_X1 _19481_ (
    .A1(_08540_),
    .A2(_11802_),
    .ZN(_11803_)
  );
  AND2_X1 _19482_ (
    .A1(_11799_),
    .A2(_11803_),
    .ZN(_11804_)
  );
  INV_X1 _19483_ (
    .A(_11804_),
    .ZN(_11805_)
  );
  AND2_X1 _19484_ (
    .A1(_11792_),
    .A2(_11805_),
    .ZN(_11806_)
  );
  INV_X1 _19485_ (
    .A(_11806_),
    .ZN(_11807_)
  );
  AND2_X1 _19486_ (
    .A1(_08571_),
    .A2(_11807_),
    .ZN(_11808_)
  );
  INV_X1 _19487_ (
    .A(_11808_),
    .ZN(_11809_)
  );
  AND2_X1 _19488_ (
    .A1(_11779_),
    .A2(_11809_),
    .ZN(_11810_)
  );
  AND2_X1 _19489_ (
    .A1(\rf[10] [16]),
    .A2(_08541_),
    .ZN(_11811_)
  );
  INV_X1 _19490_ (
    .A(_11811_),
    .ZN(_11812_)
  );
  AND2_X1 _19491_ (
    .A1(\rf[8] [16]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_11813_)
  );
  INV_X1 _19492_ (
    .A(_11813_),
    .ZN(_11814_)
  );
  AND2_X1 _19493_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_11814_),
    .ZN(_11815_)
  );
  AND2_X1 _19494_ (
    .A1(_11812_),
    .A2(_11815_),
    .ZN(_11816_)
  );
  INV_X1 _19495_ (
    .A(_11816_),
    .ZN(_11817_)
  );
  AND2_X1 _19496_ (
    .A1(\rf[14] [16]),
    .A2(_08541_),
    .ZN(_11818_)
  );
  INV_X1 _19497_ (
    .A(_11818_),
    .ZN(_11819_)
  );
  AND2_X1 _19498_ (
    .A1(\rf[12] [16]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_11820_)
  );
  INV_X1 _19499_ (
    .A(_11820_),
    .ZN(_11821_)
  );
  AND2_X1 _19500_ (
    .A1(_08542_),
    .A2(_11821_),
    .ZN(_11822_)
  );
  AND2_X1 _19501_ (
    .A1(_11819_),
    .A2(_11822_),
    .ZN(_11823_)
  );
  INV_X1 _19502_ (
    .A(_11823_),
    .ZN(_11824_)
  );
  AND2_X1 _19503_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_11824_),
    .ZN(_11825_)
  );
  AND2_X1 _19504_ (
    .A1(_11817_),
    .A2(_11825_),
    .ZN(_11826_)
  );
  INV_X1 _19505_ (
    .A(_11826_),
    .ZN(_11827_)
  );
  AND2_X1 _19506_ (
    .A1(\rf[11] [16]),
    .A2(_08541_),
    .ZN(_11828_)
  );
  INV_X1 _19507_ (
    .A(_11828_),
    .ZN(_11829_)
  );
  AND2_X1 _19508_ (
    .A1(\rf[9] [16]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_11830_)
  );
  INV_X1 _19509_ (
    .A(_11830_),
    .ZN(_11831_)
  );
  AND2_X1 _19510_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_11831_),
    .ZN(_11832_)
  );
  AND2_X1 _19511_ (
    .A1(_11829_),
    .A2(_11832_),
    .ZN(_11833_)
  );
  INV_X1 _19512_ (
    .A(_11833_),
    .ZN(_11834_)
  );
  AND2_X1 _19513_ (
    .A1(\rf[15] [16]),
    .A2(_08541_),
    .ZN(_11835_)
  );
  INV_X1 _19514_ (
    .A(_11835_),
    .ZN(_11836_)
  );
  AND2_X1 _19515_ (
    .A1(\rf[13] [16]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_11837_)
  );
  INV_X1 _19516_ (
    .A(_11837_),
    .ZN(_11838_)
  );
  AND2_X1 _19517_ (
    .A1(_08542_),
    .A2(_11838_),
    .ZN(_11839_)
  );
  AND2_X1 _19518_ (
    .A1(_11836_),
    .A2(_11839_),
    .ZN(_11840_)
  );
  INV_X1 _19519_ (
    .A(_11840_),
    .ZN(_11841_)
  );
  AND2_X1 _19520_ (
    .A1(_08540_),
    .A2(_11841_),
    .ZN(_11842_)
  );
  AND2_X1 _19521_ (
    .A1(_11834_),
    .A2(_11842_),
    .ZN(_11843_)
  );
  INV_X1 _19522_ (
    .A(_11843_),
    .ZN(_11844_)
  );
  AND2_X1 _19523_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_11844_),
    .ZN(_11845_)
  );
  AND2_X1 _19524_ (
    .A1(_11827_),
    .A2(_11845_),
    .ZN(_11846_)
  );
  INV_X1 _19525_ (
    .A(_11846_),
    .ZN(_11847_)
  );
  AND2_X1 _19526_ (
    .A1(\rf[30] [16]),
    .A2(_08542_),
    .ZN(_11848_)
  );
  INV_X1 _19527_ (
    .A(_11848_),
    .ZN(_11849_)
  );
  AND2_X1 _19528_ (
    .A1(\rf[26] [16]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11850_)
  );
  INV_X1 _19529_ (
    .A(_11850_),
    .ZN(_11851_)
  );
  AND2_X1 _19530_ (
    .A1(_08541_),
    .A2(_11851_),
    .ZN(_11852_)
  );
  AND2_X1 _19531_ (
    .A1(_11849_),
    .A2(_11852_),
    .ZN(_11853_)
  );
  INV_X1 _19532_ (
    .A(_11853_),
    .ZN(_11854_)
  );
  AND2_X1 _19533_ (
    .A1(\rf[24] [16]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11855_)
  );
  INV_X1 _19534_ (
    .A(_11855_),
    .ZN(_11856_)
  );
  AND2_X1 _19535_ (
    .A1(\rf[28] [16]),
    .A2(_08542_),
    .ZN(_11857_)
  );
  INV_X1 _19536_ (
    .A(_11857_),
    .ZN(_11858_)
  );
  AND2_X1 _19537_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11858_),
    .ZN(_11859_)
  );
  AND2_X1 _19538_ (
    .A1(_11856_),
    .A2(_11859_),
    .ZN(_11860_)
  );
  INV_X1 _19539_ (
    .A(_11860_),
    .ZN(_11861_)
  );
  AND2_X1 _19540_ (
    .A1(_11854_),
    .A2(_11861_),
    .ZN(_11862_)
  );
  MUX2_X1 _19541_ (
    .A(\rf[29] [16]),
    .B(\rf[25] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11863_)
  );
  AND2_X1 _19542_ (
    .A1(\rf[27] [16]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11864_)
  );
  MUX2_X1 _19543_ (
    .A(_11863_),
    .B(_11864_),
    .S(_08541_),
    .Z(_11865_)
  );
  MUX2_X1 _19544_ (
    .A(_11862_),
    .B(_11865_),
    .S(_08540_),
    .Z(_11866_)
  );
  INV_X1 _19545_ (
    .A(_11866_),
    .ZN(_11867_)
  );
  AND2_X1 _19546_ (
    .A1(_08571_),
    .A2(_11867_),
    .ZN(_11868_)
  );
  INV_X1 _19547_ (
    .A(_11868_),
    .ZN(_11869_)
  );
  AND2_X1 _19548_ (
    .A1(_11847_),
    .A2(_11869_),
    .ZN(_11870_)
  );
  MUX2_X1 _19549_ (
    .A(_11810_),
    .B(_11870_),
    .S(_08543_),
    .Z(_11871_)
  );
  MUX2_X1 _19550_ (
    .A(_11871_),
    .B(_11766_),
    .S(_10131_),
    .Z(_11872_)
  );
  AND2_X1 _19551_ (
    .A1(_10082_),
    .A2(_11872_),
    .ZN(_11873_)
  );
  INV_X1 _19552_ (
    .A(_11873_),
    .ZN(_11874_)
  );
  AND2_X1 _19553_ (
    .A1(_11763_),
    .A2(_11874_),
    .ZN(_11875_)
  );
  INV_X1 _19554_ (
    .A(_11875_),
    .ZN(_11876_)
  );
  MUX2_X1 _19555_ (
    .A(ex_reg_rs_msb_0[14]),
    .B(_11876_),
    .S(_10079_),
    .Z(_00081_)
  );
  AND2_X1 _19556_ (
    .A1(_08578_),
    .A2(ibuf_io_inst_0_bits_raw[17]),
    .ZN(_11877_)
  );
  AND2_X1 _19557_ (
    .A1(_09295_),
    .A2(_11877_),
    .ZN(_11878_)
  );
  INV_X1 _19558_ (
    .A(_11878_),
    .ZN(_11879_)
  );
  MUX2_X1 _19559_ (
    .A(csr_io_rw_rdata[17]),
    .B(wb_reg_wdata[17]),
    .S(_10134_),
    .Z(_11880_)
  );
  MUX2_X1 _19560_ (
    .A(div_io_resp_bits_data[17]),
    .B(_11880_),
    .S(_08649_),
    .Z(_11881_)
  );
  MUX2_X1 _19561_ (
    .A(_11881_),
    .B(io_dmem_resp_bits_data[17]),
    .S(_08631_),
    .Z(_11882_)
  );
  MUX2_X1 _19562_ (
    .A(\rf[5] [17]),
    .B(\rf[1] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11883_)
  );
  MUX2_X1 _19563_ (
    .A(\rf[7] [17]),
    .B(\rf[3] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11884_)
  );
  MUX2_X1 _19564_ (
    .A(_11883_),
    .B(_11884_),
    .S(_08541_),
    .Z(_11885_)
  );
  AND2_X1 _19565_ (
    .A1(_08540_),
    .A2(_11885_),
    .ZN(_11886_)
  );
  INV_X1 _19566_ (
    .A(_11886_),
    .ZN(_11887_)
  );
  MUX2_X1 _19567_ (
    .A(\rf[4] [17]),
    .B(\rf[0] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11888_)
  );
  MUX2_X1 _19568_ (
    .A(\rf[6] [17]),
    .B(\rf[2] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11889_)
  );
  MUX2_X1 _19569_ (
    .A(_11888_),
    .B(_11889_),
    .S(_08541_),
    .Z(_11890_)
  );
  AND2_X1 _19570_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_11890_),
    .ZN(_11891_)
  );
  INV_X1 _19571_ (
    .A(_11891_),
    .ZN(_11892_)
  );
  AND2_X1 _19572_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_11892_),
    .ZN(_11893_)
  );
  AND2_X1 _19573_ (
    .A1(_11887_),
    .A2(_11893_),
    .ZN(_11894_)
  );
  INV_X1 _19574_ (
    .A(_11894_),
    .ZN(_11895_)
  );
  AND2_X1 _19575_ (
    .A1(_08390_),
    .A2(_08542_),
    .ZN(_11896_)
  );
  INV_X1 _19576_ (
    .A(_11896_),
    .ZN(_11897_)
  );
  AND2_X1 _19577_ (
    .A1(_08291_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11898_)
  );
  INV_X1 _19578_ (
    .A(_11898_),
    .ZN(_11899_)
  );
  AND2_X1 _19579_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11899_),
    .ZN(_11900_)
  );
  AND2_X1 _19580_ (
    .A1(_11897_),
    .A2(_11900_),
    .ZN(_11901_)
  );
  INV_X1 _19581_ (
    .A(_11901_),
    .ZN(_11902_)
  );
  MUX2_X1 _19582_ (
    .A(\rf[22] [17]),
    .B(\rf[18] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11903_)
  );
  AND2_X1 _19583_ (
    .A1(_08541_),
    .A2(_11903_),
    .ZN(_11904_)
  );
  INV_X1 _19584_ (
    .A(_11904_),
    .ZN(_11905_)
  );
  AND2_X1 _19585_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_11905_),
    .ZN(_11906_)
  );
  AND2_X1 _19586_ (
    .A1(_11902_),
    .A2(_11906_),
    .ZN(_11907_)
  );
  INV_X1 _19587_ (
    .A(_11907_),
    .ZN(_11908_)
  );
  AND2_X1 _19588_ (
    .A1(_08321_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11909_)
  );
  INV_X1 _19589_ (
    .A(_11909_),
    .ZN(_11910_)
  );
  AND2_X1 _19590_ (
    .A1(_08420_),
    .A2(_08542_),
    .ZN(_11911_)
  );
  INV_X1 _19591_ (
    .A(_11911_),
    .ZN(_11912_)
  );
  AND2_X1 _19592_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11912_),
    .ZN(_11913_)
  );
  AND2_X1 _19593_ (
    .A1(_11910_),
    .A2(_11913_),
    .ZN(_11914_)
  );
  INV_X1 _19594_ (
    .A(_11914_),
    .ZN(_11915_)
  );
  MUX2_X1 _19595_ (
    .A(\rf[23] [17]),
    .B(\rf[19] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11916_)
  );
  AND2_X1 _19596_ (
    .A1(_08541_),
    .A2(_11916_),
    .ZN(_11917_)
  );
  INV_X1 _19597_ (
    .A(_11917_),
    .ZN(_11918_)
  );
  AND2_X1 _19598_ (
    .A1(_08540_),
    .A2(_11918_),
    .ZN(_11919_)
  );
  AND2_X1 _19599_ (
    .A1(_11915_),
    .A2(_11919_),
    .ZN(_11920_)
  );
  INV_X1 _19600_ (
    .A(_11920_),
    .ZN(_11921_)
  );
  AND2_X1 _19601_ (
    .A1(_11908_),
    .A2(_11921_),
    .ZN(_11922_)
  );
  INV_X1 _19602_ (
    .A(_11922_),
    .ZN(_11923_)
  );
  AND2_X1 _19603_ (
    .A1(_08571_),
    .A2(_11923_),
    .ZN(_11924_)
  );
  INV_X1 _19604_ (
    .A(_11924_),
    .ZN(_11925_)
  );
  AND2_X1 _19605_ (
    .A1(_11895_),
    .A2(_11925_),
    .ZN(_11926_)
  );
  AND2_X1 _19606_ (
    .A1(\rf[10] [17]),
    .A2(_08541_),
    .ZN(_11927_)
  );
  INV_X1 _19607_ (
    .A(_11927_),
    .ZN(_11928_)
  );
  AND2_X1 _19608_ (
    .A1(\rf[8] [17]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_11929_)
  );
  INV_X1 _19609_ (
    .A(_11929_),
    .ZN(_11930_)
  );
  AND2_X1 _19610_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_11930_),
    .ZN(_11931_)
  );
  AND2_X1 _19611_ (
    .A1(_11928_),
    .A2(_11931_),
    .ZN(_11932_)
  );
  INV_X1 _19612_ (
    .A(_11932_),
    .ZN(_11933_)
  );
  AND2_X1 _19613_ (
    .A1(\rf[14] [17]),
    .A2(_08541_),
    .ZN(_11934_)
  );
  INV_X1 _19614_ (
    .A(_11934_),
    .ZN(_11935_)
  );
  AND2_X1 _19615_ (
    .A1(\rf[12] [17]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_11936_)
  );
  INV_X1 _19616_ (
    .A(_11936_),
    .ZN(_11937_)
  );
  AND2_X1 _19617_ (
    .A1(_08542_),
    .A2(_11937_),
    .ZN(_11938_)
  );
  AND2_X1 _19618_ (
    .A1(_11935_),
    .A2(_11938_),
    .ZN(_11939_)
  );
  INV_X1 _19619_ (
    .A(_11939_),
    .ZN(_11940_)
  );
  AND2_X1 _19620_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_11940_),
    .ZN(_11941_)
  );
  AND2_X1 _19621_ (
    .A1(_11933_),
    .A2(_11941_),
    .ZN(_11942_)
  );
  INV_X1 _19622_ (
    .A(_11942_),
    .ZN(_11943_)
  );
  AND2_X1 _19623_ (
    .A1(\rf[11] [17]),
    .A2(_08541_),
    .ZN(_11944_)
  );
  INV_X1 _19624_ (
    .A(_11944_),
    .ZN(_11945_)
  );
  AND2_X1 _19625_ (
    .A1(\rf[9] [17]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_11946_)
  );
  INV_X1 _19626_ (
    .A(_11946_),
    .ZN(_11947_)
  );
  AND2_X1 _19627_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_11947_),
    .ZN(_11948_)
  );
  AND2_X1 _19628_ (
    .A1(_11945_),
    .A2(_11948_),
    .ZN(_11949_)
  );
  INV_X1 _19629_ (
    .A(_11949_),
    .ZN(_11950_)
  );
  AND2_X1 _19630_ (
    .A1(\rf[15] [17]),
    .A2(_08541_),
    .ZN(_11951_)
  );
  INV_X1 _19631_ (
    .A(_11951_),
    .ZN(_11952_)
  );
  AND2_X1 _19632_ (
    .A1(\rf[13] [17]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_11953_)
  );
  INV_X1 _19633_ (
    .A(_11953_),
    .ZN(_11954_)
  );
  AND2_X1 _19634_ (
    .A1(_08542_),
    .A2(_11954_),
    .ZN(_11955_)
  );
  AND2_X1 _19635_ (
    .A1(_11952_),
    .A2(_11955_),
    .ZN(_11956_)
  );
  INV_X1 _19636_ (
    .A(_11956_),
    .ZN(_11957_)
  );
  AND2_X1 _19637_ (
    .A1(_08540_),
    .A2(_11957_),
    .ZN(_11958_)
  );
  AND2_X1 _19638_ (
    .A1(_11950_),
    .A2(_11958_),
    .ZN(_11959_)
  );
  INV_X1 _19639_ (
    .A(_11959_),
    .ZN(_11960_)
  );
  AND2_X1 _19640_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_11960_),
    .ZN(_11961_)
  );
  AND2_X1 _19641_ (
    .A1(_11943_),
    .A2(_11961_),
    .ZN(_11962_)
  );
  INV_X1 _19642_ (
    .A(_11962_),
    .ZN(_11963_)
  );
  AND2_X1 _19643_ (
    .A1(\rf[30] [17]),
    .A2(_08542_),
    .ZN(_11964_)
  );
  INV_X1 _19644_ (
    .A(_11964_),
    .ZN(_11965_)
  );
  AND2_X1 _19645_ (
    .A1(\rf[26] [17]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11966_)
  );
  INV_X1 _19646_ (
    .A(_11966_),
    .ZN(_11967_)
  );
  AND2_X1 _19647_ (
    .A1(_08541_),
    .A2(_11967_),
    .ZN(_11968_)
  );
  AND2_X1 _19648_ (
    .A1(_11965_),
    .A2(_11968_),
    .ZN(_11969_)
  );
  INV_X1 _19649_ (
    .A(_11969_),
    .ZN(_11970_)
  );
  AND2_X1 _19650_ (
    .A1(\rf[24] [17]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11971_)
  );
  INV_X1 _19651_ (
    .A(_11971_),
    .ZN(_11972_)
  );
  AND2_X1 _19652_ (
    .A1(\rf[28] [17]),
    .A2(_08542_),
    .ZN(_11973_)
  );
  INV_X1 _19653_ (
    .A(_11973_),
    .ZN(_11974_)
  );
  AND2_X1 _19654_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_11974_),
    .ZN(_11975_)
  );
  AND2_X1 _19655_ (
    .A1(_11972_),
    .A2(_11975_),
    .ZN(_11976_)
  );
  INV_X1 _19656_ (
    .A(_11976_),
    .ZN(_11977_)
  );
  AND2_X1 _19657_ (
    .A1(_11970_),
    .A2(_11977_),
    .ZN(_11978_)
  );
  MUX2_X1 _19658_ (
    .A(\rf[29] [17]),
    .B(\rf[25] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_11979_)
  );
  AND2_X1 _19659_ (
    .A1(\rf[27] [17]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_11980_)
  );
  MUX2_X1 _19660_ (
    .A(_11979_),
    .B(_11980_),
    .S(_08541_),
    .Z(_11981_)
  );
  MUX2_X1 _19661_ (
    .A(_11978_),
    .B(_11981_),
    .S(_08540_),
    .Z(_11982_)
  );
  INV_X1 _19662_ (
    .A(_11982_),
    .ZN(_11983_)
  );
  AND2_X1 _19663_ (
    .A1(_08571_),
    .A2(_11983_),
    .ZN(_11984_)
  );
  INV_X1 _19664_ (
    .A(_11984_),
    .ZN(_11985_)
  );
  AND2_X1 _19665_ (
    .A1(_11963_),
    .A2(_11985_),
    .ZN(_11986_)
  );
  MUX2_X1 _19666_ (
    .A(_11926_),
    .B(_11986_),
    .S(_08543_),
    .Z(_11987_)
  );
  MUX2_X1 _19667_ (
    .A(_11987_),
    .B(_11882_),
    .S(_10131_),
    .Z(_11988_)
  );
  AND2_X1 _19668_ (
    .A1(_10082_),
    .A2(_11988_),
    .ZN(_11989_)
  );
  INV_X1 _19669_ (
    .A(_11989_),
    .ZN(_11990_)
  );
  AND2_X1 _19670_ (
    .A1(_11879_),
    .A2(_11990_),
    .ZN(_11991_)
  );
  INV_X1 _19671_ (
    .A(_11991_),
    .ZN(_11992_)
  );
  MUX2_X1 _19672_ (
    .A(ex_reg_rs_msb_0[15]),
    .B(_11992_),
    .S(_10079_),
    .Z(_00082_)
  );
  AND2_X1 _19673_ (
    .A1(_08578_),
    .A2(ibuf_io_inst_0_bits_raw[18]),
    .ZN(_11993_)
  );
  AND2_X1 _19674_ (
    .A1(_09295_),
    .A2(_11993_),
    .ZN(_11994_)
  );
  INV_X1 _19675_ (
    .A(_11994_),
    .ZN(_11995_)
  );
  MUX2_X1 _19676_ (
    .A(\rf[3] [18]),
    .B(\rf[2] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_11996_)
  );
  MUX2_X1 _19677_ (
    .A(\rf[7] [18]),
    .B(\rf[6] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_11997_)
  );
  MUX2_X1 _19678_ (
    .A(_11996_),
    .B(_11997_),
    .S(_08542_),
    .Z(_11998_)
  );
  INV_X1 _19679_ (
    .A(_11998_),
    .ZN(_11999_)
  );
  AND2_X1 _19680_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_11999_),
    .ZN(_12000_)
  );
  INV_X1 _19681_ (
    .A(_12000_),
    .ZN(_12001_)
  );
  MUX2_X1 _19682_ (
    .A(\rf[14] [18]),
    .B(\rf[10] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12002_)
  );
  INV_X1 _19683_ (
    .A(_12002_),
    .ZN(_12003_)
  );
  AND2_X1 _19684_ (
    .A1(_10213_),
    .A2(_12003_),
    .ZN(_12004_)
  );
  INV_X1 _19685_ (
    .A(_12004_),
    .ZN(_12005_)
  );
  MUX2_X1 _19686_ (
    .A(\rf[15] [18]),
    .B(\rf[11] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12006_)
  );
  INV_X1 _19687_ (
    .A(_12006_),
    .ZN(_12007_)
  );
  AND2_X1 _19688_ (
    .A1(_09110_),
    .A2(_12007_),
    .ZN(_12008_)
  );
  INV_X1 _19689_ (
    .A(_12008_),
    .ZN(_12009_)
  );
  AND2_X1 _19690_ (
    .A1(_12005_),
    .A2(_12009_),
    .ZN(_12010_)
  );
  AND2_X1 _19691_ (
    .A1(_12001_),
    .A2(_12010_),
    .ZN(_12011_)
  );
  AND2_X1 _19692_ (
    .A1(_08541_),
    .A2(_12011_),
    .ZN(_12012_)
  );
  INV_X1 _19693_ (
    .A(_12012_),
    .ZN(_12013_)
  );
  MUX2_X1 _19694_ (
    .A(\rf[1] [18]),
    .B(\rf[0] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_12014_)
  );
  MUX2_X1 _19695_ (
    .A(\rf[5] [18]),
    .B(\rf[4] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_12015_)
  );
  MUX2_X1 _19696_ (
    .A(_12014_),
    .B(_12015_),
    .S(_08542_),
    .Z(_12016_)
  );
  INV_X1 _19697_ (
    .A(_12016_),
    .ZN(_12017_)
  );
  AND2_X1 _19698_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_12017_),
    .ZN(_12018_)
  );
  INV_X1 _19699_ (
    .A(_12018_),
    .ZN(_12019_)
  );
  MUX2_X1 _19700_ (
    .A(\rf[13] [18]),
    .B(\rf[9] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12020_)
  );
  INV_X1 _19701_ (
    .A(_12020_),
    .ZN(_12021_)
  );
  AND2_X1 _19702_ (
    .A1(_09110_),
    .A2(_12021_),
    .ZN(_12022_)
  );
  INV_X1 _19703_ (
    .A(_12022_),
    .ZN(_12023_)
  );
  MUX2_X1 _19704_ (
    .A(\rf[12] [18]),
    .B(\rf[8] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12024_)
  );
  INV_X1 _19705_ (
    .A(_12024_),
    .ZN(_12025_)
  );
  AND2_X1 _19706_ (
    .A1(_10213_),
    .A2(_12025_),
    .ZN(_12026_)
  );
  INV_X1 _19707_ (
    .A(_12026_),
    .ZN(_12027_)
  );
  AND2_X1 _19708_ (
    .A1(_12023_),
    .A2(_12027_),
    .ZN(_12028_)
  );
  AND2_X1 _19709_ (
    .A1(_12019_),
    .A2(_12028_),
    .ZN(_12029_)
  );
  AND2_X1 _19710_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12029_),
    .ZN(_12030_)
  );
  INV_X1 _19711_ (
    .A(_12030_),
    .ZN(_12031_)
  );
  AND2_X1 _19712_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_12031_),
    .ZN(_12032_)
  );
  AND2_X1 _19713_ (
    .A1(_12013_),
    .A2(_12032_),
    .ZN(_12033_)
  );
  INV_X1 _19714_ (
    .A(_12033_),
    .ZN(_12034_)
  );
  AND2_X1 _19715_ (
    .A1(\rf[30] [18]),
    .A2(_08542_),
    .ZN(_12035_)
  );
  INV_X1 _19716_ (
    .A(_12035_),
    .ZN(_12036_)
  );
  AND2_X1 _19717_ (
    .A1(\rf[26] [18]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12037_)
  );
  INV_X1 _19718_ (
    .A(_12037_),
    .ZN(_12038_)
  );
  AND2_X1 _19719_ (
    .A1(_08541_),
    .A2(_12038_),
    .ZN(_12039_)
  );
  AND2_X1 _19720_ (
    .A1(_12036_),
    .A2(_12039_),
    .ZN(_12040_)
  );
  INV_X1 _19721_ (
    .A(_12040_),
    .ZN(_12041_)
  );
  AND2_X1 _19722_ (
    .A1(\rf[24] [18]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12042_)
  );
  INV_X1 _19723_ (
    .A(_12042_),
    .ZN(_12043_)
  );
  AND2_X1 _19724_ (
    .A1(\rf[28] [18]),
    .A2(_08542_),
    .ZN(_12044_)
  );
  INV_X1 _19725_ (
    .A(_12044_),
    .ZN(_12045_)
  );
  AND2_X1 _19726_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12045_),
    .ZN(_12046_)
  );
  AND2_X1 _19727_ (
    .A1(_12043_),
    .A2(_12046_),
    .ZN(_12047_)
  );
  INV_X1 _19728_ (
    .A(_12047_),
    .ZN(_12048_)
  );
  AND2_X1 _19729_ (
    .A1(_12041_),
    .A2(_12048_),
    .ZN(_12049_)
  );
  MUX2_X1 _19730_ (
    .A(\rf[29] [18]),
    .B(\rf[25] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12050_)
  );
  AND2_X1 _19731_ (
    .A1(\rf[27] [18]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12051_)
  );
  MUX2_X1 _19732_ (
    .A(_12050_),
    .B(_12051_),
    .S(_08541_),
    .Z(_12052_)
  );
  MUX2_X1 _19733_ (
    .A(_12049_),
    .B(_12052_),
    .S(_08540_),
    .Z(_12053_)
  );
  AND2_X1 _19734_ (
    .A1(_08391_),
    .A2(_08542_),
    .ZN(_12054_)
  );
  INV_X1 _19735_ (
    .A(_12054_),
    .ZN(_12055_)
  );
  AND2_X1 _19736_ (
    .A1(_08292_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12056_)
  );
  INV_X1 _19737_ (
    .A(_12056_),
    .ZN(_12057_)
  );
  AND2_X1 _19738_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12057_),
    .ZN(_12058_)
  );
  AND2_X1 _19739_ (
    .A1(_12055_),
    .A2(_12058_),
    .ZN(_12059_)
  );
  INV_X1 _19740_ (
    .A(_12059_),
    .ZN(_12060_)
  );
  MUX2_X1 _19741_ (
    .A(\rf[22] [18]),
    .B(\rf[18] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12061_)
  );
  AND2_X1 _19742_ (
    .A1(_08541_),
    .A2(_12061_),
    .ZN(_12062_)
  );
  INV_X1 _19743_ (
    .A(_12062_),
    .ZN(_12063_)
  );
  AND2_X1 _19744_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_12063_),
    .ZN(_12064_)
  );
  AND2_X1 _19745_ (
    .A1(_12060_),
    .A2(_12064_),
    .ZN(_12065_)
  );
  INV_X1 _19746_ (
    .A(_12065_),
    .ZN(_12066_)
  );
  AND2_X1 _19747_ (
    .A1(_08322_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12067_)
  );
  INV_X1 _19748_ (
    .A(_12067_),
    .ZN(_12068_)
  );
  AND2_X1 _19749_ (
    .A1(_08421_),
    .A2(_08542_),
    .ZN(_12069_)
  );
  INV_X1 _19750_ (
    .A(_12069_),
    .ZN(_12070_)
  );
  AND2_X1 _19751_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12070_),
    .ZN(_12071_)
  );
  AND2_X1 _19752_ (
    .A1(_12068_),
    .A2(_12071_),
    .ZN(_12072_)
  );
  INV_X1 _19753_ (
    .A(_12072_),
    .ZN(_12073_)
  );
  MUX2_X1 _19754_ (
    .A(\rf[23] [18]),
    .B(\rf[19] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12074_)
  );
  AND2_X1 _19755_ (
    .A1(_08541_),
    .A2(_12074_),
    .ZN(_12075_)
  );
  INV_X1 _19756_ (
    .A(_12075_),
    .ZN(_12076_)
  );
  AND2_X1 _19757_ (
    .A1(_08540_),
    .A2(_12076_),
    .ZN(_12077_)
  );
  AND2_X1 _19758_ (
    .A1(_12073_),
    .A2(_12077_),
    .ZN(_12078_)
  );
  INV_X1 _19759_ (
    .A(_12078_),
    .ZN(_12079_)
  );
  AND2_X1 _19760_ (
    .A1(_12066_),
    .A2(_12079_),
    .ZN(_12080_)
  );
  MUX2_X1 _19761_ (
    .A(_12053_),
    .B(_12080_),
    .S(ibuf_io_inst_0_bits_inst_rs1[3]),
    .Z(_12081_)
  );
  INV_X1 _19762_ (
    .A(_12081_),
    .ZN(_12082_)
  );
  AND2_X1 _19763_ (
    .A1(_08571_),
    .A2(_12082_),
    .ZN(_12083_)
  );
  INV_X1 _19764_ (
    .A(_12083_),
    .ZN(_12084_)
  );
  AND2_X1 _19765_ (
    .A1(_12034_),
    .A2(_12084_),
    .ZN(_12085_)
  );
  MUX2_X1 _19766_ (
    .A(csr_io_rw_rdata[18]),
    .B(wb_reg_wdata[18]),
    .S(_10134_),
    .Z(_12086_)
  );
  MUX2_X1 _19767_ (
    .A(div_io_resp_bits_data[18]),
    .B(_12086_),
    .S(_08649_),
    .Z(_12087_)
  );
  MUX2_X1 _19768_ (
    .A(_12087_),
    .B(io_dmem_resp_bits_data[18]),
    .S(_08631_),
    .Z(_12088_)
  );
  MUX2_X1 _19769_ (
    .A(_12085_),
    .B(_12088_),
    .S(_10131_),
    .Z(_12089_)
  );
  AND2_X1 _19770_ (
    .A1(_10082_),
    .A2(_12089_),
    .ZN(_12090_)
  );
  INV_X1 _19771_ (
    .A(_12090_),
    .ZN(_12091_)
  );
  AND2_X1 _19772_ (
    .A1(_11995_),
    .A2(_12091_),
    .ZN(_12092_)
  );
  INV_X1 _19773_ (
    .A(_12092_),
    .ZN(_12093_)
  );
  MUX2_X1 _19774_ (
    .A(ex_reg_rs_msb_0[16]),
    .B(_12093_),
    .S(_10079_),
    .Z(_00083_)
  );
  AND2_X1 _19775_ (
    .A1(_08578_),
    .A2(ibuf_io_inst_0_bits_raw[19]),
    .ZN(_12094_)
  );
  AND2_X1 _19776_ (
    .A1(_09295_),
    .A2(_12094_),
    .ZN(_12095_)
  );
  INV_X1 _19777_ (
    .A(_12095_),
    .ZN(_12096_)
  );
  MUX2_X1 _19778_ (
    .A(csr_io_rw_rdata[19]),
    .B(wb_reg_wdata[19]),
    .S(_10134_),
    .Z(_12097_)
  );
  MUX2_X1 _19779_ (
    .A(div_io_resp_bits_data[19]),
    .B(_12097_),
    .S(_08649_),
    .Z(_12098_)
  );
  MUX2_X1 _19780_ (
    .A(_12098_),
    .B(io_dmem_resp_bits_data[19]),
    .S(_08631_),
    .Z(_12099_)
  );
  MUX2_X1 _19781_ (
    .A(\rf[1] [19]),
    .B(\rf[0] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_12100_)
  );
  MUX2_X1 _19782_ (
    .A(\rf[5] [19]),
    .B(\rf[4] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_12101_)
  );
  MUX2_X1 _19783_ (
    .A(_12100_),
    .B(_12101_),
    .S(_08542_),
    .Z(_12102_)
  );
  INV_X1 _19784_ (
    .A(_12102_),
    .ZN(_12103_)
  );
  AND2_X1 _19785_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_12103_),
    .ZN(_12104_)
  );
  INV_X1 _19786_ (
    .A(_12104_),
    .ZN(_12105_)
  );
  MUX2_X1 _19787_ (
    .A(\rf[12] [19]),
    .B(\rf[8] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12106_)
  );
  INV_X1 _19788_ (
    .A(_12106_),
    .ZN(_12107_)
  );
  AND2_X1 _19789_ (
    .A1(_10213_),
    .A2(_12107_),
    .ZN(_12108_)
  );
  INV_X1 _19790_ (
    .A(_12108_),
    .ZN(_12109_)
  );
  MUX2_X1 _19791_ (
    .A(\rf[13] [19]),
    .B(\rf[9] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12110_)
  );
  INV_X1 _19792_ (
    .A(_12110_),
    .ZN(_12111_)
  );
  AND2_X1 _19793_ (
    .A1(_09110_),
    .A2(_12111_),
    .ZN(_12112_)
  );
  INV_X1 _19794_ (
    .A(_12112_),
    .ZN(_12113_)
  );
  AND2_X1 _19795_ (
    .A1(_12109_),
    .A2(_12113_),
    .ZN(_12114_)
  );
  AND2_X1 _19796_ (
    .A1(_12105_),
    .A2(_12114_),
    .ZN(_12115_)
  );
  AND2_X1 _19797_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12115_),
    .ZN(_12116_)
  );
  INV_X1 _19798_ (
    .A(_12116_),
    .ZN(_12117_)
  );
  MUX2_X1 _19799_ (
    .A(\rf[3] [19]),
    .B(\rf[2] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_12118_)
  );
  MUX2_X1 _19800_ (
    .A(\rf[7] [19]),
    .B(\rf[6] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_12119_)
  );
  MUX2_X1 _19801_ (
    .A(_12118_),
    .B(_12119_),
    .S(_08542_),
    .Z(_12120_)
  );
  INV_X1 _19802_ (
    .A(_12120_),
    .ZN(_12121_)
  );
  AND2_X1 _19803_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_12121_),
    .ZN(_12122_)
  );
  INV_X1 _19804_ (
    .A(_12122_),
    .ZN(_12123_)
  );
  MUX2_X1 _19805_ (
    .A(\rf[14] [19]),
    .B(\rf[10] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12124_)
  );
  INV_X1 _19806_ (
    .A(_12124_),
    .ZN(_12125_)
  );
  AND2_X1 _19807_ (
    .A1(_10213_),
    .A2(_12125_),
    .ZN(_12126_)
  );
  INV_X1 _19808_ (
    .A(_12126_),
    .ZN(_12127_)
  );
  MUX2_X1 _19809_ (
    .A(\rf[15] [19]),
    .B(\rf[11] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12128_)
  );
  INV_X1 _19810_ (
    .A(_12128_),
    .ZN(_12129_)
  );
  AND2_X1 _19811_ (
    .A1(_09110_),
    .A2(_12129_),
    .ZN(_12130_)
  );
  INV_X1 _19812_ (
    .A(_12130_),
    .ZN(_12131_)
  );
  AND2_X1 _19813_ (
    .A1(_12127_),
    .A2(_12131_),
    .ZN(_12132_)
  );
  AND2_X1 _19814_ (
    .A1(_08541_),
    .A2(_12132_),
    .ZN(_12133_)
  );
  AND2_X1 _19815_ (
    .A1(_12123_),
    .A2(_12133_),
    .ZN(_12134_)
  );
  INV_X1 _19816_ (
    .A(_12134_),
    .ZN(_12135_)
  );
  AND2_X1 _19817_ (
    .A1(\rf[30] [19]),
    .A2(_08542_),
    .ZN(_12136_)
  );
  INV_X1 _19818_ (
    .A(_12136_),
    .ZN(_12137_)
  );
  AND2_X1 _19819_ (
    .A1(\rf[26] [19]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12138_)
  );
  INV_X1 _19820_ (
    .A(_12138_),
    .ZN(_12139_)
  );
  AND2_X1 _19821_ (
    .A1(_08541_),
    .A2(_12139_),
    .ZN(_12140_)
  );
  AND2_X1 _19822_ (
    .A1(_12137_),
    .A2(_12140_),
    .ZN(_12141_)
  );
  INV_X1 _19823_ (
    .A(_12141_),
    .ZN(_12142_)
  );
  AND2_X1 _19824_ (
    .A1(\rf[24] [19]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12143_)
  );
  INV_X1 _19825_ (
    .A(_12143_),
    .ZN(_12144_)
  );
  AND2_X1 _19826_ (
    .A1(\rf[28] [19]),
    .A2(_08542_),
    .ZN(_12145_)
  );
  INV_X1 _19827_ (
    .A(_12145_),
    .ZN(_12146_)
  );
  AND2_X1 _19828_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12146_),
    .ZN(_12147_)
  );
  AND2_X1 _19829_ (
    .A1(_12144_),
    .A2(_12147_),
    .ZN(_12148_)
  );
  INV_X1 _19830_ (
    .A(_12148_),
    .ZN(_12149_)
  );
  AND2_X1 _19831_ (
    .A1(_12142_),
    .A2(_12149_),
    .ZN(_12150_)
  );
  MUX2_X1 _19832_ (
    .A(\rf[29] [19]),
    .B(\rf[25] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12151_)
  );
  AND2_X1 _19833_ (
    .A1(\rf[27] [19]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12152_)
  );
  MUX2_X1 _19834_ (
    .A(_12151_),
    .B(_12152_),
    .S(_08541_),
    .Z(_12153_)
  );
  MUX2_X1 _19835_ (
    .A(_12150_),
    .B(_12153_),
    .S(_08540_),
    .Z(_12154_)
  );
  AND2_X1 _19836_ (
    .A1(_08392_),
    .A2(_08542_),
    .ZN(_12155_)
  );
  INV_X1 _19837_ (
    .A(_12155_),
    .ZN(_12156_)
  );
  AND2_X1 _19838_ (
    .A1(_08293_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12157_)
  );
  INV_X1 _19839_ (
    .A(_12157_),
    .ZN(_12158_)
  );
  AND2_X1 _19840_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12158_),
    .ZN(_12159_)
  );
  AND2_X1 _19841_ (
    .A1(_12156_),
    .A2(_12159_),
    .ZN(_12160_)
  );
  INV_X1 _19842_ (
    .A(_12160_),
    .ZN(_12161_)
  );
  MUX2_X1 _19843_ (
    .A(\rf[22] [19]),
    .B(\rf[18] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12162_)
  );
  AND2_X1 _19844_ (
    .A1(_08541_),
    .A2(_12162_),
    .ZN(_12163_)
  );
  INV_X1 _19845_ (
    .A(_12163_),
    .ZN(_12164_)
  );
  AND2_X1 _19846_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_12164_),
    .ZN(_12165_)
  );
  AND2_X1 _19847_ (
    .A1(_12161_),
    .A2(_12165_),
    .ZN(_12166_)
  );
  INV_X1 _19848_ (
    .A(_12166_),
    .ZN(_12167_)
  );
  AND2_X1 _19849_ (
    .A1(_08323_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12168_)
  );
  INV_X1 _19850_ (
    .A(_12168_),
    .ZN(_12169_)
  );
  AND2_X1 _19851_ (
    .A1(_08422_),
    .A2(_08542_),
    .ZN(_12170_)
  );
  INV_X1 _19852_ (
    .A(_12170_),
    .ZN(_12171_)
  );
  AND2_X1 _19853_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12171_),
    .ZN(_12172_)
  );
  AND2_X1 _19854_ (
    .A1(_12169_),
    .A2(_12172_),
    .ZN(_12173_)
  );
  INV_X1 _19855_ (
    .A(_12173_),
    .ZN(_12174_)
  );
  MUX2_X1 _19856_ (
    .A(\rf[23] [19]),
    .B(\rf[19] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12175_)
  );
  AND2_X1 _19857_ (
    .A1(_08541_),
    .A2(_12175_),
    .ZN(_12176_)
  );
  INV_X1 _19858_ (
    .A(_12176_),
    .ZN(_12177_)
  );
  AND2_X1 _19859_ (
    .A1(_08540_),
    .A2(_12177_),
    .ZN(_12178_)
  );
  AND2_X1 _19860_ (
    .A1(_12174_),
    .A2(_12178_),
    .ZN(_12179_)
  );
  INV_X1 _19861_ (
    .A(_12179_),
    .ZN(_12180_)
  );
  AND2_X1 _19862_ (
    .A1(_12167_),
    .A2(_12180_),
    .ZN(_12181_)
  );
  MUX2_X1 _19863_ (
    .A(_12154_),
    .B(_12181_),
    .S(ibuf_io_inst_0_bits_inst_rs1[3]),
    .Z(_12182_)
  );
  AND2_X1 _19864_ (
    .A1(_12117_),
    .A2(_12135_),
    .ZN(_12183_)
  );
  INV_X1 _19865_ (
    .A(_12183_),
    .ZN(_12184_)
  );
  MUX2_X1 _19866_ (
    .A(_12182_),
    .B(_12184_),
    .S(ibuf_io_inst_0_bits_inst_rs1[4]),
    .Z(_12185_)
  );
  MUX2_X1 _19867_ (
    .A(_12185_),
    .B(_12099_),
    .S(_10131_),
    .Z(_12186_)
  );
  AND2_X1 _19868_ (
    .A1(_10082_),
    .A2(_12186_),
    .ZN(_12187_)
  );
  INV_X1 _19869_ (
    .A(_12187_),
    .ZN(_12188_)
  );
  AND2_X1 _19870_ (
    .A1(_12096_),
    .A2(_12188_),
    .ZN(_12189_)
  );
  INV_X1 _19871_ (
    .A(_12189_),
    .ZN(_12190_)
  );
  MUX2_X1 _19872_ (
    .A(ex_reg_rs_msb_0[17]),
    .B(_12190_),
    .S(_10079_),
    .Z(_00084_)
  );
  AND2_X1 _19873_ (
    .A1(_08578_),
    .A2(ibuf_io_inst_0_bits_raw[20]),
    .ZN(_12191_)
  );
  AND2_X1 _19874_ (
    .A1(_09295_),
    .A2(_12191_),
    .ZN(_12192_)
  );
  INV_X1 _19875_ (
    .A(_12192_),
    .ZN(_12193_)
  );
  AND2_X1 _19876_ (
    .A1(_08343_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12194_)
  );
  INV_X1 _19877_ (
    .A(_12194_),
    .ZN(_12195_)
  );
  AND2_X1 _19878_ (
    .A1(_08481_),
    .A2(_08542_),
    .ZN(_12196_)
  );
  INV_X1 _19879_ (
    .A(_12196_),
    .ZN(_12197_)
  );
  AND2_X1 _19880_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_12197_),
    .ZN(_12198_)
  );
  AND2_X1 _19881_ (
    .A1(_12195_),
    .A2(_12198_),
    .ZN(_12199_)
  );
  INV_X1 _19882_ (
    .A(_12199_),
    .ZN(_12200_)
  );
  MUX2_X1 _19883_ (
    .A(\rf[15] [20]),
    .B(\rf[11] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12201_)
  );
  AND2_X1 _19884_ (
    .A1(_08540_),
    .A2(_12201_),
    .ZN(_12202_)
  );
  INV_X1 _19885_ (
    .A(_12202_),
    .ZN(_12203_)
  );
  AND2_X1 _19886_ (
    .A1(_08541_),
    .A2(_12203_),
    .ZN(_12204_)
  );
  AND2_X1 _19887_ (
    .A1(_12200_),
    .A2(_12204_),
    .ZN(_12205_)
  );
  INV_X1 _19888_ (
    .A(_12205_),
    .ZN(_12206_)
  );
  AND2_X1 _19889_ (
    .A1(_08364_),
    .A2(_08542_),
    .ZN(_12207_)
  );
  INV_X1 _19890_ (
    .A(_12207_),
    .ZN(_12208_)
  );
  AND2_X1 _19891_ (
    .A1(_08265_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12209_)
  );
  INV_X1 _19892_ (
    .A(_12209_),
    .ZN(_12210_)
  );
  AND2_X1 _19893_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_12210_),
    .ZN(_12211_)
  );
  AND2_X1 _19894_ (
    .A1(_12208_),
    .A2(_12211_),
    .ZN(_12212_)
  );
  INV_X1 _19895_ (
    .A(_12212_),
    .ZN(_12213_)
  );
  MUX2_X1 _19896_ (
    .A(\rf[13] [20]),
    .B(\rf[9] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12214_)
  );
  AND2_X1 _19897_ (
    .A1(_08540_),
    .A2(_12214_),
    .ZN(_12215_)
  );
  INV_X1 _19898_ (
    .A(_12215_),
    .ZN(_12216_)
  );
  AND2_X1 _19899_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12216_),
    .ZN(_12217_)
  );
  AND2_X1 _19900_ (
    .A1(_12213_),
    .A2(_12217_),
    .ZN(_12218_)
  );
  INV_X1 _19901_ (
    .A(_12218_),
    .ZN(_12219_)
  );
  AND2_X1 _19902_ (
    .A1(_08543_),
    .A2(_12219_),
    .ZN(_12220_)
  );
  AND2_X1 _19903_ (
    .A1(_12206_),
    .A2(_12220_),
    .ZN(_12221_)
  );
  INV_X1 _19904_ (
    .A(_12221_),
    .ZN(_12222_)
  );
  AND2_X1 _19905_ (
    .A1(_08255_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12223_)
  );
  INV_X1 _19906_ (
    .A(_12223_),
    .ZN(_12224_)
  );
  AND2_X1 _19907_ (
    .A1(_08250_),
    .A2(_08542_),
    .ZN(_12225_)
  );
  INV_X1 _19908_ (
    .A(_12225_),
    .ZN(_12226_)
  );
  AND2_X1 _19909_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_12226_),
    .ZN(_12227_)
  );
  AND2_X1 _19910_ (
    .A1(_12224_),
    .A2(_12227_),
    .ZN(_12228_)
  );
  INV_X1 _19911_ (
    .A(_12228_),
    .ZN(_12229_)
  );
  MUX2_X1 _19912_ (
    .A(\rf[5] [20]),
    .B(\rf[1] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12230_)
  );
  AND2_X1 _19913_ (
    .A1(_08540_),
    .A2(_12230_),
    .ZN(_12231_)
  );
  INV_X1 _19914_ (
    .A(_12231_),
    .ZN(_12232_)
  );
  AND2_X1 _19915_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12232_),
    .ZN(_12233_)
  );
  AND2_X1 _19916_ (
    .A1(_12229_),
    .A2(_12233_),
    .ZN(_12234_)
  );
  INV_X1 _19917_ (
    .A(_12234_),
    .ZN(_12235_)
  );
  MUX2_X1 _19918_ (
    .A(\rf[7] [20]),
    .B(\rf[3] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12236_)
  );
  AND2_X1 _19919_ (
    .A1(_08540_),
    .A2(_12236_),
    .ZN(_12237_)
  );
  INV_X1 _19920_ (
    .A(_12237_),
    .ZN(_12238_)
  );
  AND2_X1 _19921_ (
    .A1(_08502_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12239_)
  );
  INV_X1 _19922_ (
    .A(_12239_),
    .ZN(_12240_)
  );
  AND2_X1 _19923_ (
    .A1(_08246_),
    .A2(_08542_),
    .ZN(_12241_)
  );
  INV_X1 _19924_ (
    .A(_12241_),
    .ZN(_12242_)
  );
  AND2_X1 _19925_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_12242_),
    .ZN(_12243_)
  );
  AND2_X1 _19926_ (
    .A1(_12240_),
    .A2(_12243_),
    .ZN(_12244_)
  );
  INV_X1 _19927_ (
    .A(_12244_),
    .ZN(_12245_)
  );
  AND2_X1 _19928_ (
    .A1(_12238_),
    .A2(_12245_),
    .ZN(_12246_)
  );
  AND2_X1 _19929_ (
    .A1(_08541_),
    .A2(_12246_),
    .ZN(_12247_)
  );
  INV_X1 _19930_ (
    .A(_12247_),
    .ZN(_12248_)
  );
  AND2_X1 _19931_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_12235_),
    .ZN(_12249_)
  );
  AND2_X1 _19932_ (
    .A1(_12248_),
    .A2(_12249_),
    .ZN(_12250_)
  );
  INV_X1 _19933_ (
    .A(_12250_),
    .ZN(_12251_)
  );
  AND2_X1 _19934_ (
    .A1(_12222_),
    .A2(_12251_),
    .ZN(_12252_)
  );
  MUX2_X1 _19935_ (
    .A(\rf[30] [20]),
    .B(\rf[26] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12253_)
  );
  AND2_X1 _19936_ (
    .A1(\rf[27] [20]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12254_)
  );
  MUX2_X1 _19937_ (
    .A(_12253_),
    .B(_12254_),
    .S(_08540_),
    .Z(_12255_)
  );
  INV_X1 _19938_ (
    .A(_12255_),
    .ZN(_12256_)
  );
  MUX2_X1 _19939_ (
    .A(\rf[29] [20]),
    .B(\rf[25] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12257_)
  );
  AND2_X1 _19940_ (
    .A1(_08540_),
    .A2(_12257_),
    .ZN(_12258_)
  );
  INV_X1 _19941_ (
    .A(_12258_),
    .ZN(_12259_)
  );
  MUX2_X1 _19942_ (
    .A(\rf[28] [20]),
    .B(\rf[24] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12260_)
  );
  AND2_X1 _19943_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_12260_),
    .ZN(_12261_)
  );
  INV_X1 _19944_ (
    .A(_12261_),
    .ZN(_12262_)
  );
  AND2_X1 _19945_ (
    .A1(_08541_),
    .A2(_12256_),
    .ZN(_12263_)
  );
  INV_X1 _19946_ (
    .A(_12263_),
    .ZN(_12264_)
  );
  AND2_X1 _19947_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12262_),
    .ZN(_12265_)
  );
  AND2_X1 _19948_ (
    .A1(_12259_),
    .A2(_12265_),
    .ZN(_12266_)
  );
  INV_X1 _19949_ (
    .A(_12266_),
    .ZN(_12267_)
  );
  AND2_X1 _19950_ (
    .A1(_08543_),
    .A2(_12264_),
    .ZN(_12268_)
  );
  AND2_X1 _19951_ (
    .A1(_12267_),
    .A2(_12268_),
    .ZN(_12269_)
  );
  INV_X1 _19952_ (
    .A(_12269_),
    .ZN(_12270_)
  );
  AND2_X1 _19953_ (
    .A1(_08354_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12271_)
  );
  INV_X1 _19954_ (
    .A(_12271_),
    .ZN(_12272_)
  );
  AND2_X1 _19955_ (
    .A1(_08492_),
    .A2(_08542_),
    .ZN(_12273_)
  );
  INV_X1 _19956_ (
    .A(_12273_),
    .ZN(_12274_)
  );
  AND2_X1 _19957_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_12274_),
    .ZN(_12275_)
  );
  AND2_X1 _19958_ (
    .A1(_12272_),
    .A2(_12275_),
    .ZN(_12276_)
  );
  INV_X1 _19959_ (
    .A(_12276_),
    .ZN(_12277_)
  );
  MUX2_X1 _19960_ (
    .A(\rf[23] [20]),
    .B(\rf[19] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12278_)
  );
  AND2_X1 _19961_ (
    .A1(_08540_),
    .A2(_12278_),
    .ZN(_12279_)
  );
  INV_X1 _19962_ (
    .A(_12279_),
    .ZN(_12280_)
  );
  AND2_X1 _19963_ (
    .A1(_08541_),
    .A2(_12280_),
    .ZN(_12281_)
  );
  AND2_X1 _19964_ (
    .A1(_12277_),
    .A2(_12281_),
    .ZN(_12282_)
  );
  INV_X1 _19965_ (
    .A(_12282_),
    .ZN(_12283_)
  );
  MUX2_X1 _19966_ (
    .A(\rf[21] [20]),
    .B(\rf[17] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12284_)
  );
  AND2_X1 _19967_ (
    .A1(_08540_),
    .A2(_12284_),
    .ZN(_12285_)
  );
  INV_X1 _19968_ (
    .A(_12285_),
    .ZN(_12286_)
  );
  AND2_X1 _19969_ (
    .A1(_08393_),
    .A2(_08542_),
    .ZN(_12287_)
  );
  INV_X1 _19970_ (
    .A(_12287_),
    .ZN(_12288_)
  );
  AND2_X1 _19971_ (
    .A1(_08294_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12289_)
  );
  INV_X1 _19972_ (
    .A(_12289_),
    .ZN(_12290_)
  );
  AND2_X1 _19973_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_12290_),
    .ZN(_12291_)
  );
  AND2_X1 _19974_ (
    .A1(_12288_),
    .A2(_12291_),
    .ZN(_12292_)
  );
  INV_X1 _19975_ (
    .A(_12292_),
    .ZN(_12293_)
  );
  AND2_X1 _19976_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12286_),
    .ZN(_12294_)
  );
  AND2_X1 _19977_ (
    .A1(_12293_),
    .A2(_12294_),
    .ZN(_12295_)
  );
  INV_X1 _19978_ (
    .A(_12295_),
    .ZN(_12296_)
  );
  AND2_X1 _19979_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_12283_),
    .ZN(_12297_)
  );
  AND2_X1 _19980_ (
    .A1(_12296_),
    .A2(_12297_),
    .ZN(_12298_)
  );
  INV_X1 _19981_ (
    .A(_12298_),
    .ZN(_12299_)
  );
  AND2_X1 _19982_ (
    .A1(_12270_),
    .A2(_12299_),
    .ZN(_12300_)
  );
  MUX2_X1 _19983_ (
    .A(_12252_),
    .B(_12300_),
    .S(_08571_),
    .Z(_12301_)
  );
  INV_X1 _19984_ (
    .A(_12301_),
    .ZN(_12302_)
  );
  MUX2_X1 _19985_ (
    .A(csr_io_rw_rdata[20]),
    .B(wb_reg_wdata[20]),
    .S(_10134_),
    .Z(_12303_)
  );
  MUX2_X1 _19986_ (
    .A(div_io_resp_bits_data[20]),
    .B(_12303_),
    .S(_08649_),
    .Z(_12304_)
  );
  MUX2_X1 _19987_ (
    .A(_12304_),
    .B(io_dmem_resp_bits_data[20]),
    .S(_08631_),
    .Z(_12305_)
  );
  MUX2_X1 _19988_ (
    .A(_12302_),
    .B(_12305_),
    .S(_10131_),
    .Z(_12306_)
  );
  AND2_X1 _19989_ (
    .A1(_10082_),
    .A2(_12306_),
    .ZN(_12307_)
  );
  INV_X1 _19990_ (
    .A(_12307_),
    .ZN(_12308_)
  );
  AND2_X1 _19991_ (
    .A1(_12193_),
    .A2(_12308_),
    .ZN(_12309_)
  );
  INV_X1 _19992_ (
    .A(_12309_),
    .ZN(_12310_)
  );
  MUX2_X1 _19993_ (
    .A(ex_reg_rs_msb_0[18]),
    .B(_12310_),
    .S(_10079_),
    .Z(_00085_)
  );
  AND2_X1 _19994_ (
    .A1(_08578_),
    .A2(ibuf_io_inst_0_bits_raw[21]),
    .ZN(_12311_)
  );
  AND2_X1 _19995_ (
    .A1(_09295_),
    .A2(_12311_),
    .ZN(_12312_)
  );
  INV_X1 _19996_ (
    .A(_12312_),
    .ZN(_12313_)
  );
  MUX2_X1 _19997_ (
    .A(csr_io_rw_rdata[21]),
    .B(wb_reg_wdata[21]),
    .S(_10134_),
    .Z(_12314_)
  );
  MUX2_X1 _19998_ (
    .A(div_io_resp_bits_data[21]),
    .B(_12314_),
    .S(_08649_),
    .Z(_12315_)
  );
  MUX2_X1 _19999_ (
    .A(_12315_),
    .B(io_dmem_resp_bits_data[21]),
    .S(_08631_),
    .Z(_12316_)
  );
  MUX2_X1 _20000_ (
    .A(\rf[5] [21]),
    .B(\rf[1] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12317_)
  );
  MUX2_X1 _20001_ (
    .A(\rf[7] [21]),
    .B(\rf[3] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12318_)
  );
  MUX2_X1 _20002_ (
    .A(_12317_),
    .B(_12318_),
    .S(_08541_),
    .Z(_12319_)
  );
  AND2_X1 _20003_ (
    .A1(_08540_),
    .A2(_12319_),
    .ZN(_12320_)
  );
  INV_X1 _20004_ (
    .A(_12320_),
    .ZN(_12321_)
  );
  MUX2_X1 _20005_ (
    .A(\rf[4] [21]),
    .B(\rf[0] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12322_)
  );
  MUX2_X1 _20006_ (
    .A(\rf[6] [21]),
    .B(\rf[2] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12323_)
  );
  MUX2_X1 _20007_ (
    .A(_12322_),
    .B(_12323_),
    .S(_08541_),
    .Z(_12324_)
  );
  AND2_X1 _20008_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_12324_),
    .ZN(_12325_)
  );
  INV_X1 _20009_ (
    .A(_12325_),
    .ZN(_12326_)
  );
  AND2_X1 _20010_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_12326_),
    .ZN(_12327_)
  );
  AND2_X1 _20011_ (
    .A1(_12321_),
    .A2(_12327_),
    .ZN(_12328_)
  );
  INV_X1 _20012_ (
    .A(_12328_),
    .ZN(_12329_)
  );
  AND2_X1 _20013_ (
    .A1(_08394_),
    .A2(_08542_),
    .ZN(_12330_)
  );
  INV_X1 _20014_ (
    .A(_12330_),
    .ZN(_12331_)
  );
  AND2_X1 _20015_ (
    .A1(_08295_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12332_)
  );
  INV_X1 _20016_ (
    .A(_12332_),
    .ZN(_12333_)
  );
  AND2_X1 _20017_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12333_),
    .ZN(_12334_)
  );
  AND2_X1 _20018_ (
    .A1(_12331_),
    .A2(_12334_),
    .ZN(_12335_)
  );
  INV_X1 _20019_ (
    .A(_12335_),
    .ZN(_12336_)
  );
  MUX2_X1 _20020_ (
    .A(\rf[22] [21]),
    .B(\rf[18] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12337_)
  );
  AND2_X1 _20021_ (
    .A1(_08541_),
    .A2(_12337_),
    .ZN(_12338_)
  );
  INV_X1 _20022_ (
    .A(_12338_),
    .ZN(_12339_)
  );
  AND2_X1 _20023_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_12339_),
    .ZN(_12340_)
  );
  AND2_X1 _20024_ (
    .A1(_12336_),
    .A2(_12340_),
    .ZN(_12341_)
  );
  INV_X1 _20025_ (
    .A(_12341_),
    .ZN(_12342_)
  );
  AND2_X1 _20026_ (
    .A1(_08325_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12343_)
  );
  INV_X1 _20027_ (
    .A(_12343_),
    .ZN(_12344_)
  );
  AND2_X1 _20028_ (
    .A1(_08424_),
    .A2(_08542_),
    .ZN(_12345_)
  );
  INV_X1 _20029_ (
    .A(_12345_),
    .ZN(_12346_)
  );
  AND2_X1 _20030_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12346_),
    .ZN(_12347_)
  );
  AND2_X1 _20031_ (
    .A1(_12344_),
    .A2(_12347_),
    .ZN(_12348_)
  );
  INV_X1 _20032_ (
    .A(_12348_),
    .ZN(_12349_)
  );
  MUX2_X1 _20033_ (
    .A(\rf[23] [21]),
    .B(\rf[19] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12350_)
  );
  AND2_X1 _20034_ (
    .A1(_08541_),
    .A2(_12350_),
    .ZN(_12351_)
  );
  INV_X1 _20035_ (
    .A(_12351_),
    .ZN(_12352_)
  );
  AND2_X1 _20036_ (
    .A1(_08540_),
    .A2(_12352_),
    .ZN(_12353_)
  );
  AND2_X1 _20037_ (
    .A1(_12349_),
    .A2(_12353_),
    .ZN(_12354_)
  );
  INV_X1 _20038_ (
    .A(_12354_),
    .ZN(_12355_)
  );
  AND2_X1 _20039_ (
    .A1(_12342_),
    .A2(_12355_),
    .ZN(_12356_)
  );
  INV_X1 _20040_ (
    .A(_12356_),
    .ZN(_12357_)
  );
  AND2_X1 _20041_ (
    .A1(_08571_),
    .A2(_12357_),
    .ZN(_12358_)
  );
  INV_X1 _20042_ (
    .A(_12358_),
    .ZN(_12359_)
  );
  AND2_X1 _20043_ (
    .A1(_12329_),
    .A2(_12359_),
    .ZN(_12360_)
  );
  AND2_X1 _20044_ (
    .A1(\rf[10] [21]),
    .A2(_08541_),
    .ZN(_12361_)
  );
  INV_X1 _20045_ (
    .A(_12361_),
    .ZN(_12362_)
  );
  AND2_X1 _20046_ (
    .A1(\rf[8] [21]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_12363_)
  );
  INV_X1 _20047_ (
    .A(_12363_),
    .ZN(_12364_)
  );
  AND2_X1 _20048_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_12364_),
    .ZN(_12365_)
  );
  AND2_X1 _20049_ (
    .A1(_12362_),
    .A2(_12365_),
    .ZN(_12366_)
  );
  INV_X1 _20050_ (
    .A(_12366_),
    .ZN(_12367_)
  );
  AND2_X1 _20051_ (
    .A1(\rf[14] [21]),
    .A2(_08541_),
    .ZN(_12368_)
  );
  INV_X1 _20052_ (
    .A(_12368_),
    .ZN(_12369_)
  );
  AND2_X1 _20053_ (
    .A1(\rf[12] [21]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_12370_)
  );
  INV_X1 _20054_ (
    .A(_12370_),
    .ZN(_12371_)
  );
  AND2_X1 _20055_ (
    .A1(_08542_),
    .A2(_12371_),
    .ZN(_12372_)
  );
  AND2_X1 _20056_ (
    .A1(_12369_),
    .A2(_12372_),
    .ZN(_12373_)
  );
  INV_X1 _20057_ (
    .A(_12373_),
    .ZN(_12374_)
  );
  AND2_X1 _20058_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_12374_),
    .ZN(_12375_)
  );
  AND2_X1 _20059_ (
    .A1(_12367_),
    .A2(_12375_),
    .ZN(_12376_)
  );
  INV_X1 _20060_ (
    .A(_12376_),
    .ZN(_12377_)
  );
  AND2_X1 _20061_ (
    .A1(\rf[11] [21]),
    .A2(_08541_),
    .ZN(_12378_)
  );
  INV_X1 _20062_ (
    .A(_12378_),
    .ZN(_12379_)
  );
  AND2_X1 _20063_ (
    .A1(\rf[9] [21]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_12380_)
  );
  INV_X1 _20064_ (
    .A(_12380_),
    .ZN(_12381_)
  );
  AND2_X1 _20065_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_12381_),
    .ZN(_12382_)
  );
  AND2_X1 _20066_ (
    .A1(_12379_),
    .A2(_12382_),
    .ZN(_12383_)
  );
  INV_X1 _20067_ (
    .A(_12383_),
    .ZN(_12384_)
  );
  AND2_X1 _20068_ (
    .A1(\rf[15] [21]),
    .A2(_08541_),
    .ZN(_12385_)
  );
  INV_X1 _20069_ (
    .A(_12385_),
    .ZN(_12386_)
  );
  AND2_X1 _20070_ (
    .A1(\rf[13] [21]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_12387_)
  );
  INV_X1 _20071_ (
    .A(_12387_),
    .ZN(_12388_)
  );
  AND2_X1 _20072_ (
    .A1(_08542_),
    .A2(_12388_),
    .ZN(_12389_)
  );
  AND2_X1 _20073_ (
    .A1(_12386_),
    .A2(_12389_),
    .ZN(_12390_)
  );
  INV_X1 _20074_ (
    .A(_12390_),
    .ZN(_12391_)
  );
  AND2_X1 _20075_ (
    .A1(_08540_),
    .A2(_12391_),
    .ZN(_12392_)
  );
  AND2_X1 _20076_ (
    .A1(_12384_),
    .A2(_12392_),
    .ZN(_12393_)
  );
  INV_X1 _20077_ (
    .A(_12393_),
    .ZN(_12394_)
  );
  AND2_X1 _20078_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_12394_),
    .ZN(_12395_)
  );
  AND2_X1 _20079_ (
    .A1(_12377_),
    .A2(_12395_),
    .ZN(_12396_)
  );
  INV_X1 _20080_ (
    .A(_12396_),
    .ZN(_12397_)
  );
  AND2_X1 _20081_ (
    .A1(\rf[30] [21]),
    .A2(_08542_),
    .ZN(_12398_)
  );
  INV_X1 _20082_ (
    .A(_12398_),
    .ZN(_12399_)
  );
  AND2_X1 _20083_ (
    .A1(\rf[26] [21]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12400_)
  );
  INV_X1 _20084_ (
    .A(_12400_),
    .ZN(_12401_)
  );
  AND2_X1 _20085_ (
    .A1(_08541_),
    .A2(_12401_),
    .ZN(_12402_)
  );
  AND2_X1 _20086_ (
    .A1(_12399_),
    .A2(_12402_),
    .ZN(_12403_)
  );
  INV_X1 _20087_ (
    .A(_12403_),
    .ZN(_12404_)
  );
  AND2_X1 _20088_ (
    .A1(\rf[24] [21]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12405_)
  );
  INV_X1 _20089_ (
    .A(_12405_),
    .ZN(_12406_)
  );
  AND2_X1 _20090_ (
    .A1(\rf[28] [21]),
    .A2(_08542_),
    .ZN(_12407_)
  );
  INV_X1 _20091_ (
    .A(_12407_),
    .ZN(_12408_)
  );
  AND2_X1 _20092_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12408_),
    .ZN(_12409_)
  );
  AND2_X1 _20093_ (
    .A1(_12406_),
    .A2(_12409_),
    .ZN(_12410_)
  );
  INV_X1 _20094_ (
    .A(_12410_),
    .ZN(_12411_)
  );
  AND2_X1 _20095_ (
    .A1(_12404_),
    .A2(_12411_),
    .ZN(_12412_)
  );
  MUX2_X1 _20096_ (
    .A(\rf[29] [21]),
    .B(\rf[25] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12413_)
  );
  AND2_X1 _20097_ (
    .A1(\rf[27] [21]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12414_)
  );
  MUX2_X1 _20098_ (
    .A(_12413_),
    .B(_12414_),
    .S(_08541_),
    .Z(_12415_)
  );
  MUX2_X1 _20099_ (
    .A(_12412_),
    .B(_12415_),
    .S(_08540_),
    .Z(_12416_)
  );
  INV_X1 _20100_ (
    .A(_12416_),
    .ZN(_12417_)
  );
  AND2_X1 _20101_ (
    .A1(_08571_),
    .A2(_12417_),
    .ZN(_12418_)
  );
  INV_X1 _20102_ (
    .A(_12418_),
    .ZN(_12419_)
  );
  AND2_X1 _20103_ (
    .A1(_12397_),
    .A2(_12419_),
    .ZN(_12420_)
  );
  MUX2_X1 _20104_ (
    .A(_12360_),
    .B(_12420_),
    .S(_08543_),
    .Z(_12421_)
  );
  MUX2_X1 _20105_ (
    .A(_12421_),
    .B(_12316_),
    .S(_10131_),
    .Z(_12422_)
  );
  AND2_X1 _20106_ (
    .A1(_10082_),
    .A2(_12422_),
    .ZN(_12423_)
  );
  INV_X1 _20107_ (
    .A(_12423_),
    .ZN(_12424_)
  );
  AND2_X1 _20108_ (
    .A1(_12313_),
    .A2(_12424_),
    .ZN(_12425_)
  );
  INV_X1 _20109_ (
    .A(_12425_),
    .ZN(_12426_)
  );
  MUX2_X1 _20110_ (
    .A(ex_reg_rs_msb_0[19]),
    .B(_12426_),
    .S(_10079_),
    .Z(_00086_)
  );
  AND2_X1 _20111_ (
    .A1(_08578_),
    .A2(ibuf_io_inst_0_bits_raw[22]),
    .ZN(_12427_)
  );
  AND2_X1 _20112_ (
    .A1(_09295_),
    .A2(_12427_),
    .ZN(_12428_)
  );
  INV_X1 _20113_ (
    .A(_12428_),
    .ZN(_12429_)
  );
  MUX2_X1 _20114_ (
    .A(\rf[5] [22]),
    .B(\rf[1] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12430_)
  );
  MUX2_X1 _20115_ (
    .A(\rf[7] [22]),
    .B(\rf[3] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12431_)
  );
  MUX2_X1 _20116_ (
    .A(_12430_),
    .B(_12431_),
    .S(_08541_),
    .Z(_12432_)
  );
  AND2_X1 _20117_ (
    .A1(_08540_),
    .A2(_12432_),
    .ZN(_12433_)
  );
  INV_X1 _20118_ (
    .A(_12433_),
    .ZN(_12434_)
  );
  MUX2_X1 _20119_ (
    .A(\rf[4] [22]),
    .B(\rf[0] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12435_)
  );
  MUX2_X1 _20120_ (
    .A(\rf[6] [22]),
    .B(\rf[2] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12436_)
  );
  MUX2_X1 _20121_ (
    .A(_12435_),
    .B(_12436_),
    .S(_08541_),
    .Z(_12437_)
  );
  AND2_X1 _20122_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_12437_),
    .ZN(_12438_)
  );
  INV_X1 _20123_ (
    .A(_12438_),
    .ZN(_12439_)
  );
  AND2_X1 _20124_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_12439_),
    .ZN(_12440_)
  );
  AND2_X1 _20125_ (
    .A1(_12434_),
    .A2(_12440_),
    .ZN(_12441_)
  );
  INV_X1 _20126_ (
    .A(_12441_),
    .ZN(_12442_)
  );
  AND2_X1 _20127_ (
    .A1(_08395_),
    .A2(_08542_),
    .ZN(_12443_)
  );
  INV_X1 _20128_ (
    .A(_12443_),
    .ZN(_12444_)
  );
  AND2_X1 _20129_ (
    .A1(_08296_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12445_)
  );
  INV_X1 _20130_ (
    .A(_12445_),
    .ZN(_12446_)
  );
  AND2_X1 _20131_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12446_),
    .ZN(_12447_)
  );
  AND2_X1 _20132_ (
    .A1(_12444_),
    .A2(_12447_),
    .ZN(_12448_)
  );
  INV_X1 _20133_ (
    .A(_12448_),
    .ZN(_12449_)
  );
  MUX2_X1 _20134_ (
    .A(\rf[22] [22]),
    .B(\rf[18] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12450_)
  );
  AND2_X1 _20135_ (
    .A1(_08541_),
    .A2(_12450_),
    .ZN(_12451_)
  );
  INV_X1 _20136_ (
    .A(_12451_),
    .ZN(_12452_)
  );
  AND2_X1 _20137_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_12452_),
    .ZN(_12453_)
  );
  AND2_X1 _20138_ (
    .A1(_12449_),
    .A2(_12453_),
    .ZN(_12454_)
  );
  INV_X1 _20139_ (
    .A(_12454_),
    .ZN(_12455_)
  );
  AND2_X1 _20140_ (
    .A1(_08326_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12456_)
  );
  INV_X1 _20141_ (
    .A(_12456_),
    .ZN(_12457_)
  );
  AND2_X1 _20142_ (
    .A1(_08425_),
    .A2(_08542_),
    .ZN(_12458_)
  );
  INV_X1 _20143_ (
    .A(_12458_),
    .ZN(_12459_)
  );
  AND2_X1 _20144_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12459_),
    .ZN(_12460_)
  );
  AND2_X1 _20145_ (
    .A1(_12457_),
    .A2(_12460_),
    .ZN(_12461_)
  );
  INV_X1 _20146_ (
    .A(_12461_),
    .ZN(_12462_)
  );
  MUX2_X1 _20147_ (
    .A(\rf[23] [22]),
    .B(\rf[19] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12463_)
  );
  AND2_X1 _20148_ (
    .A1(_08541_),
    .A2(_12463_),
    .ZN(_12464_)
  );
  INV_X1 _20149_ (
    .A(_12464_),
    .ZN(_12465_)
  );
  AND2_X1 _20150_ (
    .A1(_08540_),
    .A2(_12465_),
    .ZN(_12466_)
  );
  AND2_X1 _20151_ (
    .A1(_12462_),
    .A2(_12466_),
    .ZN(_12467_)
  );
  INV_X1 _20152_ (
    .A(_12467_),
    .ZN(_12468_)
  );
  AND2_X1 _20153_ (
    .A1(_12455_),
    .A2(_12468_),
    .ZN(_12469_)
  );
  INV_X1 _20154_ (
    .A(_12469_),
    .ZN(_12470_)
  );
  AND2_X1 _20155_ (
    .A1(_08571_),
    .A2(_12470_),
    .ZN(_12471_)
  );
  INV_X1 _20156_ (
    .A(_12471_),
    .ZN(_12472_)
  );
  AND2_X1 _20157_ (
    .A1(_12442_),
    .A2(_12472_),
    .ZN(_12473_)
  );
  AND2_X1 _20158_ (
    .A1(\rf[10] [22]),
    .A2(_08541_),
    .ZN(_12474_)
  );
  INV_X1 _20159_ (
    .A(_12474_),
    .ZN(_12475_)
  );
  AND2_X1 _20160_ (
    .A1(\rf[8] [22]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_12476_)
  );
  INV_X1 _20161_ (
    .A(_12476_),
    .ZN(_12477_)
  );
  AND2_X1 _20162_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_12477_),
    .ZN(_12478_)
  );
  AND2_X1 _20163_ (
    .A1(_12475_),
    .A2(_12478_),
    .ZN(_12479_)
  );
  INV_X1 _20164_ (
    .A(_12479_),
    .ZN(_12480_)
  );
  AND2_X1 _20165_ (
    .A1(\rf[14] [22]),
    .A2(_08541_),
    .ZN(_12481_)
  );
  INV_X1 _20166_ (
    .A(_12481_),
    .ZN(_12482_)
  );
  AND2_X1 _20167_ (
    .A1(\rf[12] [22]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_12483_)
  );
  INV_X1 _20168_ (
    .A(_12483_),
    .ZN(_12484_)
  );
  AND2_X1 _20169_ (
    .A1(_08542_),
    .A2(_12484_),
    .ZN(_12485_)
  );
  AND2_X1 _20170_ (
    .A1(_12482_),
    .A2(_12485_),
    .ZN(_12486_)
  );
  INV_X1 _20171_ (
    .A(_12486_),
    .ZN(_12487_)
  );
  AND2_X1 _20172_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_12487_),
    .ZN(_12488_)
  );
  AND2_X1 _20173_ (
    .A1(_12480_),
    .A2(_12488_),
    .ZN(_12489_)
  );
  INV_X1 _20174_ (
    .A(_12489_),
    .ZN(_12490_)
  );
  AND2_X1 _20175_ (
    .A1(\rf[11] [22]),
    .A2(_08541_),
    .ZN(_12491_)
  );
  INV_X1 _20176_ (
    .A(_12491_),
    .ZN(_12492_)
  );
  AND2_X1 _20177_ (
    .A1(\rf[9] [22]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_12493_)
  );
  INV_X1 _20178_ (
    .A(_12493_),
    .ZN(_12494_)
  );
  AND2_X1 _20179_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_12494_),
    .ZN(_12495_)
  );
  AND2_X1 _20180_ (
    .A1(_12492_),
    .A2(_12495_),
    .ZN(_12496_)
  );
  INV_X1 _20181_ (
    .A(_12496_),
    .ZN(_12497_)
  );
  AND2_X1 _20182_ (
    .A1(\rf[15] [22]),
    .A2(_08541_),
    .ZN(_12498_)
  );
  INV_X1 _20183_ (
    .A(_12498_),
    .ZN(_12499_)
  );
  AND2_X1 _20184_ (
    .A1(\rf[13] [22]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_12500_)
  );
  INV_X1 _20185_ (
    .A(_12500_),
    .ZN(_12501_)
  );
  AND2_X1 _20186_ (
    .A1(_08542_),
    .A2(_12501_),
    .ZN(_12502_)
  );
  AND2_X1 _20187_ (
    .A1(_12499_),
    .A2(_12502_),
    .ZN(_12503_)
  );
  INV_X1 _20188_ (
    .A(_12503_),
    .ZN(_12504_)
  );
  AND2_X1 _20189_ (
    .A1(_08540_),
    .A2(_12504_),
    .ZN(_12505_)
  );
  AND2_X1 _20190_ (
    .A1(_12497_),
    .A2(_12505_),
    .ZN(_12506_)
  );
  INV_X1 _20191_ (
    .A(_12506_),
    .ZN(_12507_)
  );
  AND2_X1 _20192_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_12507_),
    .ZN(_12508_)
  );
  AND2_X1 _20193_ (
    .A1(_12490_),
    .A2(_12508_),
    .ZN(_12509_)
  );
  INV_X1 _20194_ (
    .A(_12509_),
    .ZN(_12510_)
  );
  AND2_X1 _20195_ (
    .A1(\rf[30] [22]),
    .A2(_08542_),
    .ZN(_12511_)
  );
  INV_X1 _20196_ (
    .A(_12511_),
    .ZN(_12512_)
  );
  AND2_X1 _20197_ (
    .A1(\rf[26] [22]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12513_)
  );
  INV_X1 _20198_ (
    .A(_12513_),
    .ZN(_12514_)
  );
  AND2_X1 _20199_ (
    .A1(_08541_),
    .A2(_12514_),
    .ZN(_12515_)
  );
  AND2_X1 _20200_ (
    .A1(_12512_),
    .A2(_12515_),
    .ZN(_12516_)
  );
  INV_X1 _20201_ (
    .A(_12516_),
    .ZN(_12517_)
  );
  AND2_X1 _20202_ (
    .A1(\rf[24] [22]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12518_)
  );
  INV_X1 _20203_ (
    .A(_12518_),
    .ZN(_12519_)
  );
  AND2_X1 _20204_ (
    .A1(\rf[28] [22]),
    .A2(_08542_),
    .ZN(_12520_)
  );
  INV_X1 _20205_ (
    .A(_12520_),
    .ZN(_12521_)
  );
  AND2_X1 _20206_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12521_),
    .ZN(_12522_)
  );
  AND2_X1 _20207_ (
    .A1(_12519_),
    .A2(_12522_),
    .ZN(_12523_)
  );
  INV_X1 _20208_ (
    .A(_12523_),
    .ZN(_12524_)
  );
  AND2_X1 _20209_ (
    .A1(_12517_),
    .A2(_12524_),
    .ZN(_12525_)
  );
  MUX2_X1 _20210_ (
    .A(\rf[29] [22]),
    .B(\rf[25] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12526_)
  );
  AND2_X1 _20211_ (
    .A1(\rf[27] [22]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12527_)
  );
  MUX2_X1 _20212_ (
    .A(_12526_),
    .B(_12527_),
    .S(_08541_),
    .Z(_12528_)
  );
  MUX2_X1 _20213_ (
    .A(_12525_),
    .B(_12528_),
    .S(_08540_),
    .Z(_12529_)
  );
  INV_X1 _20214_ (
    .A(_12529_),
    .ZN(_12530_)
  );
  AND2_X1 _20215_ (
    .A1(_08571_),
    .A2(_12530_),
    .ZN(_12531_)
  );
  INV_X1 _20216_ (
    .A(_12531_),
    .ZN(_12532_)
  );
  AND2_X1 _20217_ (
    .A1(_12510_),
    .A2(_12532_),
    .ZN(_12533_)
  );
  MUX2_X1 _20218_ (
    .A(_12473_),
    .B(_12533_),
    .S(_08543_),
    .Z(_12534_)
  );
  MUX2_X1 _20219_ (
    .A(csr_io_rw_rdata[22]),
    .B(wb_reg_wdata[22]),
    .S(_10134_),
    .Z(_12535_)
  );
  MUX2_X1 _20220_ (
    .A(div_io_resp_bits_data[22]),
    .B(_12535_),
    .S(_08649_),
    .Z(_12536_)
  );
  MUX2_X1 _20221_ (
    .A(_12536_),
    .B(io_dmem_resp_bits_data[22]),
    .S(_08631_),
    .Z(_12537_)
  );
  MUX2_X1 _20222_ (
    .A(_12534_),
    .B(_12537_),
    .S(_10131_),
    .Z(_12538_)
  );
  AND2_X1 _20223_ (
    .A1(_10082_),
    .A2(_12538_),
    .ZN(_12539_)
  );
  INV_X1 _20224_ (
    .A(_12539_),
    .ZN(_12540_)
  );
  AND2_X1 _20225_ (
    .A1(_12429_),
    .A2(_12540_),
    .ZN(_12541_)
  );
  INV_X1 _20226_ (
    .A(_12541_),
    .ZN(_12542_)
  );
  MUX2_X1 _20227_ (
    .A(ex_reg_rs_msb_0[20]),
    .B(_12542_),
    .S(_10079_),
    .Z(_00087_)
  );
  AND2_X1 _20228_ (
    .A1(_08578_),
    .A2(ibuf_io_inst_0_bits_raw[23]),
    .ZN(_12543_)
  );
  AND2_X1 _20229_ (
    .A1(_09295_),
    .A2(_12543_),
    .ZN(_12544_)
  );
  INV_X1 _20230_ (
    .A(_12544_),
    .ZN(_12545_)
  );
  MUX2_X1 _20231_ (
    .A(\rf[3] [23]),
    .B(\rf[2] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_12546_)
  );
  MUX2_X1 _20232_ (
    .A(\rf[7] [23]),
    .B(\rf[6] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_12547_)
  );
  MUX2_X1 _20233_ (
    .A(_12546_),
    .B(_12547_),
    .S(_08542_),
    .Z(_12548_)
  );
  INV_X1 _20234_ (
    .A(_12548_),
    .ZN(_12549_)
  );
  AND2_X1 _20235_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_12549_),
    .ZN(_12550_)
  );
  INV_X1 _20236_ (
    .A(_12550_),
    .ZN(_12551_)
  );
  MUX2_X1 _20237_ (
    .A(\rf[15] [23]),
    .B(\rf[11] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12552_)
  );
  INV_X1 _20238_ (
    .A(_12552_),
    .ZN(_12553_)
  );
  AND2_X1 _20239_ (
    .A1(_09110_),
    .A2(_12553_),
    .ZN(_12554_)
  );
  INV_X1 _20240_ (
    .A(_12554_),
    .ZN(_12555_)
  );
  MUX2_X1 _20241_ (
    .A(\rf[14] [23]),
    .B(\rf[10] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12556_)
  );
  INV_X1 _20242_ (
    .A(_12556_),
    .ZN(_12557_)
  );
  AND2_X1 _20243_ (
    .A1(_10213_),
    .A2(_12557_),
    .ZN(_12558_)
  );
  INV_X1 _20244_ (
    .A(_12558_),
    .ZN(_12559_)
  );
  AND2_X1 _20245_ (
    .A1(_12555_),
    .A2(_12559_),
    .ZN(_12560_)
  );
  AND2_X1 _20246_ (
    .A1(_12551_),
    .A2(_12560_),
    .ZN(_12561_)
  );
  AND2_X1 _20247_ (
    .A1(_08541_),
    .A2(_12561_),
    .ZN(_12562_)
  );
  INV_X1 _20248_ (
    .A(_12562_),
    .ZN(_12563_)
  );
  MUX2_X1 _20249_ (
    .A(\rf[1] [23]),
    .B(\rf[0] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_12564_)
  );
  MUX2_X1 _20250_ (
    .A(\rf[5] [23]),
    .B(\rf[4] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_12565_)
  );
  MUX2_X1 _20251_ (
    .A(_12564_),
    .B(_12565_),
    .S(_08542_),
    .Z(_12566_)
  );
  INV_X1 _20252_ (
    .A(_12566_),
    .ZN(_12567_)
  );
  AND2_X1 _20253_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_12567_),
    .ZN(_12568_)
  );
  INV_X1 _20254_ (
    .A(_12568_),
    .ZN(_12569_)
  );
  MUX2_X1 _20255_ (
    .A(\rf[13] [23]),
    .B(\rf[9] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12570_)
  );
  INV_X1 _20256_ (
    .A(_12570_),
    .ZN(_12571_)
  );
  AND2_X1 _20257_ (
    .A1(_09110_),
    .A2(_12571_),
    .ZN(_12572_)
  );
  INV_X1 _20258_ (
    .A(_12572_),
    .ZN(_12573_)
  );
  MUX2_X1 _20259_ (
    .A(\rf[12] [23]),
    .B(\rf[8] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12574_)
  );
  INV_X1 _20260_ (
    .A(_12574_),
    .ZN(_12575_)
  );
  AND2_X1 _20261_ (
    .A1(_10213_),
    .A2(_12575_),
    .ZN(_12576_)
  );
  INV_X1 _20262_ (
    .A(_12576_),
    .ZN(_12577_)
  );
  AND2_X1 _20263_ (
    .A1(_12573_),
    .A2(_12577_),
    .ZN(_12578_)
  );
  AND2_X1 _20264_ (
    .A1(_12569_),
    .A2(_12578_),
    .ZN(_12579_)
  );
  AND2_X1 _20265_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12579_),
    .ZN(_12580_)
  );
  INV_X1 _20266_ (
    .A(_12580_),
    .ZN(_12581_)
  );
  AND2_X1 _20267_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_12581_),
    .ZN(_12582_)
  );
  AND2_X1 _20268_ (
    .A1(_12563_),
    .A2(_12582_),
    .ZN(_12583_)
  );
  INV_X1 _20269_ (
    .A(_12583_),
    .ZN(_12584_)
  );
  AND2_X1 _20270_ (
    .A1(\rf[30] [23]),
    .A2(_08542_),
    .ZN(_12585_)
  );
  INV_X1 _20271_ (
    .A(_12585_),
    .ZN(_12586_)
  );
  AND2_X1 _20272_ (
    .A1(\rf[26] [23]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12587_)
  );
  INV_X1 _20273_ (
    .A(_12587_),
    .ZN(_12588_)
  );
  AND2_X1 _20274_ (
    .A1(_08541_),
    .A2(_12588_),
    .ZN(_12589_)
  );
  AND2_X1 _20275_ (
    .A1(_12586_),
    .A2(_12589_),
    .ZN(_12590_)
  );
  INV_X1 _20276_ (
    .A(_12590_),
    .ZN(_12591_)
  );
  AND2_X1 _20277_ (
    .A1(\rf[24] [23]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12592_)
  );
  INV_X1 _20278_ (
    .A(_12592_),
    .ZN(_12593_)
  );
  AND2_X1 _20279_ (
    .A1(\rf[28] [23]),
    .A2(_08542_),
    .ZN(_12594_)
  );
  INV_X1 _20280_ (
    .A(_12594_),
    .ZN(_12595_)
  );
  AND2_X1 _20281_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12595_),
    .ZN(_12596_)
  );
  AND2_X1 _20282_ (
    .A1(_12593_),
    .A2(_12596_),
    .ZN(_12597_)
  );
  INV_X1 _20283_ (
    .A(_12597_),
    .ZN(_12598_)
  );
  AND2_X1 _20284_ (
    .A1(_12591_),
    .A2(_12598_),
    .ZN(_12599_)
  );
  MUX2_X1 _20285_ (
    .A(\rf[29] [23]),
    .B(\rf[25] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12600_)
  );
  AND2_X1 _20286_ (
    .A1(\rf[27] [23]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12601_)
  );
  MUX2_X1 _20287_ (
    .A(_12600_),
    .B(_12601_),
    .S(_08541_),
    .Z(_12602_)
  );
  MUX2_X1 _20288_ (
    .A(_12599_),
    .B(_12602_),
    .S(_08540_),
    .Z(_12603_)
  );
  AND2_X1 _20289_ (
    .A1(_08396_),
    .A2(_08542_),
    .ZN(_12604_)
  );
  INV_X1 _20290_ (
    .A(_12604_),
    .ZN(_12605_)
  );
  AND2_X1 _20291_ (
    .A1(_08297_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12606_)
  );
  INV_X1 _20292_ (
    .A(_12606_),
    .ZN(_12607_)
  );
  AND2_X1 _20293_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12607_),
    .ZN(_12608_)
  );
  AND2_X1 _20294_ (
    .A1(_12605_),
    .A2(_12608_),
    .ZN(_12609_)
  );
  INV_X1 _20295_ (
    .A(_12609_),
    .ZN(_12610_)
  );
  MUX2_X1 _20296_ (
    .A(\rf[22] [23]),
    .B(\rf[18] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12611_)
  );
  AND2_X1 _20297_ (
    .A1(_08541_),
    .A2(_12611_),
    .ZN(_12612_)
  );
  INV_X1 _20298_ (
    .A(_12612_),
    .ZN(_12613_)
  );
  AND2_X1 _20299_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_12613_),
    .ZN(_12614_)
  );
  AND2_X1 _20300_ (
    .A1(_12610_),
    .A2(_12614_),
    .ZN(_12615_)
  );
  INV_X1 _20301_ (
    .A(_12615_),
    .ZN(_12616_)
  );
  AND2_X1 _20302_ (
    .A1(_08327_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12617_)
  );
  INV_X1 _20303_ (
    .A(_12617_),
    .ZN(_12618_)
  );
  AND2_X1 _20304_ (
    .A1(_08426_),
    .A2(_08542_),
    .ZN(_12619_)
  );
  INV_X1 _20305_ (
    .A(_12619_),
    .ZN(_12620_)
  );
  AND2_X1 _20306_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12620_),
    .ZN(_12621_)
  );
  AND2_X1 _20307_ (
    .A1(_12618_),
    .A2(_12621_),
    .ZN(_12622_)
  );
  INV_X1 _20308_ (
    .A(_12622_),
    .ZN(_12623_)
  );
  MUX2_X1 _20309_ (
    .A(\rf[23] [23]),
    .B(\rf[19] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12624_)
  );
  AND2_X1 _20310_ (
    .A1(_08541_),
    .A2(_12624_),
    .ZN(_12625_)
  );
  INV_X1 _20311_ (
    .A(_12625_),
    .ZN(_12626_)
  );
  AND2_X1 _20312_ (
    .A1(_08540_),
    .A2(_12626_),
    .ZN(_12627_)
  );
  AND2_X1 _20313_ (
    .A1(_12623_),
    .A2(_12627_),
    .ZN(_12628_)
  );
  INV_X1 _20314_ (
    .A(_12628_),
    .ZN(_12629_)
  );
  AND2_X1 _20315_ (
    .A1(_12616_),
    .A2(_12629_),
    .ZN(_12630_)
  );
  MUX2_X1 _20316_ (
    .A(_12603_),
    .B(_12630_),
    .S(ibuf_io_inst_0_bits_inst_rs1[3]),
    .Z(_12631_)
  );
  INV_X1 _20317_ (
    .A(_12631_),
    .ZN(_12632_)
  );
  AND2_X1 _20318_ (
    .A1(_08571_),
    .A2(_12632_),
    .ZN(_12633_)
  );
  INV_X1 _20319_ (
    .A(_12633_),
    .ZN(_12634_)
  );
  AND2_X1 _20320_ (
    .A1(_12584_),
    .A2(_12634_),
    .ZN(_12635_)
  );
  MUX2_X1 _20321_ (
    .A(csr_io_rw_rdata[23]),
    .B(wb_reg_wdata[23]),
    .S(_10134_),
    .Z(_12636_)
  );
  MUX2_X1 _20322_ (
    .A(div_io_resp_bits_data[23]),
    .B(_12636_),
    .S(_08649_),
    .Z(_12637_)
  );
  MUX2_X1 _20323_ (
    .A(_12637_),
    .B(io_dmem_resp_bits_data[23]),
    .S(_08631_),
    .Z(_12638_)
  );
  MUX2_X1 _20324_ (
    .A(_12635_),
    .B(_12638_),
    .S(_10131_),
    .Z(_12639_)
  );
  AND2_X1 _20325_ (
    .A1(_10082_),
    .A2(_12639_),
    .ZN(_12640_)
  );
  INV_X1 _20326_ (
    .A(_12640_),
    .ZN(_12641_)
  );
  AND2_X1 _20327_ (
    .A1(_12545_),
    .A2(_12641_),
    .ZN(_12642_)
  );
  INV_X1 _20328_ (
    .A(_12642_),
    .ZN(_12643_)
  );
  MUX2_X1 _20329_ (
    .A(ex_reg_rs_msb_0[21]),
    .B(_12643_),
    .S(_10079_),
    .Z(_00088_)
  );
  AND2_X1 _20330_ (
    .A1(_08578_),
    .A2(ibuf_io_inst_0_bits_raw[24]),
    .ZN(_12644_)
  );
  AND2_X1 _20331_ (
    .A1(_09295_),
    .A2(_12644_),
    .ZN(_12645_)
  );
  INV_X1 _20332_ (
    .A(_12645_),
    .ZN(_12646_)
  );
  MUX2_X1 _20333_ (
    .A(csr_io_rw_rdata[24]),
    .B(wb_reg_wdata[24]),
    .S(_10134_),
    .Z(_12647_)
  );
  MUX2_X1 _20334_ (
    .A(div_io_resp_bits_data[24]),
    .B(_12647_),
    .S(_08649_),
    .Z(_12648_)
  );
  MUX2_X1 _20335_ (
    .A(_12648_),
    .B(io_dmem_resp_bits_data[24]),
    .S(_08631_),
    .Z(_12649_)
  );
  MUX2_X1 _20336_ (
    .A(\rf[5] [24]),
    .B(\rf[1] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12650_)
  );
  MUX2_X1 _20337_ (
    .A(\rf[7] [24]),
    .B(\rf[3] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12651_)
  );
  MUX2_X1 _20338_ (
    .A(_12650_),
    .B(_12651_),
    .S(_08541_),
    .Z(_12652_)
  );
  AND2_X1 _20339_ (
    .A1(_08540_),
    .A2(_12652_),
    .ZN(_12653_)
  );
  INV_X1 _20340_ (
    .A(_12653_),
    .ZN(_12654_)
  );
  MUX2_X1 _20341_ (
    .A(\rf[4] [24]),
    .B(\rf[0] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12655_)
  );
  MUX2_X1 _20342_ (
    .A(\rf[6] [24]),
    .B(\rf[2] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12656_)
  );
  MUX2_X1 _20343_ (
    .A(_12655_),
    .B(_12656_),
    .S(_08541_),
    .Z(_12657_)
  );
  AND2_X1 _20344_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_12657_),
    .ZN(_12658_)
  );
  INV_X1 _20345_ (
    .A(_12658_),
    .ZN(_12659_)
  );
  AND2_X1 _20346_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_12659_),
    .ZN(_12660_)
  );
  AND2_X1 _20347_ (
    .A1(_12654_),
    .A2(_12660_),
    .ZN(_12661_)
  );
  INV_X1 _20348_ (
    .A(_12661_),
    .ZN(_12662_)
  );
  AND2_X1 _20349_ (
    .A1(_08397_),
    .A2(_08542_),
    .ZN(_12663_)
  );
  INV_X1 _20350_ (
    .A(_12663_),
    .ZN(_12664_)
  );
  AND2_X1 _20351_ (
    .A1(_08298_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12665_)
  );
  INV_X1 _20352_ (
    .A(_12665_),
    .ZN(_12666_)
  );
  AND2_X1 _20353_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12666_),
    .ZN(_12667_)
  );
  AND2_X1 _20354_ (
    .A1(_12664_),
    .A2(_12667_),
    .ZN(_12668_)
  );
  INV_X1 _20355_ (
    .A(_12668_),
    .ZN(_12669_)
  );
  MUX2_X1 _20356_ (
    .A(\rf[22] [24]),
    .B(\rf[18] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12670_)
  );
  AND2_X1 _20357_ (
    .A1(_08541_),
    .A2(_12670_),
    .ZN(_12671_)
  );
  INV_X1 _20358_ (
    .A(_12671_),
    .ZN(_12672_)
  );
  AND2_X1 _20359_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_12672_),
    .ZN(_12673_)
  );
  AND2_X1 _20360_ (
    .A1(_12669_),
    .A2(_12673_),
    .ZN(_12674_)
  );
  INV_X1 _20361_ (
    .A(_12674_),
    .ZN(_12675_)
  );
  AND2_X1 _20362_ (
    .A1(_08328_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12676_)
  );
  INV_X1 _20363_ (
    .A(_12676_),
    .ZN(_12677_)
  );
  AND2_X1 _20364_ (
    .A1(_08427_),
    .A2(_08542_),
    .ZN(_12678_)
  );
  INV_X1 _20365_ (
    .A(_12678_),
    .ZN(_12679_)
  );
  AND2_X1 _20366_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12679_),
    .ZN(_12680_)
  );
  AND2_X1 _20367_ (
    .A1(_12677_),
    .A2(_12680_),
    .ZN(_12681_)
  );
  INV_X1 _20368_ (
    .A(_12681_),
    .ZN(_12682_)
  );
  MUX2_X1 _20369_ (
    .A(\rf[23] [24]),
    .B(\rf[19] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12683_)
  );
  AND2_X1 _20370_ (
    .A1(_08541_),
    .A2(_12683_),
    .ZN(_12684_)
  );
  INV_X1 _20371_ (
    .A(_12684_),
    .ZN(_12685_)
  );
  AND2_X1 _20372_ (
    .A1(_08540_),
    .A2(_12685_),
    .ZN(_12686_)
  );
  AND2_X1 _20373_ (
    .A1(_12682_),
    .A2(_12686_),
    .ZN(_12687_)
  );
  INV_X1 _20374_ (
    .A(_12687_),
    .ZN(_12688_)
  );
  AND2_X1 _20375_ (
    .A1(_12675_),
    .A2(_12688_),
    .ZN(_12689_)
  );
  INV_X1 _20376_ (
    .A(_12689_),
    .ZN(_12690_)
  );
  AND2_X1 _20377_ (
    .A1(_08571_),
    .A2(_12690_),
    .ZN(_12691_)
  );
  INV_X1 _20378_ (
    .A(_12691_),
    .ZN(_12692_)
  );
  AND2_X1 _20379_ (
    .A1(_12662_),
    .A2(_12692_),
    .ZN(_12693_)
  );
  AND2_X1 _20380_ (
    .A1(\rf[10] [24]),
    .A2(_08541_),
    .ZN(_12694_)
  );
  INV_X1 _20381_ (
    .A(_12694_),
    .ZN(_12695_)
  );
  AND2_X1 _20382_ (
    .A1(\rf[8] [24]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_12696_)
  );
  INV_X1 _20383_ (
    .A(_12696_),
    .ZN(_12697_)
  );
  AND2_X1 _20384_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_12697_),
    .ZN(_12698_)
  );
  AND2_X1 _20385_ (
    .A1(_12695_),
    .A2(_12698_),
    .ZN(_12699_)
  );
  INV_X1 _20386_ (
    .A(_12699_),
    .ZN(_12700_)
  );
  AND2_X1 _20387_ (
    .A1(\rf[14] [24]),
    .A2(_08541_),
    .ZN(_12701_)
  );
  INV_X1 _20388_ (
    .A(_12701_),
    .ZN(_12702_)
  );
  AND2_X1 _20389_ (
    .A1(\rf[12] [24]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_12703_)
  );
  INV_X1 _20390_ (
    .A(_12703_),
    .ZN(_12704_)
  );
  AND2_X1 _20391_ (
    .A1(_08542_),
    .A2(_12704_),
    .ZN(_12705_)
  );
  AND2_X1 _20392_ (
    .A1(_12702_),
    .A2(_12705_),
    .ZN(_12706_)
  );
  INV_X1 _20393_ (
    .A(_12706_),
    .ZN(_12707_)
  );
  AND2_X1 _20394_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_12707_),
    .ZN(_12708_)
  );
  AND2_X1 _20395_ (
    .A1(_12700_),
    .A2(_12708_),
    .ZN(_12709_)
  );
  INV_X1 _20396_ (
    .A(_12709_),
    .ZN(_12710_)
  );
  AND2_X1 _20397_ (
    .A1(\rf[11] [24]),
    .A2(_08541_),
    .ZN(_12711_)
  );
  INV_X1 _20398_ (
    .A(_12711_),
    .ZN(_12712_)
  );
  AND2_X1 _20399_ (
    .A1(\rf[9] [24]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_12713_)
  );
  INV_X1 _20400_ (
    .A(_12713_),
    .ZN(_12714_)
  );
  AND2_X1 _20401_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_12714_),
    .ZN(_12715_)
  );
  AND2_X1 _20402_ (
    .A1(_12712_),
    .A2(_12715_),
    .ZN(_12716_)
  );
  INV_X1 _20403_ (
    .A(_12716_),
    .ZN(_12717_)
  );
  AND2_X1 _20404_ (
    .A1(\rf[15] [24]),
    .A2(_08541_),
    .ZN(_12718_)
  );
  INV_X1 _20405_ (
    .A(_12718_),
    .ZN(_12719_)
  );
  AND2_X1 _20406_ (
    .A1(\rf[13] [24]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_12720_)
  );
  INV_X1 _20407_ (
    .A(_12720_),
    .ZN(_12721_)
  );
  AND2_X1 _20408_ (
    .A1(_08542_),
    .A2(_12721_),
    .ZN(_12722_)
  );
  AND2_X1 _20409_ (
    .A1(_12719_),
    .A2(_12722_),
    .ZN(_12723_)
  );
  INV_X1 _20410_ (
    .A(_12723_),
    .ZN(_12724_)
  );
  AND2_X1 _20411_ (
    .A1(_08540_),
    .A2(_12724_),
    .ZN(_12725_)
  );
  AND2_X1 _20412_ (
    .A1(_12717_),
    .A2(_12725_),
    .ZN(_12726_)
  );
  INV_X1 _20413_ (
    .A(_12726_),
    .ZN(_12727_)
  );
  AND2_X1 _20414_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_12727_),
    .ZN(_12728_)
  );
  AND2_X1 _20415_ (
    .A1(_12710_),
    .A2(_12728_),
    .ZN(_12729_)
  );
  INV_X1 _20416_ (
    .A(_12729_),
    .ZN(_12730_)
  );
  AND2_X1 _20417_ (
    .A1(\rf[30] [24]),
    .A2(_08542_),
    .ZN(_12731_)
  );
  INV_X1 _20418_ (
    .A(_12731_),
    .ZN(_12732_)
  );
  AND2_X1 _20419_ (
    .A1(\rf[26] [24]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12733_)
  );
  INV_X1 _20420_ (
    .A(_12733_),
    .ZN(_12734_)
  );
  AND2_X1 _20421_ (
    .A1(_08541_),
    .A2(_12734_),
    .ZN(_12735_)
  );
  AND2_X1 _20422_ (
    .A1(_12732_),
    .A2(_12735_),
    .ZN(_12736_)
  );
  INV_X1 _20423_ (
    .A(_12736_),
    .ZN(_12737_)
  );
  AND2_X1 _20424_ (
    .A1(\rf[24] [24]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12738_)
  );
  INV_X1 _20425_ (
    .A(_12738_),
    .ZN(_12739_)
  );
  AND2_X1 _20426_ (
    .A1(\rf[28] [24]),
    .A2(_08542_),
    .ZN(_12740_)
  );
  INV_X1 _20427_ (
    .A(_12740_),
    .ZN(_12741_)
  );
  AND2_X1 _20428_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12741_),
    .ZN(_12742_)
  );
  AND2_X1 _20429_ (
    .A1(_12739_),
    .A2(_12742_),
    .ZN(_12743_)
  );
  INV_X1 _20430_ (
    .A(_12743_),
    .ZN(_12744_)
  );
  AND2_X1 _20431_ (
    .A1(_12737_),
    .A2(_12744_),
    .ZN(_12745_)
  );
  MUX2_X1 _20432_ (
    .A(\rf[29] [24]),
    .B(\rf[25] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12746_)
  );
  AND2_X1 _20433_ (
    .A1(\rf[27] [24]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12747_)
  );
  MUX2_X1 _20434_ (
    .A(_12746_),
    .B(_12747_),
    .S(_08541_),
    .Z(_12748_)
  );
  MUX2_X1 _20435_ (
    .A(_12745_),
    .B(_12748_),
    .S(_08540_),
    .Z(_12749_)
  );
  INV_X1 _20436_ (
    .A(_12749_),
    .ZN(_12750_)
  );
  AND2_X1 _20437_ (
    .A1(_08571_),
    .A2(_12750_),
    .ZN(_12751_)
  );
  INV_X1 _20438_ (
    .A(_12751_),
    .ZN(_12752_)
  );
  AND2_X1 _20439_ (
    .A1(_12730_),
    .A2(_12752_),
    .ZN(_12753_)
  );
  MUX2_X1 _20440_ (
    .A(_12693_),
    .B(_12753_),
    .S(_08543_),
    .Z(_12754_)
  );
  MUX2_X1 _20441_ (
    .A(_12754_),
    .B(_12649_),
    .S(_10131_),
    .Z(_12755_)
  );
  AND2_X1 _20442_ (
    .A1(_10082_),
    .A2(_12755_),
    .ZN(_12756_)
  );
  INV_X1 _20443_ (
    .A(_12756_),
    .ZN(_12757_)
  );
  AND2_X1 _20444_ (
    .A1(_12646_),
    .A2(_12757_),
    .ZN(_12758_)
  );
  INV_X1 _20445_ (
    .A(_12758_),
    .ZN(_12759_)
  );
  MUX2_X1 _20446_ (
    .A(ex_reg_rs_msb_0[22]),
    .B(_12759_),
    .S(_10079_),
    .Z(_00089_)
  );
  AND2_X1 _20447_ (
    .A1(_08578_),
    .A2(ibuf_io_inst_0_bits_raw[25]),
    .ZN(_12760_)
  );
  AND2_X1 _20448_ (
    .A1(_09295_),
    .A2(_12760_),
    .ZN(_12761_)
  );
  INV_X1 _20449_ (
    .A(_12761_),
    .ZN(_12762_)
  );
  MUX2_X1 _20450_ (
    .A(csr_io_rw_rdata[25]),
    .B(wb_reg_wdata[25]),
    .S(_10134_),
    .Z(_12763_)
  );
  MUX2_X1 _20451_ (
    .A(div_io_resp_bits_data[25]),
    .B(_12763_),
    .S(_08649_),
    .Z(_12764_)
  );
  MUX2_X1 _20452_ (
    .A(_12764_),
    .B(io_dmem_resp_bits_data[25]),
    .S(_08631_),
    .Z(_12765_)
  );
  MUX2_X1 _20453_ (
    .A(\rf[5] [25]),
    .B(\rf[1] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12766_)
  );
  MUX2_X1 _20454_ (
    .A(\rf[7] [25]),
    .B(\rf[3] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12767_)
  );
  MUX2_X1 _20455_ (
    .A(_12766_),
    .B(_12767_),
    .S(_08541_),
    .Z(_12768_)
  );
  AND2_X1 _20456_ (
    .A1(_08540_),
    .A2(_12768_),
    .ZN(_12769_)
  );
  INV_X1 _20457_ (
    .A(_12769_),
    .ZN(_12770_)
  );
  MUX2_X1 _20458_ (
    .A(\rf[4] [25]),
    .B(\rf[0] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12771_)
  );
  MUX2_X1 _20459_ (
    .A(\rf[6] [25]),
    .B(\rf[2] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12772_)
  );
  MUX2_X1 _20460_ (
    .A(_12771_),
    .B(_12772_),
    .S(_08541_),
    .Z(_12773_)
  );
  AND2_X1 _20461_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_12773_),
    .ZN(_12774_)
  );
  INV_X1 _20462_ (
    .A(_12774_),
    .ZN(_12775_)
  );
  AND2_X1 _20463_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_12775_),
    .ZN(_12776_)
  );
  AND2_X1 _20464_ (
    .A1(_12770_),
    .A2(_12776_),
    .ZN(_12777_)
  );
  INV_X1 _20465_ (
    .A(_12777_),
    .ZN(_12778_)
  );
  AND2_X1 _20466_ (
    .A1(_08398_),
    .A2(_08542_),
    .ZN(_12779_)
  );
  INV_X1 _20467_ (
    .A(_12779_),
    .ZN(_12780_)
  );
  AND2_X1 _20468_ (
    .A1(_08299_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12781_)
  );
  INV_X1 _20469_ (
    .A(_12781_),
    .ZN(_12782_)
  );
  AND2_X1 _20470_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12782_),
    .ZN(_12783_)
  );
  AND2_X1 _20471_ (
    .A1(_12780_),
    .A2(_12783_),
    .ZN(_12784_)
  );
  INV_X1 _20472_ (
    .A(_12784_),
    .ZN(_12785_)
  );
  MUX2_X1 _20473_ (
    .A(\rf[22] [25]),
    .B(\rf[18] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12786_)
  );
  AND2_X1 _20474_ (
    .A1(_08541_),
    .A2(_12786_),
    .ZN(_12787_)
  );
  INV_X1 _20475_ (
    .A(_12787_),
    .ZN(_12788_)
  );
  AND2_X1 _20476_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_12788_),
    .ZN(_12789_)
  );
  AND2_X1 _20477_ (
    .A1(_12785_),
    .A2(_12789_),
    .ZN(_12790_)
  );
  INV_X1 _20478_ (
    .A(_12790_),
    .ZN(_12791_)
  );
  AND2_X1 _20479_ (
    .A1(_08329_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12792_)
  );
  INV_X1 _20480_ (
    .A(_12792_),
    .ZN(_12793_)
  );
  AND2_X1 _20481_ (
    .A1(_08428_),
    .A2(_08542_),
    .ZN(_12794_)
  );
  INV_X1 _20482_ (
    .A(_12794_),
    .ZN(_12795_)
  );
  AND2_X1 _20483_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12795_),
    .ZN(_12796_)
  );
  AND2_X1 _20484_ (
    .A1(_12793_),
    .A2(_12796_),
    .ZN(_12797_)
  );
  INV_X1 _20485_ (
    .A(_12797_),
    .ZN(_12798_)
  );
  MUX2_X1 _20486_ (
    .A(\rf[23] [25]),
    .B(\rf[19] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12799_)
  );
  AND2_X1 _20487_ (
    .A1(_08541_),
    .A2(_12799_),
    .ZN(_12800_)
  );
  INV_X1 _20488_ (
    .A(_12800_),
    .ZN(_12801_)
  );
  AND2_X1 _20489_ (
    .A1(_08540_),
    .A2(_12801_),
    .ZN(_12802_)
  );
  AND2_X1 _20490_ (
    .A1(_12798_),
    .A2(_12802_),
    .ZN(_12803_)
  );
  INV_X1 _20491_ (
    .A(_12803_),
    .ZN(_12804_)
  );
  AND2_X1 _20492_ (
    .A1(_12791_),
    .A2(_12804_),
    .ZN(_12805_)
  );
  INV_X1 _20493_ (
    .A(_12805_),
    .ZN(_12806_)
  );
  AND2_X1 _20494_ (
    .A1(_08571_),
    .A2(_12806_),
    .ZN(_12807_)
  );
  INV_X1 _20495_ (
    .A(_12807_),
    .ZN(_12808_)
  );
  AND2_X1 _20496_ (
    .A1(_12778_),
    .A2(_12808_),
    .ZN(_12809_)
  );
  AND2_X1 _20497_ (
    .A1(\rf[10] [25]),
    .A2(_08541_),
    .ZN(_12810_)
  );
  INV_X1 _20498_ (
    .A(_12810_),
    .ZN(_12811_)
  );
  AND2_X1 _20499_ (
    .A1(\rf[8] [25]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_12812_)
  );
  INV_X1 _20500_ (
    .A(_12812_),
    .ZN(_12813_)
  );
  AND2_X1 _20501_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_12813_),
    .ZN(_12814_)
  );
  AND2_X1 _20502_ (
    .A1(_12811_),
    .A2(_12814_),
    .ZN(_12815_)
  );
  INV_X1 _20503_ (
    .A(_12815_),
    .ZN(_12816_)
  );
  AND2_X1 _20504_ (
    .A1(\rf[14] [25]),
    .A2(_08541_),
    .ZN(_12817_)
  );
  INV_X1 _20505_ (
    .A(_12817_),
    .ZN(_12818_)
  );
  AND2_X1 _20506_ (
    .A1(\rf[12] [25]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_12819_)
  );
  INV_X1 _20507_ (
    .A(_12819_),
    .ZN(_12820_)
  );
  AND2_X1 _20508_ (
    .A1(_08542_),
    .A2(_12820_),
    .ZN(_12821_)
  );
  AND2_X1 _20509_ (
    .A1(_12818_),
    .A2(_12821_),
    .ZN(_12822_)
  );
  INV_X1 _20510_ (
    .A(_12822_),
    .ZN(_12823_)
  );
  AND2_X1 _20511_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_12823_),
    .ZN(_12824_)
  );
  AND2_X1 _20512_ (
    .A1(_12816_),
    .A2(_12824_),
    .ZN(_12825_)
  );
  INV_X1 _20513_ (
    .A(_12825_),
    .ZN(_12826_)
  );
  AND2_X1 _20514_ (
    .A1(\rf[11] [25]),
    .A2(_08541_),
    .ZN(_12827_)
  );
  INV_X1 _20515_ (
    .A(_12827_),
    .ZN(_12828_)
  );
  AND2_X1 _20516_ (
    .A1(\rf[9] [25]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_12829_)
  );
  INV_X1 _20517_ (
    .A(_12829_),
    .ZN(_12830_)
  );
  AND2_X1 _20518_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_12830_),
    .ZN(_12831_)
  );
  AND2_X1 _20519_ (
    .A1(_12828_),
    .A2(_12831_),
    .ZN(_12832_)
  );
  INV_X1 _20520_ (
    .A(_12832_),
    .ZN(_12833_)
  );
  AND2_X1 _20521_ (
    .A1(\rf[15] [25]),
    .A2(_08541_),
    .ZN(_12834_)
  );
  INV_X1 _20522_ (
    .A(_12834_),
    .ZN(_12835_)
  );
  AND2_X1 _20523_ (
    .A1(\rf[13] [25]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_12836_)
  );
  INV_X1 _20524_ (
    .A(_12836_),
    .ZN(_12837_)
  );
  AND2_X1 _20525_ (
    .A1(_08542_),
    .A2(_12837_),
    .ZN(_12838_)
  );
  AND2_X1 _20526_ (
    .A1(_12835_),
    .A2(_12838_),
    .ZN(_12839_)
  );
  INV_X1 _20527_ (
    .A(_12839_),
    .ZN(_12840_)
  );
  AND2_X1 _20528_ (
    .A1(_08540_),
    .A2(_12840_),
    .ZN(_12841_)
  );
  AND2_X1 _20529_ (
    .A1(_12833_),
    .A2(_12841_),
    .ZN(_12842_)
  );
  INV_X1 _20530_ (
    .A(_12842_),
    .ZN(_12843_)
  );
  AND2_X1 _20531_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_12843_),
    .ZN(_12844_)
  );
  AND2_X1 _20532_ (
    .A1(_12826_),
    .A2(_12844_),
    .ZN(_12845_)
  );
  INV_X1 _20533_ (
    .A(_12845_),
    .ZN(_12846_)
  );
  AND2_X1 _20534_ (
    .A1(\rf[30] [25]),
    .A2(_08542_),
    .ZN(_12847_)
  );
  INV_X1 _20535_ (
    .A(_12847_),
    .ZN(_12848_)
  );
  AND2_X1 _20536_ (
    .A1(\rf[26] [25]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12849_)
  );
  INV_X1 _20537_ (
    .A(_12849_),
    .ZN(_12850_)
  );
  AND2_X1 _20538_ (
    .A1(_08541_),
    .A2(_12850_),
    .ZN(_12851_)
  );
  AND2_X1 _20539_ (
    .A1(_12848_),
    .A2(_12851_),
    .ZN(_12852_)
  );
  INV_X1 _20540_ (
    .A(_12852_),
    .ZN(_12853_)
  );
  AND2_X1 _20541_ (
    .A1(\rf[24] [25]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12854_)
  );
  INV_X1 _20542_ (
    .A(_12854_),
    .ZN(_12855_)
  );
  AND2_X1 _20543_ (
    .A1(\rf[28] [25]),
    .A2(_08542_),
    .ZN(_12856_)
  );
  INV_X1 _20544_ (
    .A(_12856_),
    .ZN(_12857_)
  );
  AND2_X1 _20545_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12857_),
    .ZN(_12858_)
  );
  AND2_X1 _20546_ (
    .A1(_12855_),
    .A2(_12858_),
    .ZN(_12859_)
  );
  INV_X1 _20547_ (
    .A(_12859_),
    .ZN(_12860_)
  );
  AND2_X1 _20548_ (
    .A1(_12853_),
    .A2(_12860_),
    .ZN(_12861_)
  );
  MUX2_X1 _20549_ (
    .A(\rf[29] [25]),
    .B(\rf[25] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12862_)
  );
  AND2_X1 _20550_ (
    .A1(\rf[27] [25]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12863_)
  );
  MUX2_X1 _20551_ (
    .A(_12862_),
    .B(_12863_),
    .S(_08541_),
    .Z(_12864_)
  );
  MUX2_X1 _20552_ (
    .A(_12861_),
    .B(_12864_),
    .S(_08540_),
    .Z(_12865_)
  );
  INV_X1 _20553_ (
    .A(_12865_),
    .ZN(_12866_)
  );
  AND2_X1 _20554_ (
    .A1(_08571_),
    .A2(_12866_),
    .ZN(_12867_)
  );
  INV_X1 _20555_ (
    .A(_12867_),
    .ZN(_12868_)
  );
  AND2_X1 _20556_ (
    .A1(_12846_),
    .A2(_12868_),
    .ZN(_12869_)
  );
  MUX2_X1 _20557_ (
    .A(_12809_),
    .B(_12869_),
    .S(_08543_),
    .Z(_12870_)
  );
  MUX2_X1 _20558_ (
    .A(_12870_),
    .B(_12765_),
    .S(_10131_),
    .Z(_12871_)
  );
  AND2_X1 _20559_ (
    .A1(_10082_),
    .A2(_12871_),
    .ZN(_12872_)
  );
  INV_X1 _20560_ (
    .A(_12872_),
    .ZN(_12873_)
  );
  AND2_X1 _20561_ (
    .A1(_12762_),
    .A2(_12873_),
    .ZN(_12874_)
  );
  INV_X1 _20562_ (
    .A(_12874_),
    .ZN(_12875_)
  );
  MUX2_X1 _20563_ (
    .A(ex_reg_rs_msb_0[23]),
    .B(_12875_),
    .S(_10079_),
    .Z(_00090_)
  );
  AND2_X1 _20564_ (
    .A1(_08578_),
    .A2(ibuf_io_inst_0_bits_raw[26]),
    .ZN(_12876_)
  );
  AND2_X1 _20565_ (
    .A1(_09295_),
    .A2(_12876_),
    .ZN(_12877_)
  );
  INV_X1 _20566_ (
    .A(_12877_),
    .ZN(_12878_)
  );
  MUX2_X1 _20567_ (
    .A(\rf[5] [26]),
    .B(\rf[1] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12879_)
  );
  MUX2_X1 _20568_ (
    .A(\rf[7] [26]),
    .B(\rf[3] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12880_)
  );
  MUX2_X1 _20569_ (
    .A(_12879_),
    .B(_12880_),
    .S(_08541_),
    .Z(_12881_)
  );
  AND2_X1 _20570_ (
    .A1(_08540_),
    .A2(_12881_),
    .ZN(_12882_)
  );
  INV_X1 _20571_ (
    .A(_12882_),
    .ZN(_12883_)
  );
  MUX2_X1 _20572_ (
    .A(\rf[4] [26]),
    .B(\rf[0] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12884_)
  );
  MUX2_X1 _20573_ (
    .A(\rf[6] [26]),
    .B(\rf[2] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12885_)
  );
  MUX2_X1 _20574_ (
    .A(_12884_),
    .B(_12885_),
    .S(_08541_),
    .Z(_12886_)
  );
  AND2_X1 _20575_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_12886_),
    .ZN(_12887_)
  );
  INV_X1 _20576_ (
    .A(_12887_),
    .ZN(_12888_)
  );
  AND2_X1 _20577_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_12888_),
    .ZN(_12889_)
  );
  AND2_X1 _20578_ (
    .A1(_12883_),
    .A2(_12889_),
    .ZN(_12890_)
  );
  INV_X1 _20579_ (
    .A(_12890_),
    .ZN(_12891_)
  );
  AND2_X1 _20580_ (
    .A1(_08399_),
    .A2(_08542_),
    .ZN(_12892_)
  );
  INV_X1 _20581_ (
    .A(_12892_),
    .ZN(_12893_)
  );
  AND2_X1 _20582_ (
    .A1(_08300_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12894_)
  );
  INV_X1 _20583_ (
    .A(_12894_),
    .ZN(_12895_)
  );
  AND2_X1 _20584_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12895_),
    .ZN(_12896_)
  );
  AND2_X1 _20585_ (
    .A1(_12893_),
    .A2(_12896_),
    .ZN(_12897_)
  );
  INV_X1 _20586_ (
    .A(_12897_),
    .ZN(_12898_)
  );
  MUX2_X1 _20587_ (
    .A(\rf[22] [26]),
    .B(\rf[18] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12899_)
  );
  AND2_X1 _20588_ (
    .A1(_08541_),
    .A2(_12899_),
    .ZN(_12900_)
  );
  INV_X1 _20589_ (
    .A(_12900_),
    .ZN(_12901_)
  );
  AND2_X1 _20590_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_12901_),
    .ZN(_12902_)
  );
  AND2_X1 _20591_ (
    .A1(_12898_),
    .A2(_12902_),
    .ZN(_12903_)
  );
  INV_X1 _20592_ (
    .A(_12903_),
    .ZN(_12904_)
  );
  AND2_X1 _20593_ (
    .A1(_08330_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12905_)
  );
  INV_X1 _20594_ (
    .A(_12905_),
    .ZN(_12906_)
  );
  AND2_X1 _20595_ (
    .A1(_08429_),
    .A2(_08542_),
    .ZN(_12907_)
  );
  INV_X1 _20596_ (
    .A(_12907_),
    .ZN(_12908_)
  );
  AND2_X1 _20597_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12908_),
    .ZN(_12909_)
  );
  AND2_X1 _20598_ (
    .A1(_12906_),
    .A2(_12909_),
    .ZN(_12910_)
  );
  INV_X1 _20599_ (
    .A(_12910_),
    .ZN(_12911_)
  );
  MUX2_X1 _20600_ (
    .A(\rf[23] [26]),
    .B(\rf[19] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12912_)
  );
  AND2_X1 _20601_ (
    .A1(_08541_),
    .A2(_12912_),
    .ZN(_12913_)
  );
  INV_X1 _20602_ (
    .A(_12913_),
    .ZN(_12914_)
  );
  AND2_X1 _20603_ (
    .A1(_08540_),
    .A2(_12914_),
    .ZN(_12915_)
  );
  AND2_X1 _20604_ (
    .A1(_12911_),
    .A2(_12915_),
    .ZN(_12916_)
  );
  INV_X1 _20605_ (
    .A(_12916_),
    .ZN(_12917_)
  );
  AND2_X1 _20606_ (
    .A1(_12904_),
    .A2(_12917_),
    .ZN(_12918_)
  );
  INV_X1 _20607_ (
    .A(_12918_),
    .ZN(_12919_)
  );
  AND2_X1 _20608_ (
    .A1(_08571_),
    .A2(_12919_),
    .ZN(_12920_)
  );
  INV_X1 _20609_ (
    .A(_12920_),
    .ZN(_12921_)
  );
  AND2_X1 _20610_ (
    .A1(_12891_),
    .A2(_12921_),
    .ZN(_12922_)
  );
  AND2_X1 _20611_ (
    .A1(\rf[10] [26]),
    .A2(_08541_),
    .ZN(_12923_)
  );
  INV_X1 _20612_ (
    .A(_12923_),
    .ZN(_12924_)
  );
  AND2_X1 _20613_ (
    .A1(\rf[8] [26]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_12925_)
  );
  INV_X1 _20614_ (
    .A(_12925_),
    .ZN(_12926_)
  );
  AND2_X1 _20615_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_12926_),
    .ZN(_12927_)
  );
  AND2_X1 _20616_ (
    .A1(_12924_),
    .A2(_12927_),
    .ZN(_12928_)
  );
  INV_X1 _20617_ (
    .A(_12928_),
    .ZN(_12929_)
  );
  AND2_X1 _20618_ (
    .A1(\rf[14] [26]),
    .A2(_08541_),
    .ZN(_12930_)
  );
  INV_X1 _20619_ (
    .A(_12930_),
    .ZN(_12931_)
  );
  AND2_X1 _20620_ (
    .A1(\rf[12] [26]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_12932_)
  );
  INV_X1 _20621_ (
    .A(_12932_),
    .ZN(_12933_)
  );
  AND2_X1 _20622_ (
    .A1(_08542_),
    .A2(_12933_),
    .ZN(_12934_)
  );
  AND2_X1 _20623_ (
    .A1(_12931_),
    .A2(_12934_),
    .ZN(_12935_)
  );
  INV_X1 _20624_ (
    .A(_12935_),
    .ZN(_12936_)
  );
  AND2_X1 _20625_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_12936_),
    .ZN(_12937_)
  );
  AND2_X1 _20626_ (
    .A1(_12929_),
    .A2(_12937_),
    .ZN(_12938_)
  );
  INV_X1 _20627_ (
    .A(_12938_),
    .ZN(_12939_)
  );
  AND2_X1 _20628_ (
    .A1(\rf[11] [26]),
    .A2(_08541_),
    .ZN(_12940_)
  );
  INV_X1 _20629_ (
    .A(_12940_),
    .ZN(_12941_)
  );
  AND2_X1 _20630_ (
    .A1(\rf[9] [26]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_12942_)
  );
  INV_X1 _20631_ (
    .A(_12942_),
    .ZN(_12943_)
  );
  AND2_X1 _20632_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_12943_),
    .ZN(_12944_)
  );
  AND2_X1 _20633_ (
    .A1(_12941_),
    .A2(_12944_),
    .ZN(_12945_)
  );
  INV_X1 _20634_ (
    .A(_12945_),
    .ZN(_12946_)
  );
  AND2_X1 _20635_ (
    .A1(\rf[15] [26]),
    .A2(_08541_),
    .ZN(_12947_)
  );
  INV_X1 _20636_ (
    .A(_12947_),
    .ZN(_12948_)
  );
  AND2_X1 _20637_ (
    .A1(\rf[13] [26]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_12949_)
  );
  INV_X1 _20638_ (
    .A(_12949_),
    .ZN(_12950_)
  );
  AND2_X1 _20639_ (
    .A1(_08542_),
    .A2(_12950_),
    .ZN(_12951_)
  );
  AND2_X1 _20640_ (
    .A1(_12948_),
    .A2(_12951_),
    .ZN(_12952_)
  );
  INV_X1 _20641_ (
    .A(_12952_),
    .ZN(_12953_)
  );
  AND2_X1 _20642_ (
    .A1(_08540_),
    .A2(_12953_),
    .ZN(_12954_)
  );
  AND2_X1 _20643_ (
    .A1(_12946_),
    .A2(_12954_),
    .ZN(_12955_)
  );
  INV_X1 _20644_ (
    .A(_12955_),
    .ZN(_12956_)
  );
  AND2_X1 _20645_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_12956_),
    .ZN(_12957_)
  );
  AND2_X1 _20646_ (
    .A1(_12939_),
    .A2(_12957_),
    .ZN(_12958_)
  );
  INV_X1 _20647_ (
    .A(_12958_),
    .ZN(_12959_)
  );
  AND2_X1 _20648_ (
    .A1(\rf[30] [26]),
    .A2(_08542_),
    .ZN(_12960_)
  );
  INV_X1 _20649_ (
    .A(_12960_),
    .ZN(_12961_)
  );
  AND2_X1 _20650_ (
    .A1(\rf[26] [26]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12962_)
  );
  INV_X1 _20651_ (
    .A(_12962_),
    .ZN(_12963_)
  );
  AND2_X1 _20652_ (
    .A1(_08541_),
    .A2(_12963_),
    .ZN(_12964_)
  );
  AND2_X1 _20653_ (
    .A1(_12961_),
    .A2(_12964_),
    .ZN(_12965_)
  );
  INV_X1 _20654_ (
    .A(_12965_),
    .ZN(_12966_)
  );
  AND2_X1 _20655_ (
    .A1(\rf[24] [26]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12967_)
  );
  INV_X1 _20656_ (
    .A(_12967_),
    .ZN(_12968_)
  );
  AND2_X1 _20657_ (
    .A1(\rf[28] [26]),
    .A2(_08542_),
    .ZN(_12969_)
  );
  INV_X1 _20658_ (
    .A(_12969_),
    .ZN(_12970_)
  );
  AND2_X1 _20659_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_12970_),
    .ZN(_12971_)
  );
  AND2_X1 _20660_ (
    .A1(_12968_),
    .A2(_12971_),
    .ZN(_12972_)
  );
  INV_X1 _20661_ (
    .A(_12972_),
    .ZN(_12973_)
  );
  AND2_X1 _20662_ (
    .A1(_12966_),
    .A2(_12973_),
    .ZN(_12974_)
  );
  MUX2_X1 _20663_ (
    .A(\rf[29] [26]),
    .B(\rf[25] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12975_)
  );
  AND2_X1 _20664_ (
    .A1(\rf[27] [26]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_12976_)
  );
  MUX2_X1 _20665_ (
    .A(_12975_),
    .B(_12976_),
    .S(_08541_),
    .Z(_12977_)
  );
  MUX2_X1 _20666_ (
    .A(_12974_),
    .B(_12977_),
    .S(_08540_),
    .Z(_12978_)
  );
  INV_X1 _20667_ (
    .A(_12978_),
    .ZN(_12979_)
  );
  AND2_X1 _20668_ (
    .A1(_08571_),
    .A2(_12979_),
    .ZN(_12980_)
  );
  INV_X1 _20669_ (
    .A(_12980_),
    .ZN(_12981_)
  );
  AND2_X1 _20670_ (
    .A1(_12959_),
    .A2(_12981_),
    .ZN(_12982_)
  );
  MUX2_X1 _20671_ (
    .A(_12922_),
    .B(_12982_),
    .S(_08543_),
    .Z(_12983_)
  );
  MUX2_X1 _20672_ (
    .A(csr_io_rw_rdata[26]),
    .B(wb_reg_wdata[26]),
    .S(_10134_),
    .Z(_12984_)
  );
  MUX2_X1 _20673_ (
    .A(div_io_resp_bits_data[26]),
    .B(_12984_),
    .S(_08649_),
    .Z(_12985_)
  );
  MUX2_X1 _20674_ (
    .A(_12985_),
    .B(io_dmem_resp_bits_data[26]),
    .S(_08631_),
    .Z(_12986_)
  );
  MUX2_X1 _20675_ (
    .A(_12983_),
    .B(_12986_),
    .S(_10131_),
    .Z(_12987_)
  );
  AND2_X1 _20676_ (
    .A1(_10082_),
    .A2(_12987_),
    .ZN(_12988_)
  );
  INV_X1 _20677_ (
    .A(_12988_),
    .ZN(_12989_)
  );
  AND2_X1 _20678_ (
    .A1(_12878_),
    .A2(_12989_),
    .ZN(_12990_)
  );
  INV_X1 _20679_ (
    .A(_12990_),
    .ZN(_12991_)
  );
  MUX2_X1 _20680_ (
    .A(ex_reg_rs_msb_0[24]),
    .B(_12991_),
    .S(_10079_),
    .Z(_00091_)
  );
  AND2_X1 _20681_ (
    .A1(_08578_),
    .A2(ibuf_io_inst_0_bits_raw[27]),
    .ZN(_12992_)
  );
  AND2_X1 _20682_ (
    .A1(_09295_),
    .A2(_12992_),
    .ZN(_12993_)
  );
  INV_X1 _20683_ (
    .A(_12993_),
    .ZN(_12994_)
  );
  MUX2_X1 _20684_ (
    .A(\rf[5] [27]),
    .B(\rf[1] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12995_)
  );
  MUX2_X1 _20685_ (
    .A(\rf[7] [27]),
    .B(\rf[3] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_12996_)
  );
  MUX2_X1 _20686_ (
    .A(_12995_),
    .B(_12996_),
    .S(_08541_),
    .Z(_12997_)
  );
  AND2_X1 _20687_ (
    .A1(_08540_),
    .A2(_12997_),
    .ZN(_12998_)
  );
  INV_X1 _20688_ (
    .A(_12998_),
    .ZN(_12999_)
  );
  MUX2_X1 _20689_ (
    .A(\rf[4] [27]),
    .B(\rf[0] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13000_)
  );
  MUX2_X1 _20690_ (
    .A(\rf[6] [27]),
    .B(\rf[2] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13001_)
  );
  MUX2_X1 _20691_ (
    .A(_13000_),
    .B(_13001_),
    .S(_08541_),
    .Z(_13002_)
  );
  AND2_X1 _20692_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13002_),
    .ZN(_13003_)
  );
  INV_X1 _20693_ (
    .A(_13003_),
    .ZN(_13004_)
  );
  AND2_X1 _20694_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_13004_),
    .ZN(_13005_)
  );
  AND2_X1 _20695_ (
    .A1(_12999_),
    .A2(_13005_),
    .ZN(_13006_)
  );
  INV_X1 _20696_ (
    .A(_13006_),
    .ZN(_13007_)
  );
  AND2_X1 _20697_ (
    .A1(_08400_),
    .A2(_08542_),
    .ZN(_13008_)
  );
  INV_X1 _20698_ (
    .A(_13008_),
    .ZN(_13009_)
  );
  AND2_X1 _20699_ (
    .A1(_08301_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13010_)
  );
  INV_X1 _20700_ (
    .A(_13010_),
    .ZN(_13011_)
  );
  AND2_X1 _20701_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_13011_),
    .ZN(_13012_)
  );
  AND2_X1 _20702_ (
    .A1(_13009_),
    .A2(_13012_),
    .ZN(_13013_)
  );
  INV_X1 _20703_ (
    .A(_13013_),
    .ZN(_13014_)
  );
  MUX2_X1 _20704_ (
    .A(\rf[22] [27]),
    .B(\rf[18] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13015_)
  );
  AND2_X1 _20705_ (
    .A1(_08541_),
    .A2(_13015_),
    .ZN(_13016_)
  );
  INV_X1 _20706_ (
    .A(_13016_),
    .ZN(_13017_)
  );
  AND2_X1 _20707_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13017_),
    .ZN(_13018_)
  );
  AND2_X1 _20708_ (
    .A1(_13014_),
    .A2(_13018_),
    .ZN(_13019_)
  );
  INV_X1 _20709_ (
    .A(_13019_),
    .ZN(_13020_)
  );
  AND2_X1 _20710_ (
    .A1(_08331_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13021_)
  );
  INV_X1 _20711_ (
    .A(_13021_),
    .ZN(_13022_)
  );
  AND2_X1 _20712_ (
    .A1(_08430_),
    .A2(_08542_),
    .ZN(_13023_)
  );
  INV_X1 _20713_ (
    .A(_13023_),
    .ZN(_13024_)
  );
  AND2_X1 _20714_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_13024_),
    .ZN(_13025_)
  );
  AND2_X1 _20715_ (
    .A1(_13022_),
    .A2(_13025_),
    .ZN(_13026_)
  );
  INV_X1 _20716_ (
    .A(_13026_),
    .ZN(_13027_)
  );
  MUX2_X1 _20717_ (
    .A(\rf[23] [27]),
    .B(\rf[19] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13028_)
  );
  AND2_X1 _20718_ (
    .A1(_08541_),
    .A2(_13028_),
    .ZN(_13029_)
  );
  INV_X1 _20719_ (
    .A(_13029_),
    .ZN(_13030_)
  );
  AND2_X1 _20720_ (
    .A1(_08540_),
    .A2(_13030_),
    .ZN(_13031_)
  );
  AND2_X1 _20721_ (
    .A1(_13027_),
    .A2(_13031_),
    .ZN(_13032_)
  );
  INV_X1 _20722_ (
    .A(_13032_),
    .ZN(_13033_)
  );
  AND2_X1 _20723_ (
    .A1(_13020_),
    .A2(_13033_),
    .ZN(_13034_)
  );
  INV_X1 _20724_ (
    .A(_13034_),
    .ZN(_13035_)
  );
  AND2_X1 _20725_ (
    .A1(_08571_),
    .A2(_13035_),
    .ZN(_13036_)
  );
  INV_X1 _20726_ (
    .A(_13036_),
    .ZN(_13037_)
  );
  AND2_X1 _20727_ (
    .A1(_13007_),
    .A2(_13037_),
    .ZN(_13038_)
  );
  AND2_X1 _20728_ (
    .A1(\rf[10] [27]),
    .A2(_08541_),
    .ZN(_13039_)
  );
  INV_X1 _20729_ (
    .A(_13039_),
    .ZN(_13040_)
  );
  AND2_X1 _20730_ (
    .A1(\rf[8] [27]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_13041_)
  );
  INV_X1 _20731_ (
    .A(_13041_),
    .ZN(_13042_)
  );
  AND2_X1 _20732_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_13042_),
    .ZN(_13043_)
  );
  AND2_X1 _20733_ (
    .A1(_13040_),
    .A2(_13043_),
    .ZN(_13044_)
  );
  INV_X1 _20734_ (
    .A(_13044_),
    .ZN(_13045_)
  );
  AND2_X1 _20735_ (
    .A1(\rf[14] [27]),
    .A2(_08541_),
    .ZN(_13046_)
  );
  INV_X1 _20736_ (
    .A(_13046_),
    .ZN(_13047_)
  );
  AND2_X1 _20737_ (
    .A1(\rf[12] [27]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_13048_)
  );
  INV_X1 _20738_ (
    .A(_13048_),
    .ZN(_13049_)
  );
  AND2_X1 _20739_ (
    .A1(_08542_),
    .A2(_13049_),
    .ZN(_13050_)
  );
  AND2_X1 _20740_ (
    .A1(_13047_),
    .A2(_13050_),
    .ZN(_13051_)
  );
  INV_X1 _20741_ (
    .A(_13051_),
    .ZN(_13052_)
  );
  AND2_X1 _20742_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13052_),
    .ZN(_13053_)
  );
  AND2_X1 _20743_ (
    .A1(_13045_),
    .A2(_13053_),
    .ZN(_13054_)
  );
  INV_X1 _20744_ (
    .A(_13054_),
    .ZN(_13055_)
  );
  AND2_X1 _20745_ (
    .A1(\rf[11] [27]),
    .A2(_08541_),
    .ZN(_13056_)
  );
  INV_X1 _20746_ (
    .A(_13056_),
    .ZN(_13057_)
  );
  AND2_X1 _20747_ (
    .A1(\rf[9] [27]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_13058_)
  );
  INV_X1 _20748_ (
    .A(_13058_),
    .ZN(_13059_)
  );
  AND2_X1 _20749_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_13059_),
    .ZN(_13060_)
  );
  AND2_X1 _20750_ (
    .A1(_13057_),
    .A2(_13060_),
    .ZN(_13061_)
  );
  INV_X1 _20751_ (
    .A(_13061_),
    .ZN(_13062_)
  );
  AND2_X1 _20752_ (
    .A1(\rf[15] [27]),
    .A2(_08541_),
    .ZN(_13063_)
  );
  INV_X1 _20753_ (
    .A(_13063_),
    .ZN(_13064_)
  );
  AND2_X1 _20754_ (
    .A1(\rf[13] [27]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_13065_)
  );
  INV_X1 _20755_ (
    .A(_13065_),
    .ZN(_13066_)
  );
  AND2_X1 _20756_ (
    .A1(_08542_),
    .A2(_13066_),
    .ZN(_13067_)
  );
  AND2_X1 _20757_ (
    .A1(_13064_),
    .A2(_13067_),
    .ZN(_13068_)
  );
  INV_X1 _20758_ (
    .A(_13068_),
    .ZN(_13069_)
  );
  AND2_X1 _20759_ (
    .A1(_08540_),
    .A2(_13069_),
    .ZN(_13070_)
  );
  AND2_X1 _20760_ (
    .A1(_13062_),
    .A2(_13070_),
    .ZN(_13071_)
  );
  INV_X1 _20761_ (
    .A(_13071_),
    .ZN(_13072_)
  );
  AND2_X1 _20762_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_13072_),
    .ZN(_13073_)
  );
  AND2_X1 _20763_ (
    .A1(_13055_),
    .A2(_13073_),
    .ZN(_13074_)
  );
  INV_X1 _20764_ (
    .A(_13074_),
    .ZN(_13075_)
  );
  AND2_X1 _20765_ (
    .A1(\rf[30] [27]),
    .A2(_08542_),
    .ZN(_13076_)
  );
  INV_X1 _20766_ (
    .A(_13076_),
    .ZN(_13077_)
  );
  AND2_X1 _20767_ (
    .A1(\rf[26] [27]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13078_)
  );
  INV_X1 _20768_ (
    .A(_13078_),
    .ZN(_13079_)
  );
  AND2_X1 _20769_ (
    .A1(_08541_),
    .A2(_13079_),
    .ZN(_13080_)
  );
  AND2_X1 _20770_ (
    .A1(_13077_),
    .A2(_13080_),
    .ZN(_13081_)
  );
  INV_X1 _20771_ (
    .A(_13081_),
    .ZN(_13082_)
  );
  AND2_X1 _20772_ (
    .A1(\rf[24] [27]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13083_)
  );
  INV_X1 _20773_ (
    .A(_13083_),
    .ZN(_13084_)
  );
  AND2_X1 _20774_ (
    .A1(\rf[28] [27]),
    .A2(_08542_),
    .ZN(_13085_)
  );
  INV_X1 _20775_ (
    .A(_13085_),
    .ZN(_13086_)
  );
  AND2_X1 _20776_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_13086_),
    .ZN(_13087_)
  );
  AND2_X1 _20777_ (
    .A1(_13084_),
    .A2(_13087_),
    .ZN(_13088_)
  );
  INV_X1 _20778_ (
    .A(_13088_),
    .ZN(_13089_)
  );
  AND2_X1 _20779_ (
    .A1(_13082_),
    .A2(_13089_),
    .ZN(_13090_)
  );
  MUX2_X1 _20780_ (
    .A(\rf[29] [27]),
    .B(\rf[25] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13091_)
  );
  AND2_X1 _20781_ (
    .A1(\rf[27] [27]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13092_)
  );
  MUX2_X1 _20782_ (
    .A(_13091_),
    .B(_13092_),
    .S(_08541_),
    .Z(_13093_)
  );
  MUX2_X1 _20783_ (
    .A(_13090_),
    .B(_13093_),
    .S(_08540_),
    .Z(_13094_)
  );
  INV_X1 _20784_ (
    .A(_13094_),
    .ZN(_13095_)
  );
  AND2_X1 _20785_ (
    .A1(_08571_),
    .A2(_13095_),
    .ZN(_13096_)
  );
  INV_X1 _20786_ (
    .A(_13096_),
    .ZN(_13097_)
  );
  AND2_X1 _20787_ (
    .A1(_13075_),
    .A2(_13097_),
    .ZN(_13098_)
  );
  MUX2_X1 _20788_ (
    .A(_13038_),
    .B(_13098_),
    .S(_08543_),
    .Z(_13099_)
  );
  MUX2_X1 _20789_ (
    .A(csr_io_rw_rdata[27]),
    .B(wb_reg_wdata[27]),
    .S(_10134_),
    .Z(_13100_)
  );
  MUX2_X1 _20790_ (
    .A(div_io_resp_bits_data[27]),
    .B(_13100_),
    .S(_08649_),
    .Z(_13101_)
  );
  MUX2_X1 _20791_ (
    .A(_13101_),
    .B(io_dmem_resp_bits_data[27]),
    .S(_08631_),
    .Z(_13102_)
  );
  MUX2_X1 _20792_ (
    .A(_13099_),
    .B(_13102_),
    .S(_10131_),
    .Z(_13103_)
  );
  AND2_X1 _20793_ (
    .A1(_10082_),
    .A2(_13103_),
    .ZN(_13104_)
  );
  INV_X1 _20794_ (
    .A(_13104_),
    .ZN(_13105_)
  );
  AND2_X1 _20795_ (
    .A1(_12994_),
    .A2(_13105_),
    .ZN(_13106_)
  );
  INV_X1 _20796_ (
    .A(_13106_),
    .ZN(_13107_)
  );
  MUX2_X1 _20797_ (
    .A(ex_reg_rs_msb_0[25]),
    .B(_13107_),
    .S(_10079_),
    .Z(_00092_)
  );
  AND2_X1 _20798_ (
    .A1(_08578_),
    .A2(ibuf_io_inst_0_bits_raw[28]),
    .ZN(_13108_)
  );
  AND2_X1 _20799_ (
    .A1(_09295_),
    .A2(_13108_),
    .ZN(_13109_)
  );
  INV_X1 _20800_ (
    .A(_13109_),
    .ZN(_13110_)
  );
  MUX2_X1 _20801_ (
    .A(\rf[5] [28]),
    .B(\rf[1] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13111_)
  );
  MUX2_X1 _20802_ (
    .A(\rf[7] [28]),
    .B(\rf[3] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13112_)
  );
  MUX2_X1 _20803_ (
    .A(_13111_),
    .B(_13112_),
    .S(_08541_),
    .Z(_13113_)
  );
  AND2_X1 _20804_ (
    .A1(_08540_),
    .A2(_13113_),
    .ZN(_13114_)
  );
  INV_X1 _20805_ (
    .A(_13114_),
    .ZN(_13115_)
  );
  MUX2_X1 _20806_ (
    .A(\rf[4] [28]),
    .B(\rf[0] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13116_)
  );
  MUX2_X1 _20807_ (
    .A(\rf[6] [28]),
    .B(\rf[2] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13117_)
  );
  MUX2_X1 _20808_ (
    .A(_13116_),
    .B(_13117_),
    .S(_08541_),
    .Z(_13118_)
  );
  AND2_X1 _20809_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13118_),
    .ZN(_13119_)
  );
  INV_X1 _20810_ (
    .A(_13119_),
    .ZN(_13120_)
  );
  AND2_X1 _20811_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_13120_),
    .ZN(_13121_)
  );
  AND2_X1 _20812_ (
    .A1(_13115_),
    .A2(_13121_),
    .ZN(_13122_)
  );
  INV_X1 _20813_ (
    .A(_13122_),
    .ZN(_13123_)
  );
  AND2_X1 _20814_ (
    .A1(_08401_),
    .A2(_08542_),
    .ZN(_13124_)
  );
  INV_X1 _20815_ (
    .A(_13124_),
    .ZN(_13125_)
  );
  AND2_X1 _20816_ (
    .A1(_08302_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13126_)
  );
  INV_X1 _20817_ (
    .A(_13126_),
    .ZN(_13127_)
  );
  AND2_X1 _20818_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_13127_),
    .ZN(_13128_)
  );
  AND2_X1 _20819_ (
    .A1(_13125_),
    .A2(_13128_),
    .ZN(_13129_)
  );
  INV_X1 _20820_ (
    .A(_13129_),
    .ZN(_13130_)
  );
  MUX2_X1 _20821_ (
    .A(\rf[22] [28]),
    .B(\rf[18] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13131_)
  );
  AND2_X1 _20822_ (
    .A1(_08541_),
    .A2(_13131_),
    .ZN(_13132_)
  );
  INV_X1 _20823_ (
    .A(_13132_),
    .ZN(_13133_)
  );
  AND2_X1 _20824_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13133_),
    .ZN(_13134_)
  );
  AND2_X1 _20825_ (
    .A1(_13130_),
    .A2(_13134_),
    .ZN(_13135_)
  );
  INV_X1 _20826_ (
    .A(_13135_),
    .ZN(_13136_)
  );
  AND2_X1 _20827_ (
    .A1(_08332_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13137_)
  );
  INV_X1 _20828_ (
    .A(_13137_),
    .ZN(_13138_)
  );
  AND2_X1 _20829_ (
    .A1(_08431_),
    .A2(_08542_),
    .ZN(_13139_)
  );
  INV_X1 _20830_ (
    .A(_13139_),
    .ZN(_13140_)
  );
  AND2_X1 _20831_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_13140_),
    .ZN(_13141_)
  );
  AND2_X1 _20832_ (
    .A1(_13138_),
    .A2(_13141_),
    .ZN(_13142_)
  );
  INV_X1 _20833_ (
    .A(_13142_),
    .ZN(_13143_)
  );
  MUX2_X1 _20834_ (
    .A(\rf[23] [28]),
    .B(\rf[19] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13144_)
  );
  AND2_X1 _20835_ (
    .A1(_08541_),
    .A2(_13144_),
    .ZN(_13145_)
  );
  INV_X1 _20836_ (
    .A(_13145_),
    .ZN(_13146_)
  );
  AND2_X1 _20837_ (
    .A1(_08540_),
    .A2(_13146_),
    .ZN(_13147_)
  );
  AND2_X1 _20838_ (
    .A1(_13143_),
    .A2(_13147_),
    .ZN(_13148_)
  );
  INV_X1 _20839_ (
    .A(_13148_),
    .ZN(_13149_)
  );
  AND2_X1 _20840_ (
    .A1(_13136_),
    .A2(_13149_),
    .ZN(_13150_)
  );
  INV_X1 _20841_ (
    .A(_13150_),
    .ZN(_13151_)
  );
  AND2_X1 _20842_ (
    .A1(_08571_),
    .A2(_13151_),
    .ZN(_13152_)
  );
  INV_X1 _20843_ (
    .A(_13152_),
    .ZN(_13153_)
  );
  AND2_X1 _20844_ (
    .A1(_13123_),
    .A2(_13153_),
    .ZN(_13154_)
  );
  AND2_X1 _20845_ (
    .A1(\rf[10] [28]),
    .A2(_08541_),
    .ZN(_13155_)
  );
  INV_X1 _20846_ (
    .A(_13155_),
    .ZN(_13156_)
  );
  AND2_X1 _20847_ (
    .A1(\rf[8] [28]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_13157_)
  );
  INV_X1 _20848_ (
    .A(_13157_),
    .ZN(_13158_)
  );
  AND2_X1 _20849_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_13158_),
    .ZN(_13159_)
  );
  AND2_X1 _20850_ (
    .A1(_13156_),
    .A2(_13159_),
    .ZN(_13160_)
  );
  INV_X1 _20851_ (
    .A(_13160_),
    .ZN(_13161_)
  );
  AND2_X1 _20852_ (
    .A1(\rf[14] [28]),
    .A2(_08541_),
    .ZN(_13162_)
  );
  INV_X1 _20853_ (
    .A(_13162_),
    .ZN(_13163_)
  );
  AND2_X1 _20854_ (
    .A1(\rf[12] [28]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_13164_)
  );
  INV_X1 _20855_ (
    .A(_13164_),
    .ZN(_13165_)
  );
  AND2_X1 _20856_ (
    .A1(_08542_),
    .A2(_13165_),
    .ZN(_13166_)
  );
  AND2_X1 _20857_ (
    .A1(_13163_),
    .A2(_13166_),
    .ZN(_13167_)
  );
  INV_X1 _20858_ (
    .A(_13167_),
    .ZN(_13168_)
  );
  AND2_X1 _20859_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13168_),
    .ZN(_13169_)
  );
  AND2_X1 _20860_ (
    .A1(_13161_),
    .A2(_13169_),
    .ZN(_13170_)
  );
  INV_X1 _20861_ (
    .A(_13170_),
    .ZN(_13171_)
  );
  AND2_X1 _20862_ (
    .A1(\rf[11] [28]),
    .A2(_08541_),
    .ZN(_13172_)
  );
  INV_X1 _20863_ (
    .A(_13172_),
    .ZN(_13173_)
  );
  AND2_X1 _20864_ (
    .A1(\rf[9] [28]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_13174_)
  );
  INV_X1 _20865_ (
    .A(_13174_),
    .ZN(_13175_)
  );
  AND2_X1 _20866_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_13175_),
    .ZN(_13176_)
  );
  AND2_X1 _20867_ (
    .A1(_13173_),
    .A2(_13176_),
    .ZN(_13177_)
  );
  INV_X1 _20868_ (
    .A(_13177_),
    .ZN(_13178_)
  );
  AND2_X1 _20869_ (
    .A1(\rf[15] [28]),
    .A2(_08541_),
    .ZN(_13179_)
  );
  INV_X1 _20870_ (
    .A(_13179_),
    .ZN(_13180_)
  );
  AND2_X1 _20871_ (
    .A1(\rf[13] [28]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_13181_)
  );
  INV_X1 _20872_ (
    .A(_13181_),
    .ZN(_13182_)
  );
  AND2_X1 _20873_ (
    .A1(_08542_),
    .A2(_13182_),
    .ZN(_13183_)
  );
  AND2_X1 _20874_ (
    .A1(_13180_),
    .A2(_13183_),
    .ZN(_13184_)
  );
  INV_X1 _20875_ (
    .A(_13184_),
    .ZN(_13185_)
  );
  AND2_X1 _20876_ (
    .A1(_08540_),
    .A2(_13185_),
    .ZN(_13186_)
  );
  AND2_X1 _20877_ (
    .A1(_13178_),
    .A2(_13186_),
    .ZN(_13187_)
  );
  INV_X1 _20878_ (
    .A(_13187_),
    .ZN(_13188_)
  );
  AND2_X1 _20879_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_13188_),
    .ZN(_13189_)
  );
  AND2_X1 _20880_ (
    .A1(_13171_),
    .A2(_13189_),
    .ZN(_13190_)
  );
  INV_X1 _20881_ (
    .A(_13190_),
    .ZN(_13191_)
  );
  AND2_X1 _20882_ (
    .A1(\rf[30] [28]),
    .A2(_08542_),
    .ZN(_13192_)
  );
  INV_X1 _20883_ (
    .A(_13192_),
    .ZN(_13193_)
  );
  AND2_X1 _20884_ (
    .A1(\rf[26] [28]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13194_)
  );
  INV_X1 _20885_ (
    .A(_13194_),
    .ZN(_13195_)
  );
  AND2_X1 _20886_ (
    .A1(_08541_),
    .A2(_13195_),
    .ZN(_13196_)
  );
  AND2_X1 _20887_ (
    .A1(_13193_),
    .A2(_13196_),
    .ZN(_13197_)
  );
  INV_X1 _20888_ (
    .A(_13197_),
    .ZN(_13198_)
  );
  AND2_X1 _20889_ (
    .A1(\rf[24] [28]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13199_)
  );
  INV_X1 _20890_ (
    .A(_13199_),
    .ZN(_13200_)
  );
  AND2_X1 _20891_ (
    .A1(\rf[28] [28]),
    .A2(_08542_),
    .ZN(_13201_)
  );
  INV_X1 _20892_ (
    .A(_13201_),
    .ZN(_13202_)
  );
  AND2_X1 _20893_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_13202_),
    .ZN(_13203_)
  );
  AND2_X1 _20894_ (
    .A1(_13200_),
    .A2(_13203_),
    .ZN(_13204_)
  );
  INV_X1 _20895_ (
    .A(_13204_),
    .ZN(_13205_)
  );
  AND2_X1 _20896_ (
    .A1(_13198_),
    .A2(_13205_),
    .ZN(_13206_)
  );
  MUX2_X1 _20897_ (
    .A(\rf[29] [28]),
    .B(\rf[25] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13207_)
  );
  AND2_X1 _20898_ (
    .A1(\rf[27] [28]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13208_)
  );
  MUX2_X1 _20899_ (
    .A(_13207_),
    .B(_13208_),
    .S(_08541_),
    .Z(_13209_)
  );
  MUX2_X1 _20900_ (
    .A(_13206_),
    .B(_13209_),
    .S(_08540_),
    .Z(_13210_)
  );
  INV_X1 _20901_ (
    .A(_13210_),
    .ZN(_13211_)
  );
  AND2_X1 _20902_ (
    .A1(_08571_),
    .A2(_13211_),
    .ZN(_13212_)
  );
  INV_X1 _20903_ (
    .A(_13212_),
    .ZN(_13213_)
  );
  AND2_X1 _20904_ (
    .A1(_13191_),
    .A2(_13213_),
    .ZN(_13214_)
  );
  MUX2_X1 _20905_ (
    .A(_13154_),
    .B(_13214_),
    .S(_08543_),
    .Z(_13215_)
  );
  MUX2_X1 _20906_ (
    .A(csr_io_rw_rdata[28]),
    .B(wb_reg_wdata[28]),
    .S(_10134_),
    .Z(_13216_)
  );
  MUX2_X1 _20907_ (
    .A(div_io_resp_bits_data[28]),
    .B(_13216_),
    .S(_08649_),
    .Z(_13217_)
  );
  MUX2_X1 _20908_ (
    .A(_13217_),
    .B(io_dmem_resp_bits_data[28]),
    .S(_08631_),
    .Z(_13218_)
  );
  MUX2_X1 _20909_ (
    .A(_13215_),
    .B(_13218_),
    .S(_10131_),
    .Z(_13219_)
  );
  AND2_X1 _20910_ (
    .A1(_10082_),
    .A2(_13219_),
    .ZN(_13220_)
  );
  INV_X1 _20911_ (
    .A(_13220_),
    .ZN(_13221_)
  );
  AND2_X1 _20912_ (
    .A1(_13110_),
    .A2(_13221_),
    .ZN(_13222_)
  );
  INV_X1 _20913_ (
    .A(_13222_),
    .ZN(_13223_)
  );
  MUX2_X1 _20914_ (
    .A(ex_reg_rs_msb_0[26]),
    .B(_13223_),
    .S(_10079_),
    .Z(_00093_)
  );
  AND2_X1 _20915_ (
    .A1(_08578_),
    .A2(ibuf_io_inst_0_bits_raw[29]),
    .ZN(_13224_)
  );
  AND2_X1 _20916_ (
    .A1(_09295_),
    .A2(_13224_),
    .ZN(_13225_)
  );
  INV_X1 _20917_ (
    .A(_13225_),
    .ZN(_13226_)
  );
  AND2_X1 _20918_ (
    .A1(_08350_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13227_)
  );
  INV_X1 _20919_ (
    .A(_13227_),
    .ZN(_13228_)
  );
  AND2_X1 _20920_ (
    .A1(_08488_),
    .A2(_08542_),
    .ZN(_13229_)
  );
  INV_X1 _20921_ (
    .A(_13229_),
    .ZN(_13230_)
  );
  AND2_X1 _20922_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13230_),
    .ZN(_13231_)
  );
  AND2_X1 _20923_ (
    .A1(_13228_),
    .A2(_13231_),
    .ZN(_13232_)
  );
  INV_X1 _20924_ (
    .A(_13232_),
    .ZN(_13233_)
  );
  MUX2_X1 _20925_ (
    .A(\rf[15] [29]),
    .B(\rf[11] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13234_)
  );
  AND2_X1 _20926_ (
    .A1(_08540_),
    .A2(_13234_),
    .ZN(_13235_)
  );
  INV_X1 _20927_ (
    .A(_13235_),
    .ZN(_13236_)
  );
  AND2_X1 _20928_ (
    .A1(_08541_),
    .A2(_13236_),
    .ZN(_13237_)
  );
  AND2_X1 _20929_ (
    .A1(_13233_),
    .A2(_13237_),
    .ZN(_13238_)
  );
  INV_X1 _20930_ (
    .A(_13238_),
    .ZN(_13239_)
  );
  AND2_X1 _20931_ (
    .A1(_08371_),
    .A2(_08542_),
    .ZN(_13240_)
  );
  INV_X1 _20932_ (
    .A(_13240_),
    .ZN(_13241_)
  );
  AND2_X1 _20933_ (
    .A1(_08272_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13242_)
  );
  INV_X1 _20934_ (
    .A(_13242_),
    .ZN(_13243_)
  );
  AND2_X1 _20935_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13243_),
    .ZN(_13244_)
  );
  AND2_X1 _20936_ (
    .A1(_13241_),
    .A2(_13244_),
    .ZN(_13245_)
  );
  INV_X1 _20937_ (
    .A(_13245_),
    .ZN(_13246_)
  );
  MUX2_X1 _20938_ (
    .A(\rf[13] [29]),
    .B(\rf[9] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13247_)
  );
  AND2_X1 _20939_ (
    .A1(_08540_),
    .A2(_13247_),
    .ZN(_13248_)
  );
  INV_X1 _20940_ (
    .A(_13248_),
    .ZN(_13249_)
  );
  AND2_X1 _20941_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_13249_),
    .ZN(_13250_)
  );
  AND2_X1 _20942_ (
    .A1(_13246_),
    .A2(_13250_),
    .ZN(_13251_)
  );
  INV_X1 _20943_ (
    .A(_13251_),
    .ZN(_13252_)
  );
  AND2_X1 _20944_ (
    .A1(_08543_),
    .A2(_13252_),
    .ZN(_13253_)
  );
  AND2_X1 _20945_ (
    .A1(_13239_),
    .A2(_13253_),
    .ZN(_13254_)
  );
  INV_X1 _20946_ (
    .A(_13254_),
    .ZN(_13255_)
  );
  AND2_X1 _20947_ (
    .A1(_08256_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13256_)
  );
  INV_X1 _20948_ (
    .A(_13256_),
    .ZN(_13257_)
  );
  AND2_X1 _20949_ (
    .A1(_08252_),
    .A2(_08542_),
    .ZN(_13258_)
  );
  INV_X1 _20950_ (
    .A(_13258_),
    .ZN(_13259_)
  );
  AND2_X1 _20951_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13259_),
    .ZN(_13260_)
  );
  AND2_X1 _20952_ (
    .A1(_13257_),
    .A2(_13260_),
    .ZN(_13261_)
  );
  INV_X1 _20953_ (
    .A(_13261_),
    .ZN(_13262_)
  );
  MUX2_X1 _20954_ (
    .A(\rf[5] [29]),
    .B(\rf[1] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13263_)
  );
  AND2_X1 _20955_ (
    .A1(_08540_),
    .A2(_13263_),
    .ZN(_13264_)
  );
  INV_X1 _20956_ (
    .A(_13264_),
    .ZN(_13265_)
  );
  AND2_X1 _20957_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_13265_),
    .ZN(_13266_)
  );
  AND2_X1 _20958_ (
    .A1(_13262_),
    .A2(_13266_),
    .ZN(_13267_)
  );
  INV_X1 _20959_ (
    .A(_13267_),
    .ZN(_13268_)
  );
  MUX2_X1 _20960_ (
    .A(\rf[7] [29]),
    .B(\rf[3] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13269_)
  );
  AND2_X1 _20961_ (
    .A1(_08540_),
    .A2(_13269_),
    .ZN(_13270_)
  );
  INV_X1 _20962_ (
    .A(_13270_),
    .ZN(_13271_)
  );
  AND2_X1 _20963_ (
    .A1(_08503_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13272_)
  );
  INV_X1 _20964_ (
    .A(_13272_),
    .ZN(_13273_)
  );
  AND2_X1 _20965_ (
    .A1(_08247_),
    .A2(_08542_),
    .ZN(_13274_)
  );
  INV_X1 _20966_ (
    .A(_13274_),
    .ZN(_13275_)
  );
  AND2_X1 _20967_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13275_),
    .ZN(_13276_)
  );
  AND2_X1 _20968_ (
    .A1(_13273_),
    .A2(_13276_),
    .ZN(_13277_)
  );
  INV_X1 _20969_ (
    .A(_13277_),
    .ZN(_13278_)
  );
  AND2_X1 _20970_ (
    .A1(_13271_),
    .A2(_13278_),
    .ZN(_13279_)
  );
  AND2_X1 _20971_ (
    .A1(_08541_),
    .A2(_13279_),
    .ZN(_13280_)
  );
  INV_X1 _20972_ (
    .A(_13280_),
    .ZN(_13281_)
  );
  AND2_X1 _20973_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_13268_),
    .ZN(_13282_)
  );
  AND2_X1 _20974_ (
    .A1(_13281_),
    .A2(_13282_),
    .ZN(_13283_)
  );
  INV_X1 _20975_ (
    .A(_13283_),
    .ZN(_13284_)
  );
  AND2_X1 _20976_ (
    .A1(_13255_),
    .A2(_13284_),
    .ZN(_13285_)
  );
  MUX2_X1 _20977_ (
    .A(\rf[30] [29]),
    .B(\rf[26] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13286_)
  );
  AND2_X1 _20978_ (
    .A1(\rf[27] [29]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13287_)
  );
  MUX2_X1 _20979_ (
    .A(_13286_),
    .B(_13287_),
    .S(_08540_),
    .Z(_13288_)
  );
  INV_X1 _20980_ (
    .A(_13288_),
    .ZN(_13289_)
  );
  MUX2_X1 _20981_ (
    .A(\rf[29] [29]),
    .B(\rf[25] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13290_)
  );
  AND2_X1 _20982_ (
    .A1(_08540_),
    .A2(_13290_),
    .ZN(_13291_)
  );
  INV_X1 _20983_ (
    .A(_13291_),
    .ZN(_13292_)
  );
  MUX2_X1 _20984_ (
    .A(\rf[28] [29]),
    .B(\rf[24] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13293_)
  );
  AND2_X1 _20985_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13293_),
    .ZN(_13294_)
  );
  INV_X1 _20986_ (
    .A(_13294_),
    .ZN(_13295_)
  );
  AND2_X1 _20987_ (
    .A1(_08541_),
    .A2(_13289_),
    .ZN(_13296_)
  );
  INV_X1 _20988_ (
    .A(_13296_),
    .ZN(_13297_)
  );
  AND2_X1 _20989_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_13295_),
    .ZN(_13298_)
  );
  AND2_X1 _20990_ (
    .A1(_13292_),
    .A2(_13298_),
    .ZN(_13299_)
  );
  INV_X1 _20991_ (
    .A(_13299_),
    .ZN(_13300_)
  );
  AND2_X1 _20992_ (
    .A1(_08543_),
    .A2(_13297_),
    .ZN(_13301_)
  );
  AND2_X1 _20993_ (
    .A1(_13300_),
    .A2(_13301_),
    .ZN(_13302_)
  );
  INV_X1 _20994_ (
    .A(_13302_),
    .ZN(_13303_)
  );
  AND2_X1 _20995_ (
    .A1(_08355_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13304_)
  );
  INV_X1 _20996_ (
    .A(_13304_),
    .ZN(_13305_)
  );
  AND2_X1 _20997_ (
    .A1(_08493_),
    .A2(_08542_),
    .ZN(_13306_)
  );
  INV_X1 _20998_ (
    .A(_13306_),
    .ZN(_13307_)
  );
  AND2_X1 _20999_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13307_),
    .ZN(_13308_)
  );
  AND2_X1 _21000_ (
    .A1(_13305_),
    .A2(_13308_),
    .ZN(_13309_)
  );
  INV_X1 _21001_ (
    .A(_13309_),
    .ZN(_13310_)
  );
  MUX2_X1 _21002_ (
    .A(\rf[23] [29]),
    .B(\rf[19] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13311_)
  );
  AND2_X1 _21003_ (
    .A1(_08540_),
    .A2(_13311_),
    .ZN(_13312_)
  );
  INV_X1 _21004_ (
    .A(_13312_),
    .ZN(_13313_)
  );
  AND2_X1 _21005_ (
    .A1(_08541_),
    .A2(_13313_),
    .ZN(_13314_)
  );
  AND2_X1 _21006_ (
    .A1(_13310_),
    .A2(_13314_),
    .ZN(_13315_)
  );
  INV_X1 _21007_ (
    .A(_13315_),
    .ZN(_13316_)
  );
  MUX2_X1 _21008_ (
    .A(\rf[21] [29]),
    .B(\rf[17] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13317_)
  );
  AND2_X1 _21009_ (
    .A1(_08540_),
    .A2(_13317_),
    .ZN(_13318_)
  );
  INV_X1 _21010_ (
    .A(_13318_),
    .ZN(_13319_)
  );
  AND2_X1 _21011_ (
    .A1(_08402_),
    .A2(_08542_),
    .ZN(_13320_)
  );
  INV_X1 _21012_ (
    .A(_13320_),
    .ZN(_13321_)
  );
  AND2_X1 _21013_ (
    .A1(_08303_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13322_)
  );
  INV_X1 _21014_ (
    .A(_13322_),
    .ZN(_13323_)
  );
  AND2_X1 _21015_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13323_),
    .ZN(_13324_)
  );
  AND2_X1 _21016_ (
    .A1(_13321_),
    .A2(_13324_),
    .ZN(_13325_)
  );
  INV_X1 _21017_ (
    .A(_13325_),
    .ZN(_13326_)
  );
  AND2_X1 _21018_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_13319_),
    .ZN(_13327_)
  );
  AND2_X1 _21019_ (
    .A1(_13326_),
    .A2(_13327_),
    .ZN(_13328_)
  );
  INV_X1 _21020_ (
    .A(_13328_),
    .ZN(_13329_)
  );
  AND2_X1 _21021_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_13316_),
    .ZN(_13330_)
  );
  AND2_X1 _21022_ (
    .A1(_13329_),
    .A2(_13330_),
    .ZN(_13331_)
  );
  INV_X1 _21023_ (
    .A(_13331_),
    .ZN(_13332_)
  );
  AND2_X1 _21024_ (
    .A1(_13303_),
    .A2(_13332_),
    .ZN(_13333_)
  );
  MUX2_X1 _21025_ (
    .A(_13285_),
    .B(_13333_),
    .S(_08571_),
    .Z(_13334_)
  );
  INV_X1 _21026_ (
    .A(_13334_),
    .ZN(_13335_)
  );
  MUX2_X1 _21027_ (
    .A(csr_io_rw_rdata[29]),
    .B(wb_reg_wdata[29]),
    .S(_10134_),
    .Z(_13336_)
  );
  MUX2_X1 _21028_ (
    .A(div_io_resp_bits_data[29]),
    .B(_13336_),
    .S(_08649_),
    .Z(_13337_)
  );
  MUX2_X1 _21029_ (
    .A(_13337_),
    .B(io_dmem_resp_bits_data[29]),
    .S(_08631_),
    .Z(_13338_)
  );
  MUX2_X1 _21030_ (
    .A(_13335_),
    .B(_13338_),
    .S(_10131_),
    .Z(_13339_)
  );
  AND2_X1 _21031_ (
    .A1(_10082_),
    .A2(_13339_),
    .ZN(_13340_)
  );
  INV_X1 _21032_ (
    .A(_13340_),
    .ZN(_13341_)
  );
  AND2_X1 _21033_ (
    .A1(_13226_),
    .A2(_13341_),
    .ZN(_13342_)
  );
  INV_X1 _21034_ (
    .A(_13342_),
    .ZN(_13343_)
  );
  MUX2_X1 _21035_ (
    .A(ex_reg_rs_msb_0[27]),
    .B(_13343_),
    .S(_10079_),
    .Z(_00094_)
  );
  AND2_X1 _21036_ (
    .A1(_08578_),
    .A2(ibuf_io_inst_0_bits_raw[30]),
    .ZN(_13344_)
  );
  AND2_X1 _21037_ (
    .A1(_09295_),
    .A2(_13344_),
    .ZN(_13345_)
  );
  INV_X1 _21038_ (
    .A(_13345_),
    .ZN(_13346_)
  );
  MUX2_X1 _21039_ (
    .A(csr_io_rw_rdata[30]),
    .B(wb_reg_wdata[30]),
    .S(_10134_),
    .Z(_13347_)
  );
  MUX2_X1 _21040_ (
    .A(div_io_resp_bits_data[30]),
    .B(_13347_),
    .S(_08649_),
    .Z(_13348_)
  );
  MUX2_X1 _21041_ (
    .A(_13348_),
    .B(io_dmem_resp_bits_data[30]),
    .S(_08631_),
    .Z(_13349_)
  );
  MUX2_X1 _21042_ (
    .A(\rf[5] [30]),
    .B(\rf[1] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13350_)
  );
  MUX2_X1 _21043_ (
    .A(\rf[7] [30]),
    .B(\rf[3] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13351_)
  );
  MUX2_X1 _21044_ (
    .A(_13350_),
    .B(_13351_),
    .S(_08541_),
    .Z(_13352_)
  );
  AND2_X1 _21045_ (
    .A1(_08540_),
    .A2(_13352_),
    .ZN(_13353_)
  );
  INV_X1 _21046_ (
    .A(_13353_),
    .ZN(_13354_)
  );
  MUX2_X1 _21047_ (
    .A(\rf[4] [30]),
    .B(\rf[0] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13355_)
  );
  MUX2_X1 _21048_ (
    .A(\rf[6] [30]),
    .B(\rf[2] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13356_)
  );
  MUX2_X1 _21049_ (
    .A(_13355_),
    .B(_13356_),
    .S(_08541_),
    .Z(_13357_)
  );
  AND2_X1 _21050_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13357_),
    .ZN(_13358_)
  );
  INV_X1 _21051_ (
    .A(_13358_),
    .ZN(_13359_)
  );
  AND2_X1 _21052_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_13359_),
    .ZN(_13360_)
  );
  AND2_X1 _21053_ (
    .A1(_13354_),
    .A2(_13360_),
    .ZN(_13361_)
  );
  INV_X1 _21054_ (
    .A(_13361_),
    .ZN(_13362_)
  );
  AND2_X1 _21055_ (
    .A1(_08403_),
    .A2(_08542_),
    .ZN(_13363_)
  );
  INV_X1 _21056_ (
    .A(_13363_),
    .ZN(_13364_)
  );
  AND2_X1 _21057_ (
    .A1(_08304_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13365_)
  );
  INV_X1 _21058_ (
    .A(_13365_),
    .ZN(_13366_)
  );
  AND2_X1 _21059_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_13366_),
    .ZN(_13367_)
  );
  AND2_X1 _21060_ (
    .A1(_13364_),
    .A2(_13367_),
    .ZN(_13368_)
  );
  INV_X1 _21061_ (
    .A(_13368_),
    .ZN(_13369_)
  );
  MUX2_X1 _21062_ (
    .A(\rf[22] [30]),
    .B(\rf[18] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13370_)
  );
  AND2_X1 _21063_ (
    .A1(_08541_),
    .A2(_13370_),
    .ZN(_13371_)
  );
  INV_X1 _21064_ (
    .A(_13371_),
    .ZN(_13372_)
  );
  AND2_X1 _21065_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13372_),
    .ZN(_13373_)
  );
  AND2_X1 _21066_ (
    .A1(_13369_),
    .A2(_13373_),
    .ZN(_13374_)
  );
  INV_X1 _21067_ (
    .A(_13374_),
    .ZN(_13375_)
  );
  AND2_X1 _21068_ (
    .A1(_08334_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13376_)
  );
  INV_X1 _21069_ (
    .A(_13376_),
    .ZN(_13377_)
  );
  AND2_X1 _21070_ (
    .A1(_08433_),
    .A2(_08542_),
    .ZN(_13378_)
  );
  INV_X1 _21071_ (
    .A(_13378_),
    .ZN(_13379_)
  );
  AND2_X1 _21072_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_13379_),
    .ZN(_13380_)
  );
  AND2_X1 _21073_ (
    .A1(_13377_),
    .A2(_13380_),
    .ZN(_13381_)
  );
  INV_X1 _21074_ (
    .A(_13381_),
    .ZN(_13382_)
  );
  MUX2_X1 _21075_ (
    .A(\rf[23] [30]),
    .B(\rf[19] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13383_)
  );
  AND2_X1 _21076_ (
    .A1(_08541_),
    .A2(_13383_),
    .ZN(_13384_)
  );
  INV_X1 _21077_ (
    .A(_13384_),
    .ZN(_13385_)
  );
  AND2_X1 _21078_ (
    .A1(_08540_),
    .A2(_13385_),
    .ZN(_13386_)
  );
  AND2_X1 _21079_ (
    .A1(_13382_),
    .A2(_13386_),
    .ZN(_13387_)
  );
  INV_X1 _21080_ (
    .A(_13387_),
    .ZN(_13388_)
  );
  AND2_X1 _21081_ (
    .A1(_13375_),
    .A2(_13388_),
    .ZN(_13389_)
  );
  INV_X1 _21082_ (
    .A(_13389_),
    .ZN(_13390_)
  );
  AND2_X1 _21083_ (
    .A1(_08571_),
    .A2(_13390_),
    .ZN(_13391_)
  );
  INV_X1 _21084_ (
    .A(_13391_),
    .ZN(_13392_)
  );
  AND2_X1 _21085_ (
    .A1(_13362_),
    .A2(_13392_),
    .ZN(_13393_)
  );
  AND2_X1 _21086_ (
    .A1(\rf[10] [30]),
    .A2(_08541_),
    .ZN(_13394_)
  );
  INV_X1 _21087_ (
    .A(_13394_),
    .ZN(_13395_)
  );
  AND2_X1 _21088_ (
    .A1(\rf[8] [30]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_13396_)
  );
  INV_X1 _21089_ (
    .A(_13396_),
    .ZN(_13397_)
  );
  AND2_X1 _21090_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_13397_),
    .ZN(_13398_)
  );
  AND2_X1 _21091_ (
    .A1(_13395_),
    .A2(_13398_),
    .ZN(_13399_)
  );
  INV_X1 _21092_ (
    .A(_13399_),
    .ZN(_13400_)
  );
  AND2_X1 _21093_ (
    .A1(\rf[14] [30]),
    .A2(_08541_),
    .ZN(_13401_)
  );
  INV_X1 _21094_ (
    .A(_13401_),
    .ZN(_13402_)
  );
  AND2_X1 _21095_ (
    .A1(\rf[12] [30]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_13403_)
  );
  INV_X1 _21096_ (
    .A(_13403_),
    .ZN(_13404_)
  );
  AND2_X1 _21097_ (
    .A1(_08542_),
    .A2(_13404_),
    .ZN(_13405_)
  );
  AND2_X1 _21098_ (
    .A1(_13402_),
    .A2(_13405_),
    .ZN(_13406_)
  );
  INV_X1 _21099_ (
    .A(_13406_),
    .ZN(_13407_)
  );
  AND2_X1 _21100_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13407_),
    .ZN(_13408_)
  );
  AND2_X1 _21101_ (
    .A1(_13400_),
    .A2(_13408_),
    .ZN(_13409_)
  );
  INV_X1 _21102_ (
    .A(_13409_),
    .ZN(_13410_)
  );
  AND2_X1 _21103_ (
    .A1(\rf[11] [30]),
    .A2(_08541_),
    .ZN(_13411_)
  );
  INV_X1 _21104_ (
    .A(_13411_),
    .ZN(_13412_)
  );
  AND2_X1 _21105_ (
    .A1(\rf[9] [30]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_13413_)
  );
  INV_X1 _21106_ (
    .A(_13413_),
    .ZN(_13414_)
  );
  AND2_X1 _21107_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_13414_),
    .ZN(_13415_)
  );
  AND2_X1 _21108_ (
    .A1(_13412_),
    .A2(_13415_),
    .ZN(_13416_)
  );
  INV_X1 _21109_ (
    .A(_13416_),
    .ZN(_13417_)
  );
  AND2_X1 _21110_ (
    .A1(\rf[15] [30]),
    .A2(_08541_),
    .ZN(_13418_)
  );
  INV_X1 _21111_ (
    .A(_13418_),
    .ZN(_13419_)
  );
  AND2_X1 _21112_ (
    .A1(\rf[13] [30]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_13420_)
  );
  INV_X1 _21113_ (
    .A(_13420_),
    .ZN(_13421_)
  );
  AND2_X1 _21114_ (
    .A1(_08542_),
    .A2(_13421_),
    .ZN(_13422_)
  );
  AND2_X1 _21115_ (
    .A1(_13419_),
    .A2(_13422_),
    .ZN(_13423_)
  );
  INV_X1 _21116_ (
    .A(_13423_),
    .ZN(_13424_)
  );
  AND2_X1 _21117_ (
    .A1(_08540_),
    .A2(_13424_),
    .ZN(_13425_)
  );
  AND2_X1 _21118_ (
    .A1(_13417_),
    .A2(_13425_),
    .ZN(_13426_)
  );
  INV_X1 _21119_ (
    .A(_13426_),
    .ZN(_13427_)
  );
  AND2_X1 _21120_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_13427_),
    .ZN(_13428_)
  );
  AND2_X1 _21121_ (
    .A1(_13410_),
    .A2(_13428_),
    .ZN(_13429_)
  );
  INV_X1 _21122_ (
    .A(_13429_),
    .ZN(_13430_)
  );
  AND2_X1 _21123_ (
    .A1(\rf[30] [30]),
    .A2(_08542_),
    .ZN(_13431_)
  );
  INV_X1 _21124_ (
    .A(_13431_),
    .ZN(_13432_)
  );
  AND2_X1 _21125_ (
    .A1(\rf[26] [30]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13433_)
  );
  INV_X1 _21126_ (
    .A(_13433_),
    .ZN(_13434_)
  );
  AND2_X1 _21127_ (
    .A1(_08541_),
    .A2(_13434_),
    .ZN(_13435_)
  );
  AND2_X1 _21128_ (
    .A1(_13432_),
    .A2(_13435_),
    .ZN(_13436_)
  );
  INV_X1 _21129_ (
    .A(_13436_),
    .ZN(_13437_)
  );
  AND2_X1 _21130_ (
    .A1(\rf[24] [30]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13438_)
  );
  INV_X1 _21131_ (
    .A(_13438_),
    .ZN(_13439_)
  );
  AND2_X1 _21132_ (
    .A1(\rf[28] [30]),
    .A2(_08542_),
    .ZN(_13440_)
  );
  INV_X1 _21133_ (
    .A(_13440_),
    .ZN(_13441_)
  );
  AND2_X1 _21134_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_13441_),
    .ZN(_13442_)
  );
  AND2_X1 _21135_ (
    .A1(_13439_),
    .A2(_13442_),
    .ZN(_13443_)
  );
  INV_X1 _21136_ (
    .A(_13443_),
    .ZN(_13444_)
  );
  AND2_X1 _21137_ (
    .A1(_13437_),
    .A2(_13444_),
    .ZN(_13445_)
  );
  MUX2_X1 _21138_ (
    .A(\rf[29] [30]),
    .B(\rf[25] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13446_)
  );
  AND2_X1 _21139_ (
    .A1(\rf[27] [30]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13447_)
  );
  MUX2_X1 _21140_ (
    .A(_13446_),
    .B(_13447_),
    .S(_08541_),
    .Z(_13448_)
  );
  MUX2_X1 _21141_ (
    .A(_13445_),
    .B(_13448_),
    .S(_08540_),
    .Z(_13449_)
  );
  INV_X1 _21142_ (
    .A(_13449_),
    .ZN(_13450_)
  );
  AND2_X1 _21143_ (
    .A1(_08571_),
    .A2(_13450_),
    .ZN(_13451_)
  );
  INV_X1 _21144_ (
    .A(_13451_),
    .ZN(_13452_)
  );
  AND2_X1 _21145_ (
    .A1(_13430_),
    .A2(_13452_),
    .ZN(_13453_)
  );
  MUX2_X1 _21146_ (
    .A(_13393_),
    .B(_13453_),
    .S(_08543_),
    .Z(_13454_)
  );
  MUX2_X1 _21147_ (
    .A(_13454_),
    .B(_13349_),
    .S(_10131_),
    .Z(_13455_)
  );
  AND2_X1 _21148_ (
    .A1(_10082_),
    .A2(_13455_),
    .ZN(_13456_)
  );
  INV_X1 _21149_ (
    .A(_13456_),
    .ZN(_13457_)
  );
  AND2_X1 _21150_ (
    .A1(_13346_),
    .A2(_13457_),
    .ZN(_13458_)
  );
  INV_X1 _21151_ (
    .A(_13458_),
    .ZN(_13459_)
  );
  MUX2_X1 _21152_ (
    .A(ex_reg_rs_msb_0[28]),
    .B(_13459_),
    .S(_10079_),
    .Z(_00095_)
  );
  AND2_X1 _21153_ (
    .A1(_08578_),
    .A2(ibuf_io_inst_0_bits_raw[31]),
    .ZN(_13460_)
  );
  AND2_X1 _21154_ (
    .A1(_09295_),
    .A2(_13460_),
    .ZN(_13461_)
  );
  INV_X1 _21155_ (
    .A(_13461_),
    .ZN(_13462_)
  );
  MUX2_X1 _21156_ (
    .A(csr_io_rw_rdata[31]),
    .B(wb_reg_wdata[31]),
    .S(_10134_),
    .Z(_13463_)
  );
  MUX2_X1 _21157_ (
    .A(div_io_resp_bits_data[31]),
    .B(_13463_),
    .S(_08649_),
    .Z(_13464_)
  );
  MUX2_X1 _21158_ (
    .A(_13464_),
    .B(io_dmem_resp_bits_data[31]),
    .S(_08631_),
    .Z(_13465_)
  );
  MUX2_X1 _21159_ (
    .A(\rf[5] [31]),
    .B(\rf[1] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13466_)
  );
  MUX2_X1 _21160_ (
    .A(\rf[7] [31]),
    .B(\rf[3] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13467_)
  );
  MUX2_X1 _21161_ (
    .A(_13466_),
    .B(_13467_),
    .S(_08541_),
    .Z(_13468_)
  );
  AND2_X1 _21162_ (
    .A1(_08540_),
    .A2(_13468_),
    .ZN(_13469_)
  );
  INV_X1 _21163_ (
    .A(_13469_),
    .ZN(_13470_)
  );
  MUX2_X1 _21164_ (
    .A(\rf[4] [31]),
    .B(\rf[0] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13471_)
  );
  MUX2_X1 _21165_ (
    .A(\rf[6] [31]),
    .B(\rf[2] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13472_)
  );
  MUX2_X1 _21166_ (
    .A(_13471_),
    .B(_13472_),
    .S(_08541_),
    .Z(_13473_)
  );
  AND2_X1 _21167_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13473_),
    .ZN(_13474_)
  );
  INV_X1 _21168_ (
    .A(_13474_),
    .ZN(_13475_)
  );
  AND2_X1 _21169_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_13475_),
    .ZN(_13476_)
  );
  AND2_X1 _21170_ (
    .A1(_13470_),
    .A2(_13476_),
    .ZN(_13477_)
  );
  INV_X1 _21171_ (
    .A(_13477_),
    .ZN(_13478_)
  );
  AND2_X1 _21172_ (
    .A1(_08230_),
    .A2(_08542_),
    .ZN(_13479_)
  );
  INV_X1 _21173_ (
    .A(_13479_),
    .ZN(_13480_)
  );
  AND2_X1 _21174_ (
    .A1(_08232_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13481_)
  );
  INV_X1 _21175_ (
    .A(_13481_),
    .ZN(_13482_)
  );
  AND2_X1 _21176_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_13482_),
    .ZN(_13483_)
  );
  AND2_X1 _21177_ (
    .A1(_13480_),
    .A2(_13483_),
    .ZN(_13484_)
  );
  INV_X1 _21178_ (
    .A(_13484_),
    .ZN(_13485_)
  );
  MUX2_X1 _21179_ (
    .A(\rf[22] [31]),
    .B(\rf[18] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13486_)
  );
  AND2_X1 _21180_ (
    .A1(_08541_),
    .A2(_13486_),
    .ZN(_13487_)
  );
  INV_X1 _21181_ (
    .A(_13487_),
    .ZN(_13488_)
  );
  AND2_X1 _21182_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13488_),
    .ZN(_13489_)
  );
  AND2_X1 _21183_ (
    .A1(_13485_),
    .A2(_13489_),
    .ZN(_13490_)
  );
  INV_X1 _21184_ (
    .A(_13490_),
    .ZN(_13491_)
  );
  AND2_X1 _21185_ (
    .A1(_08231_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13492_)
  );
  INV_X1 _21186_ (
    .A(_13492_),
    .ZN(_13493_)
  );
  AND2_X1 _21187_ (
    .A1(_08229_),
    .A2(_08542_),
    .ZN(_13494_)
  );
  INV_X1 _21188_ (
    .A(_13494_),
    .ZN(_13495_)
  );
  AND2_X1 _21189_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_13495_),
    .ZN(_13496_)
  );
  AND2_X1 _21190_ (
    .A1(_13493_),
    .A2(_13496_),
    .ZN(_13497_)
  );
  INV_X1 _21191_ (
    .A(_13497_),
    .ZN(_13498_)
  );
  MUX2_X1 _21192_ (
    .A(\rf[23] [31]),
    .B(\rf[19] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13499_)
  );
  AND2_X1 _21193_ (
    .A1(_08541_),
    .A2(_13499_),
    .ZN(_13500_)
  );
  INV_X1 _21194_ (
    .A(_13500_),
    .ZN(_13501_)
  );
  AND2_X1 _21195_ (
    .A1(_08540_),
    .A2(_13501_),
    .ZN(_13502_)
  );
  AND2_X1 _21196_ (
    .A1(_13498_),
    .A2(_13502_),
    .ZN(_13503_)
  );
  INV_X1 _21197_ (
    .A(_13503_),
    .ZN(_13504_)
  );
  AND2_X1 _21198_ (
    .A1(_13491_),
    .A2(_13504_),
    .ZN(_13505_)
  );
  INV_X1 _21199_ (
    .A(_13505_),
    .ZN(_13506_)
  );
  AND2_X1 _21200_ (
    .A1(_08571_),
    .A2(_13506_),
    .ZN(_13507_)
  );
  INV_X1 _21201_ (
    .A(_13507_),
    .ZN(_13508_)
  );
  AND2_X1 _21202_ (
    .A1(_13478_),
    .A2(_13508_),
    .ZN(_13509_)
  );
  AND2_X1 _21203_ (
    .A1(\rf[10] [31]),
    .A2(_08541_),
    .ZN(_13510_)
  );
  INV_X1 _21204_ (
    .A(_13510_),
    .ZN(_13511_)
  );
  AND2_X1 _21205_ (
    .A1(\rf[8] [31]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_13512_)
  );
  INV_X1 _21206_ (
    .A(_13512_),
    .ZN(_13513_)
  );
  AND2_X1 _21207_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_13513_),
    .ZN(_13514_)
  );
  AND2_X1 _21208_ (
    .A1(_13511_),
    .A2(_13514_),
    .ZN(_13515_)
  );
  INV_X1 _21209_ (
    .A(_13515_),
    .ZN(_13516_)
  );
  AND2_X1 _21210_ (
    .A1(\rf[14] [31]),
    .A2(_08541_),
    .ZN(_13517_)
  );
  INV_X1 _21211_ (
    .A(_13517_),
    .ZN(_13518_)
  );
  AND2_X1 _21212_ (
    .A1(\rf[12] [31]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_13519_)
  );
  INV_X1 _21213_ (
    .A(_13519_),
    .ZN(_13520_)
  );
  AND2_X1 _21214_ (
    .A1(_08542_),
    .A2(_13520_),
    .ZN(_13521_)
  );
  AND2_X1 _21215_ (
    .A1(_13518_),
    .A2(_13521_),
    .ZN(_13522_)
  );
  INV_X1 _21216_ (
    .A(_13522_),
    .ZN(_13523_)
  );
  AND2_X1 _21217_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13523_),
    .ZN(_13524_)
  );
  AND2_X1 _21218_ (
    .A1(_13516_),
    .A2(_13524_),
    .ZN(_13525_)
  );
  INV_X1 _21219_ (
    .A(_13525_),
    .ZN(_13526_)
  );
  AND2_X1 _21220_ (
    .A1(\rf[11] [31]),
    .A2(_08541_),
    .ZN(_13527_)
  );
  INV_X1 _21221_ (
    .A(_13527_),
    .ZN(_13528_)
  );
  AND2_X1 _21222_ (
    .A1(\rf[9] [31]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_13529_)
  );
  INV_X1 _21223_ (
    .A(_13529_),
    .ZN(_13530_)
  );
  AND2_X1 _21224_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_13530_),
    .ZN(_13531_)
  );
  AND2_X1 _21225_ (
    .A1(_13528_),
    .A2(_13531_),
    .ZN(_13532_)
  );
  INV_X1 _21226_ (
    .A(_13532_),
    .ZN(_13533_)
  );
  AND2_X1 _21227_ (
    .A1(\rf[15] [31]),
    .A2(_08541_),
    .ZN(_13534_)
  );
  INV_X1 _21228_ (
    .A(_13534_),
    .ZN(_13535_)
  );
  AND2_X1 _21229_ (
    .A1(\rf[13] [31]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_13536_)
  );
  INV_X1 _21230_ (
    .A(_13536_),
    .ZN(_13537_)
  );
  AND2_X1 _21231_ (
    .A1(_08542_),
    .A2(_13537_),
    .ZN(_13538_)
  );
  AND2_X1 _21232_ (
    .A1(_13535_),
    .A2(_13538_),
    .ZN(_13539_)
  );
  INV_X1 _21233_ (
    .A(_13539_),
    .ZN(_13540_)
  );
  AND2_X1 _21234_ (
    .A1(_08540_),
    .A2(_13540_),
    .ZN(_13541_)
  );
  AND2_X1 _21235_ (
    .A1(_13533_),
    .A2(_13541_),
    .ZN(_13542_)
  );
  INV_X1 _21236_ (
    .A(_13542_),
    .ZN(_13543_)
  );
  AND2_X1 _21237_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_13543_),
    .ZN(_13544_)
  );
  AND2_X1 _21238_ (
    .A1(_13526_),
    .A2(_13544_),
    .ZN(_13545_)
  );
  INV_X1 _21239_ (
    .A(_13545_),
    .ZN(_13546_)
  );
  AND2_X1 _21240_ (
    .A1(\rf[30] [31]),
    .A2(_08542_),
    .ZN(_13547_)
  );
  INV_X1 _21241_ (
    .A(_13547_),
    .ZN(_13548_)
  );
  AND2_X1 _21242_ (
    .A1(\rf[26] [31]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13549_)
  );
  INV_X1 _21243_ (
    .A(_13549_),
    .ZN(_13550_)
  );
  AND2_X1 _21244_ (
    .A1(_08541_),
    .A2(_13550_),
    .ZN(_13551_)
  );
  AND2_X1 _21245_ (
    .A1(_13548_),
    .A2(_13551_),
    .ZN(_13552_)
  );
  INV_X1 _21246_ (
    .A(_13552_),
    .ZN(_13553_)
  );
  AND2_X1 _21247_ (
    .A1(\rf[24] [31]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13554_)
  );
  INV_X1 _21248_ (
    .A(_13554_),
    .ZN(_13555_)
  );
  AND2_X1 _21249_ (
    .A1(\rf[28] [31]),
    .A2(_08542_),
    .ZN(_13556_)
  );
  INV_X1 _21250_ (
    .A(_13556_),
    .ZN(_13557_)
  );
  AND2_X1 _21251_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_13557_),
    .ZN(_13558_)
  );
  AND2_X1 _21252_ (
    .A1(_13555_),
    .A2(_13558_),
    .ZN(_13559_)
  );
  INV_X1 _21253_ (
    .A(_13559_),
    .ZN(_13560_)
  );
  AND2_X1 _21254_ (
    .A1(_13553_),
    .A2(_13560_),
    .ZN(_13561_)
  );
  MUX2_X1 _21255_ (
    .A(\rf[29] [31]),
    .B(\rf[25] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13562_)
  );
  AND2_X1 _21256_ (
    .A1(\rf[27] [31]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13563_)
  );
  MUX2_X1 _21257_ (
    .A(_13562_),
    .B(_13563_),
    .S(_08541_),
    .Z(_13564_)
  );
  MUX2_X1 _21258_ (
    .A(_13561_),
    .B(_13564_),
    .S(_08540_),
    .Z(_13565_)
  );
  INV_X1 _21259_ (
    .A(_13565_),
    .ZN(_13566_)
  );
  AND2_X1 _21260_ (
    .A1(_08571_),
    .A2(_13566_),
    .ZN(_13567_)
  );
  INV_X1 _21261_ (
    .A(_13567_),
    .ZN(_13568_)
  );
  AND2_X1 _21262_ (
    .A1(_13546_),
    .A2(_13568_),
    .ZN(_13569_)
  );
  MUX2_X1 _21263_ (
    .A(_13509_),
    .B(_13569_),
    .S(_08543_),
    .Z(_13570_)
  );
  MUX2_X1 _21264_ (
    .A(_13570_),
    .B(_13465_),
    .S(_10131_),
    .Z(_13571_)
  );
  AND2_X1 _21265_ (
    .A1(_10082_),
    .A2(_13571_),
    .ZN(_13572_)
  );
  INV_X1 _21266_ (
    .A(_13572_),
    .ZN(_13573_)
  );
  AND2_X1 _21267_ (
    .A1(_13462_),
    .A2(_13573_),
    .ZN(_13574_)
  );
  INV_X1 _21268_ (
    .A(_13574_),
    .ZN(_13575_)
  );
  MUX2_X1 _21269_ (
    .A(ex_reg_rs_msb_0[29]),
    .B(_13575_),
    .S(_10079_),
    .Z(_00096_)
  );
  AND2_X1 _21270_ (
    .A1(_08127_),
    .A2(_09295_),
    .ZN(_13576_)
  );
  INV_X1 _21271_ (
    .A(_13576_),
    .ZN(_13577_)
  );
  MUX2_X1 _21272_ (
    .A(csr_io_rw_rdata[0]),
    .B(wb_reg_wdata[0]),
    .S(_10134_),
    .Z(_13578_)
  );
  MUX2_X1 _21273_ (
    .A(div_io_resp_bits_data[0]),
    .B(_13578_),
    .S(_08649_),
    .Z(_13579_)
  );
  MUX2_X1 _21274_ (
    .A(_13579_),
    .B(io_dmem_resp_bits_data[0]),
    .S(_08631_),
    .Z(_13580_)
  );
  INV_X1 _21275_ (
    .A(_13580_),
    .ZN(_13581_)
  );
  AND2_X1 _21276_ (
    .A1(_10131_),
    .A2(_13581_),
    .ZN(_13582_)
  );
  INV_X1 _21277_ (
    .A(_13582_),
    .ZN(_13583_)
  );
  AND2_X1 _21278_ (
    .A1(_08305_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13584_)
  );
  INV_X1 _21279_ (
    .A(_13584_),
    .ZN(_13585_)
  );
  AND2_X1 _21280_ (
    .A1(_08404_),
    .A2(_08542_),
    .ZN(_13586_)
  );
  INV_X1 _21281_ (
    .A(_13586_),
    .ZN(_13587_)
  );
  AND2_X1 _21282_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_13587_),
    .ZN(_13588_)
  );
  AND2_X1 _21283_ (
    .A1(_13585_),
    .A2(_13588_),
    .ZN(_13589_)
  );
  INV_X1 _21284_ (
    .A(_13589_),
    .ZN(_13590_)
  );
  MUX2_X1 _21285_ (
    .A(\rf[23] [0]),
    .B(\rf[19] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13591_)
  );
  AND2_X1 _21286_ (
    .A1(_08541_),
    .A2(_13591_),
    .ZN(_13592_)
  );
  INV_X1 _21287_ (
    .A(_13592_),
    .ZN(_13593_)
  );
  AND2_X1 _21288_ (
    .A1(_08540_),
    .A2(_13593_),
    .ZN(_13594_)
  );
  AND2_X1 _21289_ (
    .A1(_13590_),
    .A2(_13594_),
    .ZN(_13595_)
  );
  INV_X1 _21290_ (
    .A(_13595_),
    .ZN(_13596_)
  );
  AND2_X1 _21291_ (
    .A1(_08373_),
    .A2(_08542_),
    .ZN(_13597_)
  );
  INV_X1 _21292_ (
    .A(_13597_),
    .ZN(_13598_)
  );
  AND2_X1 _21293_ (
    .A1(_08274_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13599_)
  );
  INV_X1 _21294_ (
    .A(_13599_),
    .ZN(_13600_)
  );
  AND2_X1 _21295_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_13600_),
    .ZN(_13601_)
  );
  AND2_X1 _21296_ (
    .A1(_13598_),
    .A2(_13601_),
    .ZN(_13602_)
  );
  INV_X1 _21297_ (
    .A(_13602_),
    .ZN(_13603_)
  );
  MUX2_X1 _21298_ (
    .A(\rf[22] [0]),
    .B(\rf[18] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13604_)
  );
  AND2_X1 _21299_ (
    .A1(_08541_),
    .A2(_13604_),
    .ZN(_13605_)
  );
  INV_X1 _21300_ (
    .A(_13605_),
    .ZN(_13606_)
  );
  AND2_X1 _21301_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13606_),
    .ZN(_13607_)
  );
  AND2_X1 _21302_ (
    .A1(_13603_),
    .A2(_13607_),
    .ZN(_13608_)
  );
  INV_X1 _21303_ (
    .A(_13608_),
    .ZN(_13609_)
  );
  AND2_X1 _21304_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_13596_),
    .ZN(_13610_)
  );
  AND2_X1 _21305_ (
    .A1(_13609_),
    .A2(_13610_),
    .ZN(_13611_)
  );
  INV_X1 _21306_ (
    .A(_13611_),
    .ZN(_13612_)
  );
  AND2_X1 _21307_ (
    .A1(_08434_),
    .A2(_08542_),
    .ZN(_13613_)
  );
  INV_X1 _21308_ (
    .A(_13613_),
    .ZN(_13614_)
  );
  AND2_X1 _21309_ (
    .A1(_08504_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13615_)
  );
  INV_X1 _21310_ (
    .A(_13615_),
    .ZN(_13616_)
  );
  AND2_X1 _21311_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_13616_),
    .ZN(_13617_)
  );
  AND2_X1 _21312_ (
    .A1(_13614_),
    .A2(_13617_),
    .ZN(_13618_)
  );
  INV_X1 _21313_ (
    .A(_13618_),
    .ZN(_13619_)
  );
  MUX2_X1 _21314_ (
    .A(\rf[30] [0]),
    .B(\rf[26] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13620_)
  );
  AND2_X1 _21315_ (
    .A1(_08541_),
    .A2(_13620_),
    .ZN(_13621_)
  );
  INV_X1 _21316_ (
    .A(_13621_),
    .ZN(_13622_)
  );
  AND2_X1 _21317_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13622_),
    .ZN(_13623_)
  );
  AND2_X1 _21318_ (
    .A1(_13619_),
    .A2(_13623_),
    .ZN(_13624_)
  );
  INV_X1 _21319_ (
    .A(_13624_),
    .ZN(_13625_)
  );
  MUX2_X1 _21320_ (
    .A(\rf[29] [0]),
    .B(\rf[25] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13626_)
  );
  AND2_X1 _21321_ (
    .A1(\rf[27] [0]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13627_)
  );
  MUX2_X1 _21322_ (
    .A(_13626_),
    .B(_13627_),
    .S(_08541_),
    .Z(_13628_)
  );
  INV_X1 _21323_ (
    .A(_13628_),
    .ZN(_13629_)
  );
  AND2_X1 _21324_ (
    .A1(_08540_),
    .A2(_13629_),
    .ZN(_13630_)
  );
  INV_X1 _21325_ (
    .A(_13630_),
    .ZN(_13631_)
  );
  AND2_X1 _21326_ (
    .A1(_08543_),
    .A2(_13631_),
    .ZN(_13632_)
  );
  AND2_X1 _21327_ (
    .A1(_13625_),
    .A2(_13632_),
    .ZN(_13633_)
  );
  INV_X1 _21328_ (
    .A(_13633_),
    .ZN(_13634_)
  );
  AND2_X1 _21329_ (
    .A1(_13612_),
    .A2(_13634_),
    .ZN(_13635_)
  );
  AND2_X1 _21330_ (
    .A1(_08335_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13636_)
  );
  INV_X1 _21331_ (
    .A(_13636_),
    .ZN(_13637_)
  );
  AND2_X1 _21332_ (
    .A1(_08473_),
    .A2(_08542_),
    .ZN(_13638_)
  );
  INV_X1 _21333_ (
    .A(_13638_),
    .ZN(_13639_)
  );
  AND2_X1 _21334_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13639_),
    .ZN(_13640_)
  );
  AND2_X1 _21335_ (
    .A1(_13637_),
    .A2(_13640_),
    .ZN(_13641_)
  );
  INV_X1 _21336_ (
    .A(_13641_),
    .ZN(_13642_)
  );
  MUX2_X1 _21337_ (
    .A(\rf[15] [0]),
    .B(\rf[11] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13643_)
  );
  AND2_X1 _21338_ (
    .A1(_08540_),
    .A2(_13643_),
    .ZN(_13644_)
  );
  INV_X1 _21339_ (
    .A(_13644_),
    .ZN(_13645_)
  );
  AND2_X1 _21340_ (
    .A1(_08541_),
    .A2(_13645_),
    .ZN(_13646_)
  );
  AND2_X1 _21341_ (
    .A1(_13642_),
    .A2(_13646_),
    .ZN(_13647_)
  );
  INV_X1 _21342_ (
    .A(_13647_),
    .ZN(_13648_)
  );
  AND2_X1 _21343_ (
    .A1(_08356_),
    .A2(_08542_),
    .ZN(_13649_)
  );
  INV_X1 _21344_ (
    .A(_13649_),
    .ZN(_13650_)
  );
  AND2_X1 _21345_ (
    .A1(_08257_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13651_)
  );
  INV_X1 _21346_ (
    .A(_13651_),
    .ZN(_13652_)
  );
  AND2_X1 _21347_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13652_),
    .ZN(_13653_)
  );
  AND2_X1 _21348_ (
    .A1(_13650_),
    .A2(_13653_),
    .ZN(_13654_)
  );
  INV_X1 _21349_ (
    .A(_13654_),
    .ZN(_13655_)
  );
  MUX2_X1 _21350_ (
    .A(\rf[13] [0]),
    .B(\rf[9] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13656_)
  );
  AND2_X1 _21351_ (
    .A1(_08540_),
    .A2(_13656_),
    .ZN(_13657_)
  );
  INV_X1 _21352_ (
    .A(_13657_),
    .ZN(_13658_)
  );
  AND2_X1 _21353_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_13658_),
    .ZN(_13659_)
  );
  AND2_X1 _21354_ (
    .A1(_13655_),
    .A2(_13659_),
    .ZN(_13660_)
  );
  INV_X1 _21355_ (
    .A(_13660_),
    .ZN(_13661_)
  );
  AND2_X1 _21356_ (
    .A1(_08543_),
    .A2(_13661_),
    .ZN(_13662_)
  );
  AND2_X1 _21357_ (
    .A1(_13648_),
    .A2(_13662_),
    .ZN(_13663_)
  );
  INV_X1 _21358_ (
    .A(_13663_),
    .ZN(_13664_)
  );
  MUX2_X1 _21359_ (
    .A(\rf[6] [0]),
    .B(\rf[2] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13665_)
  );
  AND2_X1 _21360_ (
    .A1(_08541_),
    .A2(_13665_),
    .ZN(_13666_)
  );
  INV_X1 _21361_ (
    .A(_13666_),
    .ZN(_13667_)
  );
  MUX2_X1 _21362_ (
    .A(\rf[4] [0]),
    .B(\rf[0] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13668_)
  );
  AND2_X1 _21363_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_13668_),
    .ZN(_13669_)
  );
  INV_X1 _21364_ (
    .A(_13669_),
    .ZN(_13670_)
  );
  AND2_X1 _21365_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13670_),
    .ZN(_13671_)
  );
  AND2_X1 _21366_ (
    .A1(_13667_),
    .A2(_13671_),
    .ZN(_13672_)
  );
  INV_X1 _21367_ (
    .A(_13672_),
    .ZN(_13673_)
  );
  MUX2_X1 _21368_ (
    .A(\rf[7] [0]),
    .B(\rf[3] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13674_)
  );
  AND2_X1 _21369_ (
    .A1(_08541_),
    .A2(_13674_),
    .ZN(_13675_)
  );
  INV_X1 _21370_ (
    .A(_13675_),
    .ZN(_13676_)
  );
  MUX2_X1 _21371_ (
    .A(\rf[5] [0]),
    .B(\rf[1] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13677_)
  );
  AND2_X1 _21372_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_13677_),
    .ZN(_13678_)
  );
  INV_X1 _21373_ (
    .A(_13678_),
    .ZN(_13679_)
  );
  AND2_X1 _21374_ (
    .A1(_08540_),
    .A2(_13679_),
    .ZN(_13680_)
  );
  AND2_X1 _21375_ (
    .A1(_13676_),
    .A2(_13680_),
    .ZN(_13681_)
  );
  INV_X1 _21376_ (
    .A(_13681_),
    .ZN(_13682_)
  );
  AND2_X1 _21377_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_13682_),
    .ZN(_13683_)
  );
  AND2_X1 _21378_ (
    .A1(_13673_),
    .A2(_13683_),
    .ZN(_13684_)
  );
  INV_X1 _21379_ (
    .A(_13684_),
    .ZN(_13685_)
  );
  AND2_X1 _21380_ (
    .A1(_13664_),
    .A2(_13685_),
    .ZN(_13686_)
  );
  MUX2_X1 _21381_ (
    .A(_13635_),
    .B(_13686_),
    .S(ibuf_io_inst_0_bits_inst_rs1[4]),
    .Z(_13687_)
  );
  AND2_X1 _21382_ (
    .A1(_10132_),
    .A2(_13687_),
    .ZN(_13688_)
  );
  INV_X1 _21383_ (
    .A(_13688_),
    .ZN(_13689_)
  );
  AND2_X1 _21384_ (
    .A1(_09182_),
    .A2(_13583_),
    .ZN(_13690_)
  );
  AND2_X1 _21385_ (
    .A1(_13689_),
    .A2(_13690_),
    .ZN(_13691_)
  );
  INV_X1 _21386_ (
    .A(_13691_),
    .ZN(_13692_)
  );
  AND2_X1 _21387_ (
    .A1(_00028_),
    .A2(_09148_),
    .ZN(_13693_)
  );
  AND2_X1 _21388_ (
    .A1(_09177_),
    .A2(_13693_),
    .ZN(_13694_)
  );
  AND2_X1 _21389_ (
    .A1(_09146_),
    .A2(_13694_),
    .ZN(_13695_)
  );
  INV_X1 _21390_ (
    .A(_13695_),
    .ZN(_13696_)
  );
  AND2_X1 _21391_ (
    .A1(_09183_),
    .A2(_13696_),
    .ZN(_13697_)
  );
  AND2_X1 _21392_ (
    .A1(_09114_),
    .A2(_13697_),
    .ZN(_13698_)
  );
  INV_X1 _21393_ (
    .A(_13698_),
    .ZN(_13699_)
  );
  AND2_X1 _21394_ (
    .A1(_09294_),
    .A2(_13692_),
    .ZN(_13700_)
  );
  AND2_X1 _21395_ (
    .A1(_13699_),
    .A2(_13700_),
    .ZN(_13701_)
  );
  INV_X1 _21396_ (
    .A(_13701_),
    .ZN(_13702_)
  );
  AND2_X1 _21397_ (
    .A1(_13577_),
    .A2(_13702_),
    .ZN(_13703_)
  );
  MUX2_X1 _21398_ (
    .A(ex_reg_rs_lsb_0[0]),
    .B(_13703_),
    .S(_10244_),
    .Z(_00097_)
  );
  AND2_X1 _21399_ (
    .A1(_09147_),
    .A2(_09296_),
    .ZN(_13704_)
  );
  INV_X1 _21400_ (
    .A(_13704_),
    .ZN(_13705_)
  );
  AND2_X1 _21401_ (
    .A1(ibuf_io_inst_0_bits_raw[1]),
    .A2(_09295_),
    .ZN(_13706_)
  );
  INV_X1 _21402_ (
    .A(_13706_),
    .ZN(_13707_)
  );
  AND2_X1 _21403_ (
    .A1(_13705_),
    .A2(_13707_),
    .ZN(_13708_)
  );
  AND2_X1 _21404_ (
    .A1(_08336_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13709_)
  );
  INV_X1 _21405_ (
    .A(_13709_),
    .ZN(_13710_)
  );
  AND2_X1 _21406_ (
    .A1(_08474_),
    .A2(_08542_),
    .ZN(_13711_)
  );
  INV_X1 _21407_ (
    .A(_13711_),
    .ZN(_13712_)
  );
  AND2_X1 _21408_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13712_),
    .ZN(_13713_)
  );
  AND2_X1 _21409_ (
    .A1(_13710_),
    .A2(_13713_),
    .ZN(_13714_)
  );
  INV_X1 _21410_ (
    .A(_13714_),
    .ZN(_13715_)
  );
  MUX2_X1 _21411_ (
    .A(\rf[15] [1]),
    .B(\rf[11] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13716_)
  );
  AND2_X1 _21412_ (
    .A1(_08540_),
    .A2(_13716_),
    .ZN(_13717_)
  );
  INV_X1 _21413_ (
    .A(_13717_),
    .ZN(_13718_)
  );
  AND2_X1 _21414_ (
    .A1(_08541_),
    .A2(_13718_),
    .ZN(_13719_)
  );
  AND2_X1 _21415_ (
    .A1(_13715_),
    .A2(_13719_),
    .ZN(_13720_)
  );
  INV_X1 _21416_ (
    .A(_13720_),
    .ZN(_13721_)
  );
  AND2_X1 _21417_ (
    .A1(_08357_),
    .A2(_08542_),
    .ZN(_13722_)
  );
  INV_X1 _21418_ (
    .A(_13722_),
    .ZN(_13723_)
  );
  AND2_X1 _21419_ (
    .A1(_08258_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13724_)
  );
  INV_X1 _21420_ (
    .A(_13724_),
    .ZN(_13725_)
  );
  AND2_X1 _21421_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13725_),
    .ZN(_13726_)
  );
  AND2_X1 _21422_ (
    .A1(_13723_),
    .A2(_13726_),
    .ZN(_13727_)
  );
  INV_X1 _21423_ (
    .A(_13727_),
    .ZN(_13728_)
  );
  MUX2_X1 _21424_ (
    .A(\rf[13] [1]),
    .B(\rf[9] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13729_)
  );
  AND2_X1 _21425_ (
    .A1(_08540_),
    .A2(_13729_),
    .ZN(_13730_)
  );
  INV_X1 _21426_ (
    .A(_13730_),
    .ZN(_13731_)
  );
  AND2_X1 _21427_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_13731_),
    .ZN(_13732_)
  );
  AND2_X1 _21428_ (
    .A1(_13728_),
    .A2(_13732_),
    .ZN(_13733_)
  );
  INV_X1 _21429_ (
    .A(_13733_),
    .ZN(_13734_)
  );
  AND2_X1 _21430_ (
    .A1(_08543_),
    .A2(_13734_),
    .ZN(_13735_)
  );
  AND2_X1 _21431_ (
    .A1(_13721_),
    .A2(_13735_),
    .ZN(_13736_)
  );
  INV_X1 _21432_ (
    .A(_13736_),
    .ZN(_13737_)
  );
  MUX2_X1 _21433_ (
    .A(\rf[7] [1]),
    .B(\rf[3] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13738_)
  );
  AND2_X1 _21434_ (
    .A1(_08540_),
    .A2(_13738_),
    .ZN(_13739_)
  );
  INV_X1 _21435_ (
    .A(_13739_),
    .ZN(_13740_)
  );
  AND2_X1 _21436_ (
    .A1(_08501_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13741_)
  );
  INV_X1 _21437_ (
    .A(_13741_),
    .ZN(_13742_)
  );
  AND2_X1 _21438_ (
    .A1(_08245_),
    .A2(_08542_),
    .ZN(_13743_)
  );
  INV_X1 _21439_ (
    .A(_13743_),
    .ZN(_13744_)
  );
  AND2_X1 _21440_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13744_),
    .ZN(_13745_)
  );
  AND2_X1 _21441_ (
    .A1(_13742_),
    .A2(_13745_),
    .ZN(_13746_)
  );
  INV_X1 _21442_ (
    .A(_13746_),
    .ZN(_13747_)
  );
  AND2_X1 _21443_ (
    .A1(_13740_),
    .A2(_13747_),
    .ZN(_13748_)
  );
  AND2_X1 _21444_ (
    .A1(_08541_),
    .A2(_13748_),
    .ZN(_13749_)
  );
  INV_X1 _21445_ (
    .A(_13749_),
    .ZN(_13750_)
  );
  AND2_X1 _21446_ (
    .A1(_08254_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13751_)
  );
  INV_X1 _21447_ (
    .A(_13751_),
    .ZN(_13752_)
  );
  AND2_X1 _21448_ (
    .A1(_08249_),
    .A2(_08542_),
    .ZN(_13753_)
  );
  INV_X1 _21449_ (
    .A(_13753_),
    .ZN(_13754_)
  );
  AND2_X1 _21450_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13754_),
    .ZN(_13755_)
  );
  AND2_X1 _21451_ (
    .A1(_13752_),
    .A2(_13755_),
    .ZN(_13756_)
  );
  INV_X1 _21452_ (
    .A(_13756_),
    .ZN(_13757_)
  );
  MUX2_X1 _21453_ (
    .A(\rf[5] [1]),
    .B(\rf[1] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13758_)
  );
  AND2_X1 _21454_ (
    .A1(_08540_),
    .A2(_13758_),
    .ZN(_13759_)
  );
  INV_X1 _21455_ (
    .A(_13759_),
    .ZN(_13760_)
  );
  AND2_X1 _21456_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_13760_),
    .ZN(_13761_)
  );
  AND2_X1 _21457_ (
    .A1(_13757_),
    .A2(_13761_),
    .ZN(_13762_)
  );
  INV_X1 _21458_ (
    .A(_13762_),
    .ZN(_13763_)
  );
  AND2_X1 _21459_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_13763_),
    .ZN(_13764_)
  );
  AND2_X1 _21460_ (
    .A1(_13750_),
    .A2(_13764_),
    .ZN(_13765_)
  );
  INV_X1 _21461_ (
    .A(_13765_),
    .ZN(_13766_)
  );
  AND2_X1 _21462_ (
    .A1(_13737_),
    .A2(_13766_),
    .ZN(_13767_)
  );
  MUX2_X1 _21463_ (
    .A(\rf[29] [1]),
    .B(\rf[25] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13768_)
  );
  AND2_X1 _21464_ (
    .A1(_08540_),
    .A2(_13768_),
    .ZN(_13769_)
  );
  INV_X1 _21465_ (
    .A(_13769_),
    .ZN(_13770_)
  );
  MUX2_X1 _21466_ (
    .A(\rf[28] [1]),
    .B(\rf[24] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13771_)
  );
  AND2_X1 _21467_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13771_),
    .ZN(_13772_)
  );
  INV_X1 _21468_ (
    .A(_13772_),
    .ZN(_13773_)
  );
  AND2_X1 _21469_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_13773_),
    .ZN(_13774_)
  );
  AND2_X1 _21470_ (
    .A1(_13770_),
    .A2(_13774_),
    .ZN(_13775_)
  );
  INV_X1 _21471_ (
    .A(_13775_),
    .ZN(_13776_)
  );
  MUX2_X1 _21472_ (
    .A(\rf[30] [1]),
    .B(\rf[26] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13777_)
  );
  AND2_X1 _21473_ (
    .A1(\rf[27] [1]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13778_)
  );
  MUX2_X1 _21474_ (
    .A(_13777_),
    .B(_13778_),
    .S(_08540_),
    .Z(_13779_)
  );
  INV_X1 _21475_ (
    .A(_13779_),
    .ZN(_13780_)
  );
  AND2_X1 _21476_ (
    .A1(_08541_),
    .A2(_13780_),
    .ZN(_13781_)
  );
  INV_X1 _21477_ (
    .A(_13781_),
    .ZN(_13782_)
  );
  AND2_X1 _21478_ (
    .A1(_08543_),
    .A2(_13782_),
    .ZN(_13783_)
  );
  AND2_X1 _21479_ (
    .A1(_13776_),
    .A2(_13783_),
    .ZN(_13784_)
  );
  INV_X1 _21480_ (
    .A(_13784_),
    .ZN(_13785_)
  );
  AND2_X1 _21481_ (
    .A1(_08353_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13786_)
  );
  INV_X1 _21482_ (
    .A(_13786_),
    .ZN(_13787_)
  );
  AND2_X1 _21483_ (
    .A1(_08491_),
    .A2(_08542_),
    .ZN(_13788_)
  );
  INV_X1 _21484_ (
    .A(_13788_),
    .ZN(_13789_)
  );
  AND2_X1 _21485_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13789_),
    .ZN(_13790_)
  );
  AND2_X1 _21486_ (
    .A1(_13787_),
    .A2(_13790_),
    .ZN(_13791_)
  );
  INV_X1 _21487_ (
    .A(_13791_),
    .ZN(_13792_)
  );
  MUX2_X1 _21488_ (
    .A(\rf[23] [1]),
    .B(\rf[19] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13793_)
  );
  AND2_X1 _21489_ (
    .A1(_08540_),
    .A2(_13793_),
    .ZN(_13794_)
  );
  INV_X1 _21490_ (
    .A(_13794_),
    .ZN(_13795_)
  );
  AND2_X1 _21491_ (
    .A1(_08541_),
    .A2(_13795_),
    .ZN(_13796_)
  );
  AND2_X1 _21492_ (
    .A1(_13792_),
    .A2(_13796_),
    .ZN(_13797_)
  );
  INV_X1 _21493_ (
    .A(_13797_),
    .ZN(_13798_)
  );
  MUX2_X1 _21494_ (
    .A(\rf[21] [1]),
    .B(\rf[17] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_13799_)
  );
  AND2_X1 _21495_ (
    .A1(_08540_),
    .A2(_13799_),
    .ZN(_13800_)
  );
  INV_X1 _21496_ (
    .A(_13800_),
    .ZN(_13801_)
  );
  AND2_X1 _21497_ (
    .A1(_08374_),
    .A2(_08542_),
    .ZN(_13802_)
  );
  INV_X1 _21498_ (
    .A(_13802_),
    .ZN(_13803_)
  );
  AND2_X1 _21499_ (
    .A1(_08275_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_13804_)
  );
  INV_X1 _21500_ (
    .A(_13804_),
    .ZN(_13805_)
  );
  AND2_X1 _21501_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_13805_),
    .ZN(_13806_)
  );
  AND2_X1 _21502_ (
    .A1(_13803_),
    .A2(_13806_),
    .ZN(_13807_)
  );
  INV_X1 _21503_ (
    .A(_13807_),
    .ZN(_13808_)
  );
  AND2_X1 _21504_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_13801_),
    .ZN(_13809_)
  );
  AND2_X1 _21505_ (
    .A1(_13808_),
    .A2(_13809_),
    .ZN(_13810_)
  );
  INV_X1 _21506_ (
    .A(_13810_),
    .ZN(_13811_)
  );
  AND2_X1 _21507_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_13798_),
    .ZN(_13812_)
  );
  AND2_X1 _21508_ (
    .A1(_13811_),
    .A2(_13812_),
    .ZN(_13813_)
  );
  INV_X1 _21509_ (
    .A(_13813_),
    .ZN(_13814_)
  );
  AND2_X1 _21510_ (
    .A1(_13785_),
    .A2(_13814_),
    .ZN(_13815_)
  );
  MUX2_X1 _21511_ (
    .A(_13767_),
    .B(_13815_),
    .S(_08571_),
    .Z(_13816_)
  );
  INV_X1 _21512_ (
    .A(_13816_),
    .ZN(_13817_)
  );
  MUX2_X1 _21513_ (
    .A(csr_io_rw_rdata[1]),
    .B(wb_reg_wdata[1]),
    .S(_10134_),
    .Z(_13818_)
  );
  MUX2_X1 _21514_ (
    .A(div_io_resp_bits_data[1]),
    .B(_13818_),
    .S(_08649_),
    .Z(_13819_)
  );
  MUX2_X1 _21515_ (
    .A(_13819_),
    .B(io_dmem_resp_bits_data[1]),
    .S(_08631_),
    .Z(_13820_)
  );
  MUX2_X1 _21516_ (
    .A(_13817_),
    .B(_13820_),
    .S(_10131_),
    .Z(_13821_)
  );
  AND2_X1 _21517_ (
    .A1(_10082_),
    .A2(_13821_),
    .ZN(_13822_)
  );
  INV_X1 _21518_ (
    .A(_13822_),
    .ZN(_13823_)
  );
  AND2_X1 _21519_ (
    .A1(_13708_),
    .A2(_13823_),
    .ZN(_13824_)
  );
  INV_X1 _21520_ (
    .A(_13824_),
    .ZN(_13825_)
  );
  MUX2_X1 _21521_ (
    .A(ex_reg_rs_lsb_0[1]),
    .B(_13825_),
    .S(_10244_),
    .Z(_00098_)
  );
  AND2_X1 _21522_ (
    .A1(_09115_),
    .A2(_10022_),
    .ZN(_13826_)
  );
  INV_X1 _21523_ (
    .A(_13826_),
    .ZN(_13827_)
  );
  AND2_X1 _21524_ (
    .A1(_09696_),
    .A2(_13827_),
    .ZN(_13828_)
  );
  AND2_X1 _21525_ (
    .A1(_09842_),
    .A2(_13828_),
    .ZN(_13829_)
  );
  INV_X1 _21526_ (
    .A(_13829_),
    .ZN(_13830_)
  );
  MUX2_X1 _21527_ (
    .A(ex_reg_rs_bypass_1),
    .B(_13830_),
    .S(_10244_),
    .Z(_00099_)
  );
  AND2_X1 _21528_ (
    .A1(_09181_),
    .A2(_09294_),
    .ZN(_13831_)
  );
  MUX2_X1 _21529_ (
    .A(ex_reg_rs_bypass_0),
    .B(_13831_),
    .S(_10244_),
    .Z(_00100_)
  );
  AND2_X1 _21530_ (
    .A1(_08607_),
    .A2(_08623_),
    .ZN(_13832_)
  );
  AND2_X1 _21531_ (
    .A1(_08624_),
    .A2(_13832_),
    .ZN(_13833_)
  );
  INV_X1 _21532_ (
    .A(_13833_),
    .ZN(_13834_)
  );
  MUX2_X1 _21533_ (
    .A(mem_reg_raw_inst[0]),
    .B(wb_reg_raw_inst[0]),
    .S(_13833_),
    .Z(_00101_)
  );
  MUX2_X1 _21534_ (
    .A(mem_reg_raw_inst[1]),
    .B(wb_reg_raw_inst[1]),
    .S(_13833_),
    .Z(_00102_)
  );
  MUX2_X1 _21535_ (
    .A(mem_reg_raw_inst[2]),
    .B(wb_reg_raw_inst[2]),
    .S(_13833_),
    .Z(_00103_)
  );
  MUX2_X1 _21536_ (
    .A(mem_reg_raw_inst[3]),
    .B(wb_reg_raw_inst[3]),
    .S(_13833_),
    .Z(_00104_)
  );
  MUX2_X1 _21537_ (
    .A(mem_reg_raw_inst[4]),
    .B(wb_reg_raw_inst[4]),
    .S(_13833_),
    .Z(_00105_)
  );
  MUX2_X1 _21538_ (
    .A(mem_reg_raw_inst[5]),
    .B(wb_reg_raw_inst[5]),
    .S(_13833_),
    .Z(_00106_)
  );
  MUX2_X1 _21539_ (
    .A(mem_reg_raw_inst[6]),
    .B(wb_reg_raw_inst[6]),
    .S(_13833_),
    .Z(_00107_)
  );
  MUX2_X1 _21540_ (
    .A(mem_reg_raw_inst[7]),
    .B(wb_reg_raw_inst[7]),
    .S(_13833_),
    .Z(_00108_)
  );
  MUX2_X1 _21541_ (
    .A(mem_reg_raw_inst[8]),
    .B(wb_reg_raw_inst[8]),
    .S(_13833_),
    .Z(_00109_)
  );
  MUX2_X1 _21542_ (
    .A(mem_reg_raw_inst[9]),
    .B(wb_reg_raw_inst[9]),
    .S(_13833_),
    .Z(_00110_)
  );
  MUX2_X1 _21543_ (
    .A(mem_reg_raw_inst[10]),
    .B(wb_reg_raw_inst[10]),
    .S(_13833_),
    .Z(_00111_)
  );
  MUX2_X1 _21544_ (
    .A(mem_reg_raw_inst[11]),
    .B(wb_reg_raw_inst[11]),
    .S(_13833_),
    .Z(_00112_)
  );
  MUX2_X1 _21545_ (
    .A(mem_reg_raw_inst[12]),
    .B(wb_reg_raw_inst[12]),
    .S(_13833_),
    .Z(_00113_)
  );
  MUX2_X1 _21546_ (
    .A(mem_reg_raw_inst[13]),
    .B(wb_reg_raw_inst[13]),
    .S(_13833_),
    .Z(_00114_)
  );
  MUX2_X1 _21547_ (
    .A(mem_reg_raw_inst[14]),
    .B(wb_reg_raw_inst[14]),
    .S(_13833_),
    .Z(_00115_)
  );
  MUX2_X1 _21548_ (
    .A(mem_reg_raw_inst[15]),
    .B(wb_reg_raw_inst[15]),
    .S(_13833_),
    .Z(_00116_)
  );
  MUX2_X1 _21549_ (
    .A(mem_reg_rvc),
    .B(mem_reg_inst[21]),
    .S(mem_ctrl_jal),
    .Z(_13835_)
  );
  MUX2_X1 _21550_ (
    .A(_13835_),
    .B(mem_reg_inst[8]),
    .S(_10066_),
    .Z(_13836_)
  );
  INV_X1 _21551_ (
    .A(_13836_),
    .ZN(_13837_)
  );
  AND2_X1 _21552_ (
    .A1(mem_reg_pc[1]),
    .A2(_13836_),
    .ZN(_13838_)
  );
  INV_X1 _21553_ (
    .A(_13838_),
    .ZN(_13839_)
  );
  AND2_X1 _21554_ (
    .A1(_07985_),
    .A2(_13837_),
    .ZN(_13840_)
  );
  INV_X1 _21555_ (
    .A(_13840_),
    .ZN(_13841_)
  );
  AND2_X1 _21556_ (
    .A1(_13839_),
    .A2(_13841_),
    .ZN(_13842_)
  );
  MUX2_X1 _21557_ (
    .A(mem_reg_wdata[1]),
    .B(_13842_),
    .S(_08206_),
    .Z(_13843_)
  );
  INV_X1 _21558_ (
    .A(_13843_),
    .ZN(_13844_)
  );
  AND2_X1 _21559_ (
    .A1(_08599_),
    .A2(_13843_),
    .ZN(_13845_)
  );
  INV_X1 _21560_ (
    .A(_13845_),
    .ZN(_13846_)
  );
  AND2_X1 _21561_ (
    .A1(mem_ctrl_jalr),
    .A2(_13845_),
    .ZN(_13847_)
  );
  INV_X1 _21562_ (
    .A(_13847_),
    .ZN(_13848_)
  );
  AND2_X1 _21563_ (
    .A1(_08206_),
    .A2(_13846_),
    .ZN(_13849_)
  );
  INV_X1 _21564_ (
    .A(_13849_),
    .ZN(_13850_)
  );
  AND2_X1 _21565_ (
    .A1(_take_pc_mem_T),
    .A2(_13848_),
    .ZN(_13851_)
  );
  AND2_X1 _21566_ (
    .A1(_13850_),
    .A2(_13851_),
    .ZN(_13852_)
  );
  INV_X1 _21567_ (
    .A(_13852_),
    .ZN(_13853_)
  );
  MUX2_X1 _21568_ (
    .A(mem_reg_wdata[0]),
    .B(mem_reg_pc[0]),
    .S(_13852_),
    .Z(_13854_)
  );
  MUX2_X1 _21569_ (
    .A(wb_reg_wdata[0]),
    .B(_13854_),
    .S(_13834_),
    .Z(_00117_)
  );
  MUX2_X1 _21570_ (
    .A(mem_reg_wdata[1]),
    .B(_13842_),
    .S(_13852_),
    .Z(_13855_)
  );
  MUX2_X1 _21571_ (
    .A(wb_reg_wdata[1]),
    .B(_13855_),
    .S(_13834_),
    .Z(_00118_)
  );
  MUX2_X1 _21572_ (
    .A(_mem_br_target_T_6[2]),
    .B(mem_reg_inst[22]),
    .S(mem_ctrl_jal),
    .Z(_13856_)
  );
  MUX2_X1 _21573_ (
    .A(_13856_),
    .B(mem_reg_inst[9]),
    .S(_10066_),
    .Z(_13857_)
  );
  INV_X1 _21574_ (
    .A(_13857_),
    .ZN(_13858_)
  );
  AND2_X1 _21575_ (
    .A1(mem_reg_pc[2]),
    .A2(_13857_),
    .ZN(_13859_)
  );
  INV_X1 _21576_ (
    .A(_13859_),
    .ZN(_13860_)
  );
  AND2_X1 _21577_ (
    .A1(_07986_),
    .A2(_13858_),
    .ZN(_13861_)
  );
  INV_X1 _21578_ (
    .A(_13861_),
    .ZN(_13862_)
  );
  AND2_X1 _21579_ (
    .A1(_13860_),
    .A2(_13862_),
    .ZN(_13863_)
  );
  INV_X1 _21580_ (
    .A(_13863_),
    .ZN(_13864_)
  );
  AND2_X1 _21581_ (
    .A1(_13838_),
    .A2(_13863_),
    .ZN(_13865_)
  );
  INV_X1 _21582_ (
    .A(_13865_),
    .ZN(_13866_)
  );
  AND2_X1 _21583_ (
    .A1(_13839_),
    .A2(_13864_),
    .ZN(_13867_)
  );
  INV_X1 _21584_ (
    .A(_13867_),
    .ZN(_13868_)
  );
  AND2_X1 _21585_ (
    .A1(_13866_),
    .A2(_13868_),
    .ZN(_13869_)
  );
  MUX2_X1 _21586_ (
    .A(mem_reg_wdata[2]),
    .B(_13869_),
    .S(_13852_),
    .Z(_13870_)
  );
  MUX2_X1 _21587_ (
    .A(wb_reg_wdata[2]),
    .B(_13870_),
    .S(_13834_),
    .Z(_00119_)
  );
  AND2_X1 _21588_ (
    .A1(_13860_),
    .A2(_13866_),
    .ZN(_13871_)
  );
  INV_X1 _21589_ (
    .A(_13871_),
    .ZN(_13872_)
  );
  AND2_X1 _21590_ (
    .A1(mem_reg_inst[23]),
    .A2(mem_ctrl_jal),
    .ZN(_13873_)
  );
  MUX2_X1 _21591_ (
    .A(_13873_),
    .B(mem_reg_inst[10]),
    .S(_10066_),
    .Z(_13874_)
  );
  INV_X1 _21592_ (
    .A(_13874_),
    .ZN(_13875_)
  );
  AND2_X1 _21593_ (
    .A1(mem_reg_pc[3]),
    .A2(_13874_),
    .ZN(_13876_)
  );
  INV_X1 _21594_ (
    .A(_13876_),
    .ZN(_13877_)
  );
  AND2_X1 _21595_ (
    .A1(_07987_),
    .A2(_13875_),
    .ZN(_13878_)
  );
  INV_X1 _21596_ (
    .A(_13878_),
    .ZN(_13879_)
  );
  AND2_X1 _21597_ (
    .A1(_13877_),
    .A2(_13879_),
    .ZN(_13880_)
  );
  INV_X1 _21598_ (
    .A(_13880_),
    .ZN(_13881_)
  );
  AND2_X1 _21599_ (
    .A1(_13872_),
    .A2(_13880_),
    .ZN(_13882_)
  );
  INV_X1 _21600_ (
    .A(_13882_),
    .ZN(_13883_)
  );
  AND2_X1 _21601_ (
    .A1(_13871_),
    .A2(_13881_),
    .ZN(_13884_)
  );
  INV_X1 _21602_ (
    .A(_13884_),
    .ZN(_13885_)
  );
  AND2_X1 _21603_ (
    .A1(_13883_),
    .A2(_13885_),
    .ZN(_13886_)
  );
  MUX2_X1 _21604_ (
    .A(mem_reg_wdata[3]),
    .B(_13886_),
    .S(_13852_),
    .Z(_13887_)
  );
  MUX2_X1 _21605_ (
    .A(wb_reg_wdata[3]),
    .B(_13887_),
    .S(_13834_),
    .Z(_00120_)
  );
  AND2_X1 _21606_ (
    .A1(mem_reg_inst[24]),
    .A2(mem_ctrl_jal),
    .ZN(_13888_)
  );
  MUX2_X1 _21607_ (
    .A(_13888_),
    .B(mem_reg_inst[11]),
    .S(_10066_),
    .Z(_13889_)
  );
  INV_X1 _21608_ (
    .A(_13889_),
    .ZN(_13890_)
  );
  AND2_X1 _21609_ (
    .A1(mem_reg_pc[4]),
    .A2(_13889_),
    .ZN(_13891_)
  );
  INV_X1 _21610_ (
    .A(_13891_),
    .ZN(_13892_)
  );
  AND2_X1 _21611_ (
    .A1(_07988_),
    .A2(_13890_),
    .ZN(_13893_)
  );
  INV_X1 _21612_ (
    .A(_13893_),
    .ZN(_13894_)
  );
  AND2_X1 _21613_ (
    .A1(_13892_),
    .A2(_13894_),
    .ZN(_13895_)
  );
  INV_X1 _21614_ (
    .A(_13895_),
    .ZN(_13896_)
  );
  AND2_X1 _21615_ (
    .A1(_13872_),
    .A2(_13879_),
    .ZN(_13897_)
  );
  INV_X1 _21616_ (
    .A(_13897_),
    .ZN(_13898_)
  );
  AND2_X1 _21617_ (
    .A1(_13871_),
    .A2(_13877_),
    .ZN(_13899_)
  );
  INV_X1 _21618_ (
    .A(_13899_),
    .ZN(_13900_)
  );
  AND2_X1 _21619_ (
    .A1(_13877_),
    .A2(_13898_),
    .ZN(_13901_)
  );
  AND2_X1 _21620_ (
    .A1(_13879_),
    .A2(_13900_),
    .ZN(_13902_)
  );
  AND2_X1 _21621_ (
    .A1(_13895_),
    .A2(_13902_),
    .ZN(_13903_)
  );
  INV_X1 _21622_ (
    .A(_13903_),
    .ZN(_13904_)
  );
  AND2_X1 _21623_ (
    .A1(_13896_),
    .A2(_13901_),
    .ZN(_13905_)
  );
  INV_X1 _21624_ (
    .A(_13905_),
    .ZN(_13906_)
  );
  AND2_X1 _21625_ (
    .A1(_13904_),
    .A2(_13906_),
    .ZN(_13907_)
  );
  MUX2_X1 _21626_ (
    .A(mem_reg_wdata[4]),
    .B(_13907_),
    .S(_13852_),
    .Z(_13908_)
  );
  MUX2_X1 _21627_ (
    .A(wb_reg_wdata[4]),
    .B(_13908_),
    .S(_13834_),
    .Z(_00121_)
  );
  AND2_X1 _21628_ (
    .A1(wb_reg_wdata[5]),
    .A2(_13833_),
    .ZN(_13909_)
  );
  INV_X1 _21629_ (
    .A(_13909_),
    .ZN(_13910_)
  );
  AND2_X1 _21630_ (
    .A1(_13892_),
    .A2(_13904_),
    .ZN(_13911_)
  );
  INV_X1 _21631_ (
    .A(_13911_),
    .ZN(_13912_)
  );
  AND2_X1 _21632_ (
    .A1(mem_reg_inst[25]),
    .A2(_10069_),
    .ZN(_13913_)
  );
  INV_X1 _21633_ (
    .A(_13913_),
    .ZN(_13914_)
  );
  AND2_X1 _21634_ (
    .A1(mem_reg_pc[5]),
    .A2(_13913_),
    .ZN(_13915_)
  );
  INV_X1 _21635_ (
    .A(_13915_),
    .ZN(_13916_)
  );
  AND2_X1 _21636_ (
    .A1(_07990_),
    .A2(_13914_),
    .ZN(_13917_)
  );
  INV_X1 _21637_ (
    .A(_13917_),
    .ZN(_13918_)
  );
  AND2_X1 _21638_ (
    .A1(_13916_),
    .A2(_13918_),
    .ZN(_13919_)
  );
  INV_X1 _21639_ (
    .A(_13919_),
    .ZN(_13920_)
  );
  AND2_X1 _21640_ (
    .A1(_13912_),
    .A2(_13919_),
    .ZN(_13921_)
  );
  INV_X1 _21641_ (
    .A(_13921_),
    .ZN(_13922_)
  );
  AND2_X1 _21642_ (
    .A1(_13911_),
    .A2(_13920_),
    .ZN(_13923_)
  );
  INV_X1 _21643_ (
    .A(_13923_),
    .ZN(_13924_)
  );
  AND2_X1 _21644_ (
    .A1(_13922_),
    .A2(_13924_),
    .ZN(_13925_)
  );
  INV_X1 _21645_ (
    .A(_13925_),
    .ZN(_13926_)
  );
  AND2_X1 _21646_ (
    .A1(_13852_),
    .A2(_13926_),
    .ZN(_13927_)
  );
  INV_X1 _21647_ (
    .A(_13927_),
    .ZN(_13928_)
  );
  AND2_X1 _21648_ (
    .A1(_08057_),
    .A2(_13853_),
    .ZN(_13929_)
  );
  INV_X1 _21649_ (
    .A(_13929_),
    .ZN(_13930_)
  );
  AND2_X1 _21650_ (
    .A1(_13834_),
    .A2(_13930_),
    .ZN(_13931_)
  );
  AND2_X1 _21651_ (
    .A1(_13928_),
    .A2(_13931_),
    .ZN(_13932_)
  );
  INV_X1 _21652_ (
    .A(_13932_),
    .ZN(_13933_)
  );
  AND2_X1 _21653_ (
    .A1(_13910_),
    .A2(_13933_),
    .ZN(_13934_)
  );
  INV_X1 _21654_ (
    .A(_13934_),
    .ZN(_00122_)
  );
  AND2_X1 _21655_ (
    .A1(wb_reg_wdata[6]),
    .A2(_13833_),
    .ZN(_13935_)
  );
  INV_X1 _21656_ (
    .A(_13935_),
    .ZN(_13936_)
  );
  AND2_X1 _21657_ (
    .A1(_13916_),
    .A2(_13922_),
    .ZN(_13937_)
  );
  INV_X1 _21658_ (
    .A(_13937_),
    .ZN(_13938_)
  );
  AND2_X1 _21659_ (
    .A1(mem_reg_inst[26]),
    .A2(_10069_),
    .ZN(_13939_)
  );
  INV_X1 _21660_ (
    .A(_13939_),
    .ZN(_13940_)
  );
  AND2_X1 _21661_ (
    .A1(mem_reg_pc[6]),
    .A2(_13939_),
    .ZN(_13941_)
  );
  INV_X1 _21662_ (
    .A(_13941_),
    .ZN(_13942_)
  );
  AND2_X1 _21663_ (
    .A1(_07992_),
    .A2(_13940_),
    .ZN(_13943_)
  );
  INV_X1 _21664_ (
    .A(_13943_),
    .ZN(_13944_)
  );
  AND2_X1 _21665_ (
    .A1(_13942_),
    .A2(_13944_),
    .ZN(_13945_)
  );
  INV_X1 _21666_ (
    .A(_13945_),
    .ZN(_13946_)
  );
  AND2_X1 _21667_ (
    .A1(_13938_),
    .A2(_13945_),
    .ZN(_13947_)
  );
  INV_X1 _21668_ (
    .A(_13947_),
    .ZN(_13948_)
  );
  AND2_X1 _21669_ (
    .A1(_13937_),
    .A2(_13946_),
    .ZN(_13949_)
  );
  INV_X1 _21670_ (
    .A(_13949_),
    .ZN(_13950_)
  );
  AND2_X1 _21671_ (
    .A1(_13948_),
    .A2(_13950_),
    .ZN(_13951_)
  );
  INV_X1 _21672_ (
    .A(_13951_),
    .ZN(_13952_)
  );
  AND2_X1 _21673_ (
    .A1(_13852_),
    .A2(_13952_),
    .ZN(_13953_)
  );
  INV_X1 _21674_ (
    .A(_13953_),
    .ZN(_13954_)
  );
  AND2_X1 _21675_ (
    .A1(_08058_),
    .A2(_13853_),
    .ZN(_13955_)
  );
  INV_X1 _21676_ (
    .A(_13955_),
    .ZN(_13956_)
  );
  AND2_X1 _21677_ (
    .A1(_13834_),
    .A2(_13956_),
    .ZN(_13957_)
  );
  AND2_X1 _21678_ (
    .A1(_13954_),
    .A2(_13957_),
    .ZN(_13958_)
  );
  INV_X1 _21679_ (
    .A(_13958_),
    .ZN(_13959_)
  );
  AND2_X1 _21680_ (
    .A1(_13936_),
    .A2(_13959_),
    .ZN(_13960_)
  );
  INV_X1 _21681_ (
    .A(_13960_),
    .ZN(_00123_)
  );
  AND2_X1 _21682_ (
    .A1(wb_reg_wdata[7]),
    .A2(_13833_),
    .ZN(_13961_)
  );
  INV_X1 _21683_ (
    .A(_13961_),
    .ZN(_13962_)
  );
  AND2_X1 _21684_ (
    .A1(_13942_),
    .A2(_13948_),
    .ZN(_13963_)
  );
  INV_X1 _21685_ (
    .A(_13963_),
    .ZN(_13964_)
  );
  AND2_X1 _21686_ (
    .A1(mem_reg_inst[27]),
    .A2(_10069_),
    .ZN(_13965_)
  );
  INV_X1 _21687_ (
    .A(_13965_),
    .ZN(_13966_)
  );
  AND2_X1 _21688_ (
    .A1(mem_reg_pc[7]),
    .A2(_13965_),
    .ZN(_13967_)
  );
  INV_X1 _21689_ (
    .A(_13967_),
    .ZN(_13968_)
  );
  AND2_X1 _21690_ (
    .A1(_07994_),
    .A2(_13966_),
    .ZN(_13969_)
  );
  INV_X1 _21691_ (
    .A(_13969_),
    .ZN(_13970_)
  );
  AND2_X1 _21692_ (
    .A1(_13968_),
    .A2(_13970_),
    .ZN(_13971_)
  );
  INV_X1 _21693_ (
    .A(_13971_),
    .ZN(_13972_)
  );
  AND2_X1 _21694_ (
    .A1(_13964_),
    .A2(_13972_),
    .ZN(_13973_)
  );
  INV_X1 _21695_ (
    .A(_13973_),
    .ZN(_13974_)
  );
  AND2_X1 _21696_ (
    .A1(_13963_),
    .A2(_13971_),
    .ZN(_13975_)
  );
  INV_X1 _21697_ (
    .A(_13975_),
    .ZN(_13976_)
  );
  AND2_X1 _21698_ (
    .A1(_13974_),
    .A2(_13976_),
    .ZN(_13977_)
  );
  AND2_X1 _21699_ (
    .A1(_13852_),
    .A2(_13977_),
    .ZN(_13978_)
  );
  INV_X1 _21700_ (
    .A(_13978_),
    .ZN(_13979_)
  );
  AND2_X1 _21701_ (
    .A1(_08059_),
    .A2(_13853_),
    .ZN(_13980_)
  );
  INV_X1 _21702_ (
    .A(_13980_),
    .ZN(_13981_)
  );
  AND2_X1 _21703_ (
    .A1(_13834_),
    .A2(_13981_),
    .ZN(_13982_)
  );
  AND2_X1 _21704_ (
    .A1(_13979_),
    .A2(_13982_),
    .ZN(_13983_)
  );
  INV_X1 _21705_ (
    .A(_13983_),
    .ZN(_13984_)
  );
  AND2_X1 _21706_ (
    .A1(_13962_),
    .A2(_13984_),
    .ZN(_13985_)
  );
  INV_X1 _21707_ (
    .A(_13985_),
    .ZN(_00124_)
  );
  AND2_X1 _21708_ (
    .A1(mem_reg_inst[28]),
    .A2(_10069_),
    .ZN(_13986_)
  );
  INV_X1 _21709_ (
    .A(_13986_),
    .ZN(_13987_)
  );
  AND2_X1 _21710_ (
    .A1(mem_reg_pc[8]),
    .A2(_13986_),
    .ZN(_13988_)
  );
  INV_X1 _21711_ (
    .A(_13988_),
    .ZN(_13989_)
  );
  AND2_X1 _21712_ (
    .A1(_07996_),
    .A2(_13987_),
    .ZN(_13990_)
  );
  INV_X1 _21713_ (
    .A(_13990_),
    .ZN(_13991_)
  );
  AND2_X1 _21714_ (
    .A1(_13989_),
    .A2(_13991_),
    .ZN(_13992_)
  );
  INV_X1 _21715_ (
    .A(_13992_),
    .ZN(_13993_)
  );
  AND2_X1 _21716_ (
    .A1(_13963_),
    .A2(_13968_),
    .ZN(_13994_)
  );
  INV_X1 _21717_ (
    .A(_13994_),
    .ZN(_13995_)
  );
  AND2_X1 _21718_ (
    .A1(_13964_),
    .A2(_13970_),
    .ZN(_13996_)
  );
  INV_X1 _21719_ (
    .A(_13996_),
    .ZN(_13997_)
  );
  AND2_X1 _21720_ (
    .A1(_13970_),
    .A2(_13995_),
    .ZN(_13998_)
  );
  AND2_X1 _21721_ (
    .A1(_13968_),
    .A2(_13997_),
    .ZN(_13999_)
  );
  AND2_X1 _21722_ (
    .A1(_13992_),
    .A2(_13998_),
    .ZN(_14000_)
  );
  INV_X1 _21723_ (
    .A(_14000_),
    .ZN(_14001_)
  );
  AND2_X1 _21724_ (
    .A1(_13993_),
    .A2(_13999_),
    .ZN(_14002_)
  );
  INV_X1 _21725_ (
    .A(_14002_),
    .ZN(_14003_)
  );
  AND2_X1 _21726_ (
    .A1(_14001_),
    .A2(_14003_),
    .ZN(_14004_)
  );
  INV_X1 _21727_ (
    .A(_14004_),
    .ZN(_14005_)
  );
  MUX2_X1 _21728_ (
    .A(mem_reg_wdata[8]),
    .B(_14004_),
    .S(_13852_),
    .Z(_14006_)
  );
  MUX2_X1 _21729_ (
    .A(wb_reg_wdata[8]),
    .B(_14006_),
    .S(_13834_),
    .Z(_00125_)
  );
  AND2_X1 _21730_ (
    .A1(wb_reg_wdata[9]),
    .A2(_13833_),
    .ZN(_14007_)
  );
  INV_X1 _21731_ (
    .A(_14007_),
    .ZN(_14008_)
  );
  AND2_X1 _21732_ (
    .A1(_13989_),
    .A2(_14001_),
    .ZN(_14009_)
  );
  INV_X1 _21733_ (
    .A(_14009_),
    .ZN(_14010_)
  );
  AND2_X1 _21734_ (
    .A1(mem_reg_inst[29]),
    .A2(_10069_),
    .ZN(_14011_)
  );
  INV_X1 _21735_ (
    .A(_14011_),
    .ZN(_14012_)
  );
  AND2_X1 _21736_ (
    .A1(mem_reg_pc[9]),
    .A2(_14011_),
    .ZN(_14013_)
  );
  INV_X1 _21737_ (
    .A(_14013_),
    .ZN(_14014_)
  );
  AND2_X1 _21738_ (
    .A1(_07998_),
    .A2(_14012_),
    .ZN(_14015_)
  );
  INV_X1 _21739_ (
    .A(_14015_),
    .ZN(_14016_)
  );
  AND2_X1 _21740_ (
    .A1(_14014_),
    .A2(_14016_),
    .ZN(_14017_)
  );
  INV_X1 _21741_ (
    .A(_14017_),
    .ZN(_14018_)
  );
  AND2_X1 _21742_ (
    .A1(_14010_),
    .A2(_14018_),
    .ZN(_14019_)
  );
  INV_X1 _21743_ (
    .A(_14019_),
    .ZN(_14020_)
  );
  AND2_X1 _21744_ (
    .A1(_14009_),
    .A2(_14017_),
    .ZN(_14021_)
  );
  INV_X1 _21745_ (
    .A(_14021_),
    .ZN(_14022_)
  );
  AND2_X1 _21746_ (
    .A1(_14020_),
    .A2(_14022_),
    .ZN(_14023_)
  );
  AND2_X1 _21747_ (
    .A1(_13852_),
    .A2(_14023_),
    .ZN(_14024_)
  );
  INV_X1 _21748_ (
    .A(_14024_),
    .ZN(_14025_)
  );
  AND2_X1 _21749_ (
    .A1(_08061_),
    .A2(_13853_),
    .ZN(_14026_)
  );
  INV_X1 _21750_ (
    .A(_14026_),
    .ZN(_01588_)
  );
  AND2_X1 _21751_ (
    .A1(_13834_),
    .A2(_01588_),
    .ZN(_01589_)
  );
  AND2_X1 _21752_ (
    .A1(_14025_),
    .A2(_01589_),
    .ZN(_01590_)
  );
  INV_X1 _21753_ (
    .A(_01590_),
    .ZN(_01591_)
  );
  AND2_X1 _21754_ (
    .A1(_14008_),
    .A2(_01591_),
    .ZN(_01592_)
  );
  INV_X1 _21755_ (
    .A(_01592_),
    .ZN(_00126_)
  );
  AND2_X1 _21756_ (
    .A1(wb_reg_wdata[10]),
    .A2(_13833_),
    .ZN(_01593_)
  );
  INV_X1 _21757_ (
    .A(_01593_),
    .ZN(_01594_)
  );
  AND2_X1 _21758_ (
    .A1(mem_reg_inst[30]),
    .A2(_10069_),
    .ZN(_01595_)
  );
  INV_X1 _21759_ (
    .A(_01595_),
    .ZN(_01596_)
  );
  AND2_X1 _21760_ (
    .A1(mem_reg_pc[10]),
    .A2(_01595_),
    .ZN(_01597_)
  );
  INV_X1 _21761_ (
    .A(_01597_),
    .ZN(_01598_)
  );
  AND2_X1 _21762_ (
    .A1(_08000_),
    .A2(_01596_),
    .ZN(_01599_)
  );
  INV_X1 _21763_ (
    .A(_01599_),
    .ZN(_01600_)
  );
  AND2_X1 _21764_ (
    .A1(_01598_),
    .A2(_01600_),
    .ZN(_01601_)
  );
  INV_X1 _21765_ (
    .A(_01601_),
    .ZN(_01602_)
  );
  AND2_X1 _21766_ (
    .A1(_14009_),
    .A2(_14014_),
    .ZN(_01603_)
  );
  INV_X1 _21767_ (
    .A(_01603_),
    .ZN(_01604_)
  );
  AND2_X1 _21768_ (
    .A1(_14010_),
    .A2(_14016_),
    .ZN(_01605_)
  );
  INV_X1 _21769_ (
    .A(_01605_),
    .ZN(_01606_)
  );
  AND2_X1 _21770_ (
    .A1(_14016_),
    .A2(_01604_),
    .ZN(_01607_)
  );
  AND2_X1 _21771_ (
    .A1(_14014_),
    .A2(_01606_),
    .ZN(_01608_)
  );
  AND2_X1 _21772_ (
    .A1(_01601_),
    .A2(_01607_),
    .ZN(_01609_)
  );
  INV_X1 _21773_ (
    .A(_01609_),
    .ZN(_01610_)
  );
  AND2_X1 _21774_ (
    .A1(_01602_),
    .A2(_01608_),
    .ZN(_01611_)
  );
  INV_X1 _21775_ (
    .A(_01611_),
    .ZN(_01612_)
  );
  AND2_X1 _21776_ (
    .A1(_01610_),
    .A2(_01612_),
    .ZN(_01613_)
  );
  INV_X1 _21777_ (
    .A(_01613_),
    .ZN(_01614_)
  );
  AND2_X1 _21778_ (
    .A1(_13852_),
    .A2(_01614_),
    .ZN(_01615_)
  );
  INV_X1 _21779_ (
    .A(_01615_),
    .ZN(_01616_)
  );
  AND2_X1 _21780_ (
    .A1(_08062_),
    .A2(_13853_),
    .ZN(_01617_)
  );
  INV_X1 _21781_ (
    .A(_01617_),
    .ZN(_01618_)
  );
  AND2_X1 _21782_ (
    .A1(_13834_),
    .A2(_01618_),
    .ZN(_01619_)
  );
  AND2_X1 _21783_ (
    .A1(_01616_),
    .A2(_01619_),
    .ZN(_01620_)
  );
  INV_X1 _21784_ (
    .A(_01620_),
    .ZN(_01621_)
  );
  AND2_X1 _21785_ (
    .A1(_01594_),
    .A2(_01621_),
    .ZN(_01622_)
  );
  INV_X1 _21786_ (
    .A(_01622_),
    .ZN(_00127_)
  );
  AND2_X1 _21787_ (
    .A1(wb_reg_wdata[11]),
    .A2(_13833_),
    .ZN(_01623_)
  );
  INV_X1 _21788_ (
    .A(_01623_),
    .ZN(_01624_)
  );
  AND2_X1 _21789_ (
    .A1(_01598_),
    .A2(_01610_),
    .ZN(_01625_)
  );
  INV_X1 _21790_ (
    .A(_01625_),
    .ZN(_01626_)
  );
  AND2_X1 _21791_ (
    .A1(mem_reg_inst[20]),
    .A2(mem_ctrl_jal),
    .ZN(_01627_)
  );
  MUX2_X1 _21792_ (
    .A(_01627_),
    .B(mem_reg_inst[7]),
    .S(_10066_),
    .Z(_01628_)
  );
  INV_X1 _21793_ (
    .A(_01628_),
    .ZN(_01629_)
  );
  AND2_X1 _21794_ (
    .A1(mem_reg_pc[11]),
    .A2(_01628_),
    .ZN(_01630_)
  );
  INV_X1 _21795_ (
    .A(_01630_),
    .ZN(_01631_)
  );
  AND2_X1 _21796_ (
    .A1(_08002_),
    .A2(_01629_),
    .ZN(_01632_)
  );
  INV_X1 _21797_ (
    .A(_01632_),
    .ZN(_01633_)
  );
  AND2_X1 _21798_ (
    .A1(_01631_),
    .A2(_01633_),
    .ZN(_01634_)
  );
  INV_X1 _21799_ (
    .A(_01634_),
    .ZN(_01635_)
  );
  AND2_X1 _21800_ (
    .A1(_01626_),
    .A2(_01635_),
    .ZN(_01636_)
  );
  INV_X1 _21801_ (
    .A(_01636_),
    .ZN(_01637_)
  );
  AND2_X1 _21802_ (
    .A1(_01625_),
    .A2(_01634_),
    .ZN(_01638_)
  );
  INV_X1 _21803_ (
    .A(_01638_),
    .ZN(_01639_)
  );
  AND2_X1 _21804_ (
    .A1(_01637_),
    .A2(_01639_),
    .ZN(_01640_)
  );
  AND2_X1 _21805_ (
    .A1(_13852_),
    .A2(_01640_),
    .ZN(_01641_)
  );
  INV_X1 _21806_ (
    .A(_01641_),
    .ZN(_01642_)
  );
  AND2_X1 _21807_ (
    .A1(_08063_),
    .A2(_13853_),
    .ZN(_01643_)
  );
  INV_X1 _21808_ (
    .A(_01643_),
    .ZN(_01644_)
  );
  AND2_X1 _21809_ (
    .A1(_13834_),
    .A2(_01644_),
    .ZN(_01645_)
  );
  AND2_X1 _21810_ (
    .A1(_01642_),
    .A2(_01645_),
    .ZN(_01646_)
  );
  INV_X1 _21811_ (
    .A(_01646_),
    .ZN(_01647_)
  );
  AND2_X1 _21812_ (
    .A1(_01624_),
    .A2(_01647_),
    .ZN(_01648_)
  );
  INV_X1 _21813_ (
    .A(_01648_),
    .ZN(_00128_)
  );
  AND2_X1 _21814_ (
    .A1(wb_reg_wdata[12]),
    .A2(_13833_),
    .ZN(_01649_)
  );
  INV_X1 _21815_ (
    .A(_01649_),
    .ZN(_01650_)
  );
  AND2_X1 _21816_ (
    .A1(mem_reg_inst[12]),
    .A2(mem_ctrl_jal),
    .ZN(_01651_)
  );
  MUX2_X1 _21817_ (
    .A(_01651_),
    .B(mem_reg_inst[31]),
    .S(_10066_),
    .Z(_01652_)
  );
  INV_X1 _21818_ (
    .A(_01652_),
    .ZN(_01653_)
  );
  AND2_X1 _21819_ (
    .A1(mem_reg_pc[12]),
    .A2(_01652_),
    .ZN(_01654_)
  );
  INV_X1 _21820_ (
    .A(_01654_),
    .ZN(_01655_)
  );
  AND2_X1 _21821_ (
    .A1(_08004_),
    .A2(_01653_),
    .ZN(_01656_)
  );
  INV_X1 _21822_ (
    .A(_01656_),
    .ZN(_01657_)
  );
  AND2_X1 _21823_ (
    .A1(_01655_),
    .A2(_01657_),
    .ZN(_01658_)
  );
  INV_X1 _21824_ (
    .A(_01658_),
    .ZN(_01659_)
  );
  AND2_X1 _21825_ (
    .A1(_01625_),
    .A2(_01631_),
    .ZN(_01660_)
  );
  INV_X1 _21826_ (
    .A(_01660_),
    .ZN(_01661_)
  );
  AND2_X1 _21827_ (
    .A1(_01626_),
    .A2(_01633_),
    .ZN(_01662_)
  );
  INV_X1 _21828_ (
    .A(_01662_),
    .ZN(_01663_)
  );
  AND2_X1 _21829_ (
    .A1(_01633_),
    .A2(_01661_),
    .ZN(_01664_)
  );
  AND2_X1 _21830_ (
    .A1(_01631_),
    .A2(_01663_),
    .ZN(_01665_)
  );
  AND2_X1 _21831_ (
    .A1(_01658_),
    .A2(_01664_),
    .ZN(_01666_)
  );
  INV_X1 _21832_ (
    .A(_01666_),
    .ZN(_01667_)
  );
  AND2_X1 _21833_ (
    .A1(_01659_),
    .A2(_01665_),
    .ZN(_01668_)
  );
  INV_X1 _21834_ (
    .A(_01668_),
    .ZN(_01669_)
  );
  AND2_X1 _21835_ (
    .A1(_01667_),
    .A2(_01669_),
    .ZN(_01670_)
  );
  INV_X1 _21836_ (
    .A(_01670_),
    .ZN(_01671_)
  );
  AND2_X1 _21837_ (
    .A1(_13852_),
    .A2(_01671_),
    .ZN(_01672_)
  );
  INV_X1 _21838_ (
    .A(_01672_),
    .ZN(_01673_)
  );
  AND2_X1 _21839_ (
    .A1(_08064_),
    .A2(_13853_),
    .ZN(_01674_)
  );
  INV_X1 _21840_ (
    .A(_01674_),
    .ZN(_01675_)
  );
  AND2_X1 _21841_ (
    .A1(_13834_),
    .A2(_01675_),
    .ZN(_01676_)
  );
  AND2_X1 _21842_ (
    .A1(_01673_),
    .A2(_01676_),
    .ZN(_01677_)
  );
  INV_X1 _21843_ (
    .A(_01677_),
    .ZN(_01678_)
  );
  AND2_X1 _21844_ (
    .A1(_01650_),
    .A2(_01678_),
    .ZN(_01679_)
  );
  INV_X1 _21845_ (
    .A(_01679_),
    .ZN(_00129_)
  );
  AND2_X1 _21846_ (
    .A1(wb_reg_wdata[13]),
    .A2(_13833_),
    .ZN(_01680_)
  );
  INV_X1 _21847_ (
    .A(_01680_),
    .ZN(_01681_)
  );
  AND2_X1 _21848_ (
    .A1(_01655_),
    .A2(_01667_),
    .ZN(_01682_)
  );
  INV_X1 _21849_ (
    .A(_01682_),
    .ZN(_01683_)
  );
  AND2_X1 _21850_ (
    .A1(mem_reg_inst[13]),
    .A2(mem_ctrl_jal),
    .ZN(_01684_)
  );
  MUX2_X1 _21851_ (
    .A(_01684_),
    .B(mem_reg_inst[31]),
    .S(_10066_),
    .Z(_01685_)
  );
  INV_X1 _21852_ (
    .A(_01685_),
    .ZN(_01686_)
  );
  AND2_X1 _21853_ (
    .A1(mem_reg_pc[13]),
    .A2(_01685_),
    .ZN(_01687_)
  );
  INV_X1 _21854_ (
    .A(_01687_),
    .ZN(_01688_)
  );
  AND2_X1 _21855_ (
    .A1(_08006_),
    .A2(_01686_),
    .ZN(_01689_)
  );
  INV_X1 _21856_ (
    .A(_01689_),
    .ZN(_01690_)
  );
  AND2_X1 _21857_ (
    .A1(_01688_),
    .A2(_01690_),
    .ZN(_01691_)
  );
  INV_X1 _21858_ (
    .A(_01691_),
    .ZN(_01692_)
  );
  AND2_X1 _21859_ (
    .A1(_01683_),
    .A2(_01692_),
    .ZN(_01693_)
  );
  INV_X1 _21860_ (
    .A(_01693_),
    .ZN(_01694_)
  );
  AND2_X1 _21861_ (
    .A1(_01682_),
    .A2(_01691_),
    .ZN(_01695_)
  );
  INV_X1 _21862_ (
    .A(_01695_),
    .ZN(_01696_)
  );
  AND2_X1 _21863_ (
    .A1(_01694_),
    .A2(_01696_),
    .ZN(_01697_)
  );
  AND2_X1 _21864_ (
    .A1(_13852_),
    .A2(_01697_),
    .ZN(_01698_)
  );
  INV_X1 _21865_ (
    .A(_01698_),
    .ZN(_01699_)
  );
  AND2_X1 _21866_ (
    .A1(_08065_),
    .A2(_13853_),
    .ZN(_01700_)
  );
  INV_X1 _21867_ (
    .A(_01700_),
    .ZN(_01701_)
  );
  AND2_X1 _21868_ (
    .A1(_13834_),
    .A2(_01701_),
    .ZN(_01702_)
  );
  AND2_X1 _21869_ (
    .A1(_01699_),
    .A2(_01702_),
    .ZN(_01703_)
  );
  INV_X1 _21870_ (
    .A(_01703_),
    .ZN(_01704_)
  );
  AND2_X1 _21871_ (
    .A1(_01681_),
    .A2(_01704_),
    .ZN(_01705_)
  );
  INV_X1 _21872_ (
    .A(_01705_),
    .ZN(_00130_)
  );
  AND2_X1 _21873_ (
    .A1(wb_reg_wdata[14]),
    .A2(_13833_),
    .ZN(_01706_)
  );
  INV_X1 _21874_ (
    .A(_01706_),
    .ZN(_01707_)
  );
  AND2_X1 _21875_ (
    .A1(mem_reg_inst[14]),
    .A2(mem_ctrl_jal),
    .ZN(_01708_)
  );
  MUX2_X1 _21876_ (
    .A(_01708_),
    .B(mem_reg_inst[31]),
    .S(_10066_),
    .Z(_01709_)
  );
  INV_X1 _21877_ (
    .A(_01709_),
    .ZN(_01710_)
  );
  AND2_X1 _21878_ (
    .A1(mem_reg_pc[14]),
    .A2(_01709_),
    .ZN(_01711_)
  );
  INV_X1 _21879_ (
    .A(_01711_),
    .ZN(_01712_)
  );
  AND2_X1 _21880_ (
    .A1(_08008_),
    .A2(_01710_),
    .ZN(_01713_)
  );
  INV_X1 _21881_ (
    .A(_01713_),
    .ZN(_01714_)
  );
  AND2_X1 _21882_ (
    .A1(_01712_),
    .A2(_01714_),
    .ZN(_01715_)
  );
  INV_X1 _21883_ (
    .A(_01715_),
    .ZN(_01716_)
  );
  AND2_X1 _21884_ (
    .A1(_01682_),
    .A2(_01688_),
    .ZN(_01717_)
  );
  INV_X1 _21885_ (
    .A(_01717_),
    .ZN(_01718_)
  );
  AND2_X1 _21886_ (
    .A1(_01683_),
    .A2(_01690_),
    .ZN(_01719_)
  );
  INV_X1 _21887_ (
    .A(_01719_),
    .ZN(_01720_)
  );
  AND2_X1 _21888_ (
    .A1(_01690_),
    .A2(_01718_),
    .ZN(_01721_)
  );
  AND2_X1 _21889_ (
    .A1(_01688_),
    .A2(_01720_),
    .ZN(_01722_)
  );
  AND2_X1 _21890_ (
    .A1(_01715_),
    .A2(_01721_),
    .ZN(_01723_)
  );
  INV_X1 _21891_ (
    .A(_01723_),
    .ZN(_01724_)
  );
  AND2_X1 _21892_ (
    .A1(_01716_),
    .A2(_01722_),
    .ZN(_01725_)
  );
  INV_X1 _21893_ (
    .A(_01725_),
    .ZN(_01726_)
  );
  AND2_X1 _21894_ (
    .A1(_01724_),
    .A2(_01726_),
    .ZN(_01727_)
  );
  INV_X1 _21895_ (
    .A(_01727_),
    .ZN(_01728_)
  );
  AND2_X1 _21896_ (
    .A1(_13852_),
    .A2(_01728_),
    .ZN(_01729_)
  );
  INV_X1 _21897_ (
    .A(_01729_),
    .ZN(_01730_)
  );
  AND2_X1 _21898_ (
    .A1(_08066_),
    .A2(_13853_),
    .ZN(_01731_)
  );
  INV_X1 _21899_ (
    .A(_01731_),
    .ZN(_01732_)
  );
  AND2_X1 _21900_ (
    .A1(_13834_),
    .A2(_01732_),
    .ZN(_01733_)
  );
  AND2_X1 _21901_ (
    .A1(_01730_),
    .A2(_01733_),
    .ZN(_01734_)
  );
  INV_X1 _21902_ (
    .A(_01734_),
    .ZN(_01735_)
  );
  AND2_X1 _21903_ (
    .A1(_01707_),
    .A2(_01735_),
    .ZN(_01736_)
  );
  INV_X1 _21904_ (
    .A(_01736_),
    .ZN(_00131_)
  );
  AND2_X1 _21905_ (
    .A1(wb_reg_wdata[15]),
    .A2(_13833_),
    .ZN(_01737_)
  );
  INV_X1 _21906_ (
    .A(_01737_),
    .ZN(_01738_)
  );
  AND2_X1 _21907_ (
    .A1(_01712_),
    .A2(_01724_),
    .ZN(_01739_)
  );
  INV_X1 _21908_ (
    .A(_01739_),
    .ZN(_01740_)
  );
  AND2_X1 _21909_ (
    .A1(mem_reg_inst[15]),
    .A2(mem_ctrl_jal),
    .ZN(_01741_)
  );
  MUX2_X1 _21910_ (
    .A(_01741_),
    .B(mem_reg_inst[31]),
    .S(_10066_),
    .Z(_01742_)
  );
  INV_X1 _21911_ (
    .A(_01742_),
    .ZN(_01743_)
  );
  AND2_X1 _21912_ (
    .A1(mem_reg_pc[15]),
    .A2(_01742_),
    .ZN(_01744_)
  );
  INV_X1 _21913_ (
    .A(_01744_),
    .ZN(_01745_)
  );
  AND2_X1 _21914_ (
    .A1(_08010_),
    .A2(_01743_),
    .ZN(_01746_)
  );
  INV_X1 _21915_ (
    .A(_01746_),
    .ZN(_01747_)
  );
  AND2_X1 _21916_ (
    .A1(_01745_),
    .A2(_01747_),
    .ZN(_01748_)
  );
  INV_X1 _21917_ (
    .A(_01748_),
    .ZN(_01749_)
  );
  AND2_X1 _21918_ (
    .A1(_01740_),
    .A2(_01749_),
    .ZN(_01750_)
  );
  INV_X1 _21919_ (
    .A(_01750_),
    .ZN(_01751_)
  );
  AND2_X1 _21920_ (
    .A1(_01739_),
    .A2(_01748_),
    .ZN(_01752_)
  );
  INV_X1 _21921_ (
    .A(_01752_),
    .ZN(_01753_)
  );
  AND2_X1 _21922_ (
    .A1(_01751_),
    .A2(_01753_),
    .ZN(_01754_)
  );
  AND2_X1 _21923_ (
    .A1(_13852_),
    .A2(_01754_),
    .ZN(_01755_)
  );
  INV_X1 _21924_ (
    .A(_01755_),
    .ZN(_01756_)
  );
  AND2_X1 _21925_ (
    .A1(_08067_),
    .A2(_13853_),
    .ZN(_01757_)
  );
  INV_X1 _21926_ (
    .A(_01757_),
    .ZN(_01758_)
  );
  AND2_X1 _21927_ (
    .A1(_13834_),
    .A2(_01758_),
    .ZN(_01759_)
  );
  AND2_X1 _21928_ (
    .A1(_01756_),
    .A2(_01759_),
    .ZN(_01760_)
  );
  INV_X1 _21929_ (
    .A(_01760_),
    .ZN(_01761_)
  );
  AND2_X1 _21930_ (
    .A1(_01738_),
    .A2(_01761_),
    .ZN(_01762_)
  );
  INV_X1 _21931_ (
    .A(_01762_),
    .ZN(_00132_)
  );
  AND2_X1 _21932_ (
    .A1(wb_reg_wdata[16]),
    .A2(_13833_),
    .ZN(_01763_)
  );
  INV_X1 _21933_ (
    .A(_01763_),
    .ZN(_01764_)
  );
  AND2_X1 _21934_ (
    .A1(mem_reg_inst[16]),
    .A2(mem_ctrl_jal),
    .ZN(_01765_)
  );
  MUX2_X1 _21935_ (
    .A(_01765_),
    .B(mem_reg_inst[31]),
    .S(_10066_),
    .Z(_01766_)
  );
  INV_X1 _21936_ (
    .A(_01766_),
    .ZN(_01767_)
  );
  AND2_X1 _21937_ (
    .A1(mem_reg_pc[16]),
    .A2(_01766_),
    .ZN(_01768_)
  );
  INV_X1 _21938_ (
    .A(_01768_),
    .ZN(_01769_)
  );
  AND2_X1 _21939_ (
    .A1(_08012_),
    .A2(_01767_),
    .ZN(_01770_)
  );
  INV_X1 _21940_ (
    .A(_01770_),
    .ZN(_01771_)
  );
  AND2_X1 _21941_ (
    .A1(_01769_),
    .A2(_01771_),
    .ZN(_01772_)
  );
  INV_X1 _21942_ (
    .A(_01772_),
    .ZN(_01773_)
  );
  AND2_X1 _21943_ (
    .A1(_01739_),
    .A2(_01745_),
    .ZN(_01774_)
  );
  INV_X1 _21944_ (
    .A(_01774_),
    .ZN(_01775_)
  );
  AND2_X1 _21945_ (
    .A1(_01740_),
    .A2(_01747_),
    .ZN(_01776_)
  );
  INV_X1 _21946_ (
    .A(_01776_),
    .ZN(_01777_)
  );
  AND2_X1 _21947_ (
    .A1(_01747_),
    .A2(_01775_),
    .ZN(_01778_)
  );
  AND2_X1 _21948_ (
    .A1(_01745_),
    .A2(_01777_),
    .ZN(_01779_)
  );
  AND2_X1 _21949_ (
    .A1(_01772_),
    .A2(_01778_),
    .ZN(_01780_)
  );
  INV_X1 _21950_ (
    .A(_01780_),
    .ZN(_01781_)
  );
  AND2_X1 _21951_ (
    .A1(_01773_),
    .A2(_01779_),
    .ZN(_01782_)
  );
  INV_X1 _21952_ (
    .A(_01782_),
    .ZN(_01783_)
  );
  AND2_X1 _21953_ (
    .A1(_01781_),
    .A2(_01783_),
    .ZN(_01784_)
  );
  INV_X1 _21954_ (
    .A(_01784_),
    .ZN(_01785_)
  );
  AND2_X1 _21955_ (
    .A1(_13852_),
    .A2(_01785_),
    .ZN(_01786_)
  );
  INV_X1 _21956_ (
    .A(_01786_),
    .ZN(_01787_)
  );
  AND2_X1 _21957_ (
    .A1(_08068_),
    .A2(_13853_),
    .ZN(_01788_)
  );
  INV_X1 _21958_ (
    .A(_01788_),
    .ZN(_01789_)
  );
  AND2_X1 _21959_ (
    .A1(_13834_),
    .A2(_01789_),
    .ZN(_01790_)
  );
  AND2_X1 _21960_ (
    .A1(_01787_),
    .A2(_01790_),
    .ZN(_01791_)
  );
  INV_X1 _21961_ (
    .A(_01791_),
    .ZN(_01792_)
  );
  AND2_X1 _21962_ (
    .A1(_01764_),
    .A2(_01792_),
    .ZN(_01793_)
  );
  INV_X1 _21963_ (
    .A(_01793_),
    .ZN(_00133_)
  );
  AND2_X1 _21964_ (
    .A1(wb_reg_wdata[17]),
    .A2(_13833_),
    .ZN(_01794_)
  );
  INV_X1 _21965_ (
    .A(_01794_),
    .ZN(_01795_)
  );
  AND2_X1 _21966_ (
    .A1(_01769_),
    .A2(_01781_),
    .ZN(_01796_)
  );
  INV_X1 _21967_ (
    .A(_01796_),
    .ZN(_01797_)
  );
  AND2_X1 _21968_ (
    .A1(mem_reg_inst[17]),
    .A2(mem_ctrl_jal),
    .ZN(_01798_)
  );
  MUX2_X1 _21969_ (
    .A(_01798_),
    .B(mem_reg_inst[31]),
    .S(_10066_),
    .Z(_01799_)
  );
  INV_X1 _21970_ (
    .A(_01799_),
    .ZN(_01800_)
  );
  AND2_X1 _21971_ (
    .A1(mem_reg_pc[17]),
    .A2(_01799_),
    .ZN(_01801_)
  );
  INV_X1 _21972_ (
    .A(_01801_),
    .ZN(_01802_)
  );
  AND2_X1 _21973_ (
    .A1(_08014_),
    .A2(_01800_),
    .ZN(_01803_)
  );
  INV_X1 _21974_ (
    .A(_01803_),
    .ZN(_01804_)
  );
  AND2_X1 _21975_ (
    .A1(_01802_),
    .A2(_01804_),
    .ZN(_01805_)
  );
  INV_X1 _21976_ (
    .A(_01805_),
    .ZN(_01806_)
  );
  AND2_X1 _21977_ (
    .A1(_01797_),
    .A2(_01806_),
    .ZN(_01807_)
  );
  INV_X1 _21978_ (
    .A(_01807_),
    .ZN(_01808_)
  );
  AND2_X1 _21979_ (
    .A1(_01796_),
    .A2(_01805_),
    .ZN(_01809_)
  );
  INV_X1 _21980_ (
    .A(_01809_),
    .ZN(_01810_)
  );
  AND2_X1 _21981_ (
    .A1(_01808_),
    .A2(_01810_),
    .ZN(_01811_)
  );
  AND2_X1 _21982_ (
    .A1(_13852_),
    .A2(_01811_),
    .ZN(_01812_)
  );
  INV_X1 _21983_ (
    .A(_01812_),
    .ZN(_01813_)
  );
  AND2_X1 _21984_ (
    .A1(_08069_),
    .A2(_13853_),
    .ZN(_01814_)
  );
  INV_X1 _21985_ (
    .A(_01814_),
    .ZN(_01815_)
  );
  AND2_X1 _21986_ (
    .A1(_13834_),
    .A2(_01815_),
    .ZN(_01816_)
  );
  AND2_X1 _21987_ (
    .A1(_01813_),
    .A2(_01816_),
    .ZN(_01817_)
  );
  INV_X1 _21988_ (
    .A(_01817_),
    .ZN(_01818_)
  );
  AND2_X1 _21989_ (
    .A1(_01795_),
    .A2(_01818_),
    .ZN(_01819_)
  );
  INV_X1 _21990_ (
    .A(_01819_),
    .ZN(_00134_)
  );
  AND2_X1 _21991_ (
    .A1(wb_reg_wdata[18]),
    .A2(_13833_),
    .ZN(_01820_)
  );
  INV_X1 _21992_ (
    .A(_01820_),
    .ZN(_01821_)
  );
  AND2_X1 _21993_ (
    .A1(mem_reg_inst[18]),
    .A2(mem_ctrl_jal),
    .ZN(_01822_)
  );
  MUX2_X1 _21994_ (
    .A(_01822_),
    .B(mem_reg_inst[31]),
    .S(_10066_),
    .Z(_01823_)
  );
  INV_X1 _21995_ (
    .A(_01823_),
    .ZN(_01824_)
  );
  AND2_X1 _21996_ (
    .A1(mem_reg_pc[18]),
    .A2(_01823_),
    .ZN(_01825_)
  );
  INV_X1 _21997_ (
    .A(_01825_),
    .ZN(_01826_)
  );
  AND2_X1 _21998_ (
    .A1(_08016_),
    .A2(_01824_),
    .ZN(_01827_)
  );
  INV_X1 _21999_ (
    .A(_01827_),
    .ZN(_01828_)
  );
  AND2_X1 _22000_ (
    .A1(_01826_),
    .A2(_01828_),
    .ZN(_01829_)
  );
  INV_X1 _22001_ (
    .A(_01829_),
    .ZN(_01830_)
  );
  AND2_X1 _22002_ (
    .A1(_01796_),
    .A2(_01802_),
    .ZN(_01831_)
  );
  INV_X1 _22003_ (
    .A(_01831_),
    .ZN(_01832_)
  );
  AND2_X1 _22004_ (
    .A1(_01797_),
    .A2(_01804_),
    .ZN(_01833_)
  );
  INV_X1 _22005_ (
    .A(_01833_),
    .ZN(_01834_)
  );
  AND2_X1 _22006_ (
    .A1(_01804_),
    .A2(_01832_),
    .ZN(_01835_)
  );
  AND2_X1 _22007_ (
    .A1(_01802_),
    .A2(_01834_),
    .ZN(_01836_)
  );
  AND2_X1 _22008_ (
    .A1(_01829_),
    .A2(_01835_),
    .ZN(_01837_)
  );
  INV_X1 _22009_ (
    .A(_01837_),
    .ZN(_01838_)
  );
  AND2_X1 _22010_ (
    .A1(_01830_),
    .A2(_01836_),
    .ZN(_01839_)
  );
  INV_X1 _22011_ (
    .A(_01839_),
    .ZN(_01840_)
  );
  AND2_X1 _22012_ (
    .A1(_01838_),
    .A2(_01840_),
    .ZN(_01841_)
  );
  INV_X1 _22013_ (
    .A(_01841_),
    .ZN(_01842_)
  );
  AND2_X1 _22014_ (
    .A1(_13852_),
    .A2(_01842_),
    .ZN(_01843_)
  );
  INV_X1 _22015_ (
    .A(_01843_),
    .ZN(_01844_)
  );
  AND2_X1 _22016_ (
    .A1(_08070_),
    .A2(_13853_),
    .ZN(_01845_)
  );
  INV_X1 _22017_ (
    .A(_01845_),
    .ZN(_01846_)
  );
  AND2_X1 _22018_ (
    .A1(_13834_),
    .A2(_01846_),
    .ZN(_01847_)
  );
  AND2_X1 _22019_ (
    .A1(_01844_),
    .A2(_01847_),
    .ZN(_01848_)
  );
  INV_X1 _22020_ (
    .A(_01848_),
    .ZN(_01849_)
  );
  AND2_X1 _22021_ (
    .A1(_01821_),
    .A2(_01849_),
    .ZN(_01850_)
  );
  INV_X1 _22022_ (
    .A(_01850_),
    .ZN(_00135_)
  );
  AND2_X1 _22023_ (
    .A1(wb_reg_wdata[19]),
    .A2(_13833_),
    .ZN(_01851_)
  );
  INV_X1 _22024_ (
    .A(_01851_),
    .ZN(_01852_)
  );
  AND2_X1 _22025_ (
    .A1(_01826_),
    .A2(_01838_),
    .ZN(_01853_)
  );
  INV_X1 _22026_ (
    .A(_01853_),
    .ZN(_01854_)
  );
  AND2_X1 _22027_ (
    .A1(mem_reg_inst[19]),
    .A2(mem_ctrl_jal),
    .ZN(_01855_)
  );
  MUX2_X1 _22028_ (
    .A(_01855_),
    .B(mem_reg_inst[31]),
    .S(_10066_),
    .Z(_01856_)
  );
  INV_X1 _22029_ (
    .A(_01856_),
    .ZN(_01857_)
  );
  AND2_X1 _22030_ (
    .A1(mem_reg_pc[19]),
    .A2(_01856_),
    .ZN(_01858_)
  );
  INV_X1 _22031_ (
    .A(_01858_),
    .ZN(_01859_)
  );
  AND2_X1 _22032_ (
    .A1(_08018_),
    .A2(_01857_),
    .ZN(_01860_)
  );
  INV_X1 _22033_ (
    .A(_01860_),
    .ZN(_01861_)
  );
  AND2_X1 _22034_ (
    .A1(_01859_),
    .A2(_01861_),
    .ZN(_01862_)
  );
  INV_X1 _22035_ (
    .A(_01862_),
    .ZN(_01863_)
  );
  AND2_X1 _22036_ (
    .A1(_01854_),
    .A2(_01863_),
    .ZN(_01864_)
  );
  INV_X1 _22037_ (
    .A(_01864_),
    .ZN(_01865_)
  );
  AND2_X1 _22038_ (
    .A1(_01853_),
    .A2(_01862_),
    .ZN(_01866_)
  );
  INV_X1 _22039_ (
    .A(_01866_),
    .ZN(_01867_)
  );
  AND2_X1 _22040_ (
    .A1(_01865_),
    .A2(_01867_),
    .ZN(_01868_)
  );
  AND2_X1 _22041_ (
    .A1(_13852_),
    .A2(_01868_),
    .ZN(_01869_)
  );
  INV_X1 _22042_ (
    .A(_01869_),
    .ZN(_01870_)
  );
  AND2_X1 _22043_ (
    .A1(_08071_),
    .A2(_13853_),
    .ZN(_01871_)
  );
  INV_X1 _22044_ (
    .A(_01871_),
    .ZN(_01872_)
  );
  AND2_X1 _22045_ (
    .A1(_13834_),
    .A2(_01872_),
    .ZN(_01873_)
  );
  AND2_X1 _22046_ (
    .A1(_01870_),
    .A2(_01873_),
    .ZN(_01874_)
  );
  INV_X1 _22047_ (
    .A(_01874_),
    .ZN(_01875_)
  );
  AND2_X1 _22048_ (
    .A1(_01852_),
    .A2(_01875_),
    .ZN(_01876_)
  );
  INV_X1 _22049_ (
    .A(_01876_),
    .ZN(_00136_)
  );
  AND2_X1 _22050_ (
    .A1(wb_reg_wdata[20]),
    .A2(_13833_),
    .ZN(_01877_)
  );
  INV_X1 _22051_ (
    .A(_01877_),
    .ZN(_01878_)
  );
  AND2_X1 _22052_ (
    .A1(mem_reg_inst[31]),
    .A2(_10069_),
    .ZN(_01879_)
  );
  INV_X1 _22053_ (
    .A(_01879_),
    .ZN(_01880_)
  );
  AND2_X1 _22054_ (
    .A1(mem_reg_pc[20]),
    .A2(_01879_),
    .ZN(_01881_)
  );
  INV_X1 _22055_ (
    .A(_01881_),
    .ZN(_01882_)
  );
  AND2_X1 _22056_ (
    .A1(_08020_),
    .A2(_01880_),
    .ZN(_01883_)
  );
  INV_X1 _22057_ (
    .A(_01883_),
    .ZN(_01884_)
  );
  AND2_X1 _22058_ (
    .A1(_01882_),
    .A2(_01884_),
    .ZN(_01885_)
  );
  INV_X1 _22059_ (
    .A(_01885_),
    .ZN(_01886_)
  );
  AND2_X1 _22060_ (
    .A1(_01853_),
    .A2(_01859_),
    .ZN(_01887_)
  );
  INV_X1 _22061_ (
    .A(_01887_),
    .ZN(_01888_)
  );
  AND2_X1 _22062_ (
    .A1(_01854_),
    .A2(_01861_),
    .ZN(_01889_)
  );
  INV_X1 _22063_ (
    .A(_01889_),
    .ZN(_01890_)
  );
  AND2_X1 _22064_ (
    .A1(_01861_),
    .A2(_01888_),
    .ZN(_01891_)
  );
  AND2_X1 _22065_ (
    .A1(_01859_),
    .A2(_01890_),
    .ZN(_01892_)
  );
  AND2_X1 _22066_ (
    .A1(_01885_),
    .A2(_01891_),
    .ZN(_01893_)
  );
  INV_X1 _22067_ (
    .A(_01893_),
    .ZN(_01894_)
  );
  AND2_X1 _22068_ (
    .A1(_01886_),
    .A2(_01892_),
    .ZN(_01895_)
  );
  INV_X1 _22069_ (
    .A(_01895_),
    .ZN(_01896_)
  );
  AND2_X1 _22070_ (
    .A1(_01894_),
    .A2(_01896_),
    .ZN(_01897_)
  );
  INV_X1 _22071_ (
    .A(_01897_),
    .ZN(_01898_)
  );
  AND2_X1 _22072_ (
    .A1(_13852_),
    .A2(_01898_),
    .ZN(_01899_)
  );
  INV_X1 _22073_ (
    .A(_01899_),
    .ZN(_01900_)
  );
  AND2_X1 _22074_ (
    .A1(_08072_),
    .A2(_13853_),
    .ZN(_01901_)
  );
  INV_X1 _22075_ (
    .A(_01901_),
    .ZN(_01902_)
  );
  AND2_X1 _22076_ (
    .A1(_13834_),
    .A2(_01902_),
    .ZN(_01903_)
  );
  AND2_X1 _22077_ (
    .A1(_01900_),
    .A2(_01903_),
    .ZN(_01904_)
  );
  INV_X1 _22078_ (
    .A(_01904_),
    .ZN(_01905_)
  );
  AND2_X1 _22079_ (
    .A1(_01878_),
    .A2(_01905_),
    .ZN(_01906_)
  );
  INV_X1 _22080_ (
    .A(_01906_),
    .ZN(_00137_)
  );
  AND2_X1 _22081_ (
    .A1(wb_reg_wdata[21]),
    .A2(_13833_),
    .ZN(_01907_)
  );
  INV_X1 _22082_ (
    .A(_01907_),
    .ZN(_01908_)
  );
  AND2_X1 _22083_ (
    .A1(_01882_),
    .A2(_01894_),
    .ZN(_01909_)
  );
  INV_X1 _22084_ (
    .A(_01909_),
    .ZN(_01910_)
  );
  AND2_X1 _22085_ (
    .A1(mem_reg_pc[21]),
    .A2(_01879_),
    .ZN(_01911_)
  );
  INV_X1 _22086_ (
    .A(_01911_),
    .ZN(_01912_)
  );
  AND2_X1 _22087_ (
    .A1(_08022_),
    .A2(_01880_),
    .ZN(_01913_)
  );
  INV_X1 _22088_ (
    .A(_01913_),
    .ZN(_01914_)
  );
  AND2_X1 _22089_ (
    .A1(_01912_),
    .A2(_01914_),
    .ZN(_01915_)
  );
  INV_X1 _22090_ (
    .A(_01915_),
    .ZN(_01916_)
  );
  AND2_X1 _22091_ (
    .A1(_01909_),
    .A2(_01915_),
    .ZN(_01917_)
  );
  INV_X1 _22092_ (
    .A(_01917_),
    .ZN(_01918_)
  );
  AND2_X1 _22093_ (
    .A1(_01910_),
    .A2(_01916_),
    .ZN(_01919_)
  );
  INV_X1 _22094_ (
    .A(_01919_),
    .ZN(_01920_)
  );
  AND2_X1 _22095_ (
    .A1(_01918_),
    .A2(_01920_),
    .ZN(_01921_)
  );
  AND2_X1 _22096_ (
    .A1(_13852_),
    .A2(_01921_),
    .ZN(_01922_)
  );
  INV_X1 _22097_ (
    .A(_01922_),
    .ZN(_01923_)
  );
  AND2_X1 _22098_ (
    .A1(_08073_),
    .A2(_13853_),
    .ZN(_01924_)
  );
  INV_X1 _22099_ (
    .A(_01924_),
    .ZN(_01925_)
  );
  AND2_X1 _22100_ (
    .A1(_13834_),
    .A2(_01925_),
    .ZN(_01926_)
  );
  AND2_X1 _22101_ (
    .A1(_01923_),
    .A2(_01926_),
    .ZN(_01927_)
  );
  INV_X1 _22102_ (
    .A(_01927_),
    .ZN(_01928_)
  );
  AND2_X1 _22103_ (
    .A1(_01908_),
    .A2(_01928_),
    .ZN(_01929_)
  );
  INV_X1 _22104_ (
    .A(_01929_),
    .ZN(_00138_)
  );
  AND2_X1 _22105_ (
    .A1(wb_reg_wdata[22]),
    .A2(_13833_),
    .ZN(_01930_)
  );
  INV_X1 _22106_ (
    .A(_01930_),
    .ZN(_01931_)
  );
  AND2_X1 _22107_ (
    .A1(_01882_),
    .A2(_01912_),
    .ZN(_01932_)
  );
  INV_X1 _22108_ (
    .A(_01932_),
    .ZN(_01933_)
  );
  AND2_X1 _22109_ (
    .A1(_01893_),
    .A2(_01915_),
    .ZN(_01934_)
  );
  INV_X1 _22110_ (
    .A(_01934_),
    .ZN(_01935_)
  );
  AND2_X1 _22111_ (
    .A1(_01932_),
    .A2(_01935_),
    .ZN(_01936_)
  );
  INV_X1 _22112_ (
    .A(_01936_),
    .ZN(_01937_)
  );
  AND2_X1 _22113_ (
    .A1(mem_reg_pc[22]),
    .A2(_01879_),
    .ZN(_01938_)
  );
  INV_X1 _22114_ (
    .A(_01938_),
    .ZN(_01939_)
  );
  AND2_X1 _22115_ (
    .A1(_08024_),
    .A2(_01880_),
    .ZN(_01940_)
  );
  INV_X1 _22116_ (
    .A(_01940_),
    .ZN(_01941_)
  );
  AND2_X1 _22117_ (
    .A1(_01939_),
    .A2(_01941_),
    .ZN(_01942_)
  );
  INV_X1 _22118_ (
    .A(_01942_),
    .ZN(_01943_)
  );
  AND2_X1 _22119_ (
    .A1(_01937_),
    .A2(_01942_),
    .ZN(_01944_)
  );
  INV_X1 _22120_ (
    .A(_01944_),
    .ZN(_01945_)
  );
  AND2_X1 _22121_ (
    .A1(_01936_),
    .A2(_01943_),
    .ZN(_01946_)
  );
  INV_X1 _22122_ (
    .A(_01946_),
    .ZN(_01947_)
  );
  AND2_X1 _22123_ (
    .A1(_01945_),
    .A2(_01947_),
    .ZN(_01948_)
  );
  INV_X1 _22124_ (
    .A(_01948_),
    .ZN(_01949_)
  );
  AND2_X1 _22125_ (
    .A1(_13852_),
    .A2(_01949_),
    .ZN(_01950_)
  );
  INV_X1 _22126_ (
    .A(_01950_),
    .ZN(_01951_)
  );
  AND2_X1 _22127_ (
    .A1(_08074_),
    .A2(_13853_),
    .ZN(_01952_)
  );
  INV_X1 _22128_ (
    .A(_01952_),
    .ZN(_01953_)
  );
  AND2_X1 _22129_ (
    .A1(_13834_),
    .A2(_01953_),
    .ZN(_01954_)
  );
  AND2_X1 _22130_ (
    .A1(_01951_),
    .A2(_01954_),
    .ZN(_01955_)
  );
  INV_X1 _22131_ (
    .A(_01955_),
    .ZN(_01956_)
  );
  AND2_X1 _22132_ (
    .A1(_01931_),
    .A2(_01956_),
    .ZN(_01957_)
  );
  INV_X1 _22133_ (
    .A(_01957_),
    .ZN(_00139_)
  );
  AND2_X1 _22134_ (
    .A1(wb_reg_wdata[23]),
    .A2(_13833_),
    .ZN(_01958_)
  );
  INV_X1 _22135_ (
    .A(_01958_),
    .ZN(_01959_)
  );
  AND2_X1 _22136_ (
    .A1(_01939_),
    .A2(_01945_),
    .ZN(_01960_)
  );
  INV_X1 _22137_ (
    .A(_01960_),
    .ZN(_01961_)
  );
  AND2_X1 _22138_ (
    .A1(mem_reg_pc[23]),
    .A2(_01879_),
    .ZN(_01962_)
  );
  INV_X1 _22139_ (
    .A(_01962_),
    .ZN(_01963_)
  );
  AND2_X1 _22140_ (
    .A1(_08026_),
    .A2(_01880_),
    .ZN(_01964_)
  );
  INV_X1 _22141_ (
    .A(_01964_),
    .ZN(_01965_)
  );
  AND2_X1 _22142_ (
    .A1(_01963_),
    .A2(_01965_),
    .ZN(_01966_)
  );
  INV_X1 _22143_ (
    .A(_01966_),
    .ZN(_01967_)
  );
  AND2_X1 _22144_ (
    .A1(_01960_),
    .A2(_01966_),
    .ZN(_01968_)
  );
  INV_X1 _22145_ (
    .A(_01968_),
    .ZN(_01969_)
  );
  AND2_X1 _22146_ (
    .A1(_01961_),
    .A2(_01967_),
    .ZN(_01970_)
  );
  INV_X1 _22147_ (
    .A(_01970_),
    .ZN(_01971_)
  );
  AND2_X1 _22148_ (
    .A1(_01969_),
    .A2(_01971_),
    .ZN(_01972_)
  );
  AND2_X1 _22149_ (
    .A1(_13852_),
    .A2(_01972_),
    .ZN(_01973_)
  );
  INV_X1 _22150_ (
    .A(_01973_),
    .ZN(_01974_)
  );
  AND2_X1 _22151_ (
    .A1(_08075_),
    .A2(_13853_),
    .ZN(_01975_)
  );
  INV_X1 _22152_ (
    .A(_01975_),
    .ZN(_01976_)
  );
  AND2_X1 _22153_ (
    .A1(_13834_),
    .A2(_01976_),
    .ZN(_01977_)
  );
  AND2_X1 _22154_ (
    .A1(_01974_),
    .A2(_01977_),
    .ZN(_01978_)
  );
  INV_X1 _22155_ (
    .A(_01978_),
    .ZN(_01979_)
  );
  AND2_X1 _22156_ (
    .A1(_01959_),
    .A2(_01979_),
    .ZN(_01980_)
  );
  INV_X1 _22157_ (
    .A(_01980_),
    .ZN(_00140_)
  );
  AND2_X1 _22158_ (
    .A1(wb_reg_wdata[24]),
    .A2(_13833_),
    .ZN(_01981_)
  );
  INV_X1 _22159_ (
    .A(_01981_),
    .ZN(_01982_)
  );
  AND2_X1 _22160_ (
    .A1(_01942_),
    .A2(_01966_),
    .ZN(_01983_)
  );
  AND2_X1 _22161_ (
    .A1(_01934_),
    .A2(_01983_),
    .ZN(_01984_)
  );
  INV_X1 _22162_ (
    .A(_01984_),
    .ZN(_01985_)
  );
  AND2_X1 _22163_ (
    .A1(_01933_),
    .A2(_01983_),
    .ZN(_01986_)
  );
  INV_X1 _22164_ (
    .A(_01986_),
    .ZN(_01987_)
  );
  AND2_X1 _22165_ (
    .A1(_01939_),
    .A2(_01963_),
    .ZN(_01988_)
  );
  AND2_X1 _22166_ (
    .A1(_01987_),
    .A2(_01988_),
    .ZN(_01989_)
  );
  AND2_X1 _22167_ (
    .A1(_01985_),
    .A2(_01989_),
    .ZN(_01990_)
  );
  INV_X1 _22168_ (
    .A(_01990_),
    .ZN(_01991_)
  );
  AND2_X1 _22169_ (
    .A1(mem_reg_pc[24]),
    .A2(_01879_),
    .ZN(_01992_)
  );
  INV_X1 _22170_ (
    .A(_01992_),
    .ZN(_01993_)
  );
  AND2_X1 _22171_ (
    .A1(_08028_),
    .A2(_01880_),
    .ZN(_01994_)
  );
  INV_X1 _22172_ (
    .A(_01994_),
    .ZN(_01995_)
  );
  AND2_X1 _22173_ (
    .A1(_01993_),
    .A2(_01995_),
    .ZN(_01996_)
  );
  INV_X1 _22174_ (
    .A(_01996_),
    .ZN(_01997_)
  );
  AND2_X1 _22175_ (
    .A1(_01991_),
    .A2(_01996_),
    .ZN(_01998_)
  );
  INV_X1 _22176_ (
    .A(_01998_),
    .ZN(_01999_)
  );
  AND2_X1 _22177_ (
    .A1(_01990_),
    .A2(_01997_),
    .ZN(_02000_)
  );
  INV_X1 _22178_ (
    .A(_02000_),
    .ZN(_02001_)
  );
  AND2_X1 _22179_ (
    .A1(_01999_),
    .A2(_02001_),
    .ZN(_02002_)
  );
  INV_X1 _22180_ (
    .A(_02002_),
    .ZN(_02003_)
  );
  AND2_X1 _22181_ (
    .A1(_13852_),
    .A2(_02003_),
    .ZN(_02004_)
  );
  INV_X1 _22182_ (
    .A(_02004_),
    .ZN(_02005_)
  );
  AND2_X1 _22183_ (
    .A1(_08076_),
    .A2(_13853_),
    .ZN(_02006_)
  );
  INV_X1 _22184_ (
    .A(_02006_),
    .ZN(_02007_)
  );
  AND2_X1 _22185_ (
    .A1(_13834_),
    .A2(_02007_),
    .ZN(_02008_)
  );
  AND2_X1 _22186_ (
    .A1(_02005_),
    .A2(_02008_),
    .ZN(_02009_)
  );
  INV_X1 _22187_ (
    .A(_02009_),
    .ZN(_02010_)
  );
  AND2_X1 _22188_ (
    .A1(_01982_),
    .A2(_02010_),
    .ZN(_02011_)
  );
  INV_X1 _22189_ (
    .A(_02011_),
    .ZN(_00141_)
  );
  AND2_X1 _22190_ (
    .A1(wb_reg_wdata[25]),
    .A2(_13833_),
    .ZN(_02012_)
  );
  INV_X1 _22191_ (
    .A(_02012_),
    .ZN(_02013_)
  );
  AND2_X1 _22192_ (
    .A1(_01993_),
    .A2(_01999_),
    .ZN(_02014_)
  );
  INV_X1 _22193_ (
    .A(_02014_),
    .ZN(_02015_)
  );
  AND2_X1 _22194_ (
    .A1(mem_reg_pc[25]),
    .A2(_01879_),
    .ZN(_02016_)
  );
  INV_X1 _22195_ (
    .A(_02016_),
    .ZN(_02017_)
  );
  AND2_X1 _22196_ (
    .A1(_08030_),
    .A2(_01880_),
    .ZN(_02018_)
  );
  INV_X1 _22197_ (
    .A(_02018_),
    .ZN(_02019_)
  );
  AND2_X1 _22198_ (
    .A1(_02017_),
    .A2(_02019_),
    .ZN(_02020_)
  );
  INV_X1 _22199_ (
    .A(_02020_),
    .ZN(_02021_)
  );
  AND2_X1 _22200_ (
    .A1(_02014_),
    .A2(_02020_),
    .ZN(_02022_)
  );
  INV_X1 _22201_ (
    .A(_02022_),
    .ZN(_02023_)
  );
  AND2_X1 _22202_ (
    .A1(_02015_),
    .A2(_02021_),
    .ZN(_02024_)
  );
  INV_X1 _22203_ (
    .A(_02024_),
    .ZN(_02025_)
  );
  AND2_X1 _22204_ (
    .A1(_02023_),
    .A2(_02025_),
    .ZN(_02026_)
  );
  AND2_X1 _22205_ (
    .A1(_13852_),
    .A2(_02026_),
    .ZN(_02027_)
  );
  INV_X1 _22206_ (
    .A(_02027_),
    .ZN(_02028_)
  );
  AND2_X1 _22207_ (
    .A1(_08077_),
    .A2(_13853_),
    .ZN(_02029_)
  );
  INV_X1 _22208_ (
    .A(_02029_),
    .ZN(_02030_)
  );
  AND2_X1 _22209_ (
    .A1(_13834_),
    .A2(_02030_),
    .ZN(_02031_)
  );
  AND2_X1 _22210_ (
    .A1(_02028_),
    .A2(_02031_),
    .ZN(_02032_)
  );
  INV_X1 _22211_ (
    .A(_02032_),
    .ZN(_02033_)
  );
  AND2_X1 _22212_ (
    .A1(_02013_),
    .A2(_02033_),
    .ZN(_02034_)
  );
  INV_X1 _22213_ (
    .A(_02034_),
    .ZN(_00142_)
  );
  AND2_X1 _22214_ (
    .A1(wb_reg_wdata[26]),
    .A2(_13833_),
    .ZN(_02035_)
  );
  INV_X1 _22215_ (
    .A(_02035_),
    .ZN(_02036_)
  );
  AND2_X1 _22216_ (
    .A1(_01993_),
    .A2(_02017_),
    .ZN(_02037_)
  );
  INV_X1 _22217_ (
    .A(_02037_),
    .ZN(_02038_)
  );
  AND2_X1 _22218_ (
    .A1(_01998_),
    .A2(_02020_),
    .ZN(_02039_)
  );
  INV_X1 _22219_ (
    .A(_02039_),
    .ZN(_02040_)
  );
  AND2_X1 _22220_ (
    .A1(_02037_),
    .A2(_02040_),
    .ZN(_02041_)
  );
  INV_X1 _22221_ (
    .A(_02041_),
    .ZN(_02042_)
  );
  AND2_X1 _22222_ (
    .A1(mem_reg_pc[26]),
    .A2(_01879_),
    .ZN(_02043_)
  );
  INV_X1 _22223_ (
    .A(_02043_),
    .ZN(_02044_)
  );
  AND2_X1 _22224_ (
    .A1(_08032_),
    .A2(_01880_),
    .ZN(_02045_)
  );
  INV_X1 _22225_ (
    .A(_02045_),
    .ZN(_02046_)
  );
  AND2_X1 _22226_ (
    .A1(_02044_),
    .A2(_02046_),
    .ZN(_02047_)
  );
  INV_X1 _22227_ (
    .A(_02047_),
    .ZN(_02048_)
  );
  AND2_X1 _22228_ (
    .A1(_02042_),
    .A2(_02047_),
    .ZN(_02049_)
  );
  INV_X1 _22229_ (
    .A(_02049_),
    .ZN(_02050_)
  );
  AND2_X1 _22230_ (
    .A1(_02041_),
    .A2(_02048_),
    .ZN(_02051_)
  );
  INV_X1 _22231_ (
    .A(_02051_),
    .ZN(_02052_)
  );
  AND2_X1 _22232_ (
    .A1(_02050_),
    .A2(_02052_),
    .ZN(_02053_)
  );
  INV_X1 _22233_ (
    .A(_02053_),
    .ZN(_02054_)
  );
  AND2_X1 _22234_ (
    .A1(_13852_),
    .A2(_02054_),
    .ZN(_02055_)
  );
  INV_X1 _22235_ (
    .A(_02055_),
    .ZN(_02056_)
  );
  AND2_X1 _22236_ (
    .A1(_08078_),
    .A2(_13853_),
    .ZN(_02057_)
  );
  INV_X1 _22237_ (
    .A(_02057_),
    .ZN(_02058_)
  );
  AND2_X1 _22238_ (
    .A1(_13834_),
    .A2(_02058_),
    .ZN(_02059_)
  );
  AND2_X1 _22239_ (
    .A1(_02056_),
    .A2(_02059_),
    .ZN(_02060_)
  );
  INV_X1 _22240_ (
    .A(_02060_),
    .ZN(_02061_)
  );
  AND2_X1 _22241_ (
    .A1(_02036_),
    .A2(_02061_),
    .ZN(_02062_)
  );
  INV_X1 _22242_ (
    .A(_02062_),
    .ZN(_00143_)
  );
  AND2_X1 _22243_ (
    .A1(wb_reg_wdata[27]),
    .A2(_13833_),
    .ZN(_02063_)
  );
  INV_X1 _22244_ (
    .A(_02063_),
    .ZN(_02064_)
  );
  AND2_X1 _22245_ (
    .A1(_02044_),
    .A2(_02050_),
    .ZN(_02065_)
  );
  INV_X1 _22246_ (
    .A(_02065_),
    .ZN(_02066_)
  );
  AND2_X1 _22247_ (
    .A1(mem_reg_pc[27]),
    .A2(_01879_),
    .ZN(_02067_)
  );
  INV_X1 _22248_ (
    .A(_02067_),
    .ZN(_02068_)
  );
  AND2_X1 _22249_ (
    .A1(_08034_),
    .A2(_01880_),
    .ZN(_02069_)
  );
  INV_X1 _22250_ (
    .A(_02069_),
    .ZN(_02070_)
  );
  AND2_X1 _22251_ (
    .A1(_02068_),
    .A2(_02070_),
    .ZN(_02071_)
  );
  INV_X1 _22252_ (
    .A(_02071_),
    .ZN(_02072_)
  );
  AND2_X1 _22253_ (
    .A1(_02065_),
    .A2(_02071_),
    .ZN(_02073_)
  );
  INV_X1 _22254_ (
    .A(_02073_),
    .ZN(_02074_)
  );
  AND2_X1 _22255_ (
    .A1(_02066_),
    .A2(_02072_),
    .ZN(_02075_)
  );
  INV_X1 _22256_ (
    .A(_02075_),
    .ZN(_02076_)
  );
  AND2_X1 _22257_ (
    .A1(_02074_),
    .A2(_02076_),
    .ZN(_02077_)
  );
  AND2_X1 _22258_ (
    .A1(_13852_),
    .A2(_02077_),
    .ZN(_02078_)
  );
  INV_X1 _22259_ (
    .A(_02078_),
    .ZN(_02079_)
  );
  AND2_X1 _22260_ (
    .A1(_08079_),
    .A2(_13853_),
    .ZN(_02080_)
  );
  INV_X1 _22261_ (
    .A(_02080_),
    .ZN(_02081_)
  );
  AND2_X1 _22262_ (
    .A1(_13834_),
    .A2(_02081_),
    .ZN(_02082_)
  );
  AND2_X1 _22263_ (
    .A1(_02079_),
    .A2(_02082_),
    .ZN(_02083_)
  );
  INV_X1 _22264_ (
    .A(_02083_),
    .ZN(_02084_)
  );
  AND2_X1 _22265_ (
    .A1(_02064_),
    .A2(_02084_),
    .ZN(_02085_)
  );
  INV_X1 _22266_ (
    .A(_02085_),
    .ZN(_00144_)
  );
  AND2_X1 _22267_ (
    .A1(wb_reg_wdata[28]),
    .A2(_13833_),
    .ZN(_02086_)
  );
  INV_X1 _22268_ (
    .A(_02086_),
    .ZN(_02087_)
  );
  AND2_X1 _22269_ (
    .A1(_02047_),
    .A2(_02071_),
    .ZN(_02088_)
  );
  AND2_X1 _22270_ (
    .A1(_02039_),
    .A2(_02088_),
    .ZN(_02089_)
  );
  INV_X1 _22271_ (
    .A(_02089_),
    .ZN(_02090_)
  );
  AND2_X1 _22272_ (
    .A1(_02038_),
    .A2(_02088_),
    .ZN(_02091_)
  );
  INV_X1 _22273_ (
    .A(_02091_),
    .ZN(_02092_)
  );
  AND2_X1 _22274_ (
    .A1(_02044_),
    .A2(_02068_),
    .ZN(_02093_)
  );
  AND2_X1 _22275_ (
    .A1(_02092_),
    .A2(_02093_),
    .ZN(_02094_)
  );
  AND2_X1 _22276_ (
    .A1(_02090_),
    .A2(_02094_),
    .ZN(_02095_)
  );
  INV_X1 _22277_ (
    .A(_02095_),
    .ZN(_02096_)
  );
  AND2_X1 _22278_ (
    .A1(mem_reg_pc[28]),
    .A2(_01879_),
    .ZN(_02097_)
  );
  INV_X1 _22279_ (
    .A(_02097_),
    .ZN(_02098_)
  );
  AND2_X1 _22280_ (
    .A1(_08036_),
    .A2(_01880_),
    .ZN(_02099_)
  );
  INV_X1 _22281_ (
    .A(_02099_),
    .ZN(_02100_)
  );
  AND2_X1 _22282_ (
    .A1(_02098_),
    .A2(_02100_),
    .ZN(_02101_)
  );
  INV_X1 _22283_ (
    .A(_02101_),
    .ZN(_02102_)
  );
  AND2_X1 _22284_ (
    .A1(_02096_),
    .A2(_02101_),
    .ZN(_02103_)
  );
  INV_X1 _22285_ (
    .A(_02103_),
    .ZN(_02104_)
  );
  AND2_X1 _22286_ (
    .A1(_02095_),
    .A2(_02102_),
    .ZN(_02105_)
  );
  INV_X1 _22287_ (
    .A(_02105_),
    .ZN(_02106_)
  );
  AND2_X1 _22288_ (
    .A1(_02104_),
    .A2(_02106_),
    .ZN(_02107_)
  );
  INV_X1 _22289_ (
    .A(_02107_),
    .ZN(_02108_)
  );
  AND2_X1 _22290_ (
    .A1(_13852_),
    .A2(_02108_),
    .ZN(_02109_)
  );
  INV_X1 _22291_ (
    .A(_02109_),
    .ZN(_02110_)
  );
  AND2_X1 _22292_ (
    .A1(_08080_),
    .A2(_13853_),
    .ZN(_02111_)
  );
  INV_X1 _22293_ (
    .A(_02111_),
    .ZN(_02112_)
  );
  AND2_X1 _22294_ (
    .A1(_13834_),
    .A2(_02112_),
    .ZN(_02113_)
  );
  AND2_X1 _22295_ (
    .A1(_02110_),
    .A2(_02113_),
    .ZN(_02114_)
  );
  INV_X1 _22296_ (
    .A(_02114_),
    .ZN(_02115_)
  );
  AND2_X1 _22297_ (
    .A1(_02087_),
    .A2(_02115_),
    .ZN(_02116_)
  );
  INV_X1 _22298_ (
    .A(_02116_),
    .ZN(_00145_)
  );
  AND2_X1 _22299_ (
    .A1(wb_reg_wdata[29]),
    .A2(_13833_),
    .ZN(_02117_)
  );
  INV_X1 _22300_ (
    .A(_02117_),
    .ZN(_02118_)
  );
  AND2_X1 _22301_ (
    .A1(_02098_),
    .A2(_02104_),
    .ZN(_02119_)
  );
  INV_X1 _22302_ (
    .A(_02119_),
    .ZN(_02120_)
  );
  AND2_X1 _22303_ (
    .A1(mem_reg_pc[29]),
    .A2(_01879_),
    .ZN(_02121_)
  );
  INV_X1 _22304_ (
    .A(_02121_),
    .ZN(_02122_)
  );
  AND2_X1 _22305_ (
    .A1(_08038_),
    .A2(_01880_),
    .ZN(_02123_)
  );
  INV_X1 _22306_ (
    .A(_02123_),
    .ZN(_02124_)
  );
  AND2_X1 _22307_ (
    .A1(_02122_),
    .A2(_02124_),
    .ZN(_02125_)
  );
  INV_X1 _22308_ (
    .A(_02125_),
    .ZN(_02126_)
  );
  AND2_X1 _22309_ (
    .A1(_02119_),
    .A2(_02126_),
    .ZN(_02127_)
  );
  INV_X1 _22310_ (
    .A(_02127_),
    .ZN(_02128_)
  );
  AND2_X1 _22311_ (
    .A1(_02120_),
    .A2(_02125_),
    .ZN(_02129_)
  );
  INV_X1 _22312_ (
    .A(_02129_),
    .ZN(_02130_)
  );
  AND2_X1 _22313_ (
    .A1(_02128_),
    .A2(_02130_),
    .ZN(_02131_)
  );
  INV_X1 _22314_ (
    .A(_02131_),
    .ZN(_02132_)
  );
  AND2_X1 _22315_ (
    .A1(_13852_),
    .A2(_02132_),
    .ZN(_02133_)
  );
  INV_X1 _22316_ (
    .A(_02133_),
    .ZN(_02134_)
  );
  AND2_X1 _22317_ (
    .A1(_08081_),
    .A2(_13853_),
    .ZN(_02135_)
  );
  INV_X1 _22318_ (
    .A(_02135_),
    .ZN(_02136_)
  );
  AND2_X1 _22319_ (
    .A1(_13834_),
    .A2(_02136_),
    .ZN(_02137_)
  );
  AND2_X1 _22320_ (
    .A1(_02134_),
    .A2(_02137_),
    .ZN(_02138_)
  );
  INV_X1 _22321_ (
    .A(_02138_),
    .ZN(_02139_)
  );
  AND2_X1 _22322_ (
    .A1(_02118_),
    .A2(_02139_),
    .ZN(_02140_)
  );
  INV_X1 _22323_ (
    .A(_02140_),
    .ZN(_00146_)
  );
  AND2_X1 _22324_ (
    .A1(wb_reg_wdata[30]),
    .A2(_13833_),
    .ZN(_02141_)
  );
  INV_X1 _22325_ (
    .A(_02141_),
    .ZN(_02142_)
  );
  AND2_X1 _22326_ (
    .A1(mem_reg_pc[30]),
    .A2(_01879_),
    .ZN(_02143_)
  );
  INV_X1 _22327_ (
    .A(_02143_),
    .ZN(_02144_)
  );
  AND2_X1 _22328_ (
    .A1(_08040_),
    .A2(_01880_),
    .ZN(_02145_)
  );
  INV_X1 _22329_ (
    .A(_02145_),
    .ZN(_02146_)
  );
  AND2_X1 _22330_ (
    .A1(_02144_),
    .A2(_02146_),
    .ZN(_02147_)
  );
  INV_X1 _22331_ (
    .A(_02147_),
    .ZN(_02148_)
  );
  AND2_X1 _22332_ (
    .A1(_02120_),
    .A2(_02124_),
    .ZN(_02149_)
  );
  INV_X1 _22333_ (
    .A(_02149_),
    .ZN(_02150_)
  );
  AND2_X1 _22334_ (
    .A1(_02119_),
    .A2(_02122_),
    .ZN(_02151_)
  );
  INV_X1 _22335_ (
    .A(_02151_),
    .ZN(_02152_)
  );
  AND2_X1 _22336_ (
    .A1(_02122_),
    .A2(_02150_),
    .ZN(_02153_)
  );
  AND2_X1 _22337_ (
    .A1(_02124_),
    .A2(_02152_),
    .ZN(_02154_)
  );
  AND2_X1 _22338_ (
    .A1(_02147_),
    .A2(_02154_),
    .ZN(_02155_)
  );
  INV_X1 _22339_ (
    .A(_02155_),
    .ZN(_02156_)
  );
  AND2_X1 _22340_ (
    .A1(_02148_),
    .A2(_02153_),
    .ZN(_02157_)
  );
  INV_X1 _22341_ (
    .A(_02157_),
    .ZN(_02158_)
  );
  AND2_X1 _22342_ (
    .A1(_02156_),
    .A2(_02158_),
    .ZN(_02159_)
  );
  INV_X1 _22343_ (
    .A(_02159_),
    .ZN(_02160_)
  );
  AND2_X1 _22344_ (
    .A1(_13852_),
    .A2(_02160_),
    .ZN(_02161_)
  );
  INV_X1 _22345_ (
    .A(_02161_),
    .ZN(_02162_)
  );
  AND2_X1 _22346_ (
    .A1(_08082_),
    .A2(_13853_),
    .ZN(_02163_)
  );
  INV_X1 _22347_ (
    .A(_02163_),
    .ZN(_02164_)
  );
  AND2_X1 _22348_ (
    .A1(_13834_),
    .A2(_02164_),
    .ZN(_02165_)
  );
  AND2_X1 _22349_ (
    .A1(_02162_),
    .A2(_02165_),
    .ZN(_02166_)
  );
  INV_X1 _22350_ (
    .A(_02166_),
    .ZN(_02167_)
  );
  AND2_X1 _22351_ (
    .A1(_02142_),
    .A2(_02167_),
    .ZN(_02168_)
  );
  INV_X1 _22352_ (
    .A(_02168_),
    .ZN(_00147_)
  );
  AND2_X1 _22353_ (
    .A1(wb_reg_wdata[31]),
    .A2(_13833_),
    .ZN(_02169_)
  );
  INV_X1 _22354_ (
    .A(_02169_),
    .ZN(_02170_)
  );
  AND2_X1 _22355_ (
    .A1(_02144_),
    .A2(_02156_),
    .ZN(_02171_)
  );
  INV_X1 _22356_ (
    .A(_02171_),
    .ZN(_02172_)
  );
  AND2_X1 _22357_ (
    .A1(mem_reg_pc[31]),
    .A2(_01880_),
    .ZN(_02173_)
  );
  INV_X1 _22358_ (
    .A(_02173_),
    .ZN(_02174_)
  );
  AND2_X1 _22359_ (
    .A1(_08042_),
    .A2(_01879_),
    .ZN(_02175_)
  );
  INV_X1 _22360_ (
    .A(_02175_),
    .ZN(_02176_)
  );
  AND2_X1 _22361_ (
    .A1(mem_reg_pc[31]),
    .A2(_01879_),
    .ZN(_02177_)
  );
  INV_X1 _22362_ (
    .A(_02177_),
    .ZN(_02178_)
  );
  AND2_X1 _22363_ (
    .A1(_08042_),
    .A2(_01880_),
    .ZN(_02179_)
  );
  INV_X1 _22364_ (
    .A(_02179_),
    .ZN(_02180_)
  );
  AND2_X1 _22365_ (
    .A1(_02174_),
    .A2(_02176_),
    .ZN(_02181_)
  );
  AND2_X1 _22366_ (
    .A1(_02178_),
    .A2(_02180_),
    .ZN(_02182_)
  );
  AND2_X1 _22367_ (
    .A1(_02171_),
    .A2(_02182_),
    .ZN(_02183_)
  );
  INV_X1 _22368_ (
    .A(_02183_),
    .ZN(_02184_)
  );
  AND2_X1 _22369_ (
    .A1(_02172_),
    .A2(_02181_),
    .ZN(_02185_)
  );
  INV_X1 _22370_ (
    .A(_02185_),
    .ZN(_02186_)
  );
  AND2_X1 _22371_ (
    .A1(_02171_),
    .A2(_02181_),
    .ZN(_02187_)
  );
  INV_X1 _22372_ (
    .A(_02187_),
    .ZN(_02188_)
  );
  AND2_X1 _22373_ (
    .A1(_02172_),
    .A2(_02182_),
    .ZN(_02189_)
  );
  INV_X1 _22374_ (
    .A(_02189_),
    .ZN(_02190_)
  );
  AND2_X1 _22375_ (
    .A1(_02184_),
    .A2(_02186_),
    .ZN(_02191_)
  );
  AND2_X1 _22376_ (
    .A1(_02188_),
    .A2(_02190_),
    .ZN(_02192_)
  );
  AND2_X1 _22377_ (
    .A1(_13852_),
    .A2(_02191_),
    .ZN(_02193_)
  );
  INV_X1 _22378_ (
    .A(_02193_),
    .ZN(_02194_)
  );
  AND2_X1 _22379_ (
    .A1(_08083_),
    .A2(_13853_),
    .ZN(_02195_)
  );
  INV_X1 _22380_ (
    .A(_02195_),
    .ZN(_02196_)
  );
  AND2_X1 _22381_ (
    .A1(_13834_),
    .A2(_02196_),
    .ZN(_02197_)
  );
  AND2_X1 _22382_ (
    .A1(_02194_),
    .A2(_02197_),
    .ZN(_02198_)
  );
  INV_X1 _22383_ (
    .A(_02198_),
    .ZN(_02199_)
  );
  AND2_X1 _22384_ (
    .A1(_02170_),
    .A2(_02199_),
    .ZN(_02200_)
  );
  INV_X1 _22385_ (
    .A(_02200_),
    .ZN(_00148_)
  );
  AND2_X1 _22386_ (
    .A1(_09691_),
    .A2(_13829_),
    .ZN(_02201_)
  );
  AND2_X1 _22387_ (
    .A1(_ex_reg_valid_T),
    .A2(_02201_),
    .ZN(_02202_)
  );
  AND2_X1 _22388_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[4]),
    .A2(_10092_),
    .ZN(_02203_)
  );
  INV_X1 _22389_ (
    .A(_02203_),
    .ZN(_02204_)
  );
  AND2_X1 _22390_ (
    .A1(_08572_),
    .A2(_10093_),
    .ZN(_02205_)
  );
  INV_X1 _22391_ (
    .A(_02205_),
    .ZN(_02206_)
  );
  AND2_X1 _22392_ (
    .A1(_02204_),
    .A2(_02206_),
    .ZN(_02207_)
  );
  AND2_X1 _22393_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[2]),
    .A2(_10090_),
    .ZN(_02208_)
  );
  INV_X1 _22394_ (
    .A(_02208_),
    .ZN(_02209_)
  );
  AND2_X1 _22395_ (
    .A1(_08546_),
    .A2(_10091_),
    .ZN(_02210_)
  );
  INV_X1 _22396_ (
    .A(_02210_),
    .ZN(_02211_)
  );
  AND2_X1 _22397_ (
    .A1(_02209_),
    .A2(_02211_),
    .ZN(_02212_)
  );
  AND2_X1 _22398_ (
    .A1(_02207_),
    .A2(_02212_),
    .ZN(_02213_)
  );
  AND2_X1 _22399_ (
    .A1(_08545_),
    .A2(_10086_),
    .ZN(_02214_)
  );
  INV_X1 _22400_ (
    .A(_02214_),
    .ZN(_02215_)
  );
  AND2_X1 _22401_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_10085_),
    .ZN(_02216_)
  );
  INV_X1 _22402_ (
    .A(_02216_),
    .ZN(_02217_)
  );
  AND2_X1 _22403_ (
    .A1(_02215_),
    .A2(_02217_),
    .ZN(_02218_)
  );
  AND2_X1 _22404_ (
    .A1(_08544_),
    .A2(_10087_),
    .ZN(_02219_)
  );
  INV_X1 _22405_ (
    .A(_02219_),
    .ZN(_02220_)
  );
  AND2_X1 _22406_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_10088_),
    .ZN(_02221_)
  );
  INV_X1 _22407_ (
    .A(_02221_),
    .ZN(_02222_)
  );
  AND2_X1 _22408_ (
    .A1(_02220_),
    .A2(_02222_),
    .ZN(_02223_)
  );
  AND2_X1 _22409_ (
    .A1(_02218_),
    .A2(_02223_),
    .ZN(_02224_)
  );
  AND2_X1 _22410_ (
    .A1(_08547_),
    .A2(_10095_),
    .ZN(_02225_)
  );
  INV_X1 _22411_ (
    .A(_02225_),
    .ZN(_02226_)
  );
  AND2_X1 _22412_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_10094_),
    .ZN(_02227_)
  );
  INV_X1 _22413_ (
    .A(_02227_),
    .ZN(_02228_)
  );
  AND2_X1 _22414_ (
    .A1(_02226_),
    .A2(_02228_),
    .ZN(_02229_)
  );
  INV_X1 _22415_ (
    .A(_02229_),
    .ZN(_02230_)
  );
  AND2_X1 _22416_ (
    .A1(_02224_),
    .A2(_02230_),
    .ZN(_02231_)
  );
  AND2_X1 _22417_ (
    .A1(_02213_),
    .A2(_02231_),
    .ZN(_02232_)
  );
  AND2_X1 _22418_ (
    .A1(_10100_),
    .A2(_02232_),
    .ZN(_02233_)
  );
  INV_X1 _22419_ (
    .A(_02233_),
    .ZN(_02234_)
  );
  MUX2_X1 _22420_ (
    .A(\rf[7] [2]),
    .B(\rf[3] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02235_)
  );
  AND2_X1 _22421_ (
    .A1(_08545_),
    .A2(_02235_),
    .ZN(_02236_)
  );
  INV_X1 _22422_ (
    .A(_02236_),
    .ZN(_02237_)
  );
  MUX2_X1 _22423_ (
    .A(\rf[5] [2]),
    .B(\rf[1] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02238_)
  );
  AND2_X1 _22424_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02238_),
    .ZN(_02239_)
  );
  INV_X1 _22425_ (
    .A(_02239_),
    .ZN(_02240_)
  );
  AND2_X1 _22426_ (
    .A1(_08544_),
    .A2(_02240_),
    .ZN(_02241_)
  );
  AND2_X1 _22427_ (
    .A1(_02237_),
    .A2(_02241_),
    .ZN(_02242_)
  );
  INV_X1 _22428_ (
    .A(_02242_),
    .ZN(_02243_)
  );
  MUX2_X1 _22429_ (
    .A(\rf[6] [2]),
    .B(\rf[2] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02244_)
  );
  AND2_X1 _22430_ (
    .A1(_08545_),
    .A2(_02244_),
    .ZN(_02245_)
  );
  INV_X1 _22431_ (
    .A(_02245_),
    .ZN(_02246_)
  );
  MUX2_X1 _22432_ (
    .A(\rf[4] [2]),
    .B(\rf[0] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02247_)
  );
  AND2_X1 _22433_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02247_),
    .ZN(_02248_)
  );
  INV_X1 _22434_ (
    .A(_02248_),
    .ZN(_02249_)
  );
  AND2_X1 _22435_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_02249_),
    .ZN(_02250_)
  );
  AND2_X1 _22436_ (
    .A1(_02246_),
    .A2(_02250_),
    .ZN(_02251_)
  );
  INV_X1 _22437_ (
    .A(_02251_),
    .ZN(_02252_)
  );
  AND2_X1 _22438_ (
    .A1(_02243_),
    .A2(_02252_),
    .ZN(_02253_)
  );
  AND2_X1 _22439_ (
    .A1(\rf[14] [2]),
    .A2(_08545_),
    .ZN(_02254_)
  );
  INV_X1 _22440_ (
    .A(_02254_),
    .ZN(_02255_)
  );
  AND2_X1 _22441_ (
    .A1(\rf[12] [2]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_02256_)
  );
  INV_X1 _22442_ (
    .A(_02256_),
    .ZN(_02257_)
  );
  AND2_X1 _22443_ (
    .A1(_08546_),
    .A2(_02257_),
    .ZN(_02258_)
  );
  AND2_X1 _22444_ (
    .A1(_02255_),
    .A2(_02258_),
    .ZN(_02259_)
  );
  INV_X1 _22445_ (
    .A(_02259_),
    .ZN(_02260_)
  );
  AND2_X1 _22446_ (
    .A1(\rf[10] [2]),
    .A2(_08545_),
    .ZN(_02261_)
  );
  INV_X1 _22447_ (
    .A(_02261_),
    .ZN(_02262_)
  );
  AND2_X1 _22448_ (
    .A1(\rf[8] [2]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_02263_)
  );
  INV_X1 _22449_ (
    .A(_02263_),
    .ZN(_02264_)
  );
  AND2_X1 _22450_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[2]),
    .A2(_02264_),
    .ZN(_02265_)
  );
  AND2_X1 _22451_ (
    .A1(_02262_),
    .A2(_02265_),
    .ZN(_02266_)
  );
  INV_X1 _22452_ (
    .A(_02266_),
    .ZN(_02267_)
  );
  AND2_X1 _22453_ (
    .A1(_02260_),
    .A2(_02267_),
    .ZN(_02268_)
  );
  AND2_X1 _22454_ (
    .A1(\rf[15] [2]),
    .A2(_08545_),
    .ZN(_02269_)
  );
  INV_X1 _22455_ (
    .A(_02269_),
    .ZN(_02270_)
  );
  AND2_X1 _22456_ (
    .A1(\rf[13] [2]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_02271_)
  );
  INV_X1 _22457_ (
    .A(_02271_),
    .ZN(_02272_)
  );
  AND2_X1 _22458_ (
    .A1(_08546_),
    .A2(_02272_),
    .ZN(_02273_)
  );
  AND2_X1 _22459_ (
    .A1(_02270_),
    .A2(_02273_),
    .ZN(_02274_)
  );
  INV_X1 _22460_ (
    .A(_02274_),
    .ZN(_02275_)
  );
  AND2_X1 _22461_ (
    .A1(\rf[11] [2]),
    .A2(_08545_),
    .ZN(_02276_)
  );
  INV_X1 _22462_ (
    .A(_02276_),
    .ZN(_02277_)
  );
  AND2_X1 _22463_ (
    .A1(\rf[9] [2]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_02278_)
  );
  INV_X1 _22464_ (
    .A(_02278_),
    .ZN(_02279_)
  );
  AND2_X1 _22465_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[2]),
    .A2(_02279_),
    .ZN(_02280_)
  );
  AND2_X1 _22466_ (
    .A1(_02277_),
    .A2(_02280_),
    .ZN(_02281_)
  );
  INV_X1 _22467_ (
    .A(_02281_),
    .ZN(_02282_)
  );
  AND2_X1 _22468_ (
    .A1(_02275_),
    .A2(_02282_),
    .ZN(_02283_)
  );
  MUX2_X1 _22469_ (
    .A(_02268_),
    .B(_02283_),
    .S(_08544_),
    .Z(_02284_)
  );
  MUX2_X1 _22470_ (
    .A(_02253_),
    .B(_02284_),
    .S(_08547_),
    .Z(_02285_)
  );
  AND2_X1 _22471_ (
    .A1(\rf[26] [2]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02286_)
  );
  INV_X1 _22472_ (
    .A(_02286_),
    .ZN(_02287_)
  );
  AND2_X1 _22473_ (
    .A1(\rf[30] [2]),
    .A2(_08546_),
    .ZN(_02288_)
  );
  INV_X1 _22474_ (
    .A(_02288_),
    .ZN(_02289_)
  );
  AND2_X1 _22475_ (
    .A1(_08545_),
    .A2(_02289_),
    .ZN(_02290_)
  );
  AND2_X1 _22476_ (
    .A1(_02287_),
    .A2(_02290_),
    .ZN(_02291_)
  );
  INV_X1 _22477_ (
    .A(_02291_),
    .ZN(_02292_)
  );
  AND2_X1 _22478_ (
    .A1(\rf[24] [2]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02293_)
  );
  INV_X1 _22479_ (
    .A(_02293_),
    .ZN(_02294_)
  );
  AND2_X1 _22480_ (
    .A1(\rf[28] [2]),
    .A2(_08546_),
    .ZN(_02295_)
  );
  INV_X1 _22481_ (
    .A(_02295_),
    .ZN(_02296_)
  );
  AND2_X1 _22482_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02296_),
    .ZN(_02297_)
  );
  AND2_X1 _22483_ (
    .A1(_02294_),
    .A2(_02297_),
    .ZN(_02298_)
  );
  INV_X1 _22484_ (
    .A(_02298_),
    .ZN(_02299_)
  );
  AND2_X1 _22485_ (
    .A1(_02292_),
    .A2(_02299_),
    .ZN(_02300_)
  );
  MUX2_X1 _22486_ (
    .A(\rf[29] [2]),
    .B(\rf[25] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02301_)
  );
  AND2_X1 _22487_ (
    .A1(\rf[27] [2]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02302_)
  );
  MUX2_X1 _22488_ (
    .A(_02301_),
    .B(_02302_),
    .S(_08545_),
    .Z(_02303_)
  );
  MUX2_X1 _22489_ (
    .A(_02300_),
    .B(_02303_),
    .S(_08544_),
    .Z(_02304_)
  );
  AND2_X1 _22490_ (
    .A1(_08375_),
    .A2(_08546_),
    .ZN(_02305_)
  );
  INV_X1 _22491_ (
    .A(_02305_),
    .ZN(_02306_)
  );
  AND2_X1 _22492_ (
    .A1(_08276_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02307_)
  );
  INV_X1 _22493_ (
    .A(_02307_),
    .ZN(_02308_)
  );
  AND2_X1 _22494_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02308_),
    .ZN(_02309_)
  );
  AND2_X1 _22495_ (
    .A1(_02306_),
    .A2(_02309_),
    .ZN(_02310_)
  );
  INV_X1 _22496_ (
    .A(_02310_),
    .ZN(_02311_)
  );
  MUX2_X1 _22497_ (
    .A(\rf[22] [2]),
    .B(\rf[18] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02312_)
  );
  AND2_X1 _22498_ (
    .A1(_08545_),
    .A2(_02312_),
    .ZN(_02313_)
  );
  INV_X1 _22499_ (
    .A(_02313_),
    .ZN(_02314_)
  );
  AND2_X1 _22500_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_02314_),
    .ZN(_02315_)
  );
  AND2_X1 _22501_ (
    .A1(_02311_),
    .A2(_02315_),
    .ZN(_02316_)
  );
  INV_X1 _22502_ (
    .A(_02316_),
    .ZN(_02317_)
  );
  AND2_X1 _22503_ (
    .A1(_08306_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02318_)
  );
  INV_X1 _22504_ (
    .A(_02318_),
    .ZN(_02319_)
  );
  AND2_X1 _22505_ (
    .A1(_08405_),
    .A2(_08546_),
    .ZN(_02320_)
  );
  INV_X1 _22506_ (
    .A(_02320_),
    .ZN(_02321_)
  );
  AND2_X1 _22507_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02321_),
    .ZN(_02322_)
  );
  AND2_X1 _22508_ (
    .A1(_02319_),
    .A2(_02322_),
    .ZN(_02323_)
  );
  INV_X1 _22509_ (
    .A(_02323_),
    .ZN(_02324_)
  );
  MUX2_X1 _22510_ (
    .A(\rf[23] [2]),
    .B(\rf[19] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02325_)
  );
  AND2_X1 _22511_ (
    .A1(_08545_),
    .A2(_02325_),
    .ZN(_02326_)
  );
  INV_X1 _22512_ (
    .A(_02326_),
    .ZN(_02327_)
  );
  AND2_X1 _22513_ (
    .A1(_08544_),
    .A2(_02327_),
    .ZN(_02328_)
  );
  AND2_X1 _22514_ (
    .A1(_02324_),
    .A2(_02328_),
    .ZN(_02329_)
  );
  INV_X1 _22515_ (
    .A(_02329_),
    .ZN(_02330_)
  );
  AND2_X1 _22516_ (
    .A1(_02317_),
    .A2(_02330_),
    .ZN(_02331_)
  );
  MUX2_X1 _22517_ (
    .A(_02304_),
    .B(_02331_),
    .S(ibuf_io_inst_0_bits_inst_rs2[3]),
    .Z(_02332_)
  );
  MUX2_X1 _22518_ (
    .A(_02285_),
    .B(_02332_),
    .S(_08572_),
    .Z(_02333_)
  );
  MUX2_X1 _22519_ (
    .A(_02333_),
    .B(_10137_),
    .S(_02233_),
    .Z(_02334_)
  );
  MUX2_X1 _22520_ (
    .A(ex_reg_rs_msb_1[0]),
    .B(_02334_),
    .S(_02202_),
    .Z(_00149_)
  );
  MUX2_X1 _22521_ (
    .A(\rf[3] [3]),
    .B(\rf[2] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_02335_)
  );
  MUX2_X1 _22522_ (
    .A(\rf[7] [3]),
    .B(\rf[6] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_02336_)
  );
  MUX2_X1 _22523_ (
    .A(_02335_),
    .B(_02336_),
    .S(_08546_),
    .Z(_02337_)
  );
  INV_X1 _22524_ (
    .A(_02337_),
    .ZN(_02338_)
  );
  AND2_X1 _22525_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_02338_),
    .ZN(_02339_)
  );
  INV_X1 _22526_ (
    .A(_02339_),
    .ZN(_02340_)
  );
  AND2_X1 _22527_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08547_),
    .ZN(_02341_)
  );
  MUX2_X1 _22528_ (
    .A(\rf[14] [3]),
    .B(\rf[10] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02342_)
  );
  INV_X1 _22529_ (
    .A(_02342_),
    .ZN(_02343_)
  );
  AND2_X1 _22530_ (
    .A1(_02341_),
    .A2(_02343_),
    .ZN(_02344_)
  );
  INV_X1 _22531_ (
    .A(_02344_),
    .ZN(_02345_)
  );
  MUX2_X1 _22532_ (
    .A(\rf[15] [3]),
    .B(\rf[11] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02346_)
  );
  INV_X1 _22533_ (
    .A(_02346_),
    .ZN(_02347_)
  );
  AND2_X1 _22534_ (
    .A1(_09692_),
    .A2(_02347_),
    .ZN(_02348_)
  );
  INV_X1 _22535_ (
    .A(_02348_),
    .ZN(_02349_)
  );
  AND2_X1 _22536_ (
    .A1(_02345_),
    .A2(_02349_),
    .ZN(_02350_)
  );
  AND2_X1 _22537_ (
    .A1(_08545_),
    .A2(_02350_),
    .ZN(_02351_)
  );
  AND2_X1 _22538_ (
    .A1(_02340_),
    .A2(_02351_),
    .ZN(_02352_)
  );
  INV_X1 _22539_ (
    .A(_02352_),
    .ZN(_02353_)
  );
  MUX2_X1 _22540_ (
    .A(\rf[1] [3]),
    .B(\rf[0] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_02354_)
  );
  MUX2_X1 _22541_ (
    .A(\rf[5] [3]),
    .B(\rf[4] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_02355_)
  );
  MUX2_X1 _22542_ (
    .A(_02354_),
    .B(_02355_),
    .S(_08546_),
    .Z(_02356_)
  );
  INV_X1 _22543_ (
    .A(_02356_),
    .ZN(_02357_)
  );
  AND2_X1 _22544_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_02357_),
    .ZN(_02358_)
  );
  INV_X1 _22545_ (
    .A(_02358_),
    .ZN(_02359_)
  );
  MUX2_X1 _22546_ (
    .A(\rf[12] [3]),
    .B(\rf[8] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02360_)
  );
  INV_X1 _22547_ (
    .A(_02360_),
    .ZN(_02361_)
  );
  AND2_X1 _22548_ (
    .A1(_02341_),
    .A2(_02361_),
    .ZN(_02362_)
  );
  INV_X1 _22549_ (
    .A(_02362_),
    .ZN(_02363_)
  );
  MUX2_X1 _22550_ (
    .A(\rf[13] [3]),
    .B(\rf[9] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02364_)
  );
  INV_X1 _22551_ (
    .A(_02364_),
    .ZN(_02365_)
  );
  AND2_X1 _22552_ (
    .A1(_09692_),
    .A2(_02365_),
    .ZN(_02366_)
  );
  INV_X1 _22553_ (
    .A(_02366_),
    .ZN(_02367_)
  );
  AND2_X1 _22554_ (
    .A1(_02363_),
    .A2(_02367_),
    .ZN(_02368_)
  );
  AND2_X1 _22555_ (
    .A1(_02359_),
    .A2(_02368_),
    .ZN(_02369_)
  );
  AND2_X1 _22556_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02369_),
    .ZN(_02370_)
  );
  INV_X1 _22557_ (
    .A(_02370_),
    .ZN(_02371_)
  );
  AND2_X1 _22558_ (
    .A1(_02353_),
    .A2(_02371_),
    .ZN(_02372_)
  );
  AND2_X1 _22559_ (
    .A1(_08307_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02373_)
  );
  INV_X1 _22560_ (
    .A(_02373_),
    .ZN(_02374_)
  );
  AND2_X1 _22561_ (
    .A1(_08406_),
    .A2(_08546_),
    .ZN(_02375_)
  );
  INV_X1 _22562_ (
    .A(_02375_),
    .ZN(_02376_)
  );
  AND2_X1 _22563_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02376_),
    .ZN(_02377_)
  );
  AND2_X1 _22564_ (
    .A1(_02374_),
    .A2(_02377_),
    .ZN(_02378_)
  );
  INV_X1 _22565_ (
    .A(_02378_),
    .ZN(_02379_)
  );
  MUX2_X1 _22566_ (
    .A(\rf[23] [3]),
    .B(\rf[19] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02380_)
  );
  AND2_X1 _22567_ (
    .A1(_08545_),
    .A2(_02380_),
    .ZN(_02381_)
  );
  INV_X1 _22568_ (
    .A(_02381_),
    .ZN(_02382_)
  );
  AND2_X1 _22569_ (
    .A1(_08544_),
    .A2(_02382_),
    .ZN(_02383_)
  );
  AND2_X1 _22570_ (
    .A1(_02379_),
    .A2(_02383_),
    .ZN(_02384_)
  );
  INV_X1 _22571_ (
    .A(_02384_),
    .ZN(_02385_)
  );
  AND2_X1 _22572_ (
    .A1(_08376_),
    .A2(_08546_),
    .ZN(_02386_)
  );
  INV_X1 _22573_ (
    .A(_02386_),
    .ZN(_02387_)
  );
  AND2_X1 _22574_ (
    .A1(_08277_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02388_)
  );
  INV_X1 _22575_ (
    .A(_02388_),
    .ZN(_02389_)
  );
  AND2_X1 _22576_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02389_),
    .ZN(_02390_)
  );
  AND2_X1 _22577_ (
    .A1(_02387_),
    .A2(_02390_),
    .ZN(_02391_)
  );
  INV_X1 _22578_ (
    .A(_02391_),
    .ZN(_02392_)
  );
  MUX2_X1 _22579_ (
    .A(\rf[22] [3]),
    .B(\rf[18] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02393_)
  );
  AND2_X1 _22580_ (
    .A1(_08545_),
    .A2(_02393_),
    .ZN(_02394_)
  );
  INV_X1 _22581_ (
    .A(_02394_),
    .ZN(_02395_)
  );
  AND2_X1 _22582_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_02395_),
    .ZN(_02396_)
  );
  AND2_X1 _22583_ (
    .A1(_02392_),
    .A2(_02396_),
    .ZN(_02397_)
  );
  INV_X1 _22584_ (
    .A(_02397_),
    .ZN(_02398_)
  );
  AND2_X1 _22585_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_02385_),
    .ZN(_02399_)
  );
  AND2_X1 _22586_ (
    .A1(_02398_),
    .A2(_02399_),
    .ZN(_02400_)
  );
  INV_X1 _22587_ (
    .A(_02400_),
    .ZN(_02401_)
  );
  AND2_X1 _22588_ (
    .A1(_08436_),
    .A2(_08546_),
    .ZN(_02402_)
  );
  INV_X1 _22589_ (
    .A(_02402_),
    .ZN(_02403_)
  );
  AND2_X1 _22590_ (
    .A1(_08506_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02404_)
  );
  INV_X1 _22591_ (
    .A(_02404_),
    .ZN(_02405_)
  );
  AND2_X1 _22592_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02405_),
    .ZN(_02406_)
  );
  AND2_X1 _22593_ (
    .A1(_02403_),
    .A2(_02406_),
    .ZN(_02407_)
  );
  INV_X1 _22594_ (
    .A(_02407_),
    .ZN(_02408_)
  );
  MUX2_X1 _22595_ (
    .A(\rf[30] [3]),
    .B(\rf[26] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02409_)
  );
  AND2_X1 _22596_ (
    .A1(_08545_),
    .A2(_02409_),
    .ZN(_02410_)
  );
  INV_X1 _22597_ (
    .A(_02410_),
    .ZN(_02411_)
  );
  AND2_X1 _22598_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_02411_),
    .ZN(_02412_)
  );
  AND2_X1 _22599_ (
    .A1(_02408_),
    .A2(_02412_),
    .ZN(_02413_)
  );
  INV_X1 _22600_ (
    .A(_02413_),
    .ZN(_02414_)
  );
  MUX2_X1 _22601_ (
    .A(\rf[29] [3]),
    .B(\rf[25] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02415_)
  );
  AND2_X1 _22602_ (
    .A1(\rf[27] [3]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02416_)
  );
  MUX2_X1 _22603_ (
    .A(_02415_),
    .B(_02416_),
    .S(_08545_),
    .Z(_02417_)
  );
  INV_X1 _22604_ (
    .A(_02417_),
    .ZN(_02418_)
  );
  AND2_X1 _22605_ (
    .A1(_08544_),
    .A2(_02418_),
    .ZN(_02419_)
  );
  INV_X1 _22606_ (
    .A(_02419_),
    .ZN(_02420_)
  );
  AND2_X1 _22607_ (
    .A1(_08547_),
    .A2(_02420_),
    .ZN(_02421_)
  );
  AND2_X1 _22608_ (
    .A1(_02414_),
    .A2(_02421_),
    .ZN(_02422_)
  );
  INV_X1 _22609_ (
    .A(_02422_),
    .ZN(_02423_)
  );
  AND2_X1 _22610_ (
    .A1(_02401_),
    .A2(_02423_),
    .ZN(_02424_)
  );
  MUX2_X1 _22611_ (
    .A(_02372_),
    .B(_02424_),
    .S(_08572_),
    .Z(_02425_)
  );
  INV_X1 _22612_ (
    .A(_02425_),
    .ZN(_02426_)
  );
  MUX2_X1 _22613_ (
    .A(_02426_),
    .B(_10250_),
    .S(_02233_),
    .Z(_02427_)
  );
  MUX2_X1 _22614_ (
    .A(ex_reg_rs_msb_1[1]),
    .B(_02427_),
    .S(_02202_),
    .Z(_00150_)
  );
  MUX2_X1 _22615_ (
    .A(\rf[3] [4]),
    .B(\rf[2] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_02428_)
  );
  MUX2_X1 _22616_ (
    .A(\rf[7] [4]),
    .B(\rf[6] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_02429_)
  );
  MUX2_X1 _22617_ (
    .A(_02428_),
    .B(_02429_),
    .S(_08546_),
    .Z(_02430_)
  );
  INV_X1 _22618_ (
    .A(_02430_),
    .ZN(_02431_)
  );
  AND2_X1 _22619_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_02431_),
    .ZN(_02432_)
  );
  INV_X1 _22620_ (
    .A(_02432_),
    .ZN(_02433_)
  );
  MUX2_X1 _22621_ (
    .A(\rf[14] [4]),
    .B(\rf[10] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02434_)
  );
  INV_X1 _22622_ (
    .A(_02434_),
    .ZN(_02435_)
  );
  AND2_X1 _22623_ (
    .A1(_02341_),
    .A2(_02435_),
    .ZN(_02436_)
  );
  INV_X1 _22624_ (
    .A(_02436_),
    .ZN(_02437_)
  );
  MUX2_X1 _22625_ (
    .A(\rf[15] [4]),
    .B(\rf[11] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02438_)
  );
  INV_X1 _22626_ (
    .A(_02438_),
    .ZN(_02439_)
  );
  AND2_X1 _22627_ (
    .A1(_09692_),
    .A2(_02439_),
    .ZN(_02440_)
  );
  INV_X1 _22628_ (
    .A(_02440_),
    .ZN(_02441_)
  );
  AND2_X1 _22629_ (
    .A1(_02437_),
    .A2(_02441_),
    .ZN(_02442_)
  );
  AND2_X1 _22630_ (
    .A1(_08545_),
    .A2(_02442_),
    .ZN(_02443_)
  );
  AND2_X1 _22631_ (
    .A1(_02433_),
    .A2(_02443_),
    .ZN(_02444_)
  );
  INV_X1 _22632_ (
    .A(_02444_),
    .ZN(_02445_)
  );
  MUX2_X1 _22633_ (
    .A(\rf[1] [4]),
    .B(\rf[0] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_02446_)
  );
  MUX2_X1 _22634_ (
    .A(\rf[5] [4]),
    .B(\rf[4] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_02447_)
  );
  MUX2_X1 _22635_ (
    .A(_02446_),
    .B(_02447_),
    .S(_08546_),
    .Z(_02448_)
  );
  INV_X1 _22636_ (
    .A(_02448_),
    .ZN(_02449_)
  );
  AND2_X1 _22637_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_02449_),
    .ZN(_02450_)
  );
  INV_X1 _22638_ (
    .A(_02450_),
    .ZN(_02451_)
  );
  MUX2_X1 _22639_ (
    .A(\rf[12] [4]),
    .B(\rf[8] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02452_)
  );
  INV_X1 _22640_ (
    .A(_02452_),
    .ZN(_02453_)
  );
  AND2_X1 _22641_ (
    .A1(_02341_),
    .A2(_02453_),
    .ZN(_02454_)
  );
  INV_X1 _22642_ (
    .A(_02454_),
    .ZN(_02455_)
  );
  MUX2_X1 _22643_ (
    .A(\rf[13] [4]),
    .B(\rf[9] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02456_)
  );
  INV_X1 _22644_ (
    .A(_02456_),
    .ZN(_02457_)
  );
  AND2_X1 _22645_ (
    .A1(_09692_),
    .A2(_02457_),
    .ZN(_02458_)
  );
  INV_X1 _22646_ (
    .A(_02458_),
    .ZN(_02459_)
  );
  AND2_X1 _22647_ (
    .A1(_02455_),
    .A2(_02459_),
    .ZN(_02460_)
  );
  AND2_X1 _22648_ (
    .A1(_02451_),
    .A2(_02460_),
    .ZN(_02461_)
  );
  AND2_X1 _22649_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02461_),
    .ZN(_02462_)
  );
  INV_X1 _22650_ (
    .A(_02462_),
    .ZN(_02463_)
  );
  AND2_X1 _22651_ (
    .A1(_02445_),
    .A2(_02463_),
    .ZN(_02464_)
  );
  AND2_X1 _22652_ (
    .A1(_08308_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02465_)
  );
  INV_X1 _22653_ (
    .A(_02465_),
    .ZN(_02466_)
  );
  AND2_X1 _22654_ (
    .A1(_08407_),
    .A2(_08546_),
    .ZN(_02467_)
  );
  INV_X1 _22655_ (
    .A(_02467_),
    .ZN(_02468_)
  );
  AND2_X1 _22656_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02468_),
    .ZN(_02469_)
  );
  AND2_X1 _22657_ (
    .A1(_02466_),
    .A2(_02469_),
    .ZN(_02470_)
  );
  INV_X1 _22658_ (
    .A(_02470_),
    .ZN(_02471_)
  );
  MUX2_X1 _22659_ (
    .A(\rf[23] [4]),
    .B(\rf[19] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02472_)
  );
  AND2_X1 _22660_ (
    .A1(_08545_),
    .A2(_02472_),
    .ZN(_02473_)
  );
  INV_X1 _22661_ (
    .A(_02473_),
    .ZN(_02474_)
  );
  AND2_X1 _22662_ (
    .A1(_08544_),
    .A2(_02474_),
    .ZN(_02475_)
  );
  AND2_X1 _22663_ (
    .A1(_02471_),
    .A2(_02475_),
    .ZN(_02476_)
  );
  INV_X1 _22664_ (
    .A(_02476_),
    .ZN(_02477_)
  );
  AND2_X1 _22665_ (
    .A1(_08377_),
    .A2(_08546_),
    .ZN(_02478_)
  );
  INV_X1 _22666_ (
    .A(_02478_),
    .ZN(_02479_)
  );
  AND2_X1 _22667_ (
    .A1(_08278_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02480_)
  );
  INV_X1 _22668_ (
    .A(_02480_),
    .ZN(_02481_)
  );
  AND2_X1 _22669_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02481_),
    .ZN(_02482_)
  );
  AND2_X1 _22670_ (
    .A1(_02479_),
    .A2(_02482_),
    .ZN(_02483_)
  );
  INV_X1 _22671_ (
    .A(_02483_),
    .ZN(_02484_)
  );
  MUX2_X1 _22672_ (
    .A(\rf[22] [4]),
    .B(\rf[18] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02485_)
  );
  AND2_X1 _22673_ (
    .A1(_08545_),
    .A2(_02485_),
    .ZN(_02486_)
  );
  INV_X1 _22674_ (
    .A(_02486_),
    .ZN(_02487_)
  );
  AND2_X1 _22675_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_02487_),
    .ZN(_02488_)
  );
  AND2_X1 _22676_ (
    .A1(_02484_),
    .A2(_02488_),
    .ZN(_02489_)
  );
  INV_X1 _22677_ (
    .A(_02489_),
    .ZN(_02490_)
  );
  AND2_X1 _22678_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_02477_),
    .ZN(_02491_)
  );
  AND2_X1 _22679_ (
    .A1(_02490_),
    .A2(_02491_),
    .ZN(_02492_)
  );
  INV_X1 _22680_ (
    .A(_02492_),
    .ZN(_02493_)
  );
  AND2_X1 _22681_ (
    .A1(_08437_),
    .A2(_08546_),
    .ZN(_02494_)
  );
  INV_X1 _22682_ (
    .A(_02494_),
    .ZN(_02495_)
  );
  AND2_X1 _22683_ (
    .A1(_08507_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02496_)
  );
  INV_X1 _22684_ (
    .A(_02496_),
    .ZN(_02497_)
  );
  AND2_X1 _22685_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02497_),
    .ZN(_02498_)
  );
  AND2_X1 _22686_ (
    .A1(_02495_),
    .A2(_02498_),
    .ZN(_02499_)
  );
  INV_X1 _22687_ (
    .A(_02499_),
    .ZN(_02500_)
  );
  MUX2_X1 _22688_ (
    .A(\rf[30] [4]),
    .B(\rf[26] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02501_)
  );
  AND2_X1 _22689_ (
    .A1(_08545_),
    .A2(_02501_),
    .ZN(_02502_)
  );
  INV_X1 _22690_ (
    .A(_02502_),
    .ZN(_02503_)
  );
  AND2_X1 _22691_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_02503_),
    .ZN(_02504_)
  );
  AND2_X1 _22692_ (
    .A1(_02500_),
    .A2(_02504_),
    .ZN(_02505_)
  );
  INV_X1 _22693_ (
    .A(_02505_),
    .ZN(_02506_)
  );
  MUX2_X1 _22694_ (
    .A(\rf[29] [4]),
    .B(\rf[25] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02507_)
  );
  AND2_X1 _22695_ (
    .A1(\rf[27] [4]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02508_)
  );
  MUX2_X1 _22696_ (
    .A(_02507_),
    .B(_02508_),
    .S(_08545_),
    .Z(_02509_)
  );
  INV_X1 _22697_ (
    .A(_02509_),
    .ZN(_02510_)
  );
  AND2_X1 _22698_ (
    .A1(_08544_),
    .A2(_02510_),
    .ZN(_02511_)
  );
  INV_X1 _22699_ (
    .A(_02511_),
    .ZN(_02512_)
  );
  AND2_X1 _22700_ (
    .A1(_08547_),
    .A2(_02512_),
    .ZN(_02513_)
  );
  AND2_X1 _22701_ (
    .A1(_02506_),
    .A2(_02513_),
    .ZN(_02514_)
  );
  INV_X1 _22702_ (
    .A(_02514_),
    .ZN(_02515_)
  );
  AND2_X1 _22703_ (
    .A1(_02493_),
    .A2(_02515_),
    .ZN(_02516_)
  );
  MUX2_X1 _22704_ (
    .A(_02464_),
    .B(_02516_),
    .S(_08572_),
    .Z(_02517_)
  );
  INV_X1 _22705_ (
    .A(_02517_),
    .ZN(_02518_)
  );
  MUX2_X1 _22706_ (
    .A(_02518_),
    .B(_10389_),
    .S(_02233_),
    .Z(_02519_)
  );
  MUX2_X1 _22707_ (
    .A(ex_reg_rs_msb_1[2]),
    .B(_02519_),
    .S(_02202_),
    .Z(_00151_)
  );
  MUX2_X1 _22708_ (
    .A(\rf[7] [5]),
    .B(\rf[3] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02520_)
  );
  AND2_X1 _22709_ (
    .A1(_08545_),
    .A2(_02520_),
    .ZN(_02521_)
  );
  INV_X1 _22710_ (
    .A(_02521_),
    .ZN(_02522_)
  );
  MUX2_X1 _22711_ (
    .A(\rf[5] [5]),
    .B(\rf[1] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02523_)
  );
  AND2_X1 _22712_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02523_),
    .ZN(_02524_)
  );
  INV_X1 _22713_ (
    .A(_02524_),
    .ZN(_02525_)
  );
  AND2_X1 _22714_ (
    .A1(_08544_),
    .A2(_02525_),
    .ZN(_02526_)
  );
  AND2_X1 _22715_ (
    .A1(_02522_),
    .A2(_02526_),
    .ZN(_02527_)
  );
  INV_X1 _22716_ (
    .A(_02527_),
    .ZN(_02528_)
  );
  MUX2_X1 _22717_ (
    .A(\rf[6] [5]),
    .B(\rf[2] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02529_)
  );
  AND2_X1 _22718_ (
    .A1(_08545_),
    .A2(_02529_),
    .ZN(_02530_)
  );
  INV_X1 _22719_ (
    .A(_02530_),
    .ZN(_02531_)
  );
  MUX2_X1 _22720_ (
    .A(\rf[4] [5]),
    .B(\rf[0] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02532_)
  );
  AND2_X1 _22721_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02532_),
    .ZN(_02533_)
  );
  INV_X1 _22722_ (
    .A(_02533_),
    .ZN(_02534_)
  );
  AND2_X1 _22723_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_02534_),
    .ZN(_02535_)
  );
  AND2_X1 _22724_ (
    .A1(_02531_),
    .A2(_02535_),
    .ZN(_02536_)
  );
  INV_X1 _22725_ (
    .A(_02536_),
    .ZN(_02537_)
  );
  AND2_X1 _22726_ (
    .A1(_02528_),
    .A2(_02537_),
    .ZN(_02538_)
  );
  AND2_X1 _22727_ (
    .A1(\rf[14] [5]),
    .A2(_08545_),
    .ZN(_02539_)
  );
  INV_X1 _22728_ (
    .A(_02539_),
    .ZN(_02540_)
  );
  AND2_X1 _22729_ (
    .A1(\rf[12] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_02541_)
  );
  INV_X1 _22730_ (
    .A(_02541_),
    .ZN(_02542_)
  );
  AND2_X1 _22731_ (
    .A1(_08546_),
    .A2(_02542_),
    .ZN(_02543_)
  );
  AND2_X1 _22732_ (
    .A1(_02540_),
    .A2(_02543_),
    .ZN(_02544_)
  );
  INV_X1 _22733_ (
    .A(_02544_),
    .ZN(_02545_)
  );
  AND2_X1 _22734_ (
    .A1(\rf[10] [5]),
    .A2(_08545_),
    .ZN(_02546_)
  );
  INV_X1 _22735_ (
    .A(_02546_),
    .ZN(_02547_)
  );
  AND2_X1 _22736_ (
    .A1(\rf[8] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_02548_)
  );
  INV_X1 _22737_ (
    .A(_02548_),
    .ZN(_02549_)
  );
  AND2_X1 _22738_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[2]),
    .A2(_02549_),
    .ZN(_02550_)
  );
  AND2_X1 _22739_ (
    .A1(_02547_),
    .A2(_02550_),
    .ZN(_02551_)
  );
  INV_X1 _22740_ (
    .A(_02551_),
    .ZN(_02552_)
  );
  AND2_X1 _22741_ (
    .A1(_02545_),
    .A2(_02552_),
    .ZN(_02553_)
  );
  AND2_X1 _22742_ (
    .A1(\rf[15] [5]),
    .A2(_08545_),
    .ZN(_02554_)
  );
  INV_X1 _22743_ (
    .A(_02554_),
    .ZN(_02555_)
  );
  AND2_X1 _22744_ (
    .A1(\rf[13] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_02556_)
  );
  INV_X1 _22745_ (
    .A(_02556_),
    .ZN(_02557_)
  );
  AND2_X1 _22746_ (
    .A1(_08546_),
    .A2(_02557_),
    .ZN(_02558_)
  );
  AND2_X1 _22747_ (
    .A1(_02555_),
    .A2(_02558_),
    .ZN(_02559_)
  );
  INV_X1 _22748_ (
    .A(_02559_),
    .ZN(_02560_)
  );
  AND2_X1 _22749_ (
    .A1(\rf[11] [5]),
    .A2(_08545_),
    .ZN(_02561_)
  );
  INV_X1 _22750_ (
    .A(_02561_),
    .ZN(_02562_)
  );
  AND2_X1 _22751_ (
    .A1(\rf[9] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_02563_)
  );
  INV_X1 _22752_ (
    .A(_02563_),
    .ZN(_02564_)
  );
  AND2_X1 _22753_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[2]),
    .A2(_02564_),
    .ZN(_02565_)
  );
  AND2_X1 _22754_ (
    .A1(_02562_),
    .A2(_02565_),
    .ZN(_02566_)
  );
  INV_X1 _22755_ (
    .A(_02566_),
    .ZN(_02567_)
  );
  AND2_X1 _22756_ (
    .A1(_02560_),
    .A2(_02567_),
    .ZN(_02568_)
  );
  MUX2_X1 _22757_ (
    .A(_02553_),
    .B(_02568_),
    .S(_08544_),
    .Z(_02569_)
  );
  MUX2_X1 _22758_ (
    .A(_02538_),
    .B(_02569_),
    .S(_08547_),
    .Z(_02570_)
  );
  AND2_X1 _22759_ (
    .A1(\rf[30] [5]),
    .A2(_08546_),
    .ZN(_02571_)
  );
  INV_X1 _22760_ (
    .A(_02571_),
    .ZN(_02572_)
  );
  AND2_X1 _22761_ (
    .A1(\rf[26] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02573_)
  );
  INV_X1 _22762_ (
    .A(_02573_),
    .ZN(_02574_)
  );
  AND2_X1 _22763_ (
    .A1(_08545_),
    .A2(_02574_),
    .ZN(_02575_)
  );
  AND2_X1 _22764_ (
    .A1(_02572_),
    .A2(_02575_),
    .ZN(_02576_)
  );
  INV_X1 _22765_ (
    .A(_02576_),
    .ZN(_02577_)
  );
  AND2_X1 _22766_ (
    .A1(\rf[24] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02578_)
  );
  INV_X1 _22767_ (
    .A(_02578_),
    .ZN(_02579_)
  );
  AND2_X1 _22768_ (
    .A1(\rf[28] [5]),
    .A2(_08546_),
    .ZN(_02580_)
  );
  INV_X1 _22769_ (
    .A(_02580_),
    .ZN(_02581_)
  );
  AND2_X1 _22770_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02581_),
    .ZN(_02582_)
  );
  AND2_X1 _22771_ (
    .A1(_02579_),
    .A2(_02582_),
    .ZN(_02583_)
  );
  INV_X1 _22772_ (
    .A(_02583_),
    .ZN(_02584_)
  );
  AND2_X1 _22773_ (
    .A1(_02577_),
    .A2(_02584_),
    .ZN(_02585_)
  );
  MUX2_X1 _22774_ (
    .A(\rf[29] [5]),
    .B(\rf[25] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02586_)
  );
  AND2_X1 _22775_ (
    .A1(\rf[27] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02587_)
  );
  MUX2_X1 _22776_ (
    .A(_02586_),
    .B(_02587_),
    .S(_08545_),
    .Z(_02588_)
  );
  MUX2_X1 _22777_ (
    .A(_02585_),
    .B(_02588_),
    .S(_08544_),
    .Z(_02589_)
  );
  AND2_X1 _22778_ (
    .A1(_08378_),
    .A2(_08546_),
    .ZN(_02590_)
  );
  INV_X1 _22779_ (
    .A(_02590_),
    .ZN(_02591_)
  );
  AND2_X1 _22780_ (
    .A1(_08279_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02592_)
  );
  INV_X1 _22781_ (
    .A(_02592_),
    .ZN(_02593_)
  );
  AND2_X1 _22782_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02593_),
    .ZN(_02594_)
  );
  AND2_X1 _22783_ (
    .A1(_02591_),
    .A2(_02594_),
    .ZN(_02595_)
  );
  INV_X1 _22784_ (
    .A(_02595_),
    .ZN(_02596_)
  );
  MUX2_X1 _22785_ (
    .A(\rf[22] [5]),
    .B(\rf[18] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02597_)
  );
  AND2_X1 _22786_ (
    .A1(_08545_),
    .A2(_02597_),
    .ZN(_02598_)
  );
  INV_X1 _22787_ (
    .A(_02598_),
    .ZN(_02599_)
  );
  AND2_X1 _22788_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_02599_),
    .ZN(_02600_)
  );
  AND2_X1 _22789_ (
    .A1(_02596_),
    .A2(_02600_),
    .ZN(_02601_)
  );
  INV_X1 _22790_ (
    .A(_02601_),
    .ZN(_02602_)
  );
  AND2_X1 _22791_ (
    .A1(_08309_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02603_)
  );
  INV_X1 _22792_ (
    .A(_02603_),
    .ZN(_02604_)
  );
  AND2_X1 _22793_ (
    .A1(_08408_),
    .A2(_08546_),
    .ZN(_02605_)
  );
  INV_X1 _22794_ (
    .A(_02605_),
    .ZN(_02606_)
  );
  AND2_X1 _22795_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02606_),
    .ZN(_02607_)
  );
  AND2_X1 _22796_ (
    .A1(_02604_),
    .A2(_02607_),
    .ZN(_02608_)
  );
  INV_X1 _22797_ (
    .A(_02608_),
    .ZN(_02609_)
  );
  MUX2_X1 _22798_ (
    .A(\rf[23] [5]),
    .B(\rf[19] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02610_)
  );
  AND2_X1 _22799_ (
    .A1(_08545_),
    .A2(_02610_),
    .ZN(_02611_)
  );
  INV_X1 _22800_ (
    .A(_02611_),
    .ZN(_02612_)
  );
  AND2_X1 _22801_ (
    .A1(_08544_),
    .A2(_02612_),
    .ZN(_02613_)
  );
  AND2_X1 _22802_ (
    .A1(_02609_),
    .A2(_02613_),
    .ZN(_02614_)
  );
  INV_X1 _22803_ (
    .A(_02614_),
    .ZN(_02615_)
  );
  AND2_X1 _22804_ (
    .A1(_02602_),
    .A2(_02615_),
    .ZN(_02616_)
  );
  MUX2_X1 _22805_ (
    .A(_02589_),
    .B(_02616_),
    .S(ibuf_io_inst_0_bits_inst_rs2[3]),
    .Z(_02617_)
  );
  MUX2_X1 _22806_ (
    .A(_02570_),
    .B(_02617_),
    .S(_08572_),
    .Z(_02618_)
  );
  MUX2_X1 _22807_ (
    .A(_02618_),
    .B(_10505_),
    .S(_02233_),
    .Z(_02619_)
  );
  MUX2_X1 _22808_ (
    .A(ex_reg_rs_msb_1[3]),
    .B(_02619_),
    .S(_02202_),
    .Z(_00152_)
  );
  AND2_X1 _22809_ (
    .A1(_08337_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02620_)
  );
  INV_X1 _22810_ (
    .A(_02620_),
    .ZN(_02621_)
  );
  AND2_X1 _22811_ (
    .A1(_08475_),
    .A2(_08546_),
    .ZN(_02622_)
  );
  INV_X1 _22812_ (
    .A(_02622_),
    .ZN(_02623_)
  );
  AND2_X1 _22813_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_02623_),
    .ZN(_02624_)
  );
  AND2_X1 _22814_ (
    .A1(_02621_),
    .A2(_02624_),
    .ZN(_02625_)
  );
  INV_X1 _22815_ (
    .A(_02625_),
    .ZN(_02626_)
  );
  MUX2_X1 _22816_ (
    .A(\rf[15] [6]),
    .B(\rf[11] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02627_)
  );
  AND2_X1 _22817_ (
    .A1(_08544_),
    .A2(_02627_),
    .ZN(_02628_)
  );
  INV_X1 _22818_ (
    .A(_02628_),
    .ZN(_02629_)
  );
  AND2_X1 _22819_ (
    .A1(_08545_),
    .A2(_02629_),
    .ZN(_02630_)
  );
  AND2_X1 _22820_ (
    .A1(_02626_),
    .A2(_02630_),
    .ZN(_02631_)
  );
  INV_X1 _22821_ (
    .A(_02631_),
    .ZN(_02632_)
  );
  AND2_X1 _22822_ (
    .A1(_08358_),
    .A2(_08546_),
    .ZN(_02633_)
  );
  INV_X1 _22823_ (
    .A(_02633_),
    .ZN(_02634_)
  );
  AND2_X1 _22824_ (
    .A1(_08259_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02635_)
  );
  INV_X1 _22825_ (
    .A(_02635_),
    .ZN(_02636_)
  );
  AND2_X1 _22826_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_02636_),
    .ZN(_02637_)
  );
  AND2_X1 _22827_ (
    .A1(_02634_),
    .A2(_02637_),
    .ZN(_02638_)
  );
  INV_X1 _22828_ (
    .A(_02638_),
    .ZN(_02639_)
  );
  MUX2_X1 _22829_ (
    .A(\rf[13] [6]),
    .B(\rf[9] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02640_)
  );
  AND2_X1 _22830_ (
    .A1(_08544_),
    .A2(_02640_),
    .ZN(_02641_)
  );
  INV_X1 _22831_ (
    .A(_02641_),
    .ZN(_02642_)
  );
  AND2_X1 _22832_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02642_),
    .ZN(_02643_)
  );
  AND2_X1 _22833_ (
    .A1(_02639_),
    .A2(_02643_),
    .ZN(_02644_)
  );
  INV_X1 _22834_ (
    .A(_02644_),
    .ZN(_02645_)
  );
  AND2_X1 _22835_ (
    .A1(_08547_),
    .A2(_02645_),
    .ZN(_02646_)
  );
  AND2_X1 _22836_ (
    .A1(_02632_),
    .A2(_02646_),
    .ZN(_02647_)
  );
  INV_X1 _22837_ (
    .A(_02647_),
    .ZN(_02648_)
  );
  MUX2_X1 _22838_ (
    .A(\rf[6] [6]),
    .B(\rf[2] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02649_)
  );
  AND2_X1 _22839_ (
    .A1(_08545_),
    .A2(_02649_),
    .ZN(_02650_)
  );
  INV_X1 _22840_ (
    .A(_02650_),
    .ZN(_02651_)
  );
  MUX2_X1 _22841_ (
    .A(\rf[4] [6]),
    .B(\rf[0] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02652_)
  );
  AND2_X1 _22842_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02652_),
    .ZN(_02653_)
  );
  INV_X1 _22843_ (
    .A(_02653_),
    .ZN(_02654_)
  );
  AND2_X1 _22844_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_02654_),
    .ZN(_02655_)
  );
  AND2_X1 _22845_ (
    .A1(_02651_),
    .A2(_02655_),
    .ZN(_02656_)
  );
  INV_X1 _22846_ (
    .A(_02656_),
    .ZN(_02657_)
  );
  MUX2_X1 _22847_ (
    .A(\rf[7] [6]),
    .B(\rf[3] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02658_)
  );
  AND2_X1 _22848_ (
    .A1(_08545_),
    .A2(_02658_),
    .ZN(_02659_)
  );
  INV_X1 _22849_ (
    .A(_02659_),
    .ZN(_02660_)
  );
  MUX2_X1 _22850_ (
    .A(\rf[5] [6]),
    .B(\rf[1] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02661_)
  );
  AND2_X1 _22851_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02661_),
    .ZN(_02662_)
  );
  INV_X1 _22852_ (
    .A(_02662_),
    .ZN(_02663_)
  );
  AND2_X1 _22853_ (
    .A1(_08544_),
    .A2(_02663_),
    .ZN(_02664_)
  );
  AND2_X1 _22854_ (
    .A1(_02660_),
    .A2(_02664_),
    .ZN(_02665_)
  );
  INV_X1 _22855_ (
    .A(_02665_),
    .ZN(_02666_)
  );
  AND2_X1 _22856_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_02666_),
    .ZN(_02667_)
  );
  AND2_X1 _22857_ (
    .A1(_02657_),
    .A2(_02667_),
    .ZN(_02668_)
  );
  INV_X1 _22858_ (
    .A(_02668_),
    .ZN(_02669_)
  );
  AND2_X1 _22859_ (
    .A1(_02648_),
    .A2(_02669_),
    .ZN(_02670_)
  );
  AND2_X1 _22860_ (
    .A1(_08310_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02671_)
  );
  INV_X1 _22861_ (
    .A(_02671_),
    .ZN(_02672_)
  );
  AND2_X1 _22862_ (
    .A1(_08409_),
    .A2(_08546_),
    .ZN(_02673_)
  );
  INV_X1 _22863_ (
    .A(_02673_),
    .ZN(_02674_)
  );
  AND2_X1 _22864_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02674_),
    .ZN(_02675_)
  );
  AND2_X1 _22865_ (
    .A1(_02672_),
    .A2(_02675_),
    .ZN(_02676_)
  );
  INV_X1 _22866_ (
    .A(_02676_),
    .ZN(_02677_)
  );
  MUX2_X1 _22867_ (
    .A(\rf[23] [6]),
    .B(\rf[19] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02678_)
  );
  AND2_X1 _22868_ (
    .A1(_08545_),
    .A2(_02678_),
    .ZN(_02679_)
  );
  INV_X1 _22869_ (
    .A(_02679_),
    .ZN(_02680_)
  );
  AND2_X1 _22870_ (
    .A1(_08544_),
    .A2(_02680_),
    .ZN(_02681_)
  );
  AND2_X1 _22871_ (
    .A1(_02677_),
    .A2(_02681_),
    .ZN(_02682_)
  );
  INV_X1 _22872_ (
    .A(_02682_),
    .ZN(_02683_)
  );
  AND2_X1 _22873_ (
    .A1(_08379_),
    .A2(_08546_),
    .ZN(_02684_)
  );
  INV_X1 _22874_ (
    .A(_02684_),
    .ZN(_02685_)
  );
  AND2_X1 _22875_ (
    .A1(_08280_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02686_)
  );
  INV_X1 _22876_ (
    .A(_02686_),
    .ZN(_02687_)
  );
  AND2_X1 _22877_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02687_),
    .ZN(_02688_)
  );
  AND2_X1 _22878_ (
    .A1(_02685_),
    .A2(_02688_),
    .ZN(_02689_)
  );
  INV_X1 _22879_ (
    .A(_02689_),
    .ZN(_02690_)
  );
  MUX2_X1 _22880_ (
    .A(\rf[22] [6]),
    .B(\rf[18] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02691_)
  );
  AND2_X1 _22881_ (
    .A1(_08545_),
    .A2(_02691_),
    .ZN(_02692_)
  );
  INV_X1 _22882_ (
    .A(_02692_),
    .ZN(_02693_)
  );
  AND2_X1 _22883_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_02693_),
    .ZN(_02694_)
  );
  AND2_X1 _22884_ (
    .A1(_02690_),
    .A2(_02694_),
    .ZN(_02695_)
  );
  INV_X1 _22885_ (
    .A(_02695_),
    .ZN(_02696_)
  );
  AND2_X1 _22886_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_02683_),
    .ZN(_02697_)
  );
  AND2_X1 _22887_ (
    .A1(_02696_),
    .A2(_02697_),
    .ZN(_02698_)
  );
  INV_X1 _22888_ (
    .A(_02698_),
    .ZN(_02699_)
  );
  AND2_X1 _22889_ (
    .A1(_08438_),
    .A2(_08546_),
    .ZN(_02700_)
  );
  INV_X1 _22890_ (
    .A(_02700_),
    .ZN(_02701_)
  );
  AND2_X1 _22891_ (
    .A1(_08508_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02702_)
  );
  INV_X1 _22892_ (
    .A(_02702_),
    .ZN(_02703_)
  );
  AND2_X1 _22893_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02703_),
    .ZN(_02704_)
  );
  AND2_X1 _22894_ (
    .A1(_02701_),
    .A2(_02704_),
    .ZN(_02705_)
  );
  INV_X1 _22895_ (
    .A(_02705_),
    .ZN(_02706_)
  );
  MUX2_X1 _22896_ (
    .A(\rf[30] [6]),
    .B(\rf[26] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02707_)
  );
  AND2_X1 _22897_ (
    .A1(_08545_),
    .A2(_02707_),
    .ZN(_02708_)
  );
  INV_X1 _22898_ (
    .A(_02708_),
    .ZN(_02709_)
  );
  AND2_X1 _22899_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_02709_),
    .ZN(_02710_)
  );
  AND2_X1 _22900_ (
    .A1(_02706_),
    .A2(_02710_),
    .ZN(_02711_)
  );
  INV_X1 _22901_ (
    .A(_02711_),
    .ZN(_02712_)
  );
  MUX2_X1 _22902_ (
    .A(\rf[29] [6]),
    .B(\rf[25] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02713_)
  );
  AND2_X1 _22903_ (
    .A1(\rf[27] [6]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02714_)
  );
  MUX2_X1 _22904_ (
    .A(_02713_),
    .B(_02714_),
    .S(_08545_),
    .Z(_02715_)
  );
  INV_X1 _22905_ (
    .A(_02715_),
    .ZN(_02716_)
  );
  AND2_X1 _22906_ (
    .A1(_08544_),
    .A2(_02716_),
    .ZN(_02717_)
  );
  INV_X1 _22907_ (
    .A(_02717_),
    .ZN(_02718_)
  );
  AND2_X1 _22908_ (
    .A1(_08547_),
    .A2(_02718_),
    .ZN(_02719_)
  );
  AND2_X1 _22909_ (
    .A1(_02712_),
    .A2(_02719_),
    .ZN(_02720_)
  );
  INV_X1 _22910_ (
    .A(_02720_),
    .ZN(_02721_)
  );
  AND2_X1 _22911_ (
    .A1(_02699_),
    .A2(_02721_),
    .ZN(_02722_)
  );
  MUX2_X1 _22912_ (
    .A(_02670_),
    .B(_02722_),
    .S(_08572_),
    .Z(_02723_)
  );
  INV_X1 _22913_ (
    .A(_02723_),
    .ZN(_02724_)
  );
  MUX2_X1 _22914_ (
    .A(_02724_),
    .B(_10620_),
    .S(_02233_),
    .Z(_02725_)
  );
  MUX2_X1 _22915_ (
    .A(ex_reg_rs_msb_1[4]),
    .B(_02725_),
    .S(_02202_),
    .Z(_00153_)
  );
  MUX2_X1 _22916_ (
    .A(\rf[1] [7]),
    .B(\rf[0] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_02726_)
  );
  MUX2_X1 _22917_ (
    .A(\rf[5] [7]),
    .B(\rf[4] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_02727_)
  );
  MUX2_X1 _22918_ (
    .A(_02726_),
    .B(_02727_),
    .S(_08546_),
    .Z(_02728_)
  );
  INV_X1 _22919_ (
    .A(_02728_),
    .ZN(_02729_)
  );
  AND2_X1 _22920_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_02729_),
    .ZN(_02730_)
  );
  INV_X1 _22921_ (
    .A(_02730_),
    .ZN(_02731_)
  );
  MUX2_X1 _22922_ (
    .A(\rf[12] [7]),
    .B(\rf[8] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02732_)
  );
  INV_X1 _22923_ (
    .A(_02732_),
    .ZN(_02733_)
  );
  AND2_X1 _22924_ (
    .A1(_02341_),
    .A2(_02733_),
    .ZN(_02734_)
  );
  INV_X1 _22925_ (
    .A(_02734_),
    .ZN(_02735_)
  );
  MUX2_X1 _22926_ (
    .A(\rf[13] [7]),
    .B(\rf[9] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02736_)
  );
  INV_X1 _22927_ (
    .A(_02736_),
    .ZN(_02737_)
  );
  AND2_X1 _22928_ (
    .A1(_09692_),
    .A2(_02737_),
    .ZN(_02738_)
  );
  INV_X1 _22929_ (
    .A(_02738_),
    .ZN(_02739_)
  );
  AND2_X1 _22930_ (
    .A1(_02735_),
    .A2(_02739_),
    .ZN(_02740_)
  );
  AND2_X1 _22931_ (
    .A1(_02731_),
    .A2(_02740_),
    .ZN(_02741_)
  );
  MUX2_X1 _22932_ (
    .A(\rf[3] [7]),
    .B(\rf[2] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_02742_)
  );
  MUX2_X1 _22933_ (
    .A(\rf[7] [7]),
    .B(\rf[6] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_02743_)
  );
  MUX2_X1 _22934_ (
    .A(_02742_),
    .B(_02743_),
    .S(_08546_),
    .Z(_02744_)
  );
  INV_X1 _22935_ (
    .A(_02744_),
    .ZN(_02745_)
  );
  AND2_X1 _22936_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_02745_),
    .ZN(_02746_)
  );
  INV_X1 _22937_ (
    .A(_02746_),
    .ZN(_02747_)
  );
  MUX2_X1 _22938_ (
    .A(\rf[15] [7]),
    .B(\rf[11] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02748_)
  );
  INV_X1 _22939_ (
    .A(_02748_),
    .ZN(_02749_)
  );
  AND2_X1 _22940_ (
    .A1(_09692_),
    .A2(_02749_),
    .ZN(_02750_)
  );
  INV_X1 _22941_ (
    .A(_02750_),
    .ZN(_02751_)
  );
  MUX2_X1 _22942_ (
    .A(\rf[14] [7]),
    .B(\rf[10] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02752_)
  );
  INV_X1 _22943_ (
    .A(_02752_),
    .ZN(_02753_)
  );
  AND2_X1 _22944_ (
    .A1(_02341_),
    .A2(_02753_),
    .ZN(_02754_)
  );
  INV_X1 _22945_ (
    .A(_02754_),
    .ZN(_02755_)
  );
  AND2_X1 _22946_ (
    .A1(_02751_),
    .A2(_02755_),
    .ZN(_02756_)
  );
  AND2_X1 _22947_ (
    .A1(_02747_),
    .A2(_02756_),
    .ZN(_02757_)
  );
  MUX2_X1 _22948_ (
    .A(_02741_),
    .B(_02757_),
    .S(_08545_),
    .Z(_02758_)
  );
  AND2_X1 _22949_ (
    .A1(_08311_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02759_)
  );
  INV_X1 _22950_ (
    .A(_02759_),
    .ZN(_02760_)
  );
  AND2_X1 _22951_ (
    .A1(_08410_),
    .A2(_08546_),
    .ZN(_02761_)
  );
  INV_X1 _22952_ (
    .A(_02761_),
    .ZN(_02762_)
  );
  AND2_X1 _22953_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02762_),
    .ZN(_02763_)
  );
  AND2_X1 _22954_ (
    .A1(_02760_),
    .A2(_02763_),
    .ZN(_02764_)
  );
  INV_X1 _22955_ (
    .A(_02764_),
    .ZN(_02765_)
  );
  MUX2_X1 _22956_ (
    .A(\rf[23] [7]),
    .B(\rf[19] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02766_)
  );
  AND2_X1 _22957_ (
    .A1(_08545_),
    .A2(_02766_),
    .ZN(_02767_)
  );
  INV_X1 _22958_ (
    .A(_02767_),
    .ZN(_02768_)
  );
  AND2_X1 _22959_ (
    .A1(_08544_),
    .A2(_02768_),
    .ZN(_02769_)
  );
  AND2_X1 _22960_ (
    .A1(_02765_),
    .A2(_02769_),
    .ZN(_02770_)
  );
  INV_X1 _22961_ (
    .A(_02770_),
    .ZN(_02771_)
  );
  AND2_X1 _22962_ (
    .A1(_08380_),
    .A2(_08546_),
    .ZN(_02772_)
  );
  INV_X1 _22963_ (
    .A(_02772_),
    .ZN(_02773_)
  );
  AND2_X1 _22964_ (
    .A1(_08281_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02774_)
  );
  INV_X1 _22965_ (
    .A(_02774_),
    .ZN(_02775_)
  );
  AND2_X1 _22966_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02775_),
    .ZN(_02776_)
  );
  AND2_X1 _22967_ (
    .A1(_02773_),
    .A2(_02776_),
    .ZN(_02777_)
  );
  INV_X1 _22968_ (
    .A(_02777_),
    .ZN(_02778_)
  );
  MUX2_X1 _22969_ (
    .A(\rf[22] [7]),
    .B(\rf[18] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02779_)
  );
  AND2_X1 _22970_ (
    .A1(_08545_),
    .A2(_02779_),
    .ZN(_02780_)
  );
  INV_X1 _22971_ (
    .A(_02780_),
    .ZN(_02781_)
  );
  AND2_X1 _22972_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_02781_),
    .ZN(_02782_)
  );
  AND2_X1 _22973_ (
    .A1(_02778_),
    .A2(_02782_),
    .ZN(_02783_)
  );
  INV_X1 _22974_ (
    .A(_02783_),
    .ZN(_02784_)
  );
  AND2_X1 _22975_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_02771_),
    .ZN(_02785_)
  );
  AND2_X1 _22976_ (
    .A1(_02784_),
    .A2(_02785_),
    .ZN(_02786_)
  );
  INV_X1 _22977_ (
    .A(_02786_),
    .ZN(_02787_)
  );
  AND2_X1 _22978_ (
    .A1(_08439_),
    .A2(_08546_),
    .ZN(_02788_)
  );
  INV_X1 _22979_ (
    .A(_02788_),
    .ZN(_02789_)
  );
  AND2_X1 _22980_ (
    .A1(_08509_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02790_)
  );
  INV_X1 _22981_ (
    .A(_02790_),
    .ZN(_02791_)
  );
  AND2_X1 _22982_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02791_),
    .ZN(_02792_)
  );
  AND2_X1 _22983_ (
    .A1(_02789_),
    .A2(_02792_),
    .ZN(_02793_)
  );
  INV_X1 _22984_ (
    .A(_02793_),
    .ZN(_02794_)
  );
  MUX2_X1 _22985_ (
    .A(\rf[30] [7]),
    .B(\rf[26] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02795_)
  );
  AND2_X1 _22986_ (
    .A1(_08545_),
    .A2(_02795_),
    .ZN(_02796_)
  );
  INV_X1 _22987_ (
    .A(_02796_),
    .ZN(_02797_)
  );
  AND2_X1 _22988_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_02797_),
    .ZN(_02798_)
  );
  AND2_X1 _22989_ (
    .A1(_02794_),
    .A2(_02798_),
    .ZN(_02799_)
  );
  INV_X1 _22990_ (
    .A(_02799_),
    .ZN(_02800_)
  );
  MUX2_X1 _22991_ (
    .A(\rf[29] [7]),
    .B(\rf[25] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02801_)
  );
  AND2_X1 _22992_ (
    .A1(\rf[27] [7]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02802_)
  );
  MUX2_X1 _22993_ (
    .A(_02801_),
    .B(_02802_),
    .S(_08545_),
    .Z(_02803_)
  );
  INV_X1 _22994_ (
    .A(_02803_),
    .ZN(_02804_)
  );
  AND2_X1 _22995_ (
    .A1(_08544_),
    .A2(_02804_),
    .ZN(_02805_)
  );
  INV_X1 _22996_ (
    .A(_02805_),
    .ZN(_02806_)
  );
  AND2_X1 _22997_ (
    .A1(_08547_),
    .A2(_02806_),
    .ZN(_02807_)
  );
  AND2_X1 _22998_ (
    .A1(_02800_),
    .A2(_02807_),
    .ZN(_02808_)
  );
  INV_X1 _22999_ (
    .A(_02808_),
    .ZN(_02809_)
  );
  AND2_X1 _23000_ (
    .A1(_02787_),
    .A2(_02809_),
    .ZN(_02810_)
  );
  INV_X1 _23001_ (
    .A(_02810_),
    .ZN(_02811_)
  );
  MUX2_X1 _23002_ (
    .A(_02758_),
    .B(_02811_),
    .S(_08572_),
    .Z(_02812_)
  );
  MUX2_X1 _23003_ (
    .A(_02812_),
    .B(_10733_),
    .S(_02233_),
    .Z(_02813_)
  );
  MUX2_X1 _23004_ (
    .A(ex_reg_rs_msb_1[5]),
    .B(_02813_),
    .S(_02202_),
    .Z(_00154_)
  );
  AND2_X1 _23005_ (
    .A1(_08338_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02814_)
  );
  INV_X1 _23006_ (
    .A(_02814_),
    .ZN(_02815_)
  );
  AND2_X1 _23007_ (
    .A1(_08476_),
    .A2(_08546_),
    .ZN(_02816_)
  );
  INV_X1 _23008_ (
    .A(_02816_),
    .ZN(_02817_)
  );
  AND2_X1 _23009_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_02817_),
    .ZN(_02818_)
  );
  AND2_X1 _23010_ (
    .A1(_02815_),
    .A2(_02818_),
    .ZN(_02819_)
  );
  INV_X1 _23011_ (
    .A(_02819_),
    .ZN(_02820_)
  );
  MUX2_X1 _23012_ (
    .A(\rf[15] [8]),
    .B(\rf[11] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02821_)
  );
  AND2_X1 _23013_ (
    .A1(_08544_),
    .A2(_02821_),
    .ZN(_02822_)
  );
  INV_X1 _23014_ (
    .A(_02822_),
    .ZN(_02823_)
  );
  AND2_X1 _23015_ (
    .A1(_08545_),
    .A2(_02823_),
    .ZN(_02824_)
  );
  AND2_X1 _23016_ (
    .A1(_02820_),
    .A2(_02824_),
    .ZN(_02825_)
  );
  INV_X1 _23017_ (
    .A(_02825_),
    .ZN(_02826_)
  );
  AND2_X1 _23018_ (
    .A1(_08359_),
    .A2(_08546_),
    .ZN(_02827_)
  );
  INV_X1 _23019_ (
    .A(_02827_),
    .ZN(_02828_)
  );
  AND2_X1 _23020_ (
    .A1(_08260_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02829_)
  );
  INV_X1 _23021_ (
    .A(_02829_),
    .ZN(_02830_)
  );
  AND2_X1 _23022_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_02830_),
    .ZN(_02831_)
  );
  AND2_X1 _23023_ (
    .A1(_02828_),
    .A2(_02831_),
    .ZN(_02832_)
  );
  INV_X1 _23024_ (
    .A(_02832_),
    .ZN(_02833_)
  );
  MUX2_X1 _23025_ (
    .A(\rf[13] [8]),
    .B(\rf[9] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02834_)
  );
  AND2_X1 _23026_ (
    .A1(_08544_),
    .A2(_02834_),
    .ZN(_02835_)
  );
  INV_X1 _23027_ (
    .A(_02835_),
    .ZN(_02836_)
  );
  AND2_X1 _23028_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02836_),
    .ZN(_02837_)
  );
  AND2_X1 _23029_ (
    .A1(_02833_),
    .A2(_02837_),
    .ZN(_02838_)
  );
  INV_X1 _23030_ (
    .A(_02838_),
    .ZN(_02839_)
  );
  AND2_X1 _23031_ (
    .A1(_08547_),
    .A2(_02839_),
    .ZN(_02840_)
  );
  AND2_X1 _23032_ (
    .A1(_02826_),
    .A2(_02840_),
    .ZN(_02841_)
  );
  INV_X1 _23033_ (
    .A(_02841_),
    .ZN(_02842_)
  );
  MUX2_X1 _23034_ (
    .A(\rf[6] [8]),
    .B(\rf[2] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02843_)
  );
  AND2_X1 _23035_ (
    .A1(_08545_),
    .A2(_02843_),
    .ZN(_02844_)
  );
  INV_X1 _23036_ (
    .A(_02844_),
    .ZN(_02845_)
  );
  MUX2_X1 _23037_ (
    .A(\rf[4] [8]),
    .B(\rf[0] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02846_)
  );
  AND2_X1 _23038_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02846_),
    .ZN(_02847_)
  );
  INV_X1 _23039_ (
    .A(_02847_),
    .ZN(_02848_)
  );
  AND2_X1 _23040_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_02848_),
    .ZN(_02849_)
  );
  AND2_X1 _23041_ (
    .A1(_02845_),
    .A2(_02849_),
    .ZN(_02850_)
  );
  INV_X1 _23042_ (
    .A(_02850_),
    .ZN(_02851_)
  );
  MUX2_X1 _23043_ (
    .A(\rf[7] [8]),
    .B(\rf[3] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02852_)
  );
  AND2_X1 _23044_ (
    .A1(_08545_),
    .A2(_02852_),
    .ZN(_02853_)
  );
  INV_X1 _23045_ (
    .A(_02853_),
    .ZN(_02854_)
  );
  MUX2_X1 _23046_ (
    .A(\rf[5] [8]),
    .B(\rf[1] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02855_)
  );
  AND2_X1 _23047_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02855_),
    .ZN(_02856_)
  );
  INV_X1 _23048_ (
    .A(_02856_),
    .ZN(_02857_)
  );
  AND2_X1 _23049_ (
    .A1(_08544_),
    .A2(_02857_),
    .ZN(_02858_)
  );
  AND2_X1 _23050_ (
    .A1(_02854_),
    .A2(_02858_),
    .ZN(_02859_)
  );
  INV_X1 _23051_ (
    .A(_02859_),
    .ZN(_02860_)
  );
  AND2_X1 _23052_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_02860_),
    .ZN(_02861_)
  );
  AND2_X1 _23053_ (
    .A1(_02851_),
    .A2(_02861_),
    .ZN(_02862_)
  );
  INV_X1 _23054_ (
    .A(_02862_),
    .ZN(_02863_)
  );
  AND2_X1 _23055_ (
    .A1(_02842_),
    .A2(_02863_),
    .ZN(_02864_)
  );
  AND2_X1 _23056_ (
    .A1(_08312_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02865_)
  );
  INV_X1 _23057_ (
    .A(_02865_),
    .ZN(_02866_)
  );
  AND2_X1 _23058_ (
    .A1(_08411_),
    .A2(_08546_),
    .ZN(_02867_)
  );
  INV_X1 _23059_ (
    .A(_02867_),
    .ZN(_02868_)
  );
  AND2_X1 _23060_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02868_),
    .ZN(_02869_)
  );
  AND2_X1 _23061_ (
    .A1(_02866_),
    .A2(_02869_),
    .ZN(_02870_)
  );
  INV_X1 _23062_ (
    .A(_02870_),
    .ZN(_02871_)
  );
  MUX2_X1 _23063_ (
    .A(\rf[23] [8]),
    .B(\rf[19] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02872_)
  );
  AND2_X1 _23064_ (
    .A1(_08545_),
    .A2(_02872_),
    .ZN(_02873_)
  );
  INV_X1 _23065_ (
    .A(_02873_),
    .ZN(_02874_)
  );
  AND2_X1 _23066_ (
    .A1(_08544_),
    .A2(_02874_),
    .ZN(_02875_)
  );
  AND2_X1 _23067_ (
    .A1(_02871_),
    .A2(_02875_),
    .ZN(_02876_)
  );
  INV_X1 _23068_ (
    .A(_02876_),
    .ZN(_02877_)
  );
  AND2_X1 _23069_ (
    .A1(_08381_),
    .A2(_08546_),
    .ZN(_02878_)
  );
  INV_X1 _23070_ (
    .A(_02878_),
    .ZN(_02879_)
  );
  AND2_X1 _23071_ (
    .A1(_08282_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02880_)
  );
  INV_X1 _23072_ (
    .A(_02880_),
    .ZN(_02881_)
  );
  AND2_X1 _23073_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02881_),
    .ZN(_02882_)
  );
  AND2_X1 _23074_ (
    .A1(_02879_),
    .A2(_02882_),
    .ZN(_02883_)
  );
  INV_X1 _23075_ (
    .A(_02883_),
    .ZN(_02884_)
  );
  MUX2_X1 _23076_ (
    .A(\rf[22] [8]),
    .B(\rf[18] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02885_)
  );
  AND2_X1 _23077_ (
    .A1(_08545_),
    .A2(_02885_),
    .ZN(_02886_)
  );
  INV_X1 _23078_ (
    .A(_02886_),
    .ZN(_02887_)
  );
  AND2_X1 _23079_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_02887_),
    .ZN(_02888_)
  );
  AND2_X1 _23080_ (
    .A1(_02884_),
    .A2(_02888_),
    .ZN(_02889_)
  );
  INV_X1 _23081_ (
    .A(_02889_),
    .ZN(_02890_)
  );
  AND2_X1 _23082_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_02877_),
    .ZN(_02891_)
  );
  AND2_X1 _23083_ (
    .A1(_02890_),
    .A2(_02891_),
    .ZN(_02892_)
  );
  INV_X1 _23084_ (
    .A(_02892_),
    .ZN(_02893_)
  );
  AND2_X1 _23085_ (
    .A1(_08440_),
    .A2(_08546_),
    .ZN(_02894_)
  );
  INV_X1 _23086_ (
    .A(_02894_),
    .ZN(_02895_)
  );
  AND2_X1 _23087_ (
    .A1(_08510_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02896_)
  );
  INV_X1 _23088_ (
    .A(_02896_),
    .ZN(_02897_)
  );
  AND2_X1 _23089_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02897_),
    .ZN(_02898_)
  );
  AND2_X1 _23090_ (
    .A1(_02895_),
    .A2(_02898_),
    .ZN(_02899_)
  );
  INV_X1 _23091_ (
    .A(_02899_),
    .ZN(_02900_)
  );
  MUX2_X1 _23092_ (
    .A(\rf[30] [8]),
    .B(\rf[26] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02901_)
  );
  AND2_X1 _23093_ (
    .A1(_08545_),
    .A2(_02901_),
    .ZN(_02902_)
  );
  INV_X1 _23094_ (
    .A(_02902_),
    .ZN(_02903_)
  );
  AND2_X1 _23095_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_02903_),
    .ZN(_02904_)
  );
  AND2_X1 _23096_ (
    .A1(_02900_),
    .A2(_02904_),
    .ZN(_02905_)
  );
  INV_X1 _23097_ (
    .A(_02905_),
    .ZN(_02906_)
  );
  MUX2_X1 _23098_ (
    .A(\rf[29] [8]),
    .B(\rf[25] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02907_)
  );
  AND2_X1 _23099_ (
    .A1(\rf[27] [8]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02908_)
  );
  MUX2_X1 _23100_ (
    .A(_02907_),
    .B(_02908_),
    .S(_08545_),
    .Z(_02909_)
  );
  INV_X1 _23101_ (
    .A(_02909_),
    .ZN(_02910_)
  );
  AND2_X1 _23102_ (
    .A1(_08544_),
    .A2(_02910_),
    .ZN(_02911_)
  );
  INV_X1 _23103_ (
    .A(_02911_),
    .ZN(_02912_)
  );
  AND2_X1 _23104_ (
    .A1(_08547_),
    .A2(_02912_),
    .ZN(_02913_)
  );
  AND2_X1 _23105_ (
    .A1(_02906_),
    .A2(_02913_),
    .ZN(_02914_)
  );
  INV_X1 _23106_ (
    .A(_02914_),
    .ZN(_02915_)
  );
  AND2_X1 _23107_ (
    .A1(_02893_),
    .A2(_02915_),
    .ZN(_02916_)
  );
  MUX2_X1 _23108_ (
    .A(_02864_),
    .B(_02916_),
    .S(_08572_),
    .Z(_02917_)
  );
  INV_X1 _23109_ (
    .A(_02917_),
    .ZN(_02918_)
  );
  MUX2_X1 _23110_ (
    .A(_02918_),
    .B(_10846_),
    .S(_02233_),
    .Z(_02919_)
  );
  MUX2_X1 _23111_ (
    .A(ex_reg_rs_msb_1[6]),
    .B(_02919_),
    .S(_02202_),
    .Z(_00155_)
  );
  AND2_X1 _23112_ (
    .A1(_08339_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02920_)
  );
  INV_X1 _23113_ (
    .A(_02920_),
    .ZN(_02921_)
  );
  AND2_X1 _23114_ (
    .A1(_08477_),
    .A2(_08546_),
    .ZN(_02922_)
  );
  INV_X1 _23115_ (
    .A(_02922_),
    .ZN(_02923_)
  );
  AND2_X1 _23116_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_02923_),
    .ZN(_02924_)
  );
  AND2_X1 _23117_ (
    .A1(_02921_),
    .A2(_02924_),
    .ZN(_02925_)
  );
  INV_X1 _23118_ (
    .A(_02925_),
    .ZN(_02926_)
  );
  MUX2_X1 _23119_ (
    .A(\rf[15] [9]),
    .B(\rf[11] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02927_)
  );
  AND2_X1 _23120_ (
    .A1(_08544_),
    .A2(_02927_),
    .ZN(_02928_)
  );
  INV_X1 _23121_ (
    .A(_02928_),
    .ZN(_02929_)
  );
  AND2_X1 _23122_ (
    .A1(_08545_),
    .A2(_02929_),
    .ZN(_02930_)
  );
  AND2_X1 _23123_ (
    .A1(_02926_),
    .A2(_02930_),
    .ZN(_02931_)
  );
  INV_X1 _23124_ (
    .A(_02931_),
    .ZN(_02932_)
  );
  AND2_X1 _23125_ (
    .A1(_08360_),
    .A2(_08546_),
    .ZN(_02933_)
  );
  INV_X1 _23126_ (
    .A(_02933_),
    .ZN(_02934_)
  );
  AND2_X1 _23127_ (
    .A1(_08261_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02935_)
  );
  INV_X1 _23128_ (
    .A(_02935_),
    .ZN(_02936_)
  );
  AND2_X1 _23129_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_02936_),
    .ZN(_02937_)
  );
  AND2_X1 _23130_ (
    .A1(_02934_),
    .A2(_02937_),
    .ZN(_02938_)
  );
  INV_X1 _23131_ (
    .A(_02938_),
    .ZN(_02939_)
  );
  MUX2_X1 _23132_ (
    .A(\rf[13] [9]),
    .B(\rf[9] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02940_)
  );
  AND2_X1 _23133_ (
    .A1(_08544_),
    .A2(_02940_),
    .ZN(_02941_)
  );
  INV_X1 _23134_ (
    .A(_02941_),
    .ZN(_02942_)
  );
  AND2_X1 _23135_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02942_),
    .ZN(_02943_)
  );
  AND2_X1 _23136_ (
    .A1(_02939_),
    .A2(_02943_),
    .ZN(_02944_)
  );
  INV_X1 _23137_ (
    .A(_02944_),
    .ZN(_02945_)
  );
  AND2_X1 _23138_ (
    .A1(_08547_),
    .A2(_02945_),
    .ZN(_02946_)
  );
  AND2_X1 _23139_ (
    .A1(_02932_),
    .A2(_02946_),
    .ZN(_02947_)
  );
  INV_X1 _23140_ (
    .A(_02947_),
    .ZN(_02948_)
  );
  MUX2_X1 _23141_ (
    .A(\rf[6] [9]),
    .B(\rf[2] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02949_)
  );
  AND2_X1 _23142_ (
    .A1(_08545_),
    .A2(_02949_),
    .ZN(_02950_)
  );
  INV_X1 _23143_ (
    .A(_02950_),
    .ZN(_02951_)
  );
  MUX2_X1 _23144_ (
    .A(\rf[4] [9]),
    .B(\rf[0] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02952_)
  );
  AND2_X1 _23145_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02952_),
    .ZN(_02953_)
  );
  INV_X1 _23146_ (
    .A(_02953_),
    .ZN(_02954_)
  );
  AND2_X1 _23147_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_02954_),
    .ZN(_02955_)
  );
  AND2_X1 _23148_ (
    .A1(_02951_),
    .A2(_02955_),
    .ZN(_02956_)
  );
  INV_X1 _23149_ (
    .A(_02956_),
    .ZN(_02957_)
  );
  MUX2_X1 _23150_ (
    .A(\rf[7] [9]),
    .B(\rf[3] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02958_)
  );
  AND2_X1 _23151_ (
    .A1(_08545_),
    .A2(_02958_),
    .ZN(_02959_)
  );
  INV_X1 _23152_ (
    .A(_02959_),
    .ZN(_02960_)
  );
  MUX2_X1 _23153_ (
    .A(\rf[5] [9]),
    .B(\rf[1] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02961_)
  );
  AND2_X1 _23154_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02961_),
    .ZN(_02962_)
  );
  INV_X1 _23155_ (
    .A(_02962_),
    .ZN(_02963_)
  );
  AND2_X1 _23156_ (
    .A1(_08544_),
    .A2(_02963_),
    .ZN(_02964_)
  );
  AND2_X1 _23157_ (
    .A1(_02960_),
    .A2(_02964_),
    .ZN(_02965_)
  );
  INV_X1 _23158_ (
    .A(_02965_),
    .ZN(_02966_)
  );
  AND2_X1 _23159_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_02966_),
    .ZN(_02967_)
  );
  AND2_X1 _23160_ (
    .A1(_02957_),
    .A2(_02967_),
    .ZN(_02968_)
  );
  INV_X1 _23161_ (
    .A(_02968_),
    .ZN(_02969_)
  );
  AND2_X1 _23162_ (
    .A1(_02948_),
    .A2(_02969_),
    .ZN(_02970_)
  );
  AND2_X1 _23163_ (
    .A1(_08313_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02971_)
  );
  INV_X1 _23164_ (
    .A(_02971_),
    .ZN(_02972_)
  );
  AND2_X1 _23165_ (
    .A1(_08412_),
    .A2(_08546_),
    .ZN(_02973_)
  );
  INV_X1 _23166_ (
    .A(_02973_),
    .ZN(_02974_)
  );
  AND2_X1 _23167_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02974_),
    .ZN(_02975_)
  );
  AND2_X1 _23168_ (
    .A1(_02972_),
    .A2(_02975_),
    .ZN(_02976_)
  );
  INV_X1 _23169_ (
    .A(_02976_),
    .ZN(_02977_)
  );
  MUX2_X1 _23170_ (
    .A(\rf[23] [9]),
    .B(\rf[19] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02978_)
  );
  AND2_X1 _23171_ (
    .A1(_08545_),
    .A2(_02978_),
    .ZN(_02979_)
  );
  INV_X1 _23172_ (
    .A(_02979_),
    .ZN(_02980_)
  );
  AND2_X1 _23173_ (
    .A1(_08544_),
    .A2(_02980_),
    .ZN(_02981_)
  );
  AND2_X1 _23174_ (
    .A1(_02977_),
    .A2(_02981_),
    .ZN(_02982_)
  );
  INV_X1 _23175_ (
    .A(_02982_),
    .ZN(_02983_)
  );
  AND2_X1 _23176_ (
    .A1(_08382_),
    .A2(_08546_),
    .ZN(_02984_)
  );
  INV_X1 _23177_ (
    .A(_02984_),
    .ZN(_02985_)
  );
  AND2_X1 _23178_ (
    .A1(_08283_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02986_)
  );
  INV_X1 _23179_ (
    .A(_02986_),
    .ZN(_02987_)
  );
  AND2_X1 _23180_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02987_),
    .ZN(_02988_)
  );
  AND2_X1 _23181_ (
    .A1(_02985_),
    .A2(_02988_),
    .ZN(_02989_)
  );
  INV_X1 _23182_ (
    .A(_02989_),
    .ZN(_02990_)
  );
  MUX2_X1 _23183_ (
    .A(\rf[22] [9]),
    .B(\rf[18] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_02991_)
  );
  AND2_X1 _23184_ (
    .A1(_08545_),
    .A2(_02991_),
    .ZN(_02992_)
  );
  INV_X1 _23185_ (
    .A(_02992_),
    .ZN(_02993_)
  );
  AND2_X1 _23186_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_02993_),
    .ZN(_02994_)
  );
  AND2_X1 _23187_ (
    .A1(_02990_),
    .A2(_02994_),
    .ZN(_02995_)
  );
  INV_X1 _23188_ (
    .A(_02995_),
    .ZN(_02996_)
  );
  AND2_X1 _23189_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_02983_),
    .ZN(_02997_)
  );
  AND2_X1 _23190_ (
    .A1(_02996_),
    .A2(_02997_),
    .ZN(_02998_)
  );
  INV_X1 _23191_ (
    .A(_02998_),
    .ZN(_02999_)
  );
  AND2_X1 _23192_ (
    .A1(_08441_),
    .A2(_08546_),
    .ZN(_03000_)
  );
  INV_X1 _23193_ (
    .A(_03000_),
    .ZN(_03001_)
  );
  AND2_X1 _23194_ (
    .A1(_08511_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03002_)
  );
  INV_X1 _23195_ (
    .A(_03002_),
    .ZN(_03003_)
  );
  AND2_X1 _23196_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03003_),
    .ZN(_03004_)
  );
  AND2_X1 _23197_ (
    .A1(_03001_),
    .A2(_03004_),
    .ZN(_03005_)
  );
  INV_X1 _23198_ (
    .A(_03005_),
    .ZN(_03006_)
  );
  MUX2_X1 _23199_ (
    .A(\rf[30] [9]),
    .B(\rf[26] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03007_)
  );
  AND2_X1 _23200_ (
    .A1(_08545_),
    .A2(_03007_),
    .ZN(_03008_)
  );
  INV_X1 _23201_ (
    .A(_03008_),
    .ZN(_03009_)
  );
  AND2_X1 _23202_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03009_),
    .ZN(_03010_)
  );
  AND2_X1 _23203_ (
    .A1(_03006_),
    .A2(_03010_),
    .ZN(_03011_)
  );
  INV_X1 _23204_ (
    .A(_03011_),
    .ZN(_03012_)
  );
  MUX2_X1 _23205_ (
    .A(\rf[29] [9]),
    .B(\rf[25] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03013_)
  );
  AND2_X1 _23206_ (
    .A1(\rf[27] [9]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03014_)
  );
  MUX2_X1 _23207_ (
    .A(_03013_),
    .B(_03014_),
    .S(_08545_),
    .Z(_03015_)
  );
  INV_X1 _23208_ (
    .A(_03015_),
    .ZN(_03016_)
  );
  AND2_X1 _23209_ (
    .A1(_08544_),
    .A2(_03016_),
    .ZN(_03017_)
  );
  INV_X1 _23210_ (
    .A(_03017_),
    .ZN(_03018_)
  );
  AND2_X1 _23211_ (
    .A1(_08547_),
    .A2(_03018_),
    .ZN(_03019_)
  );
  AND2_X1 _23212_ (
    .A1(_03012_),
    .A2(_03019_),
    .ZN(_03020_)
  );
  INV_X1 _23213_ (
    .A(_03020_),
    .ZN(_03021_)
  );
  AND2_X1 _23214_ (
    .A1(_02999_),
    .A2(_03021_),
    .ZN(_03022_)
  );
  MUX2_X1 _23215_ (
    .A(_02970_),
    .B(_03022_),
    .S(_08572_),
    .Z(_03023_)
  );
  INV_X1 _23216_ (
    .A(_03023_),
    .ZN(_03024_)
  );
  MUX2_X1 _23217_ (
    .A(_03024_),
    .B(_10956_),
    .S(_02233_),
    .Z(_03025_)
  );
  MUX2_X1 _23218_ (
    .A(ex_reg_rs_msb_1[7]),
    .B(_03025_),
    .S(_02202_),
    .Z(_00156_)
  );
  MUX2_X1 _23219_ (
    .A(\rf[3] [10]),
    .B(\rf[2] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_03026_)
  );
  MUX2_X1 _23220_ (
    .A(\rf[7] [10]),
    .B(\rf[6] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_03027_)
  );
  MUX2_X1 _23221_ (
    .A(_03026_),
    .B(_03027_),
    .S(_08546_),
    .Z(_03028_)
  );
  INV_X1 _23222_ (
    .A(_03028_),
    .ZN(_03029_)
  );
  AND2_X1 _23223_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_03029_),
    .ZN(_03030_)
  );
  INV_X1 _23224_ (
    .A(_03030_),
    .ZN(_03031_)
  );
  MUX2_X1 _23225_ (
    .A(\rf[15] [10]),
    .B(\rf[11] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03032_)
  );
  INV_X1 _23226_ (
    .A(_03032_),
    .ZN(_03033_)
  );
  AND2_X1 _23227_ (
    .A1(_09692_),
    .A2(_03033_),
    .ZN(_03034_)
  );
  INV_X1 _23228_ (
    .A(_03034_),
    .ZN(_03035_)
  );
  MUX2_X1 _23229_ (
    .A(\rf[14] [10]),
    .B(\rf[10] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03036_)
  );
  INV_X1 _23230_ (
    .A(_03036_),
    .ZN(_03037_)
  );
  AND2_X1 _23231_ (
    .A1(_02341_),
    .A2(_03037_),
    .ZN(_03038_)
  );
  INV_X1 _23232_ (
    .A(_03038_),
    .ZN(_03039_)
  );
  AND2_X1 _23233_ (
    .A1(_03035_),
    .A2(_03039_),
    .ZN(_03040_)
  );
  AND2_X1 _23234_ (
    .A1(_03031_),
    .A2(_03040_),
    .ZN(_03041_)
  );
  MUX2_X1 _23235_ (
    .A(\rf[1] [10]),
    .B(\rf[0] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_03042_)
  );
  MUX2_X1 _23236_ (
    .A(\rf[5] [10]),
    .B(\rf[4] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_03043_)
  );
  MUX2_X1 _23237_ (
    .A(_03042_),
    .B(_03043_),
    .S(_08546_),
    .Z(_03044_)
  );
  INV_X1 _23238_ (
    .A(_03044_),
    .ZN(_03045_)
  );
  AND2_X1 _23239_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_03045_),
    .ZN(_03046_)
  );
  INV_X1 _23240_ (
    .A(_03046_),
    .ZN(_03047_)
  );
  MUX2_X1 _23241_ (
    .A(\rf[12] [10]),
    .B(\rf[8] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03048_)
  );
  INV_X1 _23242_ (
    .A(_03048_),
    .ZN(_03049_)
  );
  AND2_X1 _23243_ (
    .A1(_02341_),
    .A2(_03049_),
    .ZN(_03050_)
  );
  INV_X1 _23244_ (
    .A(_03050_),
    .ZN(_03051_)
  );
  MUX2_X1 _23245_ (
    .A(\rf[13] [10]),
    .B(\rf[9] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03052_)
  );
  INV_X1 _23246_ (
    .A(_03052_),
    .ZN(_03053_)
  );
  AND2_X1 _23247_ (
    .A1(_09692_),
    .A2(_03053_),
    .ZN(_03054_)
  );
  INV_X1 _23248_ (
    .A(_03054_),
    .ZN(_03055_)
  );
  AND2_X1 _23249_ (
    .A1(_03051_),
    .A2(_03055_),
    .ZN(_03056_)
  );
  AND2_X1 _23250_ (
    .A1(_03047_),
    .A2(_03056_),
    .ZN(_03057_)
  );
  AND2_X1 _23251_ (
    .A1(\rf[30] [10]),
    .A2(_08546_),
    .ZN(_03058_)
  );
  INV_X1 _23252_ (
    .A(_03058_),
    .ZN(_03059_)
  );
  AND2_X1 _23253_ (
    .A1(\rf[26] [10]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03060_)
  );
  INV_X1 _23254_ (
    .A(_03060_),
    .ZN(_03061_)
  );
  AND2_X1 _23255_ (
    .A1(_08545_),
    .A2(_03061_),
    .ZN(_03062_)
  );
  AND2_X1 _23256_ (
    .A1(_03059_),
    .A2(_03062_),
    .ZN(_03063_)
  );
  INV_X1 _23257_ (
    .A(_03063_),
    .ZN(_03064_)
  );
  AND2_X1 _23258_ (
    .A1(\rf[24] [10]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03065_)
  );
  INV_X1 _23259_ (
    .A(_03065_),
    .ZN(_03066_)
  );
  AND2_X1 _23260_ (
    .A1(\rf[28] [10]),
    .A2(_08546_),
    .ZN(_03067_)
  );
  INV_X1 _23261_ (
    .A(_03067_),
    .ZN(_03068_)
  );
  AND2_X1 _23262_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03068_),
    .ZN(_03069_)
  );
  AND2_X1 _23263_ (
    .A1(_03066_),
    .A2(_03069_),
    .ZN(_03070_)
  );
  INV_X1 _23264_ (
    .A(_03070_),
    .ZN(_03071_)
  );
  AND2_X1 _23265_ (
    .A1(_03064_),
    .A2(_03071_),
    .ZN(_03072_)
  );
  MUX2_X1 _23266_ (
    .A(\rf[29] [10]),
    .B(\rf[25] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03073_)
  );
  AND2_X1 _23267_ (
    .A1(\rf[27] [10]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03074_)
  );
  MUX2_X1 _23268_ (
    .A(_03073_),
    .B(_03074_),
    .S(_08545_),
    .Z(_03075_)
  );
  MUX2_X1 _23269_ (
    .A(_03072_),
    .B(_03075_),
    .S(_08544_),
    .Z(_03076_)
  );
  AND2_X1 _23270_ (
    .A1(_08383_),
    .A2(_08546_),
    .ZN(_03077_)
  );
  INV_X1 _23271_ (
    .A(_03077_),
    .ZN(_03078_)
  );
  AND2_X1 _23272_ (
    .A1(_08284_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03079_)
  );
  INV_X1 _23273_ (
    .A(_03079_),
    .ZN(_03080_)
  );
  AND2_X1 _23274_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03080_),
    .ZN(_03081_)
  );
  AND2_X1 _23275_ (
    .A1(_03078_),
    .A2(_03081_),
    .ZN(_03082_)
  );
  INV_X1 _23276_ (
    .A(_03082_),
    .ZN(_03083_)
  );
  MUX2_X1 _23277_ (
    .A(\rf[22] [10]),
    .B(\rf[18] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03084_)
  );
  AND2_X1 _23278_ (
    .A1(_08545_),
    .A2(_03084_),
    .ZN(_03085_)
  );
  INV_X1 _23279_ (
    .A(_03085_),
    .ZN(_03086_)
  );
  AND2_X1 _23280_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03086_),
    .ZN(_03087_)
  );
  AND2_X1 _23281_ (
    .A1(_03083_),
    .A2(_03087_),
    .ZN(_03088_)
  );
  INV_X1 _23282_ (
    .A(_03088_),
    .ZN(_03089_)
  );
  AND2_X1 _23283_ (
    .A1(_08314_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03090_)
  );
  INV_X1 _23284_ (
    .A(_03090_),
    .ZN(_03091_)
  );
  AND2_X1 _23285_ (
    .A1(_08413_),
    .A2(_08546_),
    .ZN(_03092_)
  );
  INV_X1 _23286_ (
    .A(_03092_),
    .ZN(_03093_)
  );
  AND2_X1 _23287_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03093_),
    .ZN(_03094_)
  );
  AND2_X1 _23288_ (
    .A1(_03091_),
    .A2(_03094_),
    .ZN(_03095_)
  );
  INV_X1 _23289_ (
    .A(_03095_),
    .ZN(_03096_)
  );
  MUX2_X1 _23290_ (
    .A(\rf[23] [10]),
    .B(\rf[19] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03097_)
  );
  AND2_X1 _23291_ (
    .A1(_08545_),
    .A2(_03097_),
    .ZN(_03098_)
  );
  INV_X1 _23292_ (
    .A(_03098_),
    .ZN(_03099_)
  );
  AND2_X1 _23293_ (
    .A1(_08544_),
    .A2(_03099_),
    .ZN(_03100_)
  );
  AND2_X1 _23294_ (
    .A1(_03096_),
    .A2(_03100_),
    .ZN(_03101_)
  );
  INV_X1 _23295_ (
    .A(_03101_),
    .ZN(_03102_)
  );
  AND2_X1 _23296_ (
    .A1(_03089_),
    .A2(_03102_),
    .ZN(_03103_)
  );
  MUX2_X1 _23297_ (
    .A(_03076_),
    .B(_03103_),
    .S(ibuf_io_inst_0_bits_inst_rs2[3]),
    .Z(_03104_)
  );
  MUX2_X1 _23298_ (
    .A(_03041_),
    .B(_03057_),
    .S(ibuf_io_inst_0_bits_inst_rs2[1]),
    .Z(_03105_)
  );
  MUX2_X1 _23299_ (
    .A(_03104_),
    .B(_03105_),
    .S(ibuf_io_inst_0_bits_inst_rs2[4]),
    .Z(_03106_)
  );
  MUX2_X1 _23300_ (
    .A(_03106_),
    .B(_11066_),
    .S(_02233_),
    .Z(_03107_)
  );
  MUX2_X1 _23301_ (
    .A(ex_reg_rs_msb_1[8]),
    .B(_03107_),
    .S(_02202_),
    .Z(_00157_)
  );
  AND2_X1 _23302_ (
    .A1(_08340_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03108_)
  );
  INV_X1 _23303_ (
    .A(_03108_),
    .ZN(_03109_)
  );
  AND2_X1 _23304_ (
    .A1(_08478_),
    .A2(_08546_),
    .ZN(_03110_)
  );
  INV_X1 _23305_ (
    .A(_03110_),
    .ZN(_03111_)
  );
  AND2_X1 _23306_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03111_),
    .ZN(_03112_)
  );
  AND2_X1 _23307_ (
    .A1(_03109_),
    .A2(_03112_),
    .ZN(_03113_)
  );
  INV_X1 _23308_ (
    .A(_03113_),
    .ZN(_03114_)
  );
  MUX2_X1 _23309_ (
    .A(\rf[15] [11]),
    .B(\rf[11] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03115_)
  );
  AND2_X1 _23310_ (
    .A1(_08544_),
    .A2(_03115_),
    .ZN(_03116_)
  );
  INV_X1 _23311_ (
    .A(_03116_),
    .ZN(_03117_)
  );
  AND2_X1 _23312_ (
    .A1(_08545_),
    .A2(_03117_),
    .ZN(_03118_)
  );
  AND2_X1 _23313_ (
    .A1(_03114_),
    .A2(_03118_),
    .ZN(_03119_)
  );
  INV_X1 _23314_ (
    .A(_03119_),
    .ZN(_03120_)
  );
  AND2_X1 _23315_ (
    .A1(_08361_),
    .A2(_08546_),
    .ZN(_03121_)
  );
  INV_X1 _23316_ (
    .A(_03121_),
    .ZN(_03122_)
  );
  AND2_X1 _23317_ (
    .A1(_08262_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03123_)
  );
  INV_X1 _23318_ (
    .A(_03123_),
    .ZN(_03124_)
  );
  AND2_X1 _23319_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03124_),
    .ZN(_03125_)
  );
  AND2_X1 _23320_ (
    .A1(_03122_),
    .A2(_03125_),
    .ZN(_03126_)
  );
  INV_X1 _23321_ (
    .A(_03126_),
    .ZN(_03127_)
  );
  MUX2_X1 _23322_ (
    .A(\rf[13] [11]),
    .B(\rf[9] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03128_)
  );
  AND2_X1 _23323_ (
    .A1(_08544_),
    .A2(_03128_),
    .ZN(_03129_)
  );
  INV_X1 _23324_ (
    .A(_03129_),
    .ZN(_03130_)
  );
  AND2_X1 _23325_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03130_),
    .ZN(_03131_)
  );
  AND2_X1 _23326_ (
    .A1(_03127_),
    .A2(_03131_),
    .ZN(_03132_)
  );
  INV_X1 _23327_ (
    .A(_03132_),
    .ZN(_03133_)
  );
  AND2_X1 _23328_ (
    .A1(_08547_),
    .A2(_03133_),
    .ZN(_03134_)
  );
  AND2_X1 _23329_ (
    .A1(_03120_),
    .A2(_03134_),
    .ZN(_03135_)
  );
  INV_X1 _23330_ (
    .A(_03135_),
    .ZN(_03136_)
  );
  MUX2_X1 _23331_ (
    .A(\rf[6] [11]),
    .B(\rf[2] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03137_)
  );
  AND2_X1 _23332_ (
    .A1(_08545_),
    .A2(_03137_),
    .ZN(_03138_)
  );
  INV_X1 _23333_ (
    .A(_03138_),
    .ZN(_03139_)
  );
  MUX2_X1 _23334_ (
    .A(\rf[4] [11]),
    .B(\rf[0] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03140_)
  );
  AND2_X1 _23335_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03140_),
    .ZN(_03141_)
  );
  INV_X1 _23336_ (
    .A(_03141_),
    .ZN(_03142_)
  );
  AND2_X1 _23337_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03142_),
    .ZN(_03143_)
  );
  AND2_X1 _23338_ (
    .A1(_03139_),
    .A2(_03143_),
    .ZN(_03144_)
  );
  INV_X1 _23339_ (
    .A(_03144_),
    .ZN(_03145_)
  );
  MUX2_X1 _23340_ (
    .A(\rf[7] [11]),
    .B(\rf[3] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03146_)
  );
  AND2_X1 _23341_ (
    .A1(_08545_),
    .A2(_03146_),
    .ZN(_03147_)
  );
  INV_X1 _23342_ (
    .A(_03147_),
    .ZN(_03148_)
  );
  MUX2_X1 _23343_ (
    .A(\rf[5] [11]),
    .B(\rf[1] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03149_)
  );
  AND2_X1 _23344_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03149_),
    .ZN(_03150_)
  );
  INV_X1 _23345_ (
    .A(_03150_),
    .ZN(_03151_)
  );
  AND2_X1 _23346_ (
    .A1(_08544_),
    .A2(_03151_),
    .ZN(_03152_)
  );
  AND2_X1 _23347_ (
    .A1(_03148_),
    .A2(_03152_),
    .ZN(_03153_)
  );
  INV_X1 _23348_ (
    .A(_03153_),
    .ZN(_03154_)
  );
  AND2_X1 _23349_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_03154_),
    .ZN(_03155_)
  );
  AND2_X1 _23350_ (
    .A1(_03145_),
    .A2(_03155_),
    .ZN(_03156_)
  );
  INV_X1 _23351_ (
    .A(_03156_),
    .ZN(_03157_)
  );
  AND2_X1 _23352_ (
    .A1(_03136_),
    .A2(_03157_),
    .ZN(_03158_)
  );
  AND2_X1 _23353_ (
    .A1(_08315_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03159_)
  );
  INV_X1 _23354_ (
    .A(_03159_),
    .ZN(_03160_)
  );
  AND2_X1 _23355_ (
    .A1(_08414_),
    .A2(_08546_),
    .ZN(_03161_)
  );
  INV_X1 _23356_ (
    .A(_03161_),
    .ZN(_03162_)
  );
  AND2_X1 _23357_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03162_),
    .ZN(_03163_)
  );
  AND2_X1 _23358_ (
    .A1(_03160_),
    .A2(_03163_),
    .ZN(_03164_)
  );
  INV_X1 _23359_ (
    .A(_03164_),
    .ZN(_03165_)
  );
  MUX2_X1 _23360_ (
    .A(\rf[23] [11]),
    .B(\rf[19] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03166_)
  );
  AND2_X1 _23361_ (
    .A1(_08545_),
    .A2(_03166_),
    .ZN(_03167_)
  );
  INV_X1 _23362_ (
    .A(_03167_),
    .ZN(_03168_)
  );
  AND2_X1 _23363_ (
    .A1(_08544_),
    .A2(_03168_),
    .ZN(_03169_)
  );
  AND2_X1 _23364_ (
    .A1(_03165_),
    .A2(_03169_),
    .ZN(_03170_)
  );
  INV_X1 _23365_ (
    .A(_03170_),
    .ZN(_03171_)
  );
  AND2_X1 _23366_ (
    .A1(_08384_),
    .A2(_08546_),
    .ZN(_03172_)
  );
  INV_X1 _23367_ (
    .A(_03172_),
    .ZN(_03173_)
  );
  AND2_X1 _23368_ (
    .A1(_08285_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03174_)
  );
  INV_X1 _23369_ (
    .A(_03174_),
    .ZN(_03175_)
  );
  AND2_X1 _23370_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03175_),
    .ZN(_03176_)
  );
  AND2_X1 _23371_ (
    .A1(_03173_),
    .A2(_03176_),
    .ZN(_03177_)
  );
  INV_X1 _23372_ (
    .A(_03177_),
    .ZN(_03178_)
  );
  MUX2_X1 _23373_ (
    .A(\rf[22] [11]),
    .B(\rf[18] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03179_)
  );
  AND2_X1 _23374_ (
    .A1(_08545_),
    .A2(_03179_),
    .ZN(_03180_)
  );
  INV_X1 _23375_ (
    .A(_03180_),
    .ZN(_03181_)
  );
  AND2_X1 _23376_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03181_),
    .ZN(_03182_)
  );
  AND2_X1 _23377_ (
    .A1(_03178_),
    .A2(_03182_),
    .ZN(_03183_)
  );
  INV_X1 _23378_ (
    .A(_03183_),
    .ZN(_03184_)
  );
  AND2_X1 _23379_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_03171_),
    .ZN(_03185_)
  );
  AND2_X1 _23380_ (
    .A1(_03184_),
    .A2(_03185_),
    .ZN(_03186_)
  );
  INV_X1 _23381_ (
    .A(_03186_),
    .ZN(_03187_)
  );
  AND2_X1 _23382_ (
    .A1(_08442_),
    .A2(_08546_),
    .ZN(_03188_)
  );
  INV_X1 _23383_ (
    .A(_03188_),
    .ZN(_03189_)
  );
  AND2_X1 _23384_ (
    .A1(_08512_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03190_)
  );
  INV_X1 _23385_ (
    .A(_03190_),
    .ZN(_03191_)
  );
  AND2_X1 _23386_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03191_),
    .ZN(_03192_)
  );
  AND2_X1 _23387_ (
    .A1(_03189_),
    .A2(_03192_),
    .ZN(_03193_)
  );
  INV_X1 _23388_ (
    .A(_03193_),
    .ZN(_03194_)
  );
  MUX2_X1 _23389_ (
    .A(\rf[30] [11]),
    .B(\rf[26] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03195_)
  );
  AND2_X1 _23390_ (
    .A1(_08545_),
    .A2(_03195_),
    .ZN(_03196_)
  );
  INV_X1 _23391_ (
    .A(_03196_),
    .ZN(_03197_)
  );
  AND2_X1 _23392_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03197_),
    .ZN(_03198_)
  );
  AND2_X1 _23393_ (
    .A1(_03194_),
    .A2(_03198_),
    .ZN(_03199_)
  );
  INV_X1 _23394_ (
    .A(_03199_),
    .ZN(_03200_)
  );
  MUX2_X1 _23395_ (
    .A(\rf[29] [11]),
    .B(\rf[25] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03201_)
  );
  AND2_X1 _23396_ (
    .A1(\rf[27] [11]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03202_)
  );
  MUX2_X1 _23397_ (
    .A(_03201_),
    .B(_03202_),
    .S(_08545_),
    .Z(_03203_)
  );
  INV_X1 _23398_ (
    .A(_03203_),
    .ZN(_03204_)
  );
  AND2_X1 _23399_ (
    .A1(_08544_),
    .A2(_03204_),
    .ZN(_03205_)
  );
  INV_X1 _23400_ (
    .A(_03205_),
    .ZN(_03206_)
  );
  AND2_X1 _23401_ (
    .A1(_08547_),
    .A2(_03206_),
    .ZN(_03207_)
  );
  AND2_X1 _23402_ (
    .A1(_03200_),
    .A2(_03207_),
    .ZN(_03208_)
  );
  INV_X1 _23403_ (
    .A(_03208_),
    .ZN(_03209_)
  );
  AND2_X1 _23404_ (
    .A1(_03187_),
    .A2(_03209_),
    .ZN(_03210_)
  );
  MUX2_X1 _23405_ (
    .A(_03158_),
    .B(_03210_),
    .S(_08572_),
    .Z(_03211_)
  );
  INV_X1 _23406_ (
    .A(_03211_),
    .ZN(_03212_)
  );
  MUX2_X1 _23407_ (
    .A(_03212_),
    .B(_11205_),
    .S(_02233_),
    .Z(_03213_)
  );
  MUX2_X1 _23408_ (
    .A(ex_reg_rs_msb_1[9]),
    .B(_03213_),
    .S(_02202_),
    .Z(_00158_)
  );
  MUX2_X1 _23409_ (
    .A(\rf[7] [12]),
    .B(\rf[3] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03214_)
  );
  AND2_X1 _23410_ (
    .A1(_08545_),
    .A2(_03214_),
    .ZN(_03215_)
  );
  INV_X1 _23411_ (
    .A(_03215_),
    .ZN(_03216_)
  );
  MUX2_X1 _23412_ (
    .A(\rf[5] [12]),
    .B(\rf[1] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03217_)
  );
  AND2_X1 _23413_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03217_),
    .ZN(_03218_)
  );
  INV_X1 _23414_ (
    .A(_03218_),
    .ZN(_03219_)
  );
  AND2_X1 _23415_ (
    .A1(_08544_),
    .A2(_03219_),
    .ZN(_03220_)
  );
  AND2_X1 _23416_ (
    .A1(_03216_),
    .A2(_03220_),
    .ZN(_03221_)
  );
  INV_X1 _23417_ (
    .A(_03221_),
    .ZN(_03222_)
  );
  MUX2_X1 _23418_ (
    .A(\rf[6] [12]),
    .B(\rf[2] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03223_)
  );
  AND2_X1 _23419_ (
    .A1(_08545_),
    .A2(_03223_),
    .ZN(_03224_)
  );
  INV_X1 _23420_ (
    .A(_03224_),
    .ZN(_03225_)
  );
  MUX2_X1 _23421_ (
    .A(\rf[4] [12]),
    .B(\rf[0] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03226_)
  );
  AND2_X1 _23422_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03226_),
    .ZN(_03227_)
  );
  INV_X1 _23423_ (
    .A(_03227_),
    .ZN(_03228_)
  );
  AND2_X1 _23424_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03228_),
    .ZN(_03229_)
  );
  AND2_X1 _23425_ (
    .A1(_03225_),
    .A2(_03229_),
    .ZN(_03230_)
  );
  INV_X1 _23426_ (
    .A(_03230_),
    .ZN(_03231_)
  );
  AND2_X1 _23427_ (
    .A1(_03222_),
    .A2(_03231_),
    .ZN(_03232_)
  );
  AND2_X1 _23428_ (
    .A1(\rf[14] [12]),
    .A2(_08545_),
    .ZN(_03233_)
  );
  INV_X1 _23429_ (
    .A(_03233_),
    .ZN(_03234_)
  );
  AND2_X1 _23430_ (
    .A1(\rf[12] [12]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_03235_)
  );
  INV_X1 _23431_ (
    .A(_03235_),
    .ZN(_03236_)
  );
  AND2_X1 _23432_ (
    .A1(_08546_),
    .A2(_03236_),
    .ZN(_03237_)
  );
  AND2_X1 _23433_ (
    .A1(_03234_),
    .A2(_03237_),
    .ZN(_03238_)
  );
  INV_X1 _23434_ (
    .A(_03238_),
    .ZN(_03239_)
  );
  AND2_X1 _23435_ (
    .A1(\rf[10] [12]),
    .A2(_08545_),
    .ZN(_03240_)
  );
  INV_X1 _23436_ (
    .A(_03240_),
    .ZN(_03241_)
  );
  AND2_X1 _23437_ (
    .A1(\rf[8] [12]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_03242_)
  );
  INV_X1 _23438_ (
    .A(_03242_),
    .ZN(_03243_)
  );
  AND2_X1 _23439_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[2]),
    .A2(_03243_),
    .ZN(_03244_)
  );
  AND2_X1 _23440_ (
    .A1(_03241_),
    .A2(_03244_),
    .ZN(_03245_)
  );
  INV_X1 _23441_ (
    .A(_03245_),
    .ZN(_03246_)
  );
  AND2_X1 _23442_ (
    .A1(_03239_),
    .A2(_03246_),
    .ZN(_03247_)
  );
  AND2_X1 _23443_ (
    .A1(\rf[15] [12]),
    .A2(_08545_),
    .ZN(_03248_)
  );
  INV_X1 _23444_ (
    .A(_03248_),
    .ZN(_03249_)
  );
  AND2_X1 _23445_ (
    .A1(\rf[13] [12]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_03250_)
  );
  INV_X1 _23446_ (
    .A(_03250_),
    .ZN(_03251_)
  );
  AND2_X1 _23447_ (
    .A1(_08546_),
    .A2(_03251_),
    .ZN(_03252_)
  );
  AND2_X1 _23448_ (
    .A1(_03249_),
    .A2(_03252_),
    .ZN(_03253_)
  );
  INV_X1 _23449_ (
    .A(_03253_),
    .ZN(_03254_)
  );
  AND2_X1 _23450_ (
    .A1(\rf[11] [12]),
    .A2(_08545_),
    .ZN(_03255_)
  );
  INV_X1 _23451_ (
    .A(_03255_),
    .ZN(_03256_)
  );
  AND2_X1 _23452_ (
    .A1(\rf[9] [12]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_03257_)
  );
  INV_X1 _23453_ (
    .A(_03257_),
    .ZN(_03258_)
  );
  AND2_X1 _23454_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[2]),
    .A2(_03258_),
    .ZN(_03259_)
  );
  AND2_X1 _23455_ (
    .A1(_03256_),
    .A2(_03259_),
    .ZN(_03260_)
  );
  INV_X1 _23456_ (
    .A(_03260_),
    .ZN(_03261_)
  );
  AND2_X1 _23457_ (
    .A1(_03254_),
    .A2(_03261_),
    .ZN(_03262_)
  );
  MUX2_X1 _23458_ (
    .A(_03247_),
    .B(_03262_),
    .S(_08544_),
    .Z(_03263_)
  );
  MUX2_X1 _23459_ (
    .A(_03232_),
    .B(_03263_),
    .S(_08547_),
    .Z(_03264_)
  );
  AND2_X1 _23460_ (
    .A1(\rf[30] [12]),
    .A2(_08546_),
    .ZN(_03265_)
  );
  INV_X1 _23461_ (
    .A(_03265_),
    .ZN(_03266_)
  );
  AND2_X1 _23462_ (
    .A1(\rf[26] [12]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03267_)
  );
  INV_X1 _23463_ (
    .A(_03267_),
    .ZN(_03268_)
  );
  AND2_X1 _23464_ (
    .A1(_08545_),
    .A2(_03268_),
    .ZN(_03269_)
  );
  AND2_X1 _23465_ (
    .A1(_03266_),
    .A2(_03269_),
    .ZN(_03270_)
  );
  INV_X1 _23466_ (
    .A(_03270_),
    .ZN(_03271_)
  );
  AND2_X1 _23467_ (
    .A1(\rf[24] [12]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03272_)
  );
  INV_X1 _23468_ (
    .A(_03272_),
    .ZN(_03273_)
  );
  AND2_X1 _23469_ (
    .A1(\rf[28] [12]),
    .A2(_08546_),
    .ZN(_03274_)
  );
  INV_X1 _23470_ (
    .A(_03274_),
    .ZN(_03275_)
  );
  AND2_X1 _23471_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03275_),
    .ZN(_03276_)
  );
  AND2_X1 _23472_ (
    .A1(_03273_),
    .A2(_03276_),
    .ZN(_03277_)
  );
  INV_X1 _23473_ (
    .A(_03277_),
    .ZN(_03278_)
  );
  AND2_X1 _23474_ (
    .A1(_03271_),
    .A2(_03278_),
    .ZN(_03279_)
  );
  MUX2_X1 _23475_ (
    .A(\rf[29] [12]),
    .B(\rf[25] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03280_)
  );
  AND2_X1 _23476_ (
    .A1(\rf[27] [12]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03281_)
  );
  MUX2_X1 _23477_ (
    .A(_03280_),
    .B(_03281_),
    .S(_08545_),
    .Z(_03282_)
  );
  MUX2_X1 _23478_ (
    .A(_03279_),
    .B(_03282_),
    .S(_08544_),
    .Z(_03283_)
  );
  AND2_X1 _23479_ (
    .A1(_08385_),
    .A2(_08546_),
    .ZN(_03284_)
  );
  INV_X1 _23480_ (
    .A(_03284_),
    .ZN(_03285_)
  );
  AND2_X1 _23481_ (
    .A1(_08286_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03286_)
  );
  INV_X1 _23482_ (
    .A(_03286_),
    .ZN(_03287_)
  );
  AND2_X1 _23483_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03287_),
    .ZN(_03288_)
  );
  AND2_X1 _23484_ (
    .A1(_03285_),
    .A2(_03288_),
    .ZN(_03289_)
  );
  INV_X1 _23485_ (
    .A(_03289_),
    .ZN(_03290_)
  );
  MUX2_X1 _23486_ (
    .A(\rf[22] [12]),
    .B(\rf[18] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03291_)
  );
  AND2_X1 _23487_ (
    .A1(_08545_),
    .A2(_03291_),
    .ZN(_03292_)
  );
  INV_X1 _23488_ (
    .A(_03292_),
    .ZN(_03293_)
  );
  AND2_X1 _23489_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03293_),
    .ZN(_03294_)
  );
  AND2_X1 _23490_ (
    .A1(_03290_),
    .A2(_03294_),
    .ZN(_03295_)
  );
  INV_X1 _23491_ (
    .A(_03295_),
    .ZN(_03296_)
  );
  AND2_X1 _23492_ (
    .A1(_08316_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03297_)
  );
  INV_X1 _23493_ (
    .A(_03297_),
    .ZN(_03298_)
  );
  AND2_X1 _23494_ (
    .A1(_08415_),
    .A2(_08546_),
    .ZN(_03299_)
  );
  INV_X1 _23495_ (
    .A(_03299_),
    .ZN(_03300_)
  );
  AND2_X1 _23496_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03300_),
    .ZN(_03301_)
  );
  AND2_X1 _23497_ (
    .A1(_03298_),
    .A2(_03301_),
    .ZN(_03302_)
  );
  INV_X1 _23498_ (
    .A(_03302_),
    .ZN(_03303_)
  );
  MUX2_X1 _23499_ (
    .A(\rf[23] [12]),
    .B(\rf[19] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03304_)
  );
  AND2_X1 _23500_ (
    .A1(_08545_),
    .A2(_03304_),
    .ZN(_03305_)
  );
  INV_X1 _23501_ (
    .A(_03305_),
    .ZN(_03306_)
  );
  AND2_X1 _23502_ (
    .A1(_08544_),
    .A2(_03306_),
    .ZN(_03307_)
  );
  AND2_X1 _23503_ (
    .A1(_03303_),
    .A2(_03307_),
    .ZN(_03308_)
  );
  INV_X1 _23504_ (
    .A(_03308_),
    .ZN(_03309_)
  );
  AND2_X1 _23505_ (
    .A1(_03296_),
    .A2(_03309_),
    .ZN(_03310_)
  );
  MUX2_X1 _23506_ (
    .A(_03283_),
    .B(_03310_),
    .S(ibuf_io_inst_0_bits_inst_rs2[3]),
    .Z(_03311_)
  );
  MUX2_X1 _23507_ (
    .A(_03264_),
    .B(_03311_),
    .S(_08572_),
    .Z(_03312_)
  );
  MUX2_X1 _23508_ (
    .A(_03312_),
    .B(_11315_),
    .S(_02233_),
    .Z(_03313_)
  );
  MUX2_X1 _23509_ (
    .A(ex_reg_rs_msb_1[10]),
    .B(_03313_),
    .S(_02202_),
    .Z(_00159_)
  );
  MUX2_X1 _23510_ (
    .A(\rf[7] [13]),
    .B(\rf[3] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03314_)
  );
  AND2_X1 _23511_ (
    .A1(_08545_),
    .A2(_03314_),
    .ZN(_03315_)
  );
  INV_X1 _23512_ (
    .A(_03315_),
    .ZN(_03316_)
  );
  MUX2_X1 _23513_ (
    .A(\rf[5] [13]),
    .B(\rf[1] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03317_)
  );
  AND2_X1 _23514_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03317_),
    .ZN(_03318_)
  );
  INV_X1 _23515_ (
    .A(_03318_),
    .ZN(_03319_)
  );
  AND2_X1 _23516_ (
    .A1(_08544_),
    .A2(_03319_),
    .ZN(_03320_)
  );
  AND2_X1 _23517_ (
    .A1(_03316_),
    .A2(_03320_),
    .ZN(_03321_)
  );
  INV_X1 _23518_ (
    .A(_03321_),
    .ZN(_03322_)
  );
  MUX2_X1 _23519_ (
    .A(\rf[6] [13]),
    .B(\rf[2] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03323_)
  );
  AND2_X1 _23520_ (
    .A1(_08545_),
    .A2(_03323_),
    .ZN(_03324_)
  );
  INV_X1 _23521_ (
    .A(_03324_),
    .ZN(_03325_)
  );
  MUX2_X1 _23522_ (
    .A(\rf[4] [13]),
    .B(\rf[0] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03326_)
  );
  AND2_X1 _23523_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03326_),
    .ZN(_03327_)
  );
  INV_X1 _23524_ (
    .A(_03327_),
    .ZN(_03328_)
  );
  AND2_X1 _23525_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03328_),
    .ZN(_03329_)
  );
  AND2_X1 _23526_ (
    .A1(_03325_),
    .A2(_03329_),
    .ZN(_03330_)
  );
  INV_X1 _23527_ (
    .A(_03330_),
    .ZN(_03331_)
  );
  AND2_X1 _23528_ (
    .A1(_03322_),
    .A2(_03331_),
    .ZN(_03332_)
  );
  AND2_X1 _23529_ (
    .A1(\rf[14] [13]),
    .A2(_08545_),
    .ZN(_03333_)
  );
  INV_X1 _23530_ (
    .A(_03333_),
    .ZN(_03334_)
  );
  AND2_X1 _23531_ (
    .A1(\rf[12] [13]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_03335_)
  );
  INV_X1 _23532_ (
    .A(_03335_),
    .ZN(_03336_)
  );
  AND2_X1 _23533_ (
    .A1(_08546_),
    .A2(_03336_),
    .ZN(_03337_)
  );
  AND2_X1 _23534_ (
    .A1(_03334_),
    .A2(_03337_),
    .ZN(_03338_)
  );
  INV_X1 _23535_ (
    .A(_03338_),
    .ZN(_03339_)
  );
  AND2_X1 _23536_ (
    .A1(\rf[10] [13]),
    .A2(_08545_),
    .ZN(_03340_)
  );
  INV_X1 _23537_ (
    .A(_03340_),
    .ZN(_03341_)
  );
  AND2_X1 _23538_ (
    .A1(\rf[8] [13]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_03342_)
  );
  INV_X1 _23539_ (
    .A(_03342_),
    .ZN(_03343_)
  );
  AND2_X1 _23540_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[2]),
    .A2(_03343_),
    .ZN(_03344_)
  );
  AND2_X1 _23541_ (
    .A1(_03341_),
    .A2(_03344_),
    .ZN(_03345_)
  );
  INV_X1 _23542_ (
    .A(_03345_),
    .ZN(_03346_)
  );
  AND2_X1 _23543_ (
    .A1(_03339_),
    .A2(_03346_),
    .ZN(_03347_)
  );
  AND2_X1 _23544_ (
    .A1(\rf[15] [13]),
    .A2(_08545_),
    .ZN(_03348_)
  );
  INV_X1 _23545_ (
    .A(_03348_),
    .ZN(_03349_)
  );
  AND2_X1 _23546_ (
    .A1(\rf[13] [13]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_03350_)
  );
  INV_X1 _23547_ (
    .A(_03350_),
    .ZN(_03351_)
  );
  AND2_X1 _23548_ (
    .A1(_08546_),
    .A2(_03351_),
    .ZN(_03352_)
  );
  AND2_X1 _23549_ (
    .A1(_03349_),
    .A2(_03352_),
    .ZN(_03353_)
  );
  INV_X1 _23550_ (
    .A(_03353_),
    .ZN(_03354_)
  );
  AND2_X1 _23551_ (
    .A1(\rf[11] [13]),
    .A2(_08545_),
    .ZN(_03355_)
  );
  INV_X1 _23552_ (
    .A(_03355_),
    .ZN(_03356_)
  );
  AND2_X1 _23553_ (
    .A1(\rf[9] [13]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_03357_)
  );
  INV_X1 _23554_ (
    .A(_03357_),
    .ZN(_03358_)
  );
  AND2_X1 _23555_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[2]),
    .A2(_03358_),
    .ZN(_03359_)
  );
  AND2_X1 _23556_ (
    .A1(_03356_),
    .A2(_03359_),
    .ZN(_03360_)
  );
  INV_X1 _23557_ (
    .A(_03360_),
    .ZN(_03361_)
  );
  AND2_X1 _23558_ (
    .A1(_03354_),
    .A2(_03361_),
    .ZN(_03362_)
  );
  MUX2_X1 _23559_ (
    .A(_03347_),
    .B(_03362_),
    .S(_08544_),
    .Z(_03363_)
  );
  MUX2_X1 _23560_ (
    .A(_03332_),
    .B(_03363_),
    .S(_08547_),
    .Z(_03364_)
  );
  AND2_X1 _23561_ (
    .A1(\rf[30] [13]),
    .A2(_08546_),
    .ZN(_03365_)
  );
  INV_X1 _23562_ (
    .A(_03365_),
    .ZN(_03366_)
  );
  AND2_X1 _23563_ (
    .A1(\rf[26] [13]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03367_)
  );
  INV_X1 _23564_ (
    .A(_03367_),
    .ZN(_03368_)
  );
  AND2_X1 _23565_ (
    .A1(_08545_),
    .A2(_03368_),
    .ZN(_03369_)
  );
  AND2_X1 _23566_ (
    .A1(_03366_),
    .A2(_03369_),
    .ZN(_03370_)
  );
  INV_X1 _23567_ (
    .A(_03370_),
    .ZN(_03371_)
  );
  AND2_X1 _23568_ (
    .A1(\rf[24] [13]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03372_)
  );
  INV_X1 _23569_ (
    .A(_03372_),
    .ZN(_03373_)
  );
  AND2_X1 _23570_ (
    .A1(\rf[28] [13]),
    .A2(_08546_),
    .ZN(_03374_)
  );
  INV_X1 _23571_ (
    .A(_03374_),
    .ZN(_03375_)
  );
  AND2_X1 _23572_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03375_),
    .ZN(_03376_)
  );
  AND2_X1 _23573_ (
    .A1(_03373_),
    .A2(_03376_),
    .ZN(_03377_)
  );
  INV_X1 _23574_ (
    .A(_03377_),
    .ZN(_03378_)
  );
  AND2_X1 _23575_ (
    .A1(_03371_),
    .A2(_03378_),
    .ZN(_03379_)
  );
  MUX2_X1 _23576_ (
    .A(\rf[29] [13]),
    .B(\rf[25] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03380_)
  );
  AND2_X1 _23577_ (
    .A1(\rf[27] [13]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03381_)
  );
  MUX2_X1 _23578_ (
    .A(_03380_),
    .B(_03381_),
    .S(_08545_),
    .Z(_03382_)
  );
  MUX2_X1 _23579_ (
    .A(_03379_),
    .B(_03382_),
    .S(_08544_),
    .Z(_03383_)
  );
  AND2_X1 _23580_ (
    .A1(_08386_),
    .A2(_08546_),
    .ZN(_03384_)
  );
  INV_X1 _23581_ (
    .A(_03384_),
    .ZN(_03385_)
  );
  AND2_X1 _23582_ (
    .A1(_08287_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03386_)
  );
  INV_X1 _23583_ (
    .A(_03386_),
    .ZN(_03387_)
  );
  AND2_X1 _23584_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03387_),
    .ZN(_03388_)
  );
  AND2_X1 _23585_ (
    .A1(_03385_),
    .A2(_03388_),
    .ZN(_03389_)
  );
  INV_X1 _23586_ (
    .A(_03389_),
    .ZN(_03390_)
  );
  MUX2_X1 _23587_ (
    .A(\rf[22] [13]),
    .B(\rf[18] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03391_)
  );
  AND2_X1 _23588_ (
    .A1(_08545_),
    .A2(_03391_),
    .ZN(_03392_)
  );
  INV_X1 _23589_ (
    .A(_03392_),
    .ZN(_03393_)
  );
  AND2_X1 _23590_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03393_),
    .ZN(_03394_)
  );
  AND2_X1 _23591_ (
    .A1(_03390_),
    .A2(_03394_),
    .ZN(_03395_)
  );
  INV_X1 _23592_ (
    .A(_03395_),
    .ZN(_03396_)
  );
  AND2_X1 _23593_ (
    .A1(_08317_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03397_)
  );
  INV_X1 _23594_ (
    .A(_03397_),
    .ZN(_03398_)
  );
  AND2_X1 _23595_ (
    .A1(_08416_),
    .A2(_08546_),
    .ZN(_03399_)
  );
  INV_X1 _23596_ (
    .A(_03399_),
    .ZN(_03400_)
  );
  AND2_X1 _23597_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03400_),
    .ZN(_03401_)
  );
  AND2_X1 _23598_ (
    .A1(_03398_),
    .A2(_03401_),
    .ZN(_03402_)
  );
  INV_X1 _23599_ (
    .A(_03402_),
    .ZN(_03403_)
  );
  MUX2_X1 _23600_ (
    .A(\rf[23] [13]),
    .B(\rf[19] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03404_)
  );
  AND2_X1 _23601_ (
    .A1(_08545_),
    .A2(_03404_),
    .ZN(_03405_)
  );
  INV_X1 _23602_ (
    .A(_03405_),
    .ZN(_03406_)
  );
  AND2_X1 _23603_ (
    .A1(_08544_),
    .A2(_03406_),
    .ZN(_03407_)
  );
  AND2_X1 _23604_ (
    .A1(_03403_),
    .A2(_03407_),
    .ZN(_03408_)
  );
  INV_X1 _23605_ (
    .A(_03408_),
    .ZN(_03409_)
  );
  AND2_X1 _23606_ (
    .A1(_03396_),
    .A2(_03409_),
    .ZN(_03410_)
  );
  MUX2_X1 _23607_ (
    .A(_03383_),
    .B(_03410_),
    .S(ibuf_io_inst_0_bits_inst_rs2[3]),
    .Z(_03411_)
  );
  MUX2_X1 _23608_ (
    .A(_03364_),
    .B(_03411_),
    .S(_08572_),
    .Z(_03412_)
  );
  MUX2_X1 _23609_ (
    .A(_03412_),
    .B(_11428_),
    .S(_02233_),
    .Z(_03413_)
  );
  MUX2_X1 _23610_ (
    .A(ex_reg_rs_msb_1[11]),
    .B(_03413_),
    .S(_02202_),
    .Z(_00160_)
  );
  AND2_X1 _23611_ (
    .A1(_08341_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03414_)
  );
  INV_X1 _23612_ (
    .A(_03414_),
    .ZN(_03415_)
  );
  AND2_X1 _23613_ (
    .A1(_08479_),
    .A2(_08546_),
    .ZN(_03416_)
  );
  INV_X1 _23614_ (
    .A(_03416_),
    .ZN(_03417_)
  );
  AND2_X1 _23615_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03417_),
    .ZN(_03418_)
  );
  AND2_X1 _23616_ (
    .A1(_03415_),
    .A2(_03418_),
    .ZN(_03419_)
  );
  INV_X1 _23617_ (
    .A(_03419_),
    .ZN(_03420_)
  );
  MUX2_X1 _23618_ (
    .A(\rf[15] [14]),
    .B(\rf[11] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03421_)
  );
  AND2_X1 _23619_ (
    .A1(_08544_),
    .A2(_03421_),
    .ZN(_03422_)
  );
  INV_X1 _23620_ (
    .A(_03422_),
    .ZN(_03423_)
  );
  AND2_X1 _23621_ (
    .A1(_08545_),
    .A2(_03423_),
    .ZN(_03424_)
  );
  AND2_X1 _23622_ (
    .A1(_03420_),
    .A2(_03424_),
    .ZN(_03425_)
  );
  INV_X1 _23623_ (
    .A(_03425_),
    .ZN(_03426_)
  );
  AND2_X1 _23624_ (
    .A1(_08362_),
    .A2(_08546_),
    .ZN(_03427_)
  );
  INV_X1 _23625_ (
    .A(_03427_),
    .ZN(_03428_)
  );
  AND2_X1 _23626_ (
    .A1(_08263_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03429_)
  );
  INV_X1 _23627_ (
    .A(_03429_),
    .ZN(_03430_)
  );
  AND2_X1 _23628_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03430_),
    .ZN(_03431_)
  );
  AND2_X1 _23629_ (
    .A1(_03428_),
    .A2(_03431_),
    .ZN(_03432_)
  );
  INV_X1 _23630_ (
    .A(_03432_),
    .ZN(_03433_)
  );
  MUX2_X1 _23631_ (
    .A(\rf[13] [14]),
    .B(\rf[9] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03434_)
  );
  AND2_X1 _23632_ (
    .A1(_08544_),
    .A2(_03434_),
    .ZN(_03435_)
  );
  INV_X1 _23633_ (
    .A(_03435_),
    .ZN(_03436_)
  );
  AND2_X1 _23634_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03436_),
    .ZN(_03437_)
  );
  AND2_X1 _23635_ (
    .A1(_03433_),
    .A2(_03437_),
    .ZN(_03438_)
  );
  INV_X1 _23636_ (
    .A(_03438_),
    .ZN(_03439_)
  );
  AND2_X1 _23637_ (
    .A1(_08547_),
    .A2(_03439_),
    .ZN(_03440_)
  );
  AND2_X1 _23638_ (
    .A1(_03426_),
    .A2(_03440_),
    .ZN(_03441_)
  );
  INV_X1 _23639_ (
    .A(_03441_),
    .ZN(_03442_)
  );
  MUX2_X1 _23640_ (
    .A(\rf[6] [14]),
    .B(\rf[2] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03443_)
  );
  AND2_X1 _23641_ (
    .A1(_08545_),
    .A2(_03443_),
    .ZN(_03444_)
  );
  INV_X1 _23642_ (
    .A(_03444_),
    .ZN(_03445_)
  );
  MUX2_X1 _23643_ (
    .A(\rf[4] [14]),
    .B(\rf[0] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03446_)
  );
  AND2_X1 _23644_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03446_),
    .ZN(_03447_)
  );
  INV_X1 _23645_ (
    .A(_03447_),
    .ZN(_03448_)
  );
  AND2_X1 _23646_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03448_),
    .ZN(_03449_)
  );
  AND2_X1 _23647_ (
    .A1(_03445_),
    .A2(_03449_),
    .ZN(_03450_)
  );
  INV_X1 _23648_ (
    .A(_03450_),
    .ZN(_03451_)
  );
  MUX2_X1 _23649_ (
    .A(\rf[7] [14]),
    .B(\rf[3] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03452_)
  );
  AND2_X1 _23650_ (
    .A1(_08545_),
    .A2(_03452_),
    .ZN(_03453_)
  );
  INV_X1 _23651_ (
    .A(_03453_),
    .ZN(_03454_)
  );
  MUX2_X1 _23652_ (
    .A(\rf[5] [14]),
    .B(\rf[1] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03455_)
  );
  AND2_X1 _23653_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03455_),
    .ZN(_03456_)
  );
  INV_X1 _23654_ (
    .A(_03456_),
    .ZN(_03457_)
  );
  AND2_X1 _23655_ (
    .A1(_08544_),
    .A2(_03457_),
    .ZN(_03458_)
  );
  AND2_X1 _23656_ (
    .A1(_03454_),
    .A2(_03458_),
    .ZN(_03459_)
  );
  INV_X1 _23657_ (
    .A(_03459_),
    .ZN(_03460_)
  );
  AND2_X1 _23658_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_03460_),
    .ZN(_03461_)
  );
  AND2_X1 _23659_ (
    .A1(_03451_),
    .A2(_03461_),
    .ZN(_03462_)
  );
  INV_X1 _23660_ (
    .A(_03462_),
    .ZN(_03463_)
  );
  AND2_X1 _23661_ (
    .A1(_03442_),
    .A2(_03463_),
    .ZN(_03464_)
  );
  AND2_X1 _23662_ (
    .A1(_08318_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03465_)
  );
  INV_X1 _23663_ (
    .A(_03465_),
    .ZN(_03466_)
  );
  AND2_X1 _23664_ (
    .A1(_08417_),
    .A2(_08546_),
    .ZN(_03467_)
  );
  INV_X1 _23665_ (
    .A(_03467_),
    .ZN(_03468_)
  );
  AND2_X1 _23666_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03468_),
    .ZN(_03469_)
  );
  AND2_X1 _23667_ (
    .A1(_03466_),
    .A2(_03469_),
    .ZN(_03470_)
  );
  INV_X1 _23668_ (
    .A(_03470_),
    .ZN(_03471_)
  );
  MUX2_X1 _23669_ (
    .A(\rf[23] [14]),
    .B(\rf[19] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03472_)
  );
  AND2_X1 _23670_ (
    .A1(_08545_),
    .A2(_03472_),
    .ZN(_03473_)
  );
  INV_X1 _23671_ (
    .A(_03473_),
    .ZN(_03474_)
  );
  AND2_X1 _23672_ (
    .A1(_08544_),
    .A2(_03474_),
    .ZN(_03475_)
  );
  AND2_X1 _23673_ (
    .A1(_03471_),
    .A2(_03475_),
    .ZN(_03476_)
  );
  INV_X1 _23674_ (
    .A(_03476_),
    .ZN(_03477_)
  );
  AND2_X1 _23675_ (
    .A1(_08387_),
    .A2(_08546_),
    .ZN(_03478_)
  );
  INV_X1 _23676_ (
    .A(_03478_),
    .ZN(_03479_)
  );
  AND2_X1 _23677_ (
    .A1(_08288_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03480_)
  );
  INV_X1 _23678_ (
    .A(_03480_),
    .ZN(_03481_)
  );
  AND2_X1 _23679_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03481_),
    .ZN(_03482_)
  );
  AND2_X1 _23680_ (
    .A1(_03479_),
    .A2(_03482_),
    .ZN(_03483_)
  );
  INV_X1 _23681_ (
    .A(_03483_),
    .ZN(_03484_)
  );
  MUX2_X1 _23682_ (
    .A(\rf[22] [14]),
    .B(\rf[18] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03485_)
  );
  AND2_X1 _23683_ (
    .A1(_08545_),
    .A2(_03485_),
    .ZN(_03486_)
  );
  INV_X1 _23684_ (
    .A(_03486_),
    .ZN(_03487_)
  );
  AND2_X1 _23685_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03487_),
    .ZN(_03488_)
  );
  AND2_X1 _23686_ (
    .A1(_03484_),
    .A2(_03488_),
    .ZN(_03489_)
  );
  INV_X1 _23687_ (
    .A(_03489_),
    .ZN(_03490_)
  );
  AND2_X1 _23688_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_03477_),
    .ZN(_03491_)
  );
  AND2_X1 _23689_ (
    .A1(_03490_),
    .A2(_03491_),
    .ZN(_03492_)
  );
  INV_X1 _23690_ (
    .A(_03492_),
    .ZN(_03493_)
  );
  AND2_X1 _23691_ (
    .A1(_08445_),
    .A2(_08546_),
    .ZN(_03494_)
  );
  INV_X1 _23692_ (
    .A(_03494_),
    .ZN(_03495_)
  );
  AND2_X1 _23693_ (
    .A1(_08515_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03496_)
  );
  INV_X1 _23694_ (
    .A(_03496_),
    .ZN(_03497_)
  );
  AND2_X1 _23695_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03497_),
    .ZN(_03498_)
  );
  AND2_X1 _23696_ (
    .A1(_03495_),
    .A2(_03498_),
    .ZN(_03499_)
  );
  INV_X1 _23697_ (
    .A(_03499_),
    .ZN(_03500_)
  );
  MUX2_X1 _23698_ (
    .A(\rf[30] [14]),
    .B(\rf[26] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03501_)
  );
  AND2_X1 _23699_ (
    .A1(_08545_),
    .A2(_03501_),
    .ZN(_03502_)
  );
  INV_X1 _23700_ (
    .A(_03502_),
    .ZN(_03503_)
  );
  AND2_X1 _23701_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03503_),
    .ZN(_03504_)
  );
  AND2_X1 _23702_ (
    .A1(_03500_),
    .A2(_03504_),
    .ZN(_03505_)
  );
  INV_X1 _23703_ (
    .A(_03505_),
    .ZN(_03506_)
  );
  MUX2_X1 _23704_ (
    .A(\rf[29] [14]),
    .B(\rf[25] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03507_)
  );
  AND2_X1 _23705_ (
    .A1(\rf[27] [14]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03508_)
  );
  MUX2_X1 _23706_ (
    .A(_03507_),
    .B(_03508_),
    .S(_08545_),
    .Z(_03509_)
  );
  INV_X1 _23707_ (
    .A(_03509_),
    .ZN(_03510_)
  );
  AND2_X1 _23708_ (
    .A1(_08544_),
    .A2(_03510_),
    .ZN(_03511_)
  );
  INV_X1 _23709_ (
    .A(_03511_),
    .ZN(_03512_)
  );
  AND2_X1 _23710_ (
    .A1(_08547_),
    .A2(_03512_),
    .ZN(_03513_)
  );
  AND2_X1 _23711_ (
    .A1(_03506_),
    .A2(_03513_),
    .ZN(_03514_)
  );
  INV_X1 _23712_ (
    .A(_03514_),
    .ZN(_03515_)
  );
  AND2_X1 _23713_ (
    .A1(_03493_),
    .A2(_03515_),
    .ZN(_03516_)
  );
  MUX2_X1 _23714_ (
    .A(_03464_),
    .B(_03516_),
    .S(_08572_),
    .Z(_03517_)
  );
  INV_X1 _23715_ (
    .A(_03517_),
    .ZN(_03518_)
  );
  MUX2_X1 _23716_ (
    .A(_03518_),
    .B(_11541_),
    .S(_02233_),
    .Z(_03519_)
  );
  MUX2_X1 _23717_ (
    .A(ex_reg_rs_msb_1[12]),
    .B(_03519_),
    .S(_02202_),
    .Z(_00161_)
  );
  MUX2_X1 _23718_ (
    .A(\rf[7] [15]),
    .B(\rf[3] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03520_)
  );
  AND2_X1 _23719_ (
    .A1(_08545_),
    .A2(_03520_),
    .ZN(_03521_)
  );
  INV_X1 _23720_ (
    .A(_03521_),
    .ZN(_03522_)
  );
  MUX2_X1 _23721_ (
    .A(\rf[5] [15]),
    .B(\rf[1] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03523_)
  );
  AND2_X1 _23722_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03523_),
    .ZN(_03524_)
  );
  INV_X1 _23723_ (
    .A(_03524_),
    .ZN(_03525_)
  );
  AND2_X1 _23724_ (
    .A1(_08544_),
    .A2(_03525_),
    .ZN(_03526_)
  );
  AND2_X1 _23725_ (
    .A1(_03522_),
    .A2(_03526_),
    .ZN(_03527_)
  );
  INV_X1 _23726_ (
    .A(_03527_),
    .ZN(_03528_)
  );
  MUX2_X1 _23727_ (
    .A(\rf[6] [15]),
    .B(\rf[2] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03529_)
  );
  AND2_X1 _23728_ (
    .A1(_08545_),
    .A2(_03529_),
    .ZN(_03530_)
  );
  INV_X1 _23729_ (
    .A(_03530_),
    .ZN(_03531_)
  );
  MUX2_X1 _23730_ (
    .A(\rf[4] [15]),
    .B(\rf[0] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03532_)
  );
  AND2_X1 _23731_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03532_),
    .ZN(_03533_)
  );
  INV_X1 _23732_ (
    .A(_03533_),
    .ZN(_03534_)
  );
  AND2_X1 _23733_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03534_),
    .ZN(_03535_)
  );
  AND2_X1 _23734_ (
    .A1(_03531_),
    .A2(_03535_),
    .ZN(_03536_)
  );
  INV_X1 _23735_ (
    .A(_03536_),
    .ZN(_03537_)
  );
  AND2_X1 _23736_ (
    .A1(_03528_),
    .A2(_03537_),
    .ZN(_03538_)
  );
  AND2_X1 _23737_ (
    .A1(\rf[14] [15]),
    .A2(_08545_),
    .ZN(_03539_)
  );
  INV_X1 _23738_ (
    .A(_03539_),
    .ZN(_03540_)
  );
  AND2_X1 _23739_ (
    .A1(\rf[12] [15]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_03541_)
  );
  INV_X1 _23740_ (
    .A(_03541_),
    .ZN(_03542_)
  );
  AND2_X1 _23741_ (
    .A1(_08546_),
    .A2(_03542_),
    .ZN(_03543_)
  );
  AND2_X1 _23742_ (
    .A1(_03540_),
    .A2(_03543_),
    .ZN(_03544_)
  );
  INV_X1 _23743_ (
    .A(_03544_),
    .ZN(_03545_)
  );
  AND2_X1 _23744_ (
    .A1(\rf[10] [15]),
    .A2(_08545_),
    .ZN(_03546_)
  );
  INV_X1 _23745_ (
    .A(_03546_),
    .ZN(_03547_)
  );
  AND2_X1 _23746_ (
    .A1(\rf[8] [15]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_03548_)
  );
  INV_X1 _23747_ (
    .A(_03548_),
    .ZN(_03549_)
  );
  AND2_X1 _23748_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[2]),
    .A2(_03549_),
    .ZN(_03550_)
  );
  AND2_X1 _23749_ (
    .A1(_03547_),
    .A2(_03550_),
    .ZN(_03551_)
  );
  INV_X1 _23750_ (
    .A(_03551_),
    .ZN(_03552_)
  );
  AND2_X1 _23751_ (
    .A1(_03545_),
    .A2(_03552_),
    .ZN(_03553_)
  );
  AND2_X1 _23752_ (
    .A1(\rf[15] [15]),
    .A2(_08545_),
    .ZN(_03554_)
  );
  INV_X1 _23753_ (
    .A(_03554_),
    .ZN(_03555_)
  );
  AND2_X1 _23754_ (
    .A1(\rf[13] [15]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_03556_)
  );
  INV_X1 _23755_ (
    .A(_03556_),
    .ZN(_03557_)
  );
  AND2_X1 _23756_ (
    .A1(_08546_),
    .A2(_03557_),
    .ZN(_03558_)
  );
  AND2_X1 _23757_ (
    .A1(_03555_),
    .A2(_03558_),
    .ZN(_03559_)
  );
  INV_X1 _23758_ (
    .A(_03559_),
    .ZN(_03560_)
  );
  AND2_X1 _23759_ (
    .A1(\rf[11] [15]),
    .A2(_08545_),
    .ZN(_03561_)
  );
  INV_X1 _23760_ (
    .A(_03561_),
    .ZN(_03562_)
  );
  AND2_X1 _23761_ (
    .A1(\rf[9] [15]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_03563_)
  );
  INV_X1 _23762_ (
    .A(_03563_),
    .ZN(_03564_)
  );
  AND2_X1 _23763_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[2]),
    .A2(_03564_),
    .ZN(_03565_)
  );
  AND2_X1 _23764_ (
    .A1(_03562_),
    .A2(_03565_),
    .ZN(_03566_)
  );
  INV_X1 _23765_ (
    .A(_03566_),
    .ZN(_03567_)
  );
  AND2_X1 _23766_ (
    .A1(_03560_),
    .A2(_03567_),
    .ZN(_03568_)
  );
  MUX2_X1 _23767_ (
    .A(_03553_),
    .B(_03568_),
    .S(_08544_),
    .Z(_03569_)
  );
  MUX2_X1 _23768_ (
    .A(_03538_),
    .B(_03569_),
    .S(_08547_),
    .Z(_03570_)
  );
  AND2_X1 _23769_ (
    .A1(\rf[30] [15]),
    .A2(_08546_),
    .ZN(_03571_)
  );
  INV_X1 _23770_ (
    .A(_03571_),
    .ZN(_03572_)
  );
  AND2_X1 _23771_ (
    .A1(\rf[26] [15]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03573_)
  );
  INV_X1 _23772_ (
    .A(_03573_),
    .ZN(_03574_)
  );
  AND2_X1 _23773_ (
    .A1(_08545_),
    .A2(_03574_),
    .ZN(_03575_)
  );
  AND2_X1 _23774_ (
    .A1(_03572_),
    .A2(_03575_),
    .ZN(_03576_)
  );
  INV_X1 _23775_ (
    .A(_03576_),
    .ZN(_03577_)
  );
  AND2_X1 _23776_ (
    .A1(\rf[24] [15]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03578_)
  );
  INV_X1 _23777_ (
    .A(_03578_),
    .ZN(_03579_)
  );
  AND2_X1 _23778_ (
    .A1(\rf[28] [15]),
    .A2(_08546_),
    .ZN(_03580_)
  );
  INV_X1 _23779_ (
    .A(_03580_),
    .ZN(_03581_)
  );
  AND2_X1 _23780_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03581_),
    .ZN(_03582_)
  );
  AND2_X1 _23781_ (
    .A1(_03579_),
    .A2(_03582_),
    .ZN(_03583_)
  );
  INV_X1 _23782_ (
    .A(_03583_),
    .ZN(_03584_)
  );
  AND2_X1 _23783_ (
    .A1(_03577_),
    .A2(_03584_),
    .ZN(_03585_)
  );
  MUX2_X1 _23784_ (
    .A(\rf[29] [15]),
    .B(\rf[25] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03586_)
  );
  AND2_X1 _23785_ (
    .A1(\rf[27] [15]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03587_)
  );
  MUX2_X1 _23786_ (
    .A(_03586_),
    .B(_03587_),
    .S(_08545_),
    .Z(_03588_)
  );
  MUX2_X1 _23787_ (
    .A(_03585_),
    .B(_03588_),
    .S(_08544_),
    .Z(_03589_)
  );
  AND2_X1 _23788_ (
    .A1(_08388_),
    .A2(_08546_),
    .ZN(_03590_)
  );
  INV_X1 _23789_ (
    .A(_03590_),
    .ZN(_03591_)
  );
  AND2_X1 _23790_ (
    .A1(_08289_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03592_)
  );
  INV_X1 _23791_ (
    .A(_03592_),
    .ZN(_03593_)
  );
  AND2_X1 _23792_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03593_),
    .ZN(_03594_)
  );
  AND2_X1 _23793_ (
    .A1(_03591_),
    .A2(_03594_),
    .ZN(_03595_)
  );
  INV_X1 _23794_ (
    .A(_03595_),
    .ZN(_03596_)
  );
  MUX2_X1 _23795_ (
    .A(\rf[22] [15]),
    .B(\rf[18] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03597_)
  );
  AND2_X1 _23796_ (
    .A1(_08545_),
    .A2(_03597_),
    .ZN(_03598_)
  );
  INV_X1 _23797_ (
    .A(_03598_),
    .ZN(_03599_)
  );
  AND2_X1 _23798_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03599_),
    .ZN(_03600_)
  );
  AND2_X1 _23799_ (
    .A1(_03596_),
    .A2(_03600_),
    .ZN(_03601_)
  );
  INV_X1 _23800_ (
    .A(_03601_),
    .ZN(_03602_)
  );
  AND2_X1 _23801_ (
    .A1(_08319_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03603_)
  );
  INV_X1 _23802_ (
    .A(_03603_),
    .ZN(_03604_)
  );
  AND2_X1 _23803_ (
    .A1(_08418_),
    .A2(_08546_),
    .ZN(_03605_)
  );
  INV_X1 _23804_ (
    .A(_03605_),
    .ZN(_03606_)
  );
  AND2_X1 _23805_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03606_),
    .ZN(_03607_)
  );
  AND2_X1 _23806_ (
    .A1(_03604_),
    .A2(_03607_),
    .ZN(_03608_)
  );
  INV_X1 _23807_ (
    .A(_03608_),
    .ZN(_03609_)
  );
  MUX2_X1 _23808_ (
    .A(\rf[23] [15]),
    .B(\rf[19] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03610_)
  );
  AND2_X1 _23809_ (
    .A1(_08545_),
    .A2(_03610_),
    .ZN(_03611_)
  );
  INV_X1 _23810_ (
    .A(_03611_),
    .ZN(_03612_)
  );
  AND2_X1 _23811_ (
    .A1(_08544_),
    .A2(_03612_),
    .ZN(_03613_)
  );
  AND2_X1 _23812_ (
    .A1(_03609_),
    .A2(_03613_),
    .ZN(_03614_)
  );
  INV_X1 _23813_ (
    .A(_03614_),
    .ZN(_03615_)
  );
  AND2_X1 _23814_ (
    .A1(_03602_),
    .A2(_03615_),
    .ZN(_03616_)
  );
  MUX2_X1 _23815_ (
    .A(_03589_),
    .B(_03616_),
    .S(ibuf_io_inst_0_bits_inst_rs2[3]),
    .Z(_03617_)
  );
  MUX2_X1 _23816_ (
    .A(_03570_),
    .B(_03617_),
    .S(_08572_),
    .Z(_03618_)
  );
  MUX2_X1 _23817_ (
    .A(_03618_),
    .B(_11656_),
    .S(_02233_),
    .Z(_03619_)
  );
  MUX2_X1 _23818_ (
    .A(ex_reg_rs_msb_1[13]),
    .B(_03619_),
    .S(_02202_),
    .Z(_00162_)
  );
  MUX2_X1 _23819_ (
    .A(\rf[1] [16]),
    .B(\rf[0] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_03620_)
  );
  MUX2_X1 _23820_ (
    .A(\rf[5] [16]),
    .B(\rf[4] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_03621_)
  );
  MUX2_X1 _23821_ (
    .A(_03620_),
    .B(_03621_),
    .S(_08546_),
    .Z(_03622_)
  );
  INV_X1 _23822_ (
    .A(_03622_),
    .ZN(_03623_)
  );
  AND2_X1 _23823_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_03623_),
    .ZN(_03624_)
  );
  INV_X1 _23824_ (
    .A(_03624_),
    .ZN(_03625_)
  );
  MUX2_X1 _23825_ (
    .A(\rf[12] [16]),
    .B(\rf[8] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03626_)
  );
  INV_X1 _23826_ (
    .A(_03626_),
    .ZN(_03627_)
  );
  AND2_X1 _23827_ (
    .A1(_02341_),
    .A2(_03627_),
    .ZN(_03628_)
  );
  INV_X1 _23828_ (
    .A(_03628_),
    .ZN(_03629_)
  );
  MUX2_X1 _23829_ (
    .A(\rf[13] [16]),
    .B(\rf[9] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03630_)
  );
  INV_X1 _23830_ (
    .A(_03630_),
    .ZN(_03631_)
  );
  AND2_X1 _23831_ (
    .A1(_09692_),
    .A2(_03631_),
    .ZN(_03632_)
  );
  INV_X1 _23832_ (
    .A(_03632_),
    .ZN(_03633_)
  );
  AND2_X1 _23833_ (
    .A1(_03629_),
    .A2(_03633_),
    .ZN(_03634_)
  );
  AND2_X1 _23834_ (
    .A1(_03625_),
    .A2(_03634_),
    .ZN(_03635_)
  );
  MUX2_X1 _23835_ (
    .A(\rf[3] [16]),
    .B(\rf[2] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_03636_)
  );
  MUX2_X1 _23836_ (
    .A(\rf[7] [16]),
    .B(\rf[6] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_03637_)
  );
  MUX2_X1 _23837_ (
    .A(_03636_),
    .B(_03637_),
    .S(_08546_),
    .Z(_03638_)
  );
  INV_X1 _23838_ (
    .A(_03638_),
    .ZN(_03639_)
  );
  AND2_X1 _23839_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_03639_),
    .ZN(_03640_)
  );
  INV_X1 _23840_ (
    .A(_03640_),
    .ZN(_03641_)
  );
  MUX2_X1 _23841_ (
    .A(\rf[14] [16]),
    .B(\rf[10] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03642_)
  );
  INV_X1 _23842_ (
    .A(_03642_),
    .ZN(_03643_)
  );
  AND2_X1 _23843_ (
    .A1(_02341_),
    .A2(_03643_),
    .ZN(_03644_)
  );
  INV_X1 _23844_ (
    .A(_03644_),
    .ZN(_03645_)
  );
  MUX2_X1 _23845_ (
    .A(\rf[15] [16]),
    .B(\rf[11] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03646_)
  );
  INV_X1 _23846_ (
    .A(_03646_),
    .ZN(_03647_)
  );
  AND2_X1 _23847_ (
    .A1(_09692_),
    .A2(_03647_),
    .ZN(_03648_)
  );
  INV_X1 _23848_ (
    .A(_03648_),
    .ZN(_03649_)
  );
  AND2_X1 _23849_ (
    .A1(_03645_),
    .A2(_03649_),
    .ZN(_03650_)
  );
  AND2_X1 _23850_ (
    .A1(_03641_),
    .A2(_03650_),
    .ZN(_03651_)
  );
  MUX2_X1 _23851_ (
    .A(_03635_),
    .B(_03651_),
    .S(_08545_),
    .Z(_03652_)
  );
  AND2_X1 _23852_ (
    .A1(_08320_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03653_)
  );
  INV_X1 _23853_ (
    .A(_03653_),
    .ZN(_03654_)
  );
  AND2_X1 _23854_ (
    .A1(_08419_),
    .A2(_08546_),
    .ZN(_03655_)
  );
  INV_X1 _23855_ (
    .A(_03655_),
    .ZN(_03656_)
  );
  AND2_X1 _23856_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03656_),
    .ZN(_03657_)
  );
  AND2_X1 _23857_ (
    .A1(_03654_),
    .A2(_03657_),
    .ZN(_03658_)
  );
  INV_X1 _23858_ (
    .A(_03658_),
    .ZN(_03659_)
  );
  MUX2_X1 _23859_ (
    .A(\rf[23] [16]),
    .B(\rf[19] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03660_)
  );
  AND2_X1 _23860_ (
    .A1(_08545_),
    .A2(_03660_),
    .ZN(_03661_)
  );
  INV_X1 _23861_ (
    .A(_03661_),
    .ZN(_03662_)
  );
  AND2_X1 _23862_ (
    .A1(_08544_),
    .A2(_03662_),
    .ZN(_03663_)
  );
  AND2_X1 _23863_ (
    .A1(_03659_),
    .A2(_03663_),
    .ZN(_03664_)
  );
  INV_X1 _23864_ (
    .A(_03664_),
    .ZN(_03665_)
  );
  AND2_X1 _23865_ (
    .A1(_08389_),
    .A2(_08546_),
    .ZN(_03666_)
  );
  INV_X1 _23866_ (
    .A(_03666_),
    .ZN(_03667_)
  );
  AND2_X1 _23867_ (
    .A1(_08290_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03668_)
  );
  INV_X1 _23868_ (
    .A(_03668_),
    .ZN(_03669_)
  );
  AND2_X1 _23869_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03669_),
    .ZN(_03670_)
  );
  AND2_X1 _23870_ (
    .A1(_03667_),
    .A2(_03670_),
    .ZN(_03671_)
  );
  INV_X1 _23871_ (
    .A(_03671_),
    .ZN(_03672_)
  );
  MUX2_X1 _23872_ (
    .A(\rf[22] [16]),
    .B(\rf[18] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03673_)
  );
  AND2_X1 _23873_ (
    .A1(_08545_),
    .A2(_03673_),
    .ZN(_03674_)
  );
  INV_X1 _23874_ (
    .A(_03674_),
    .ZN(_03675_)
  );
  AND2_X1 _23875_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03675_),
    .ZN(_03676_)
  );
  AND2_X1 _23876_ (
    .A1(_03672_),
    .A2(_03676_),
    .ZN(_03677_)
  );
  INV_X1 _23877_ (
    .A(_03677_),
    .ZN(_03678_)
  );
  AND2_X1 _23878_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_03665_),
    .ZN(_03679_)
  );
  AND2_X1 _23879_ (
    .A1(_03678_),
    .A2(_03679_),
    .ZN(_03680_)
  );
  INV_X1 _23880_ (
    .A(_03680_),
    .ZN(_03681_)
  );
  AND2_X1 _23881_ (
    .A1(_08446_),
    .A2(_08546_),
    .ZN(_03682_)
  );
  INV_X1 _23882_ (
    .A(_03682_),
    .ZN(_03683_)
  );
  AND2_X1 _23883_ (
    .A1(_08516_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03684_)
  );
  INV_X1 _23884_ (
    .A(_03684_),
    .ZN(_03685_)
  );
  AND2_X1 _23885_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03685_),
    .ZN(_03686_)
  );
  AND2_X1 _23886_ (
    .A1(_03683_),
    .A2(_03686_),
    .ZN(_03687_)
  );
  INV_X1 _23887_ (
    .A(_03687_),
    .ZN(_03688_)
  );
  MUX2_X1 _23888_ (
    .A(\rf[30] [16]),
    .B(\rf[26] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03689_)
  );
  AND2_X1 _23889_ (
    .A1(_08545_),
    .A2(_03689_),
    .ZN(_03690_)
  );
  INV_X1 _23890_ (
    .A(_03690_),
    .ZN(_03691_)
  );
  AND2_X1 _23891_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03691_),
    .ZN(_03692_)
  );
  AND2_X1 _23892_ (
    .A1(_03688_),
    .A2(_03692_),
    .ZN(_03693_)
  );
  INV_X1 _23893_ (
    .A(_03693_),
    .ZN(_03694_)
  );
  MUX2_X1 _23894_ (
    .A(\rf[29] [16]),
    .B(\rf[25] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03695_)
  );
  AND2_X1 _23895_ (
    .A1(\rf[27] [16]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03696_)
  );
  MUX2_X1 _23896_ (
    .A(_03695_),
    .B(_03696_),
    .S(_08545_),
    .Z(_03697_)
  );
  INV_X1 _23897_ (
    .A(_03697_),
    .ZN(_03698_)
  );
  AND2_X1 _23898_ (
    .A1(_08544_),
    .A2(_03698_),
    .ZN(_03699_)
  );
  INV_X1 _23899_ (
    .A(_03699_),
    .ZN(_03700_)
  );
  AND2_X1 _23900_ (
    .A1(_08547_),
    .A2(_03700_),
    .ZN(_03701_)
  );
  AND2_X1 _23901_ (
    .A1(_03694_),
    .A2(_03701_),
    .ZN(_03702_)
  );
  INV_X1 _23902_ (
    .A(_03702_),
    .ZN(_03703_)
  );
  AND2_X1 _23903_ (
    .A1(_03681_),
    .A2(_03703_),
    .ZN(_03704_)
  );
  INV_X1 _23904_ (
    .A(_03704_),
    .ZN(_03705_)
  );
  MUX2_X1 _23905_ (
    .A(_03652_),
    .B(_03705_),
    .S(_08572_),
    .Z(_03706_)
  );
  MUX2_X1 _23906_ (
    .A(_03706_),
    .B(_11766_),
    .S(_02233_),
    .Z(_03707_)
  );
  MUX2_X1 _23907_ (
    .A(ex_reg_rs_msb_1[14]),
    .B(_03707_),
    .S(_02202_),
    .Z(_00163_)
  );
  MUX2_X1 _23908_ (
    .A(\rf[1] [17]),
    .B(\rf[0] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_03708_)
  );
  MUX2_X1 _23909_ (
    .A(\rf[5] [17]),
    .B(\rf[4] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_03709_)
  );
  MUX2_X1 _23910_ (
    .A(_03708_),
    .B(_03709_),
    .S(_08546_),
    .Z(_03710_)
  );
  INV_X1 _23911_ (
    .A(_03710_),
    .ZN(_03711_)
  );
  AND2_X1 _23912_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_03711_),
    .ZN(_03712_)
  );
  INV_X1 _23913_ (
    .A(_03712_),
    .ZN(_03713_)
  );
  MUX2_X1 _23914_ (
    .A(\rf[12] [17]),
    .B(\rf[8] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03714_)
  );
  INV_X1 _23915_ (
    .A(_03714_),
    .ZN(_03715_)
  );
  AND2_X1 _23916_ (
    .A1(_02341_),
    .A2(_03715_),
    .ZN(_03716_)
  );
  INV_X1 _23917_ (
    .A(_03716_),
    .ZN(_03717_)
  );
  MUX2_X1 _23918_ (
    .A(\rf[13] [17]),
    .B(\rf[9] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03718_)
  );
  INV_X1 _23919_ (
    .A(_03718_),
    .ZN(_03719_)
  );
  AND2_X1 _23920_ (
    .A1(_09692_),
    .A2(_03719_),
    .ZN(_03720_)
  );
  INV_X1 _23921_ (
    .A(_03720_),
    .ZN(_03721_)
  );
  AND2_X1 _23922_ (
    .A1(_03717_),
    .A2(_03721_),
    .ZN(_03722_)
  );
  AND2_X1 _23923_ (
    .A1(_03713_),
    .A2(_03722_),
    .ZN(_03723_)
  );
  MUX2_X1 _23924_ (
    .A(\rf[3] [17]),
    .B(\rf[2] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_03724_)
  );
  MUX2_X1 _23925_ (
    .A(\rf[7] [17]),
    .B(\rf[6] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_03725_)
  );
  MUX2_X1 _23926_ (
    .A(_03724_),
    .B(_03725_),
    .S(_08546_),
    .Z(_03726_)
  );
  INV_X1 _23927_ (
    .A(_03726_),
    .ZN(_03727_)
  );
  AND2_X1 _23928_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_03727_),
    .ZN(_03728_)
  );
  INV_X1 _23929_ (
    .A(_03728_),
    .ZN(_03729_)
  );
  MUX2_X1 _23930_ (
    .A(\rf[14] [17]),
    .B(\rf[10] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03730_)
  );
  INV_X1 _23931_ (
    .A(_03730_),
    .ZN(_03731_)
  );
  AND2_X1 _23932_ (
    .A1(_02341_),
    .A2(_03731_),
    .ZN(_03732_)
  );
  INV_X1 _23933_ (
    .A(_03732_),
    .ZN(_03733_)
  );
  MUX2_X1 _23934_ (
    .A(\rf[15] [17]),
    .B(\rf[11] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03734_)
  );
  INV_X1 _23935_ (
    .A(_03734_),
    .ZN(_03735_)
  );
  AND2_X1 _23936_ (
    .A1(_09692_),
    .A2(_03735_),
    .ZN(_03736_)
  );
  INV_X1 _23937_ (
    .A(_03736_),
    .ZN(_03737_)
  );
  AND2_X1 _23938_ (
    .A1(_03733_),
    .A2(_03737_),
    .ZN(_03738_)
  );
  AND2_X1 _23939_ (
    .A1(_03729_),
    .A2(_03738_),
    .ZN(_03739_)
  );
  MUX2_X1 _23940_ (
    .A(_03723_),
    .B(_03739_),
    .S(_08545_),
    .Z(_03740_)
  );
  AND2_X1 _23941_ (
    .A1(_08321_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03741_)
  );
  INV_X1 _23942_ (
    .A(_03741_),
    .ZN(_03742_)
  );
  AND2_X1 _23943_ (
    .A1(_08420_),
    .A2(_08546_),
    .ZN(_03743_)
  );
  INV_X1 _23944_ (
    .A(_03743_),
    .ZN(_03744_)
  );
  AND2_X1 _23945_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03744_),
    .ZN(_03745_)
  );
  AND2_X1 _23946_ (
    .A1(_03742_),
    .A2(_03745_),
    .ZN(_03746_)
  );
  INV_X1 _23947_ (
    .A(_03746_),
    .ZN(_03747_)
  );
  MUX2_X1 _23948_ (
    .A(\rf[23] [17]),
    .B(\rf[19] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03748_)
  );
  AND2_X1 _23949_ (
    .A1(_08545_),
    .A2(_03748_),
    .ZN(_03749_)
  );
  INV_X1 _23950_ (
    .A(_03749_),
    .ZN(_03750_)
  );
  AND2_X1 _23951_ (
    .A1(_08544_),
    .A2(_03750_),
    .ZN(_03751_)
  );
  AND2_X1 _23952_ (
    .A1(_03747_),
    .A2(_03751_),
    .ZN(_03752_)
  );
  INV_X1 _23953_ (
    .A(_03752_),
    .ZN(_03753_)
  );
  AND2_X1 _23954_ (
    .A1(_08390_),
    .A2(_08546_),
    .ZN(_03754_)
  );
  INV_X1 _23955_ (
    .A(_03754_),
    .ZN(_03755_)
  );
  AND2_X1 _23956_ (
    .A1(_08291_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03756_)
  );
  INV_X1 _23957_ (
    .A(_03756_),
    .ZN(_03757_)
  );
  AND2_X1 _23958_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03757_),
    .ZN(_03758_)
  );
  AND2_X1 _23959_ (
    .A1(_03755_),
    .A2(_03758_),
    .ZN(_03759_)
  );
  INV_X1 _23960_ (
    .A(_03759_),
    .ZN(_03760_)
  );
  MUX2_X1 _23961_ (
    .A(\rf[22] [17]),
    .B(\rf[18] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03761_)
  );
  AND2_X1 _23962_ (
    .A1(_08545_),
    .A2(_03761_),
    .ZN(_03762_)
  );
  INV_X1 _23963_ (
    .A(_03762_),
    .ZN(_03763_)
  );
  AND2_X1 _23964_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03763_),
    .ZN(_03764_)
  );
  AND2_X1 _23965_ (
    .A1(_03760_),
    .A2(_03764_),
    .ZN(_03765_)
  );
  INV_X1 _23966_ (
    .A(_03765_),
    .ZN(_03766_)
  );
  AND2_X1 _23967_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_03753_),
    .ZN(_03767_)
  );
  AND2_X1 _23968_ (
    .A1(_03766_),
    .A2(_03767_),
    .ZN(_03768_)
  );
  INV_X1 _23969_ (
    .A(_03768_),
    .ZN(_03769_)
  );
  AND2_X1 _23970_ (
    .A1(_08447_),
    .A2(_08546_),
    .ZN(_03770_)
  );
  INV_X1 _23971_ (
    .A(_03770_),
    .ZN(_03771_)
  );
  AND2_X1 _23972_ (
    .A1(_08517_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03772_)
  );
  INV_X1 _23973_ (
    .A(_03772_),
    .ZN(_03773_)
  );
  AND2_X1 _23974_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03773_),
    .ZN(_03774_)
  );
  AND2_X1 _23975_ (
    .A1(_03771_),
    .A2(_03774_),
    .ZN(_03775_)
  );
  INV_X1 _23976_ (
    .A(_03775_),
    .ZN(_03776_)
  );
  MUX2_X1 _23977_ (
    .A(\rf[30] [17]),
    .B(\rf[26] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03777_)
  );
  AND2_X1 _23978_ (
    .A1(_08545_),
    .A2(_03777_),
    .ZN(_03778_)
  );
  INV_X1 _23979_ (
    .A(_03778_),
    .ZN(_03779_)
  );
  AND2_X1 _23980_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03779_),
    .ZN(_03780_)
  );
  AND2_X1 _23981_ (
    .A1(_03776_),
    .A2(_03780_),
    .ZN(_03781_)
  );
  INV_X1 _23982_ (
    .A(_03781_),
    .ZN(_03782_)
  );
  MUX2_X1 _23983_ (
    .A(\rf[29] [17]),
    .B(\rf[25] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03783_)
  );
  AND2_X1 _23984_ (
    .A1(\rf[27] [17]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03784_)
  );
  MUX2_X1 _23985_ (
    .A(_03783_),
    .B(_03784_),
    .S(_08545_),
    .Z(_03785_)
  );
  INV_X1 _23986_ (
    .A(_03785_),
    .ZN(_03786_)
  );
  AND2_X1 _23987_ (
    .A1(_08544_),
    .A2(_03786_),
    .ZN(_03787_)
  );
  INV_X1 _23988_ (
    .A(_03787_),
    .ZN(_03788_)
  );
  AND2_X1 _23989_ (
    .A1(_08547_),
    .A2(_03788_),
    .ZN(_03789_)
  );
  AND2_X1 _23990_ (
    .A1(_03782_),
    .A2(_03789_),
    .ZN(_03790_)
  );
  INV_X1 _23991_ (
    .A(_03790_),
    .ZN(_03791_)
  );
  AND2_X1 _23992_ (
    .A1(_03769_),
    .A2(_03791_),
    .ZN(_03792_)
  );
  INV_X1 _23993_ (
    .A(_03792_),
    .ZN(_03793_)
  );
  MUX2_X1 _23994_ (
    .A(_03740_),
    .B(_03793_),
    .S(_08572_),
    .Z(_03794_)
  );
  MUX2_X1 _23995_ (
    .A(_03794_),
    .B(_11882_),
    .S(_02233_),
    .Z(_03795_)
  );
  MUX2_X1 _23996_ (
    .A(ex_reg_rs_msb_1[15]),
    .B(_03795_),
    .S(_02202_),
    .Z(_00164_)
  );
  AND2_X1 _23997_ (
    .A1(_08342_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03796_)
  );
  INV_X1 _23998_ (
    .A(_03796_),
    .ZN(_03797_)
  );
  AND2_X1 _23999_ (
    .A1(_08480_),
    .A2(_08546_),
    .ZN(_03798_)
  );
  INV_X1 _24000_ (
    .A(_03798_),
    .ZN(_03799_)
  );
  AND2_X1 _24001_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03799_),
    .ZN(_03800_)
  );
  AND2_X1 _24002_ (
    .A1(_03797_),
    .A2(_03800_),
    .ZN(_03801_)
  );
  INV_X1 _24003_ (
    .A(_03801_),
    .ZN(_03802_)
  );
  MUX2_X1 _24004_ (
    .A(\rf[15] [18]),
    .B(\rf[11] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03803_)
  );
  AND2_X1 _24005_ (
    .A1(_08544_),
    .A2(_03803_),
    .ZN(_03804_)
  );
  INV_X1 _24006_ (
    .A(_03804_),
    .ZN(_03805_)
  );
  AND2_X1 _24007_ (
    .A1(_08545_),
    .A2(_03805_),
    .ZN(_03806_)
  );
  AND2_X1 _24008_ (
    .A1(_03802_),
    .A2(_03806_),
    .ZN(_03807_)
  );
  INV_X1 _24009_ (
    .A(_03807_),
    .ZN(_03808_)
  );
  AND2_X1 _24010_ (
    .A1(_08363_),
    .A2(_08546_),
    .ZN(_03809_)
  );
  INV_X1 _24011_ (
    .A(_03809_),
    .ZN(_03810_)
  );
  AND2_X1 _24012_ (
    .A1(_08264_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03811_)
  );
  INV_X1 _24013_ (
    .A(_03811_),
    .ZN(_03812_)
  );
  AND2_X1 _24014_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03812_),
    .ZN(_03813_)
  );
  AND2_X1 _24015_ (
    .A1(_03810_),
    .A2(_03813_),
    .ZN(_03814_)
  );
  INV_X1 _24016_ (
    .A(_03814_),
    .ZN(_03815_)
  );
  MUX2_X1 _24017_ (
    .A(\rf[13] [18]),
    .B(\rf[9] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03816_)
  );
  AND2_X1 _24018_ (
    .A1(_08544_),
    .A2(_03816_),
    .ZN(_03817_)
  );
  INV_X1 _24019_ (
    .A(_03817_),
    .ZN(_03818_)
  );
  AND2_X1 _24020_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03818_),
    .ZN(_03819_)
  );
  AND2_X1 _24021_ (
    .A1(_03815_),
    .A2(_03819_),
    .ZN(_03820_)
  );
  INV_X1 _24022_ (
    .A(_03820_),
    .ZN(_03821_)
  );
  AND2_X1 _24023_ (
    .A1(_08547_),
    .A2(_03821_),
    .ZN(_03822_)
  );
  AND2_X1 _24024_ (
    .A1(_03808_),
    .A2(_03822_),
    .ZN(_03823_)
  );
  INV_X1 _24025_ (
    .A(_03823_),
    .ZN(_03824_)
  );
  MUX2_X1 _24026_ (
    .A(\rf[6] [18]),
    .B(\rf[2] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03825_)
  );
  AND2_X1 _24027_ (
    .A1(_08545_),
    .A2(_03825_),
    .ZN(_03826_)
  );
  INV_X1 _24028_ (
    .A(_03826_),
    .ZN(_03827_)
  );
  MUX2_X1 _24029_ (
    .A(\rf[4] [18]),
    .B(\rf[0] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03828_)
  );
  AND2_X1 _24030_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03828_),
    .ZN(_03829_)
  );
  INV_X1 _24031_ (
    .A(_03829_),
    .ZN(_03830_)
  );
  AND2_X1 _24032_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03830_),
    .ZN(_03831_)
  );
  AND2_X1 _24033_ (
    .A1(_03827_),
    .A2(_03831_),
    .ZN(_03832_)
  );
  INV_X1 _24034_ (
    .A(_03832_),
    .ZN(_03833_)
  );
  MUX2_X1 _24035_ (
    .A(\rf[7] [18]),
    .B(\rf[3] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03834_)
  );
  AND2_X1 _24036_ (
    .A1(_08545_),
    .A2(_03834_),
    .ZN(_03835_)
  );
  INV_X1 _24037_ (
    .A(_03835_),
    .ZN(_03836_)
  );
  MUX2_X1 _24038_ (
    .A(\rf[5] [18]),
    .B(\rf[1] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03837_)
  );
  AND2_X1 _24039_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03837_),
    .ZN(_03838_)
  );
  INV_X1 _24040_ (
    .A(_03838_),
    .ZN(_03839_)
  );
  AND2_X1 _24041_ (
    .A1(_08544_),
    .A2(_03839_),
    .ZN(_03840_)
  );
  AND2_X1 _24042_ (
    .A1(_03836_),
    .A2(_03840_),
    .ZN(_03841_)
  );
  INV_X1 _24043_ (
    .A(_03841_),
    .ZN(_03842_)
  );
  AND2_X1 _24044_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_03842_),
    .ZN(_03843_)
  );
  AND2_X1 _24045_ (
    .A1(_03833_),
    .A2(_03843_),
    .ZN(_03844_)
  );
  INV_X1 _24046_ (
    .A(_03844_),
    .ZN(_03845_)
  );
  AND2_X1 _24047_ (
    .A1(_03824_),
    .A2(_03845_),
    .ZN(_03846_)
  );
  AND2_X1 _24048_ (
    .A1(_08322_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03847_)
  );
  INV_X1 _24049_ (
    .A(_03847_),
    .ZN(_03848_)
  );
  AND2_X1 _24050_ (
    .A1(_08421_),
    .A2(_08546_),
    .ZN(_03849_)
  );
  INV_X1 _24051_ (
    .A(_03849_),
    .ZN(_03850_)
  );
  AND2_X1 _24052_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03850_),
    .ZN(_03851_)
  );
  AND2_X1 _24053_ (
    .A1(_03848_),
    .A2(_03851_),
    .ZN(_03852_)
  );
  INV_X1 _24054_ (
    .A(_03852_),
    .ZN(_03853_)
  );
  MUX2_X1 _24055_ (
    .A(\rf[23] [18]),
    .B(\rf[19] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03854_)
  );
  AND2_X1 _24056_ (
    .A1(_08545_),
    .A2(_03854_),
    .ZN(_03855_)
  );
  INV_X1 _24057_ (
    .A(_03855_),
    .ZN(_03856_)
  );
  AND2_X1 _24058_ (
    .A1(_08544_),
    .A2(_03856_),
    .ZN(_03857_)
  );
  AND2_X1 _24059_ (
    .A1(_03853_),
    .A2(_03857_),
    .ZN(_03858_)
  );
  INV_X1 _24060_ (
    .A(_03858_),
    .ZN(_03859_)
  );
  AND2_X1 _24061_ (
    .A1(_08391_),
    .A2(_08546_),
    .ZN(_03860_)
  );
  INV_X1 _24062_ (
    .A(_03860_),
    .ZN(_03861_)
  );
  AND2_X1 _24063_ (
    .A1(_08292_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03862_)
  );
  INV_X1 _24064_ (
    .A(_03862_),
    .ZN(_03863_)
  );
  AND2_X1 _24065_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03863_),
    .ZN(_03864_)
  );
  AND2_X1 _24066_ (
    .A1(_03861_),
    .A2(_03864_),
    .ZN(_03865_)
  );
  INV_X1 _24067_ (
    .A(_03865_),
    .ZN(_03866_)
  );
  MUX2_X1 _24068_ (
    .A(\rf[22] [18]),
    .B(\rf[18] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03867_)
  );
  AND2_X1 _24069_ (
    .A1(_08545_),
    .A2(_03867_),
    .ZN(_03868_)
  );
  INV_X1 _24070_ (
    .A(_03868_),
    .ZN(_03869_)
  );
  AND2_X1 _24071_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03869_),
    .ZN(_03870_)
  );
  AND2_X1 _24072_ (
    .A1(_03866_),
    .A2(_03870_),
    .ZN(_03871_)
  );
  INV_X1 _24073_ (
    .A(_03871_),
    .ZN(_03872_)
  );
  AND2_X1 _24074_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_03859_),
    .ZN(_03873_)
  );
  AND2_X1 _24075_ (
    .A1(_03872_),
    .A2(_03873_),
    .ZN(_03874_)
  );
  INV_X1 _24076_ (
    .A(_03874_),
    .ZN(_03875_)
  );
  AND2_X1 _24077_ (
    .A1(_08448_),
    .A2(_08546_),
    .ZN(_03876_)
  );
  INV_X1 _24078_ (
    .A(_03876_),
    .ZN(_03877_)
  );
  AND2_X1 _24079_ (
    .A1(_08518_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03878_)
  );
  INV_X1 _24080_ (
    .A(_03878_),
    .ZN(_03879_)
  );
  AND2_X1 _24081_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03879_),
    .ZN(_03880_)
  );
  AND2_X1 _24082_ (
    .A1(_03877_),
    .A2(_03880_),
    .ZN(_03881_)
  );
  INV_X1 _24083_ (
    .A(_03881_),
    .ZN(_03882_)
  );
  MUX2_X1 _24084_ (
    .A(\rf[30] [18]),
    .B(\rf[26] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03883_)
  );
  AND2_X1 _24085_ (
    .A1(_08545_),
    .A2(_03883_),
    .ZN(_03884_)
  );
  INV_X1 _24086_ (
    .A(_03884_),
    .ZN(_03885_)
  );
  AND2_X1 _24087_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03885_),
    .ZN(_03886_)
  );
  AND2_X1 _24088_ (
    .A1(_03882_),
    .A2(_03886_),
    .ZN(_03887_)
  );
  INV_X1 _24089_ (
    .A(_03887_),
    .ZN(_03888_)
  );
  MUX2_X1 _24090_ (
    .A(\rf[29] [18]),
    .B(\rf[25] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03889_)
  );
  AND2_X1 _24091_ (
    .A1(\rf[27] [18]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03890_)
  );
  MUX2_X1 _24092_ (
    .A(_03889_),
    .B(_03890_),
    .S(_08545_),
    .Z(_03891_)
  );
  INV_X1 _24093_ (
    .A(_03891_),
    .ZN(_03892_)
  );
  AND2_X1 _24094_ (
    .A1(_08544_),
    .A2(_03892_),
    .ZN(_03893_)
  );
  INV_X1 _24095_ (
    .A(_03893_),
    .ZN(_03894_)
  );
  AND2_X1 _24096_ (
    .A1(_08547_),
    .A2(_03894_),
    .ZN(_03895_)
  );
  AND2_X1 _24097_ (
    .A1(_03888_),
    .A2(_03895_),
    .ZN(_03896_)
  );
  INV_X1 _24098_ (
    .A(_03896_),
    .ZN(_03897_)
  );
  AND2_X1 _24099_ (
    .A1(_03875_),
    .A2(_03897_),
    .ZN(_03898_)
  );
  MUX2_X1 _24100_ (
    .A(_03846_),
    .B(_03898_),
    .S(_08572_),
    .Z(_03899_)
  );
  INV_X1 _24101_ (
    .A(_03899_),
    .ZN(_03900_)
  );
  MUX2_X1 _24102_ (
    .A(_03900_),
    .B(_12088_),
    .S(_02233_),
    .Z(_03901_)
  );
  MUX2_X1 _24103_ (
    .A(ex_reg_rs_msb_1[16]),
    .B(_03901_),
    .S(_02202_),
    .Z(_00165_)
  );
  MUX2_X1 _24104_ (
    .A(\rf[7] [19]),
    .B(\rf[3] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03902_)
  );
  AND2_X1 _24105_ (
    .A1(_08545_),
    .A2(_03902_),
    .ZN(_03903_)
  );
  INV_X1 _24106_ (
    .A(_03903_),
    .ZN(_03904_)
  );
  MUX2_X1 _24107_ (
    .A(\rf[5] [19]),
    .B(\rf[1] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03905_)
  );
  AND2_X1 _24108_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03905_),
    .ZN(_03906_)
  );
  INV_X1 _24109_ (
    .A(_03906_),
    .ZN(_03907_)
  );
  AND2_X1 _24110_ (
    .A1(_08544_),
    .A2(_03907_),
    .ZN(_03908_)
  );
  AND2_X1 _24111_ (
    .A1(_03904_),
    .A2(_03908_),
    .ZN(_03909_)
  );
  INV_X1 _24112_ (
    .A(_03909_),
    .ZN(_03910_)
  );
  MUX2_X1 _24113_ (
    .A(\rf[6] [19]),
    .B(\rf[2] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03911_)
  );
  AND2_X1 _24114_ (
    .A1(_08545_),
    .A2(_03911_),
    .ZN(_03912_)
  );
  INV_X1 _24115_ (
    .A(_03912_),
    .ZN(_03913_)
  );
  MUX2_X1 _24116_ (
    .A(\rf[4] [19]),
    .B(\rf[0] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03914_)
  );
  AND2_X1 _24117_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03914_),
    .ZN(_03915_)
  );
  INV_X1 _24118_ (
    .A(_03915_),
    .ZN(_03916_)
  );
  AND2_X1 _24119_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03916_),
    .ZN(_03917_)
  );
  AND2_X1 _24120_ (
    .A1(_03913_),
    .A2(_03917_),
    .ZN(_03918_)
  );
  INV_X1 _24121_ (
    .A(_03918_),
    .ZN(_03919_)
  );
  AND2_X1 _24122_ (
    .A1(_03910_),
    .A2(_03919_),
    .ZN(_03920_)
  );
  AND2_X1 _24123_ (
    .A1(\rf[14] [19]),
    .A2(_08545_),
    .ZN(_03921_)
  );
  INV_X1 _24124_ (
    .A(_03921_),
    .ZN(_03922_)
  );
  AND2_X1 _24125_ (
    .A1(\rf[12] [19]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_03923_)
  );
  INV_X1 _24126_ (
    .A(_03923_),
    .ZN(_03924_)
  );
  AND2_X1 _24127_ (
    .A1(_08546_),
    .A2(_03924_),
    .ZN(_03925_)
  );
  AND2_X1 _24128_ (
    .A1(_03922_),
    .A2(_03925_),
    .ZN(_03926_)
  );
  INV_X1 _24129_ (
    .A(_03926_),
    .ZN(_03927_)
  );
  AND2_X1 _24130_ (
    .A1(\rf[10] [19]),
    .A2(_08545_),
    .ZN(_03928_)
  );
  INV_X1 _24131_ (
    .A(_03928_),
    .ZN(_03929_)
  );
  AND2_X1 _24132_ (
    .A1(\rf[8] [19]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_03930_)
  );
  INV_X1 _24133_ (
    .A(_03930_),
    .ZN(_03931_)
  );
  AND2_X1 _24134_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[2]),
    .A2(_03931_),
    .ZN(_03932_)
  );
  AND2_X1 _24135_ (
    .A1(_03929_),
    .A2(_03932_),
    .ZN(_03933_)
  );
  INV_X1 _24136_ (
    .A(_03933_),
    .ZN(_03934_)
  );
  AND2_X1 _24137_ (
    .A1(_03927_),
    .A2(_03934_),
    .ZN(_03935_)
  );
  AND2_X1 _24138_ (
    .A1(\rf[15] [19]),
    .A2(_08545_),
    .ZN(_03936_)
  );
  INV_X1 _24139_ (
    .A(_03936_),
    .ZN(_03937_)
  );
  AND2_X1 _24140_ (
    .A1(\rf[13] [19]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_03938_)
  );
  INV_X1 _24141_ (
    .A(_03938_),
    .ZN(_03939_)
  );
  AND2_X1 _24142_ (
    .A1(_08546_),
    .A2(_03939_),
    .ZN(_03940_)
  );
  AND2_X1 _24143_ (
    .A1(_03937_),
    .A2(_03940_),
    .ZN(_03941_)
  );
  INV_X1 _24144_ (
    .A(_03941_),
    .ZN(_03942_)
  );
  AND2_X1 _24145_ (
    .A1(\rf[11] [19]),
    .A2(_08545_),
    .ZN(_03943_)
  );
  INV_X1 _24146_ (
    .A(_03943_),
    .ZN(_03944_)
  );
  AND2_X1 _24147_ (
    .A1(\rf[9] [19]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_03945_)
  );
  INV_X1 _24148_ (
    .A(_03945_),
    .ZN(_03946_)
  );
  AND2_X1 _24149_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[2]),
    .A2(_03946_),
    .ZN(_03947_)
  );
  AND2_X1 _24150_ (
    .A1(_03944_),
    .A2(_03947_),
    .ZN(_03948_)
  );
  INV_X1 _24151_ (
    .A(_03948_),
    .ZN(_03949_)
  );
  AND2_X1 _24152_ (
    .A1(_03942_),
    .A2(_03949_),
    .ZN(_03950_)
  );
  MUX2_X1 _24153_ (
    .A(_03935_),
    .B(_03950_),
    .S(_08544_),
    .Z(_03951_)
  );
  MUX2_X1 _24154_ (
    .A(_03920_),
    .B(_03951_),
    .S(_08547_),
    .Z(_03952_)
  );
  AND2_X1 _24155_ (
    .A1(\rf[30] [19]),
    .A2(_08546_),
    .ZN(_03953_)
  );
  INV_X1 _24156_ (
    .A(_03953_),
    .ZN(_03954_)
  );
  AND2_X1 _24157_ (
    .A1(\rf[26] [19]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03955_)
  );
  INV_X1 _24158_ (
    .A(_03955_),
    .ZN(_03956_)
  );
  AND2_X1 _24159_ (
    .A1(_08545_),
    .A2(_03956_),
    .ZN(_03957_)
  );
  AND2_X1 _24160_ (
    .A1(_03954_),
    .A2(_03957_),
    .ZN(_03958_)
  );
  INV_X1 _24161_ (
    .A(_03958_),
    .ZN(_03959_)
  );
  AND2_X1 _24162_ (
    .A1(\rf[24] [19]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03960_)
  );
  INV_X1 _24163_ (
    .A(_03960_),
    .ZN(_03961_)
  );
  AND2_X1 _24164_ (
    .A1(\rf[28] [19]),
    .A2(_08546_),
    .ZN(_03962_)
  );
  INV_X1 _24165_ (
    .A(_03962_),
    .ZN(_03963_)
  );
  AND2_X1 _24166_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03963_),
    .ZN(_03964_)
  );
  AND2_X1 _24167_ (
    .A1(_03961_),
    .A2(_03964_),
    .ZN(_03965_)
  );
  INV_X1 _24168_ (
    .A(_03965_),
    .ZN(_03966_)
  );
  AND2_X1 _24169_ (
    .A1(_03959_),
    .A2(_03966_),
    .ZN(_03967_)
  );
  MUX2_X1 _24170_ (
    .A(\rf[29] [19]),
    .B(\rf[25] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03968_)
  );
  AND2_X1 _24171_ (
    .A1(\rf[27] [19]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03969_)
  );
  MUX2_X1 _24172_ (
    .A(_03968_),
    .B(_03969_),
    .S(_08545_),
    .Z(_03970_)
  );
  MUX2_X1 _24173_ (
    .A(_03967_),
    .B(_03970_),
    .S(_08544_),
    .Z(_03971_)
  );
  AND2_X1 _24174_ (
    .A1(_08392_),
    .A2(_08546_),
    .ZN(_03972_)
  );
  INV_X1 _24175_ (
    .A(_03972_),
    .ZN(_03973_)
  );
  AND2_X1 _24176_ (
    .A1(_08293_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03974_)
  );
  INV_X1 _24177_ (
    .A(_03974_),
    .ZN(_03975_)
  );
  AND2_X1 _24178_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03975_),
    .ZN(_03976_)
  );
  AND2_X1 _24179_ (
    .A1(_03973_),
    .A2(_03976_),
    .ZN(_03977_)
  );
  INV_X1 _24180_ (
    .A(_03977_),
    .ZN(_03978_)
  );
  MUX2_X1 _24181_ (
    .A(\rf[22] [19]),
    .B(\rf[18] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03979_)
  );
  AND2_X1 _24182_ (
    .A1(_08545_),
    .A2(_03979_),
    .ZN(_03980_)
  );
  INV_X1 _24183_ (
    .A(_03980_),
    .ZN(_03981_)
  );
  AND2_X1 _24184_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03981_),
    .ZN(_03982_)
  );
  AND2_X1 _24185_ (
    .A1(_03978_),
    .A2(_03982_),
    .ZN(_03983_)
  );
  INV_X1 _24186_ (
    .A(_03983_),
    .ZN(_03984_)
  );
  AND2_X1 _24187_ (
    .A1(_08323_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03985_)
  );
  INV_X1 _24188_ (
    .A(_03985_),
    .ZN(_03986_)
  );
  AND2_X1 _24189_ (
    .A1(_08422_),
    .A2(_08546_),
    .ZN(_03987_)
  );
  INV_X1 _24190_ (
    .A(_03987_),
    .ZN(_03988_)
  );
  AND2_X1 _24191_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03988_),
    .ZN(_03989_)
  );
  AND2_X1 _24192_ (
    .A1(_03986_),
    .A2(_03989_),
    .ZN(_03990_)
  );
  INV_X1 _24193_ (
    .A(_03990_),
    .ZN(_03991_)
  );
  MUX2_X1 _24194_ (
    .A(\rf[23] [19]),
    .B(\rf[19] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03992_)
  );
  AND2_X1 _24195_ (
    .A1(_08545_),
    .A2(_03992_),
    .ZN(_03993_)
  );
  INV_X1 _24196_ (
    .A(_03993_),
    .ZN(_03994_)
  );
  AND2_X1 _24197_ (
    .A1(_08544_),
    .A2(_03994_),
    .ZN(_03995_)
  );
  AND2_X1 _24198_ (
    .A1(_03991_),
    .A2(_03995_),
    .ZN(_03996_)
  );
  INV_X1 _24199_ (
    .A(_03996_),
    .ZN(_03997_)
  );
  AND2_X1 _24200_ (
    .A1(_03984_),
    .A2(_03997_),
    .ZN(_03998_)
  );
  MUX2_X1 _24201_ (
    .A(_03971_),
    .B(_03998_),
    .S(ibuf_io_inst_0_bits_inst_rs2[3]),
    .Z(_03999_)
  );
  MUX2_X1 _24202_ (
    .A(_03952_),
    .B(_03999_),
    .S(_08572_),
    .Z(_04000_)
  );
  MUX2_X1 _24203_ (
    .A(_04000_),
    .B(_12099_),
    .S(_02233_),
    .Z(_04001_)
  );
  MUX2_X1 _24204_ (
    .A(ex_reg_rs_msb_1[17]),
    .B(_04001_),
    .S(_02202_),
    .Z(_00166_)
  );
  AND2_X1 _24205_ (
    .A1(_08343_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04002_)
  );
  INV_X1 _24206_ (
    .A(_04002_),
    .ZN(_04003_)
  );
  AND2_X1 _24207_ (
    .A1(_08481_),
    .A2(_08546_),
    .ZN(_04004_)
  );
  INV_X1 _24208_ (
    .A(_04004_),
    .ZN(_04005_)
  );
  AND2_X1 _24209_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04005_),
    .ZN(_04006_)
  );
  AND2_X1 _24210_ (
    .A1(_04003_),
    .A2(_04006_),
    .ZN(_04007_)
  );
  INV_X1 _24211_ (
    .A(_04007_),
    .ZN(_04008_)
  );
  MUX2_X1 _24212_ (
    .A(\rf[15] [20]),
    .B(\rf[11] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04009_)
  );
  AND2_X1 _24213_ (
    .A1(_08544_),
    .A2(_04009_),
    .ZN(_04010_)
  );
  INV_X1 _24214_ (
    .A(_04010_),
    .ZN(_04011_)
  );
  AND2_X1 _24215_ (
    .A1(_08545_),
    .A2(_04011_),
    .ZN(_04012_)
  );
  AND2_X1 _24216_ (
    .A1(_04008_),
    .A2(_04012_),
    .ZN(_04013_)
  );
  INV_X1 _24217_ (
    .A(_04013_),
    .ZN(_04014_)
  );
  AND2_X1 _24218_ (
    .A1(_08364_),
    .A2(_08546_),
    .ZN(_04015_)
  );
  INV_X1 _24219_ (
    .A(_04015_),
    .ZN(_04016_)
  );
  AND2_X1 _24220_ (
    .A1(_08265_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04017_)
  );
  INV_X1 _24221_ (
    .A(_04017_),
    .ZN(_04018_)
  );
  AND2_X1 _24222_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04018_),
    .ZN(_04019_)
  );
  AND2_X1 _24223_ (
    .A1(_04016_),
    .A2(_04019_),
    .ZN(_04020_)
  );
  INV_X1 _24224_ (
    .A(_04020_),
    .ZN(_04021_)
  );
  MUX2_X1 _24225_ (
    .A(\rf[13] [20]),
    .B(\rf[9] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04022_)
  );
  AND2_X1 _24226_ (
    .A1(_08544_),
    .A2(_04022_),
    .ZN(_04023_)
  );
  INV_X1 _24227_ (
    .A(_04023_),
    .ZN(_04024_)
  );
  AND2_X1 _24228_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04024_),
    .ZN(_04025_)
  );
  AND2_X1 _24229_ (
    .A1(_04021_),
    .A2(_04025_),
    .ZN(_04026_)
  );
  INV_X1 _24230_ (
    .A(_04026_),
    .ZN(_04027_)
  );
  AND2_X1 _24231_ (
    .A1(_08547_),
    .A2(_04027_),
    .ZN(_04028_)
  );
  AND2_X1 _24232_ (
    .A1(_04014_),
    .A2(_04028_),
    .ZN(_04029_)
  );
  INV_X1 _24233_ (
    .A(_04029_),
    .ZN(_04030_)
  );
  MUX2_X1 _24234_ (
    .A(\rf[6] [20]),
    .B(\rf[2] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04031_)
  );
  AND2_X1 _24235_ (
    .A1(_08545_),
    .A2(_04031_),
    .ZN(_04032_)
  );
  INV_X1 _24236_ (
    .A(_04032_),
    .ZN(_04033_)
  );
  MUX2_X1 _24237_ (
    .A(\rf[4] [20]),
    .B(\rf[0] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04034_)
  );
  AND2_X1 _24238_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04034_),
    .ZN(_04035_)
  );
  INV_X1 _24239_ (
    .A(_04035_),
    .ZN(_04036_)
  );
  AND2_X1 _24240_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04036_),
    .ZN(_04037_)
  );
  AND2_X1 _24241_ (
    .A1(_04033_),
    .A2(_04037_),
    .ZN(_04038_)
  );
  INV_X1 _24242_ (
    .A(_04038_),
    .ZN(_04039_)
  );
  MUX2_X1 _24243_ (
    .A(\rf[7] [20]),
    .B(\rf[3] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04040_)
  );
  AND2_X1 _24244_ (
    .A1(_08545_),
    .A2(_04040_),
    .ZN(_04041_)
  );
  INV_X1 _24245_ (
    .A(_04041_),
    .ZN(_04042_)
  );
  MUX2_X1 _24246_ (
    .A(\rf[5] [20]),
    .B(\rf[1] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04043_)
  );
  AND2_X1 _24247_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04043_),
    .ZN(_04044_)
  );
  INV_X1 _24248_ (
    .A(_04044_),
    .ZN(_04045_)
  );
  AND2_X1 _24249_ (
    .A1(_08544_),
    .A2(_04045_),
    .ZN(_04046_)
  );
  AND2_X1 _24250_ (
    .A1(_04042_),
    .A2(_04046_),
    .ZN(_04047_)
  );
  INV_X1 _24251_ (
    .A(_04047_),
    .ZN(_04048_)
  );
  AND2_X1 _24252_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_04048_),
    .ZN(_04049_)
  );
  AND2_X1 _24253_ (
    .A1(_04039_),
    .A2(_04049_),
    .ZN(_04050_)
  );
  INV_X1 _24254_ (
    .A(_04050_),
    .ZN(_04051_)
  );
  AND2_X1 _24255_ (
    .A1(_04030_),
    .A2(_04051_),
    .ZN(_04052_)
  );
  AND2_X1 _24256_ (
    .A1(_08324_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04053_)
  );
  INV_X1 _24257_ (
    .A(_04053_),
    .ZN(_04054_)
  );
  AND2_X1 _24258_ (
    .A1(_08423_),
    .A2(_08546_),
    .ZN(_04055_)
  );
  INV_X1 _24259_ (
    .A(_04055_),
    .ZN(_04056_)
  );
  AND2_X1 _24260_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04056_),
    .ZN(_04057_)
  );
  AND2_X1 _24261_ (
    .A1(_04054_),
    .A2(_04057_),
    .ZN(_04058_)
  );
  INV_X1 _24262_ (
    .A(_04058_),
    .ZN(_04059_)
  );
  MUX2_X1 _24263_ (
    .A(\rf[23] [20]),
    .B(\rf[19] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04060_)
  );
  AND2_X1 _24264_ (
    .A1(_08545_),
    .A2(_04060_),
    .ZN(_04061_)
  );
  INV_X1 _24265_ (
    .A(_04061_),
    .ZN(_04062_)
  );
  AND2_X1 _24266_ (
    .A1(_08544_),
    .A2(_04062_),
    .ZN(_04063_)
  );
  AND2_X1 _24267_ (
    .A1(_04059_),
    .A2(_04063_),
    .ZN(_04064_)
  );
  INV_X1 _24268_ (
    .A(_04064_),
    .ZN(_04065_)
  );
  AND2_X1 _24269_ (
    .A1(_08393_),
    .A2(_08546_),
    .ZN(_04066_)
  );
  INV_X1 _24270_ (
    .A(_04066_),
    .ZN(_04067_)
  );
  AND2_X1 _24271_ (
    .A1(_08294_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04068_)
  );
  INV_X1 _24272_ (
    .A(_04068_),
    .ZN(_04069_)
  );
  AND2_X1 _24273_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04069_),
    .ZN(_04070_)
  );
  AND2_X1 _24274_ (
    .A1(_04067_),
    .A2(_04070_),
    .ZN(_04071_)
  );
  INV_X1 _24275_ (
    .A(_04071_),
    .ZN(_04072_)
  );
  MUX2_X1 _24276_ (
    .A(\rf[22] [20]),
    .B(\rf[18] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04073_)
  );
  AND2_X1 _24277_ (
    .A1(_08545_),
    .A2(_04073_),
    .ZN(_04074_)
  );
  INV_X1 _24278_ (
    .A(_04074_),
    .ZN(_04075_)
  );
  AND2_X1 _24279_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04075_),
    .ZN(_04076_)
  );
  AND2_X1 _24280_ (
    .A1(_04072_),
    .A2(_04076_),
    .ZN(_04077_)
  );
  INV_X1 _24281_ (
    .A(_04077_),
    .ZN(_04078_)
  );
  AND2_X1 _24282_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_04065_),
    .ZN(_04079_)
  );
  AND2_X1 _24283_ (
    .A1(_04078_),
    .A2(_04079_),
    .ZN(_04080_)
  );
  INV_X1 _24284_ (
    .A(_04080_),
    .ZN(_04081_)
  );
  AND2_X1 _24285_ (
    .A1(_08449_),
    .A2(_08546_),
    .ZN(_04082_)
  );
  INV_X1 _24286_ (
    .A(_04082_),
    .ZN(_04083_)
  );
  AND2_X1 _24287_ (
    .A1(_08519_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04084_)
  );
  INV_X1 _24288_ (
    .A(_04084_),
    .ZN(_04085_)
  );
  AND2_X1 _24289_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04085_),
    .ZN(_04086_)
  );
  AND2_X1 _24290_ (
    .A1(_04083_),
    .A2(_04086_),
    .ZN(_04087_)
  );
  INV_X1 _24291_ (
    .A(_04087_),
    .ZN(_04088_)
  );
  MUX2_X1 _24292_ (
    .A(\rf[30] [20]),
    .B(\rf[26] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04089_)
  );
  AND2_X1 _24293_ (
    .A1(_08545_),
    .A2(_04089_),
    .ZN(_04090_)
  );
  INV_X1 _24294_ (
    .A(_04090_),
    .ZN(_04091_)
  );
  AND2_X1 _24295_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04091_),
    .ZN(_04092_)
  );
  AND2_X1 _24296_ (
    .A1(_04088_),
    .A2(_04092_),
    .ZN(_04093_)
  );
  INV_X1 _24297_ (
    .A(_04093_),
    .ZN(_04094_)
  );
  MUX2_X1 _24298_ (
    .A(\rf[29] [20]),
    .B(\rf[25] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04095_)
  );
  AND2_X1 _24299_ (
    .A1(\rf[27] [20]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04096_)
  );
  MUX2_X1 _24300_ (
    .A(_04095_),
    .B(_04096_),
    .S(_08545_),
    .Z(_04097_)
  );
  INV_X1 _24301_ (
    .A(_04097_),
    .ZN(_04098_)
  );
  AND2_X1 _24302_ (
    .A1(_08544_),
    .A2(_04098_),
    .ZN(_04099_)
  );
  INV_X1 _24303_ (
    .A(_04099_),
    .ZN(_04100_)
  );
  AND2_X1 _24304_ (
    .A1(_08547_),
    .A2(_04100_),
    .ZN(_04101_)
  );
  AND2_X1 _24305_ (
    .A1(_04094_),
    .A2(_04101_),
    .ZN(_04102_)
  );
  INV_X1 _24306_ (
    .A(_04102_),
    .ZN(_04103_)
  );
  AND2_X1 _24307_ (
    .A1(_04081_),
    .A2(_04103_),
    .ZN(_04104_)
  );
  MUX2_X1 _24308_ (
    .A(_04052_),
    .B(_04104_),
    .S(_08572_),
    .Z(_04105_)
  );
  INV_X1 _24309_ (
    .A(_04105_),
    .ZN(_04106_)
  );
  MUX2_X1 _24310_ (
    .A(_04106_),
    .B(_12305_),
    .S(_02233_),
    .Z(_04107_)
  );
  MUX2_X1 _24311_ (
    .A(ex_reg_rs_msb_1[18]),
    .B(_04107_),
    .S(_02202_),
    .Z(_00167_)
  );
  AND2_X1 _24312_ (
    .A1(_08344_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04108_)
  );
  INV_X1 _24313_ (
    .A(_04108_),
    .ZN(_04109_)
  );
  AND2_X1 _24314_ (
    .A1(_08482_),
    .A2(_08546_),
    .ZN(_04110_)
  );
  INV_X1 _24315_ (
    .A(_04110_),
    .ZN(_04111_)
  );
  AND2_X1 _24316_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04111_),
    .ZN(_04112_)
  );
  AND2_X1 _24317_ (
    .A1(_04109_),
    .A2(_04112_),
    .ZN(_04113_)
  );
  INV_X1 _24318_ (
    .A(_04113_),
    .ZN(_04114_)
  );
  MUX2_X1 _24319_ (
    .A(\rf[15] [21]),
    .B(\rf[11] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04115_)
  );
  AND2_X1 _24320_ (
    .A1(_08544_),
    .A2(_04115_),
    .ZN(_04116_)
  );
  INV_X1 _24321_ (
    .A(_04116_),
    .ZN(_04117_)
  );
  AND2_X1 _24322_ (
    .A1(_08545_),
    .A2(_04117_),
    .ZN(_04118_)
  );
  AND2_X1 _24323_ (
    .A1(_04114_),
    .A2(_04118_),
    .ZN(_04119_)
  );
  INV_X1 _24324_ (
    .A(_04119_),
    .ZN(_04120_)
  );
  AND2_X1 _24325_ (
    .A1(_08365_),
    .A2(_08546_),
    .ZN(_04121_)
  );
  INV_X1 _24326_ (
    .A(_04121_),
    .ZN(_04122_)
  );
  AND2_X1 _24327_ (
    .A1(_08266_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04123_)
  );
  INV_X1 _24328_ (
    .A(_04123_),
    .ZN(_04124_)
  );
  AND2_X1 _24329_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04124_),
    .ZN(_04125_)
  );
  AND2_X1 _24330_ (
    .A1(_04122_),
    .A2(_04125_),
    .ZN(_04126_)
  );
  INV_X1 _24331_ (
    .A(_04126_),
    .ZN(_04127_)
  );
  MUX2_X1 _24332_ (
    .A(\rf[13] [21]),
    .B(\rf[9] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04128_)
  );
  AND2_X1 _24333_ (
    .A1(_08544_),
    .A2(_04128_),
    .ZN(_04129_)
  );
  INV_X1 _24334_ (
    .A(_04129_),
    .ZN(_04130_)
  );
  AND2_X1 _24335_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04130_),
    .ZN(_04131_)
  );
  AND2_X1 _24336_ (
    .A1(_04127_),
    .A2(_04131_),
    .ZN(_04132_)
  );
  INV_X1 _24337_ (
    .A(_04132_),
    .ZN(_04133_)
  );
  AND2_X1 _24338_ (
    .A1(_08547_),
    .A2(_04133_),
    .ZN(_04134_)
  );
  AND2_X1 _24339_ (
    .A1(_04120_),
    .A2(_04134_),
    .ZN(_04135_)
  );
  INV_X1 _24340_ (
    .A(_04135_),
    .ZN(_04136_)
  );
  MUX2_X1 _24341_ (
    .A(\rf[6] [21]),
    .B(\rf[2] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04137_)
  );
  AND2_X1 _24342_ (
    .A1(_08545_),
    .A2(_04137_),
    .ZN(_04138_)
  );
  INV_X1 _24343_ (
    .A(_04138_),
    .ZN(_04139_)
  );
  MUX2_X1 _24344_ (
    .A(\rf[4] [21]),
    .B(\rf[0] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04140_)
  );
  AND2_X1 _24345_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04140_),
    .ZN(_04141_)
  );
  INV_X1 _24346_ (
    .A(_04141_),
    .ZN(_04142_)
  );
  AND2_X1 _24347_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04142_),
    .ZN(_04143_)
  );
  AND2_X1 _24348_ (
    .A1(_04139_),
    .A2(_04143_),
    .ZN(_04144_)
  );
  INV_X1 _24349_ (
    .A(_04144_),
    .ZN(_04145_)
  );
  MUX2_X1 _24350_ (
    .A(\rf[7] [21]),
    .B(\rf[3] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04146_)
  );
  AND2_X1 _24351_ (
    .A1(_08545_),
    .A2(_04146_),
    .ZN(_04147_)
  );
  INV_X1 _24352_ (
    .A(_04147_),
    .ZN(_04148_)
  );
  MUX2_X1 _24353_ (
    .A(\rf[5] [21]),
    .B(\rf[1] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04149_)
  );
  AND2_X1 _24354_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04149_),
    .ZN(_04150_)
  );
  INV_X1 _24355_ (
    .A(_04150_),
    .ZN(_04151_)
  );
  AND2_X1 _24356_ (
    .A1(_08544_),
    .A2(_04151_),
    .ZN(_04152_)
  );
  AND2_X1 _24357_ (
    .A1(_04148_),
    .A2(_04152_),
    .ZN(_04153_)
  );
  INV_X1 _24358_ (
    .A(_04153_),
    .ZN(_04154_)
  );
  AND2_X1 _24359_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_04154_),
    .ZN(_04155_)
  );
  AND2_X1 _24360_ (
    .A1(_04145_),
    .A2(_04155_),
    .ZN(_04156_)
  );
  INV_X1 _24361_ (
    .A(_04156_),
    .ZN(_04157_)
  );
  AND2_X1 _24362_ (
    .A1(_04136_),
    .A2(_04157_),
    .ZN(_04158_)
  );
  AND2_X1 _24363_ (
    .A1(_08325_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04159_)
  );
  INV_X1 _24364_ (
    .A(_04159_),
    .ZN(_04160_)
  );
  AND2_X1 _24365_ (
    .A1(_08424_),
    .A2(_08546_),
    .ZN(_04161_)
  );
  INV_X1 _24366_ (
    .A(_04161_),
    .ZN(_04162_)
  );
  AND2_X1 _24367_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04162_),
    .ZN(_04163_)
  );
  AND2_X1 _24368_ (
    .A1(_04160_),
    .A2(_04163_),
    .ZN(_04164_)
  );
  INV_X1 _24369_ (
    .A(_04164_),
    .ZN(_04165_)
  );
  MUX2_X1 _24370_ (
    .A(\rf[23] [21]),
    .B(\rf[19] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04166_)
  );
  AND2_X1 _24371_ (
    .A1(_08545_),
    .A2(_04166_),
    .ZN(_04167_)
  );
  INV_X1 _24372_ (
    .A(_04167_),
    .ZN(_04168_)
  );
  AND2_X1 _24373_ (
    .A1(_08544_),
    .A2(_04168_),
    .ZN(_04169_)
  );
  AND2_X1 _24374_ (
    .A1(_04165_),
    .A2(_04169_),
    .ZN(_04170_)
  );
  INV_X1 _24375_ (
    .A(_04170_),
    .ZN(_04171_)
  );
  AND2_X1 _24376_ (
    .A1(_08394_),
    .A2(_08546_),
    .ZN(_04172_)
  );
  INV_X1 _24377_ (
    .A(_04172_),
    .ZN(_04173_)
  );
  AND2_X1 _24378_ (
    .A1(_08295_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04174_)
  );
  INV_X1 _24379_ (
    .A(_04174_),
    .ZN(_04175_)
  );
  AND2_X1 _24380_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04175_),
    .ZN(_04176_)
  );
  AND2_X1 _24381_ (
    .A1(_04173_),
    .A2(_04176_),
    .ZN(_04177_)
  );
  INV_X1 _24382_ (
    .A(_04177_),
    .ZN(_04178_)
  );
  MUX2_X1 _24383_ (
    .A(\rf[22] [21]),
    .B(\rf[18] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04179_)
  );
  AND2_X1 _24384_ (
    .A1(_08545_),
    .A2(_04179_),
    .ZN(_04180_)
  );
  INV_X1 _24385_ (
    .A(_04180_),
    .ZN(_04181_)
  );
  AND2_X1 _24386_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04181_),
    .ZN(_04182_)
  );
  AND2_X1 _24387_ (
    .A1(_04178_),
    .A2(_04182_),
    .ZN(_04183_)
  );
  INV_X1 _24388_ (
    .A(_04183_),
    .ZN(_04184_)
  );
  AND2_X1 _24389_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_04171_),
    .ZN(_04185_)
  );
  AND2_X1 _24390_ (
    .A1(_04184_),
    .A2(_04185_),
    .ZN(_04186_)
  );
  INV_X1 _24391_ (
    .A(_04186_),
    .ZN(_04187_)
  );
  AND2_X1 _24392_ (
    .A1(_08450_),
    .A2(_08546_),
    .ZN(_04188_)
  );
  INV_X1 _24393_ (
    .A(_04188_),
    .ZN(_04189_)
  );
  AND2_X1 _24394_ (
    .A1(_08520_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04190_)
  );
  INV_X1 _24395_ (
    .A(_04190_),
    .ZN(_04191_)
  );
  AND2_X1 _24396_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04191_),
    .ZN(_04192_)
  );
  AND2_X1 _24397_ (
    .A1(_04189_),
    .A2(_04192_),
    .ZN(_04193_)
  );
  INV_X1 _24398_ (
    .A(_04193_),
    .ZN(_04194_)
  );
  MUX2_X1 _24399_ (
    .A(\rf[30] [21]),
    .B(\rf[26] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04195_)
  );
  AND2_X1 _24400_ (
    .A1(_08545_),
    .A2(_04195_),
    .ZN(_04196_)
  );
  INV_X1 _24401_ (
    .A(_04196_),
    .ZN(_04197_)
  );
  AND2_X1 _24402_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04197_),
    .ZN(_04198_)
  );
  AND2_X1 _24403_ (
    .A1(_04194_),
    .A2(_04198_),
    .ZN(_04199_)
  );
  INV_X1 _24404_ (
    .A(_04199_),
    .ZN(_04200_)
  );
  MUX2_X1 _24405_ (
    .A(\rf[29] [21]),
    .B(\rf[25] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04201_)
  );
  AND2_X1 _24406_ (
    .A1(\rf[27] [21]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04202_)
  );
  MUX2_X1 _24407_ (
    .A(_04201_),
    .B(_04202_),
    .S(_08545_),
    .Z(_04203_)
  );
  INV_X1 _24408_ (
    .A(_04203_),
    .ZN(_04204_)
  );
  AND2_X1 _24409_ (
    .A1(_08544_),
    .A2(_04204_),
    .ZN(_04205_)
  );
  INV_X1 _24410_ (
    .A(_04205_),
    .ZN(_04206_)
  );
  AND2_X1 _24411_ (
    .A1(_08547_),
    .A2(_04206_),
    .ZN(_04207_)
  );
  AND2_X1 _24412_ (
    .A1(_04200_),
    .A2(_04207_),
    .ZN(_04208_)
  );
  INV_X1 _24413_ (
    .A(_04208_),
    .ZN(_04209_)
  );
  AND2_X1 _24414_ (
    .A1(_04187_),
    .A2(_04209_),
    .ZN(_04210_)
  );
  MUX2_X1 _24415_ (
    .A(_04158_),
    .B(_04210_),
    .S(_08572_),
    .Z(_04211_)
  );
  INV_X1 _24416_ (
    .A(_04211_),
    .ZN(_04212_)
  );
  MUX2_X1 _24417_ (
    .A(_04212_),
    .B(_12316_),
    .S(_02233_),
    .Z(_04213_)
  );
  MUX2_X1 _24418_ (
    .A(ex_reg_rs_msb_1[19]),
    .B(_04213_),
    .S(_02202_),
    .Z(_00168_)
  );
  AND2_X1 _24419_ (
    .A1(_08345_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04214_)
  );
  INV_X1 _24420_ (
    .A(_04214_),
    .ZN(_04215_)
  );
  AND2_X1 _24421_ (
    .A1(_08483_),
    .A2(_08546_),
    .ZN(_04216_)
  );
  INV_X1 _24422_ (
    .A(_04216_),
    .ZN(_04217_)
  );
  AND2_X1 _24423_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04217_),
    .ZN(_04218_)
  );
  AND2_X1 _24424_ (
    .A1(_04215_),
    .A2(_04218_),
    .ZN(_04219_)
  );
  INV_X1 _24425_ (
    .A(_04219_),
    .ZN(_04220_)
  );
  MUX2_X1 _24426_ (
    .A(\rf[15] [22]),
    .B(\rf[11] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04221_)
  );
  AND2_X1 _24427_ (
    .A1(_08544_),
    .A2(_04221_),
    .ZN(_04222_)
  );
  INV_X1 _24428_ (
    .A(_04222_),
    .ZN(_04223_)
  );
  AND2_X1 _24429_ (
    .A1(_08545_),
    .A2(_04223_),
    .ZN(_04224_)
  );
  AND2_X1 _24430_ (
    .A1(_04220_),
    .A2(_04224_),
    .ZN(_04225_)
  );
  INV_X1 _24431_ (
    .A(_04225_),
    .ZN(_04226_)
  );
  AND2_X1 _24432_ (
    .A1(_08366_),
    .A2(_08546_),
    .ZN(_04227_)
  );
  INV_X1 _24433_ (
    .A(_04227_),
    .ZN(_04228_)
  );
  AND2_X1 _24434_ (
    .A1(_08267_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04229_)
  );
  INV_X1 _24435_ (
    .A(_04229_),
    .ZN(_04230_)
  );
  AND2_X1 _24436_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04230_),
    .ZN(_04231_)
  );
  AND2_X1 _24437_ (
    .A1(_04228_),
    .A2(_04231_),
    .ZN(_04232_)
  );
  INV_X1 _24438_ (
    .A(_04232_),
    .ZN(_04233_)
  );
  MUX2_X1 _24439_ (
    .A(\rf[13] [22]),
    .B(\rf[9] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04234_)
  );
  AND2_X1 _24440_ (
    .A1(_08544_),
    .A2(_04234_),
    .ZN(_04235_)
  );
  INV_X1 _24441_ (
    .A(_04235_),
    .ZN(_04236_)
  );
  AND2_X1 _24442_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04236_),
    .ZN(_04237_)
  );
  AND2_X1 _24443_ (
    .A1(_04233_),
    .A2(_04237_),
    .ZN(_04238_)
  );
  INV_X1 _24444_ (
    .A(_04238_),
    .ZN(_04239_)
  );
  AND2_X1 _24445_ (
    .A1(_08547_),
    .A2(_04239_),
    .ZN(_04240_)
  );
  AND2_X1 _24446_ (
    .A1(_04226_),
    .A2(_04240_),
    .ZN(_04241_)
  );
  INV_X1 _24447_ (
    .A(_04241_),
    .ZN(_04242_)
  );
  MUX2_X1 _24448_ (
    .A(\rf[6] [22]),
    .B(\rf[2] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04243_)
  );
  AND2_X1 _24449_ (
    .A1(_08545_),
    .A2(_04243_),
    .ZN(_04244_)
  );
  INV_X1 _24450_ (
    .A(_04244_),
    .ZN(_04245_)
  );
  MUX2_X1 _24451_ (
    .A(\rf[4] [22]),
    .B(\rf[0] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04246_)
  );
  AND2_X1 _24452_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04246_),
    .ZN(_04247_)
  );
  INV_X1 _24453_ (
    .A(_04247_),
    .ZN(_04248_)
  );
  AND2_X1 _24454_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04248_),
    .ZN(_04249_)
  );
  AND2_X1 _24455_ (
    .A1(_04245_),
    .A2(_04249_),
    .ZN(_04250_)
  );
  INV_X1 _24456_ (
    .A(_04250_),
    .ZN(_04251_)
  );
  MUX2_X1 _24457_ (
    .A(\rf[7] [22]),
    .B(\rf[3] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04252_)
  );
  AND2_X1 _24458_ (
    .A1(_08545_),
    .A2(_04252_),
    .ZN(_04253_)
  );
  INV_X1 _24459_ (
    .A(_04253_),
    .ZN(_04254_)
  );
  MUX2_X1 _24460_ (
    .A(\rf[5] [22]),
    .B(\rf[1] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04255_)
  );
  AND2_X1 _24461_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04255_),
    .ZN(_04256_)
  );
  INV_X1 _24462_ (
    .A(_04256_),
    .ZN(_04257_)
  );
  AND2_X1 _24463_ (
    .A1(_08544_),
    .A2(_04257_),
    .ZN(_04258_)
  );
  AND2_X1 _24464_ (
    .A1(_04254_),
    .A2(_04258_),
    .ZN(_04259_)
  );
  INV_X1 _24465_ (
    .A(_04259_),
    .ZN(_04260_)
  );
  AND2_X1 _24466_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_04260_),
    .ZN(_04261_)
  );
  AND2_X1 _24467_ (
    .A1(_04251_),
    .A2(_04261_),
    .ZN(_04262_)
  );
  INV_X1 _24468_ (
    .A(_04262_),
    .ZN(_04263_)
  );
  AND2_X1 _24469_ (
    .A1(_04242_),
    .A2(_04263_),
    .ZN(_04264_)
  );
  AND2_X1 _24470_ (
    .A1(_08326_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04265_)
  );
  INV_X1 _24471_ (
    .A(_04265_),
    .ZN(_04266_)
  );
  AND2_X1 _24472_ (
    .A1(_08425_),
    .A2(_08546_),
    .ZN(_04267_)
  );
  INV_X1 _24473_ (
    .A(_04267_),
    .ZN(_04268_)
  );
  AND2_X1 _24474_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04268_),
    .ZN(_04269_)
  );
  AND2_X1 _24475_ (
    .A1(_04266_),
    .A2(_04269_),
    .ZN(_04270_)
  );
  INV_X1 _24476_ (
    .A(_04270_),
    .ZN(_04271_)
  );
  MUX2_X1 _24477_ (
    .A(\rf[23] [22]),
    .B(\rf[19] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04272_)
  );
  AND2_X1 _24478_ (
    .A1(_08545_),
    .A2(_04272_),
    .ZN(_04273_)
  );
  INV_X1 _24479_ (
    .A(_04273_),
    .ZN(_04274_)
  );
  AND2_X1 _24480_ (
    .A1(_08544_),
    .A2(_04274_),
    .ZN(_04275_)
  );
  AND2_X1 _24481_ (
    .A1(_04271_),
    .A2(_04275_),
    .ZN(_04276_)
  );
  INV_X1 _24482_ (
    .A(_04276_),
    .ZN(_04277_)
  );
  AND2_X1 _24483_ (
    .A1(_08395_),
    .A2(_08546_),
    .ZN(_04278_)
  );
  INV_X1 _24484_ (
    .A(_04278_),
    .ZN(_04279_)
  );
  AND2_X1 _24485_ (
    .A1(_08296_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04280_)
  );
  INV_X1 _24486_ (
    .A(_04280_),
    .ZN(_04281_)
  );
  AND2_X1 _24487_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04281_),
    .ZN(_04282_)
  );
  AND2_X1 _24488_ (
    .A1(_04279_),
    .A2(_04282_),
    .ZN(_04283_)
  );
  INV_X1 _24489_ (
    .A(_04283_),
    .ZN(_04284_)
  );
  MUX2_X1 _24490_ (
    .A(\rf[22] [22]),
    .B(\rf[18] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04285_)
  );
  AND2_X1 _24491_ (
    .A1(_08545_),
    .A2(_04285_),
    .ZN(_04286_)
  );
  INV_X1 _24492_ (
    .A(_04286_),
    .ZN(_04287_)
  );
  AND2_X1 _24493_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04287_),
    .ZN(_04288_)
  );
  AND2_X1 _24494_ (
    .A1(_04284_),
    .A2(_04288_),
    .ZN(_04289_)
  );
  INV_X1 _24495_ (
    .A(_04289_),
    .ZN(_04290_)
  );
  AND2_X1 _24496_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_04277_),
    .ZN(_04291_)
  );
  AND2_X1 _24497_ (
    .A1(_04290_),
    .A2(_04291_),
    .ZN(_04292_)
  );
  INV_X1 _24498_ (
    .A(_04292_),
    .ZN(_04293_)
  );
  AND2_X1 _24499_ (
    .A1(_08451_),
    .A2(_08546_),
    .ZN(_04294_)
  );
  INV_X1 _24500_ (
    .A(_04294_),
    .ZN(_04295_)
  );
  AND2_X1 _24501_ (
    .A1(_08521_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04296_)
  );
  INV_X1 _24502_ (
    .A(_04296_),
    .ZN(_04297_)
  );
  AND2_X1 _24503_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04297_),
    .ZN(_04298_)
  );
  AND2_X1 _24504_ (
    .A1(_04295_),
    .A2(_04298_),
    .ZN(_04299_)
  );
  INV_X1 _24505_ (
    .A(_04299_),
    .ZN(_04300_)
  );
  MUX2_X1 _24506_ (
    .A(\rf[30] [22]),
    .B(\rf[26] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04301_)
  );
  AND2_X1 _24507_ (
    .A1(_08545_),
    .A2(_04301_),
    .ZN(_04302_)
  );
  INV_X1 _24508_ (
    .A(_04302_),
    .ZN(_04303_)
  );
  AND2_X1 _24509_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04303_),
    .ZN(_04304_)
  );
  AND2_X1 _24510_ (
    .A1(_04300_),
    .A2(_04304_),
    .ZN(_04305_)
  );
  INV_X1 _24511_ (
    .A(_04305_),
    .ZN(_04306_)
  );
  MUX2_X1 _24512_ (
    .A(\rf[29] [22]),
    .B(\rf[25] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04307_)
  );
  AND2_X1 _24513_ (
    .A1(\rf[27] [22]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04308_)
  );
  MUX2_X1 _24514_ (
    .A(_04307_),
    .B(_04308_),
    .S(_08545_),
    .Z(_04309_)
  );
  INV_X1 _24515_ (
    .A(_04309_),
    .ZN(_04310_)
  );
  AND2_X1 _24516_ (
    .A1(_08544_),
    .A2(_04310_),
    .ZN(_04311_)
  );
  INV_X1 _24517_ (
    .A(_04311_),
    .ZN(_04312_)
  );
  AND2_X1 _24518_ (
    .A1(_08547_),
    .A2(_04312_),
    .ZN(_04313_)
  );
  AND2_X1 _24519_ (
    .A1(_04306_),
    .A2(_04313_),
    .ZN(_04314_)
  );
  INV_X1 _24520_ (
    .A(_04314_),
    .ZN(_04315_)
  );
  AND2_X1 _24521_ (
    .A1(_04293_),
    .A2(_04315_),
    .ZN(_04316_)
  );
  MUX2_X1 _24522_ (
    .A(_04264_),
    .B(_04316_),
    .S(_08572_),
    .Z(_04317_)
  );
  INV_X1 _24523_ (
    .A(_04317_),
    .ZN(_04318_)
  );
  MUX2_X1 _24524_ (
    .A(_04318_),
    .B(_12537_),
    .S(_02233_),
    .Z(_04319_)
  );
  MUX2_X1 _24525_ (
    .A(ex_reg_rs_msb_1[20]),
    .B(_04319_),
    .S(_02202_),
    .Z(_00169_)
  );
  MUX2_X1 _24526_ (
    .A(\rf[3] [23]),
    .B(\rf[2] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_04320_)
  );
  MUX2_X1 _24527_ (
    .A(\rf[7] [23]),
    .B(\rf[6] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_04321_)
  );
  MUX2_X1 _24528_ (
    .A(_04320_),
    .B(_04321_),
    .S(_08546_),
    .Z(_04322_)
  );
  INV_X1 _24529_ (
    .A(_04322_),
    .ZN(_04323_)
  );
  AND2_X1 _24530_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_04323_),
    .ZN(_04324_)
  );
  INV_X1 _24531_ (
    .A(_04324_),
    .ZN(_04325_)
  );
  MUX2_X1 _24532_ (
    .A(\rf[14] [23]),
    .B(\rf[10] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04326_)
  );
  INV_X1 _24533_ (
    .A(_04326_),
    .ZN(_04327_)
  );
  AND2_X1 _24534_ (
    .A1(_02341_),
    .A2(_04327_),
    .ZN(_04328_)
  );
  INV_X1 _24535_ (
    .A(_04328_),
    .ZN(_04329_)
  );
  MUX2_X1 _24536_ (
    .A(\rf[15] [23]),
    .B(\rf[11] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04330_)
  );
  INV_X1 _24537_ (
    .A(_04330_),
    .ZN(_04331_)
  );
  AND2_X1 _24538_ (
    .A1(_09692_),
    .A2(_04331_),
    .ZN(_04332_)
  );
  INV_X1 _24539_ (
    .A(_04332_),
    .ZN(_04333_)
  );
  AND2_X1 _24540_ (
    .A1(_04329_),
    .A2(_04333_),
    .ZN(_04334_)
  );
  AND2_X1 _24541_ (
    .A1(_04325_),
    .A2(_04334_),
    .ZN(_04335_)
  );
  MUX2_X1 _24542_ (
    .A(\rf[1] [23]),
    .B(\rf[0] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_04336_)
  );
  MUX2_X1 _24543_ (
    .A(\rf[5] [23]),
    .B(\rf[4] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_04337_)
  );
  MUX2_X1 _24544_ (
    .A(_04336_),
    .B(_04337_),
    .S(_08546_),
    .Z(_04338_)
  );
  INV_X1 _24545_ (
    .A(_04338_),
    .ZN(_04339_)
  );
  AND2_X1 _24546_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_04339_),
    .ZN(_04340_)
  );
  INV_X1 _24547_ (
    .A(_04340_),
    .ZN(_04341_)
  );
  MUX2_X1 _24548_ (
    .A(\rf[12] [23]),
    .B(\rf[8] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04342_)
  );
  INV_X1 _24549_ (
    .A(_04342_),
    .ZN(_04343_)
  );
  AND2_X1 _24550_ (
    .A1(_02341_),
    .A2(_04343_),
    .ZN(_04344_)
  );
  INV_X1 _24551_ (
    .A(_04344_),
    .ZN(_04345_)
  );
  MUX2_X1 _24552_ (
    .A(\rf[13] [23]),
    .B(\rf[9] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04346_)
  );
  INV_X1 _24553_ (
    .A(_04346_),
    .ZN(_04347_)
  );
  AND2_X1 _24554_ (
    .A1(_09692_),
    .A2(_04347_),
    .ZN(_04348_)
  );
  INV_X1 _24555_ (
    .A(_04348_),
    .ZN(_04349_)
  );
  AND2_X1 _24556_ (
    .A1(_04345_),
    .A2(_04349_),
    .ZN(_04350_)
  );
  AND2_X1 _24557_ (
    .A1(_04341_),
    .A2(_04350_),
    .ZN(_04351_)
  );
  AND2_X1 _24558_ (
    .A1(\rf[30] [23]),
    .A2(_08546_),
    .ZN(_04352_)
  );
  INV_X1 _24559_ (
    .A(_04352_),
    .ZN(_04353_)
  );
  AND2_X1 _24560_ (
    .A1(\rf[26] [23]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04354_)
  );
  INV_X1 _24561_ (
    .A(_04354_),
    .ZN(_04355_)
  );
  AND2_X1 _24562_ (
    .A1(_08545_),
    .A2(_04355_),
    .ZN(_04356_)
  );
  AND2_X1 _24563_ (
    .A1(_04353_),
    .A2(_04356_),
    .ZN(_04357_)
  );
  INV_X1 _24564_ (
    .A(_04357_),
    .ZN(_04358_)
  );
  AND2_X1 _24565_ (
    .A1(\rf[24] [23]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04359_)
  );
  INV_X1 _24566_ (
    .A(_04359_),
    .ZN(_04360_)
  );
  AND2_X1 _24567_ (
    .A1(\rf[28] [23]),
    .A2(_08546_),
    .ZN(_04361_)
  );
  INV_X1 _24568_ (
    .A(_04361_),
    .ZN(_04362_)
  );
  AND2_X1 _24569_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04362_),
    .ZN(_04363_)
  );
  AND2_X1 _24570_ (
    .A1(_04360_),
    .A2(_04363_),
    .ZN(_04364_)
  );
  INV_X1 _24571_ (
    .A(_04364_),
    .ZN(_04365_)
  );
  AND2_X1 _24572_ (
    .A1(_04358_),
    .A2(_04365_),
    .ZN(_04366_)
  );
  MUX2_X1 _24573_ (
    .A(\rf[29] [23]),
    .B(\rf[25] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04367_)
  );
  AND2_X1 _24574_ (
    .A1(\rf[27] [23]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04368_)
  );
  MUX2_X1 _24575_ (
    .A(_04367_),
    .B(_04368_),
    .S(_08545_),
    .Z(_04369_)
  );
  MUX2_X1 _24576_ (
    .A(_04366_),
    .B(_04369_),
    .S(_08544_),
    .Z(_04370_)
  );
  AND2_X1 _24577_ (
    .A1(_08396_),
    .A2(_08546_),
    .ZN(_04371_)
  );
  INV_X1 _24578_ (
    .A(_04371_),
    .ZN(_04372_)
  );
  AND2_X1 _24579_ (
    .A1(_08297_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04373_)
  );
  INV_X1 _24580_ (
    .A(_04373_),
    .ZN(_04374_)
  );
  AND2_X1 _24581_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04374_),
    .ZN(_04375_)
  );
  AND2_X1 _24582_ (
    .A1(_04372_),
    .A2(_04375_),
    .ZN(_04376_)
  );
  INV_X1 _24583_ (
    .A(_04376_),
    .ZN(_04377_)
  );
  MUX2_X1 _24584_ (
    .A(\rf[22] [23]),
    .B(\rf[18] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04378_)
  );
  AND2_X1 _24585_ (
    .A1(_08545_),
    .A2(_04378_),
    .ZN(_04379_)
  );
  INV_X1 _24586_ (
    .A(_04379_),
    .ZN(_04380_)
  );
  AND2_X1 _24587_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04380_),
    .ZN(_04381_)
  );
  AND2_X1 _24588_ (
    .A1(_04377_),
    .A2(_04381_),
    .ZN(_04382_)
  );
  INV_X1 _24589_ (
    .A(_04382_),
    .ZN(_04383_)
  );
  AND2_X1 _24590_ (
    .A1(_08327_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04384_)
  );
  INV_X1 _24591_ (
    .A(_04384_),
    .ZN(_04385_)
  );
  AND2_X1 _24592_ (
    .A1(_08426_),
    .A2(_08546_),
    .ZN(_04386_)
  );
  INV_X1 _24593_ (
    .A(_04386_),
    .ZN(_04387_)
  );
  AND2_X1 _24594_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04387_),
    .ZN(_04388_)
  );
  AND2_X1 _24595_ (
    .A1(_04385_),
    .A2(_04388_),
    .ZN(_04389_)
  );
  INV_X1 _24596_ (
    .A(_04389_),
    .ZN(_04390_)
  );
  MUX2_X1 _24597_ (
    .A(\rf[23] [23]),
    .B(\rf[19] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04391_)
  );
  AND2_X1 _24598_ (
    .A1(_08545_),
    .A2(_04391_),
    .ZN(_04392_)
  );
  INV_X1 _24599_ (
    .A(_04392_),
    .ZN(_04393_)
  );
  AND2_X1 _24600_ (
    .A1(_08544_),
    .A2(_04393_),
    .ZN(_04394_)
  );
  AND2_X1 _24601_ (
    .A1(_04390_),
    .A2(_04394_),
    .ZN(_04395_)
  );
  INV_X1 _24602_ (
    .A(_04395_),
    .ZN(_04396_)
  );
  AND2_X1 _24603_ (
    .A1(_04383_),
    .A2(_04396_),
    .ZN(_04397_)
  );
  MUX2_X1 _24604_ (
    .A(_04370_),
    .B(_04397_),
    .S(ibuf_io_inst_0_bits_inst_rs2[3]),
    .Z(_04398_)
  );
  MUX2_X1 _24605_ (
    .A(_04335_),
    .B(_04351_),
    .S(ibuf_io_inst_0_bits_inst_rs2[1]),
    .Z(_04399_)
  );
  MUX2_X1 _24606_ (
    .A(_04398_),
    .B(_04399_),
    .S(ibuf_io_inst_0_bits_inst_rs2[4]),
    .Z(_04400_)
  );
  MUX2_X1 _24607_ (
    .A(_04400_),
    .B(_12638_),
    .S(_02233_),
    .Z(_04401_)
  );
  MUX2_X1 _24608_ (
    .A(ex_reg_rs_msb_1[21]),
    .B(_04401_),
    .S(_02202_),
    .Z(_00170_)
  );
  AND2_X1 _24609_ (
    .A1(_08346_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04402_)
  );
  INV_X1 _24610_ (
    .A(_04402_),
    .ZN(_04403_)
  );
  AND2_X1 _24611_ (
    .A1(_08484_),
    .A2(_08546_),
    .ZN(_04404_)
  );
  INV_X1 _24612_ (
    .A(_04404_),
    .ZN(_04405_)
  );
  AND2_X1 _24613_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04405_),
    .ZN(_04406_)
  );
  AND2_X1 _24614_ (
    .A1(_04403_),
    .A2(_04406_),
    .ZN(_04407_)
  );
  INV_X1 _24615_ (
    .A(_04407_),
    .ZN(_04408_)
  );
  MUX2_X1 _24616_ (
    .A(\rf[15] [24]),
    .B(\rf[11] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04409_)
  );
  AND2_X1 _24617_ (
    .A1(_08544_),
    .A2(_04409_),
    .ZN(_04410_)
  );
  INV_X1 _24618_ (
    .A(_04410_),
    .ZN(_04411_)
  );
  AND2_X1 _24619_ (
    .A1(_08545_),
    .A2(_04411_),
    .ZN(_04412_)
  );
  AND2_X1 _24620_ (
    .A1(_04408_),
    .A2(_04412_),
    .ZN(_04413_)
  );
  INV_X1 _24621_ (
    .A(_04413_),
    .ZN(_04414_)
  );
  AND2_X1 _24622_ (
    .A1(_08367_),
    .A2(_08546_),
    .ZN(_04415_)
  );
  INV_X1 _24623_ (
    .A(_04415_),
    .ZN(_04416_)
  );
  AND2_X1 _24624_ (
    .A1(_08268_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04417_)
  );
  INV_X1 _24625_ (
    .A(_04417_),
    .ZN(_04418_)
  );
  AND2_X1 _24626_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04418_),
    .ZN(_04419_)
  );
  AND2_X1 _24627_ (
    .A1(_04416_),
    .A2(_04419_),
    .ZN(_04420_)
  );
  INV_X1 _24628_ (
    .A(_04420_),
    .ZN(_04421_)
  );
  MUX2_X1 _24629_ (
    .A(\rf[13] [24]),
    .B(\rf[9] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04422_)
  );
  AND2_X1 _24630_ (
    .A1(_08544_),
    .A2(_04422_),
    .ZN(_04423_)
  );
  INV_X1 _24631_ (
    .A(_04423_),
    .ZN(_04424_)
  );
  AND2_X1 _24632_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04424_),
    .ZN(_04425_)
  );
  AND2_X1 _24633_ (
    .A1(_04421_),
    .A2(_04425_),
    .ZN(_04426_)
  );
  INV_X1 _24634_ (
    .A(_04426_),
    .ZN(_04427_)
  );
  AND2_X1 _24635_ (
    .A1(_08547_),
    .A2(_04427_),
    .ZN(_04428_)
  );
  AND2_X1 _24636_ (
    .A1(_04414_),
    .A2(_04428_),
    .ZN(_04429_)
  );
  INV_X1 _24637_ (
    .A(_04429_),
    .ZN(_04430_)
  );
  MUX2_X1 _24638_ (
    .A(\rf[6] [24]),
    .B(\rf[2] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04431_)
  );
  AND2_X1 _24639_ (
    .A1(_08545_),
    .A2(_04431_),
    .ZN(_04432_)
  );
  INV_X1 _24640_ (
    .A(_04432_),
    .ZN(_04433_)
  );
  MUX2_X1 _24641_ (
    .A(\rf[4] [24]),
    .B(\rf[0] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04434_)
  );
  AND2_X1 _24642_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04434_),
    .ZN(_04435_)
  );
  INV_X1 _24643_ (
    .A(_04435_),
    .ZN(_04436_)
  );
  AND2_X1 _24644_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04436_),
    .ZN(_04437_)
  );
  AND2_X1 _24645_ (
    .A1(_04433_),
    .A2(_04437_),
    .ZN(_04438_)
  );
  INV_X1 _24646_ (
    .A(_04438_),
    .ZN(_04439_)
  );
  MUX2_X1 _24647_ (
    .A(\rf[7] [24]),
    .B(\rf[3] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04440_)
  );
  AND2_X1 _24648_ (
    .A1(_08545_),
    .A2(_04440_),
    .ZN(_04441_)
  );
  INV_X1 _24649_ (
    .A(_04441_),
    .ZN(_04442_)
  );
  MUX2_X1 _24650_ (
    .A(\rf[5] [24]),
    .B(\rf[1] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04443_)
  );
  AND2_X1 _24651_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04443_),
    .ZN(_04444_)
  );
  INV_X1 _24652_ (
    .A(_04444_),
    .ZN(_04445_)
  );
  AND2_X1 _24653_ (
    .A1(_08544_),
    .A2(_04445_),
    .ZN(_04446_)
  );
  AND2_X1 _24654_ (
    .A1(_04442_),
    .A2(_04446_),
    .ZN(_04447_)
  );
  INV_X1 _24655_ (
    .A(_04447_),
    .ZN(_04448_)
  );
  AND2_X1 _24656_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_04448_),
    .ZN(_04449_)
  );
  AND2_X1 _24657_ (
    .A1(_04439_),
    .A2(_04449_),
    .ZN(_04450_)
  );
  INV_X1 _24658_ (
    .A(_04450_),
    .ZN(_04451_)
  );
  AND2_X1 _24659_ (
    .A1(_04430_),
    .A2(_04451_),
    .ZN(_04452_)
  );
  AND2_X1 _24660_ (
    .A1(_08328_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04453_)
  );
  INV_X1 _24661_ (
    .A(_04453_),
    .ZN(_04454_)
  );
  AND2_X1 _24662_ (
    .A1(_08427_),
    .A2(_08546_),
    .ZN(_04455_)
  );
  INV_X1 _24663_ (
    .A(_04455_),
    .ZN(_04456_)
  );
  AND2_X1 _24664_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04456_),
    .ZN(_04457_)
  );
  AND2_X1 _24665_ (
    .A1(_04454_),
    .A2(_04457_),
    .ZN(_04458_)
  );
  INV_X1 _24666_ (
    .A(_04458_),
    .ZN(_04459_)
  );
  MUX2_X1 _24667_ (
    .A(\rf[23] [24]),
    .B(\rf[19] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04460_)
  );
  AND2_X1 _24668_ (
    .A1(_08545_),
    .A2(_04460_),
    .ZN(_04461_)
  );
  INV_X1 _24669_ (
    .A(_04461_),
    .ZN(_04462_)
  );
  AND2_X1 _24670_ (
    .A1(_08544_),
    .A2(_04462_),
    .ZN(_04463_)
  );
  AND2_X1 _24671_ (
    .A1(_04459_),
    .A2(_04463_),
    .ZN(_04464_)
  );
  INV_X1 _24672_ (
    .A(_04464_),
    .ZN(_04465_)
  );
  AND2_X1 _24673_ (
    .A1(_08397_),
    .A2(_08546_),
    .ZN(_04466_)
  );
  INV_X1 _24674_ (
    .A(_04466_),
    .ZN(_04467_)
  );
  AND2_X1 _24675_ (
    .A1(_08298_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04468_)
  );
  INV_X1 _24676_ (
    .A(_04468_),
    .ZN(_04469_)
  );
  AND2_X1 _24677_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04469_),
    .ZN(_04470_)
  );
  AND2_X1 _24678_ (
    .A1(_04467_),
    .A2(_04470_),
    .ZN(_04471_)
  );
  INV_X1 _24679_ (
    .A(_04471_),
    .ZN(_04472_)
  );
  MUX2_X1 _24680_ (
    .A(\rf[22] [24]),
    .B(\rf[18] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04473_)
  );
  AND2_X1 _24681_ (
    .A1(_08545_),
    .A2(_04473_),
    .ZN(_04474_)
  );
  INV_X1 _24682_ (
    .A(_04474_),
    .ZN(_04475_)
  );
  AND2_X1 _24683_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04475_),
    .ZN(_04476_)
  );
  AND2_X1 _24684_ (
    .A1(_04472_),
    .A2(_04476_),
    .ZN(_04477_)
  );
  INV_X1 _24685_ (
    .A(_04477_),
    .ZN(_04478_)
  );
  AND2_X1 _24686_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_04465_),
    .ZN(_04479_)
  );
  AND2_X1 _24687_ (
    .A1(_04478_),
    .A2(_04479_),
    .ZN(_04480_)
  );
  INV_X1 _24688_ (
    .A(_04480_),
    .ZN(_04481_)
  );
  AND2_X1 _24689_ (
    .A1(_08452_),
    .A2(_08546_),
    .ZN(_04482_)
  );
  INV_X1 _24690_ (
    .A(_04482_),
    .ZN(_04483_)
  );
  AND2_X1 _24691_ (
    .A1(_08522_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04484_)
  );
  INV_X1 _24692_ (
    .A(_04484_),
    .ZN(_04485_)
  );
  AND2_X1 _24693_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04485_),
    .ZN(_04486_)
  );
  AND2_X1 _24694_ (
    .A1(_04483_),
    .A2(_04486_),
    .ZN(_04487_)
  );
  INV_X1 _24695_ (
    .A(_04487_),
    .ZN(_04488_)
  );
  MUX2_X1 _24696_ (
    .A(\rf[30] [24]),
    .B(\rf[26] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04489_)
  );
  AND2_X1 _24697_ (
    .A1(_08545_),
    .A2(_04489_),
    .ZN(_04490_)
  );
  INV_X1 _24698_ (
    .A(_04490_),
    .ZN(_04491_)
  );
  AND2_X1 _24699_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04491_),
    .ZN(_04492_)
  );
  AND2_X1 _24700_ (
    .A1(_04488_),
    .A2(_04492_),
    .ZN(_04493_)
  );
  INV_X1 _24701_ (
    .A(_04493_),
    .ZN(_04494_)
  );
  MUX2_X1 _24702_ (
    .A(\rf[29] [24]),
    .B(\rf[25] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04495_)
  );
  AND2_X1 _24703_ (
    .A1(\rf[27] [24]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04496_)
  );
  MUX2_X1 _24704_ (
    .A(_04495_),
    .B(_04496_),
    .S(_08545_),
    .Z(_04497_)
  );
  INV_X1 _24705_ (
    .A(_04497_),
    .ZN(_04498_)
  );
  AND2_X1 _24706_ (
    .A1(_08544_),
    .A2(_04498_),
    .ZN(_04499_)
  );
  INV_X1 _24707_ (
    .A(_04499_),
    .ZN(_04500_)
  );
  AND2_X1 _24708_ (
    .A1(_08547_),
    .A2(_04500_),
    .ZN(_04501_)
  );
  AND2_X1 _24709_ (
    .A1(_04494_),
    .A2(_04501_),
    .ZN(_04502_)
  );
  INV_X1 _24710_ (
    .A(_04502_),
    .ZN(_04503_)
  );
  AND2_X1 _24711_ (
    .A1(_04481_),
    .A2(_04503_),
    .ZN(_04504_)
  );
  MUX2_X1 _24712_ (
    .A(_04452_),
    .B(_04504_),
    .S(_08572_),
    .Z(_04505_)
  );
  INV_X1 _24713_ (
    .A(_04505_),
    .ZN(_04506_)
  );
  MUX2_X1 _24714_ (
    .A(_04506_),
    .B(_12649_),
    .S(_02233_),
    .Z(_04507_)
  );
  MUX2_X1 _24715_ (
    .A(ex_reg_rs_msb_1[22]),
    .B(_04507_),
    .S(_02202_),
    .Z(_00171_)
  );
  AND2_X1 _24716_ (
    .A1(_08347_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04508_)
  );
  INV_X1 _24717_ (
    .A(_04508_),
    .ZN(_04509_)
  );
  AND2_X1 _24718_ (
    .A1(_08485_),
    .A2(_08546_),
    .ZN(_04510_)
  );
  INV_X1 _24719_ (
    .A(_04510_),
    .ZN(_04511_)
  );
  AND2_X1 _24720_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04511_),
    .ZN(_04512_)
  );
  AND2_X1 _24721_ (
    .A1(_04509_),
    .A2(_04512_),
    .ZN(_04513_)
  );
  INV_X1 _24722_ (
    .A(_04513_),
    .ZN(_04514_)
  );
  MUX2_X1 _24723_ (
    .A(\rf[15] [25]),
    .B(\rf[11] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04515_)
  );
  AND2_X1 _24724_ (
    .A1(_08544_),
    .A2(_04515_),
    .ZN(_04516_)
  );
  INV_X1 _24725_ (
    .A(_04516_),
    .ZN(_04517_)
  );
  AND2_X1 _24726_ (
    .A1(_08545_),
    .A2(_04517_),
    .ZN(_04518_)
  );
  AND2_X1 _24727_ (
    .A1(_04514_),
    .A2(_04518_),
    .ZN(_04519_)
  );
  INV_X1 _24728_ (
    .A(_04519_),
    .ZN(_04520_)
  );
  AND2_X1 _24729_ (
    .A1(_08368_),
    .A2(_08546_),
    .ZN(_04521_)
  );
  INV_X1 _24730_ (
    .A(_04521_),
    .ZN(_04522_)
  );
  AND2_X1 _24731_ (
    .A1(_08269_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04523_)
  );
  INV_X1 _24732_ (
    .A(_04523_),
    .ZN(_04524_)
  );
  AND2_X1 _24733_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04524_),
    .ZN(_04525_)
  );
  AND2_X1 _24734_ (
    .A1(_04522_),
    .A2(_04525_),
    .ZN(_04526_)
  );
  INV_X1 _24735_ (
    .A(_04526_),
    .ZN(_04527_)
  );
  MUX2_X1 _24736_ (
    .A(\rf[13] [25]),
    .B(\rf[9] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04528_)
  );
  AND2_X1 _24737_ (
    .A1(_08544_),
    .A2(_04528_),
    .ZN(_04529_)
  );
  INV_X1 _24738_ (
    .A(_04529_),
    .ZN(_04530_)
  );
  AND2_X1 _24739_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04530_),
    .ZN(_04531_)
  );
  AND2_X1 _24740_ (
    .A1(_04527_),
    .A2(_04531_),
    .ZN(_04532_)
  );
  INV_X1 _24741_ (
    .A(_04532_),
    .ZN(_04533_)
  );
  AND2_X1 _24742_ (
    .A1(_08547_),
    .A2(_04533_),
    .ZN(_04534_)
  );
  AND2_X1 _24743_ (
    .A1(_04520_),
    .A2(_04534_),
    .ZN(_04535_)
  );
  INV_X1 _24744_ (
    .A(_04535_),
    .ZN(_04536_)
  );
  MUX2_X1 _24745_ (
    .A(\rf[6] [25]),
    .B(\rf[2] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04537_)
  );
  AND2_X1 _24746_ (
    .A1(_08545_),
    .A2(_04537_),
    .ZN(_04538_)
  );
  INV_X1 _24747_ (
    .A(_04538_),
    .ZN(_04539_)
  );
  MUX2_X1 _24748_ (
    .A(\rf[4] [25]),
    .B(\rf[0] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04540_)
  );
  AND2_X1 _24749_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04540_),
    .ZN(_04541_)
  );
  INV_X1 _24750_ (
    .A(_04541_),
    .ZN(_04542_)
  );
  AND2_X1 _24751_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04542_),
    .ZN(_04543_)
  );
  AND2_X1 _24752_ (
    .A1(_04539_),
    .A2(_04543_),
    .ZN(_04544_)
  );
  INV_X1 _24753_ (
    .A(_04544_),
    .ZN(_04545_)
  );
  MUX2_X1 _24754_ (
    .A(\rf[7] [25]),
    .B(\rf[3] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04546_)
  );
  AND2_X1 _24755_ (
    .A1(_08545_),
    .A2(_04546_),
    .ZN(_04547_)
  );
  INV_X1 _24756_ (
    .A(_04547_),
    .ZN(_04548_)
  );
  MUX2_X1 _24757_ (
    .A(\rf[5] [25]),
    .B(\rf[1] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04549_)
  );
  AND2_X1 _24758_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04549_),
    .ZN(_04550_)
  );
  INV_X1 _24759_ (
    .A(_04550_),
    .ZN(_04551_)
  );
  AND2_X1 _24760_ (
    .A1(_08544_),
    .A2(_04551_),
    .ZN(_04552_)
  );
  AND2_X1 _24761_ (
    .A1(_04548_),
    .A2(_04552_),
    .ZN(_04553_)
  );
  INV_X1 _24762_ (
    .A(_04553_),
    .ZN(_04554_)
  );
  AND2_X1 _24763_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_04554_),
    .ZN(_04555_)
  );
  AND2_X1 _24764_ (
    .A1(_04545_),
    .A2(_04555_),
    .ZN(_04556_)
  );
  INV_X1 _24765_ (
    .A(_04556_),
    .ZN(_04557_)
  );
  AND2_X1 _24766_ (
    .A1(_04536_),
    .A2(_04557_),
    .ZN(_04558_)
  );
  AND2_X1 _24767_ (
    .A1(_08329_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04559_)
  );
  INV_X1 _24768_ (
    .A(_04559_),
    .ZN(_04560_)
  );
  AND2_X1 _24769_ (
    .A1(_08428_),
    .A2(_08546_),
    .ZN(_04561_)
  );
  INV_X1 _24770_ (
    .A(_04561_),
    .ZN(_04562_)
  );
  AND2_X1 _24771_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04562_),
    .ZN(_04563_)
  );
  AND2_X1 _24772_ (
    .A1(_04560_),
    .A2(_04563_),
    .ZN(_04564_)
  );
  INV_X1 _24773_ (
    .A(_04564_),
    .ZN(_04565_)
  );
  MUX2_X1 _24774_ (
    .A(\rf[23] [25]),
    .B(\rf[19] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04566_)
  );
  AND2_X1 _24775_ (
    .A1(_08545_),
    .A2(_04566_),
    .ZN(_04567_)
  );
  INV_X1 _24776_ (
    .A(_04567_),
    .ZN(_04568_)
  );
  AND2_X1 _24777_ (
    .A1(_08544_),
    .A2(_04568_),
    .ZN(_04569_)
  );
  AND2_X1 _24778_ (
    .A1(_04565_),
    .A2(_04569_),
    .ZN(_04570_)
  );
  INV_X1 _24779_ (
    .A(_04570_),
    .ZN(_04571_)
  );
  AND2_X1 _24780_ (
    .A1(_08398_),
    .A2(_08546_),
    .ZN(_04572_)
  );
  INV_X1 _24781_ (
    .A(_04572_),
    .ZN(_04573_)
  );
  AND2_X1 _24782_ (
    .A1(_08299_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04574_)
  );
  INV_X1 _24783_ (
    .A(_04574_),
    .ZN(_04575_)
  );
  AND2_X1 _24784_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04575_),
    .ZN(_04576_)
  );
  AND2_X1 _24785_ (
    .A1(_04573_),
    .A2(_04576_),
    .ZN(_04577_)
  );
  INV_X1 _24786_ (
    .A(_04577_),
    .ZN(_04578_)
  );
  MUX2_X1 _24787_ (
    .A(\rf[22] [25]),
    .B(\rf[18] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04579_)
  );
  AND2_X1 _24788_ (
    .A1(_08545_),
    .A2(_04579_),
    .ZN(_04580_)
  );
  INV_X1 _24789_ (
    .A(_04580_),
    .ZN(_04581_)
  );
  AND2_X1 _24790_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04581_),
    .ZN(_04582_)
  );
  AND2_X1 _24791_ (
    .A1(_04578_),
    .A2(_04582_),
    .ZN(_04583_)
  );
  INV_X1 _24792_ (
    .A(_04583_),
    .ZN(_04584_)
  );
  AND2_X1 _24793_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_04571_),
    .ZN(_04585_)
  );
  AND2_X1 _24794_ (
    .A1(_04584_),
    .A2(_04585_),
    .ZN(_04586_)
  );
  INV_X1 _24795_ (
    .A(_04586_),
    .ZN(_04587_)
  );
  AND2_X1 _24796_ (
    .A1(_08453_),
    .A2(_08546_),
    .ZN(_04588_)
  );
  INV_X1 _24797_ (
    .A(_04588_),
    .ZN(_04589_)
  );
  AND2_X1 _24798_ (
    .A1(_08523_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04590_)
  );
  INV_X1 _24799_ (
    .A(_04590_),
    .ZN(_04591_)
  );
  AND2_X1 _24800_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04591_),
    .ZN(_04592_)
  );
  AND2_X1 _24801_ (
    .A1(_04589_),
    .A2(_04592_),
    .ZN(_04593_)
  );
  INV_X1 _24802_ (
    .A(_04593_),
    .ZN(_04594_)
  );
  MUX2_X1 _24803_ (
    .A(\rf[30] [25]),
    .B(\rf[26] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04595_)
  );
  AND2_X1 _24804_ (
    .A1(_08545_),
    .A2(_04595_),
    .ZN(_04596_)
  );
  INV_X1 _24805_ (
    .A(_04596_),
    .ZN(_04597_)
  );
  AND2_X1 _24806_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04597_),
    .ZN(_04598_)
  );
  AND2_X1 _24807_ (
    .A1(_04594_),
    .A2(_04598_),
    .ZN(_04599_)
  );
  INV_X1 _24808_ (
    .A(_04599_),
    .ZN(_04600_)
  );
  MUX2_X1 _24809_ (
    .A(\rf[29] [25]),
    .B(\rf[25] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04601_)
  );
  AND2_X1 _24810_ (
    .A1(\rf[27] [25]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04602_)
  );
  MUX2_X1 _24811_ (
    .A(_04601_),
    .B(_04602_),
    .S(_08545_),
    .Z(_04603_)
  );
  INV_X1 _24812_ (
    .A(_04603_),
    .ZN(_04604_)
  );
  AND2_X1 _24813_ (
    .A1(_08544_),
    .A2(_04604_),
    .ZN(_04605_)
  );
  INV_X1 _24814_ (
    .A(_04605_),
    .ZN(_04606_)
  );
  AND2_X1 _24815_ (
    .A1(_08547_),
    .A2(_04606_),
    .ZN(_04607_)
  );
  AND2_X1 _24816_ (
    .A1(_04600_),
    .A2(_04607_),
    .ZN(_04608_)
  );
  INV_X1 _24817_ (
    .A(_04608_),
    .ZN(_04609_)
  );
  AND2_X1 _24818_ (
    .A1(_04587_),
    .A2(_04609_),
    .ZN(_04610_)
  );
  MUX2_X1 _24819_ (
    .A(_04558_),
    .B(_04610_),
    .S(_08572_),
    .Z(_04611_)
  );
  INV_X1 _24820_ (
    .A(_04611_),
    .ZN(_04612_)
  );
  MUX2_X1 _24821_ (
    .A(_04612_),
    .B(_12765_),
    .S(_02233_),
    .Z(_04613_)
  );
  MUX2_X1 _24822_ (
    .A(ex_reg_rs_msb_1[23]),
    .B(_04613_),
    .S(_02202_),
    .Z(_00172_)
  );
  MUX2_X1 _24823_ (
    .A(\rf[1] [26]),
    .B(\rf[0] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_04614_)
  );
  MUX2_X1 _24824_ (
    .A(\rf[5] [26]),
    .B(\rf[4] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_04615_)
  );
  MUX2_X1 _24825_ (
    .A(_04614_),
    .B(_04615_),
    .S(_08546_),
    .Z(_04616_)
  );
  INV_X1 _24826_ (
    .A(_04616_),
    .ZN(_04617_)
  );
  AND2_X1 _24827_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_04617_),
    .ZN(_04618_)
  );
  INV_X1 _24828_ (
    .A(_04618_),
    .ZN(_04619_)
  );
  MUX2_X1 _24829_ (
    .A(\rf[13] [26]),
    .B(\rf[9] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04620_)
  );
  INV_X1 _24830_ (
    .A(_04620_),
    .ZN(_04621_)
  );
  AND2_X1 _24831_ (
    .A1(_09692_),
    .A2(_04621_),
    .ZN(_04622_)
  );
  INV_X1 _24832_ (
    .A(_04622_),
    .ZN(_04623_)
  );
  MUX2_X1 _24833_ (
    .A(\rf[12] [26]),
    .B(\rf[8] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04624_)
  );
  INV_X1 _24834_ (
    .A(_04624_),
    .ZN(_04625_)
  );
  AND2_X1 _24835_ (
    .A1(_02341_),
    .A2(_04625_),
    .ZN(_04626_)
  );
  INV_X1 _24836_ (
    .A(_04626_),
    .ZN(_04627_)
  );
  AND2_X1 _24837_ (
    .A1(_04623_),
    .A2(_04627_),
    .ZN(_04628_)
  );
  AND2_X1 _24838_ (
    .A1(_04619_),
    .A2(_04628_),
    .ZN(_04629_)
  );
  MUX2_X1 _24839_ (
    .A(\rf[3] [26]),
    .B(\rf[2] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_04630_)
  );
  MUX2_X1 _24840_ (
    .A(\rf[7] [26]),
    .B(\rf[6] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_04631_)
  );
  MUX2_X1 _24841_ (
    .A(_04630_),
    .B(_04631_),
    .S(_08546_),
    .Z(_04632_)
  );
  INV_X1 _24842_ (
    .A(_04632_),
    .ZN(_04633_)
  );
  AND2_X1 _24843_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_04633_),
    .ZN(_04634_)
  );
  INV_X1 _24844_ (
    .A(_04634_),
    .ZN(_04635_)
  );
  MUX2_X1 _24845_ (
    .A(\rf[14] [26]),
    .B(\rf[10] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04636_)
  );
  INV_X1 _24846_ (
    .A(_04636_),
    .ZN(_04637_)
  );
  AND2_X1 _24847_ (
    .A1(_02341_),
    .A2(_04637_),
    .ZN(_04638_)
  );
  INV_X1 _24848_ (
    .A(_04638_),
    .ZN(_04639_)
  );
  MUX2_X1 _24849_ (
    .A(\rf[15] [26]),
    .B(\rf[11] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04640_)
  );
  INV_X1 _24850_ (
    .A(_04640_),
    .ZN(_04641_)
  );
  AND2_X1 _24851_ (
    .A1(_09692_),
    .A2(_04641_),
    .ZN(_04642_)
  );
  INV_X1 _24852_ (
    .A(_04642_),
    .ZN(_04643_)
  );
  AND2_X1 _24853_ (
    .A1(_04639_),
    .A2(_04643_),
    .ZN(_04644_)
  );
  AND2_X1 _24854_ (
    .A1(_04635_),
    .A2(_04644_),
    .ZN(_04645_)
  );
  MUX2_X1 _24855_ (
    .A(_04629_),
    .B(_04645_),
    .S(_08545_),
    .Z(_04646_)
  );
  AND2_X1 _24856_ (
    .A1(_08330_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04647_)
  );
  INV_X1 _24857_ (
    .A(_04647_),
    .ZN(_04648_)
  );
  AND2_X1 _24858_ (
    .A1(_08429_),
    .A2(_08546_),
    .ZN(_04649_)
  );
  INV_X1 _24859_ (
    .A(_04649_),
    .ZN(_04650_)
  );
  AND2_X1 _24860_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04650_),
    .ZN(_04651_)
  );
  AND2_X1 _24861_ (
    .A1(_04648_),
    .A2(_04651_),
    .ZN(_04652_)
  );
  INV_X1 _24862_ (
    .A(_04652_),
    .ZN(_04653_)
  );
  MUX2_X1 _24863_ (
    .A(\rf[23] [26]),
    .B(\rf[19] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04654_)
  );
  AND2_X1 _24864_ (
    .A1(_08545_),
    .A2(_04654_),
    .ZN(_04655_)
  );
  INV_X1 _24865_ (
    .A(_04655_),
    .ZN(_04656_)
  );
  AND2_X1 _24866_ (
    .A1(_08544_),
    .A2(_04656_),
    .ZN(_04657_)
  );
  AND2_X1 _24867_ (
    .A1(_04653_),
    .A2(_04657_),
    .ZN(_04658_)
  );
  INV_X1 _24868_ (
    .A(_04658_),
    .ZN(_04659_)
  );
  AND2_X1 _24869_ (
    .A1(_08399_),
    .A2(_08546_),
    .ZN(_04660_)
  );
  INV_X1 _24870_ (
    .A(_04660_),
    .ZN(_04661_)
  );
  AND2_X1 _24871_ (
    .A1(_08300_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04662_)
  );
  INV_X1 _24872_ (
    .A(_04662_),
    .ZN(_04663_)
  );
  AND2_X1 _24873_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04663_),
    .ZN(_04664_)
  );
  AND2_X1 _24874_ (
    .A1(_04661_),
    .A2(_04664_),
    .ZN(_04665_)
  );
  INV_X1 _24875_ (
    .A(_04665_),
    .ZN(_04666_)
  );
  MUX2_X1 _24876_ (
    .A(\rf[22] [26]),
    .B(\rf[18] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04667_)
  );
  AND2_X1 _24877_ (
    .A1(_08545_),
    .A2(_04667_),
    .ZN(_04668_)
  );
  INV_X1 _24878_ (
    .A(_04668_),
    .ZN(_04669_)
  );
  AND2_X1 _24879_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04669_),
    .ZN(_04670_)
  );
  AND2_X1 _24880_ (
    .A1(_04666_),
    .A2(_04670_),
    .ZN(_04671_)
  );
  INV_X1 _24881_ (
    .A(_04671_),
    .ZN(_04672_)
  );
  AND2_X1 _24882_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_04659_),
    .ZN(_04673_)
  );
  AND2_X1 _24883_ (
    .A1(_04672_),
    .A2(_04673_),
    .ZN(_04674_)
  );
  INV_X1 _24884_ (
    .A(_04674_),
    .ZN(_04675_)
  );
  AND2_X1 _24885_ (
    .A1(_08454_),
    .A2(_08546_),
    .ZN(_04676_)
  );
  INV_X1 _24886_ (
    .A(_04676_),
    .ZN(_04677_)
  );
  AND2_X1 _24887_ (
    .A1(_08524_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04678_)
  );
  INV_X1 _24888_ (
    .A(_04678_),
    .ZN(_04679_)
  );
  AND2_X1 _24889_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04679_),
    .ZN(_04680_)
  );
  AND2_X1 _24890_ (
    .A1(_04677_),
    .A2(_04680_),
    .ZN(_04681_)
  );
  INV_X1 _24891_ (
    .A(_04681_),
    .ZN(_04682_)
  );
  MUX2_X1 _24892_ (
    .A(\rf[30] [26]),
    .B(\rf[26] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04683_)
  );
  AND2_X1 _24893_ (
    .A1(_08545_),
    .A2(_04683_),
    .ZN(_04684_)
  );
  INV_X1 _24894_ (
    .A(_04684_),
    .ZN(_04685_)
  );
  AND2_X1 _24895_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04685_),
    .ZN(_04686_)
  );
  AND2_X1 _24896_ (
    .A1(_04682_),
    .A2(_04686_),
    .ZN(_04687_)
  );
  INV_X1 _24897_ (
    .A(_04687_),
    .ZN(_04688_)
  );
  MUX2_X1 _24898_ (
    .A(\rf[29] [26]),
    .B(\rf[25] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04689_)
  );
  AND2_X1 _24899_ (
    .A1(\rf[27] [26]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04690_)
  );
  MUX2_X1 _24900_ (
    .A(_04689_),
    .B(_04690_),
    .S(_08545_),
    .Z(_04691_)
  );
  INV_X1 _24901_ (
    .A(_04691_),
    .ZN(_04692_)
  );
  AND2_X1 _24902_ (
    .A1(_08544_),
    .A2(_04692_),
    .ZN(_04693_)
  );
  INV_X1 _24903_ (
    .A(_04693_),
    .ZN(_04694_)
  );
  AND2_X1 _24904_ (
    .A1(_08547_),
    .A2(_04694_),
    .ZN(_04695_)
  );
  AND2_X1 _24905_ (
    .A1(_04688_),
    .A2(_04695_),
    .ZN(_04696_)
  );
  INV_X1 _24906_ (
    .A(_04696_),
    .ZN(_04697_)
  );
  AND2_X1 _24907_ (
    .A1(_04675_),
    .A2(_04697_),
    .ZN(_04698_)
  );
  INV_X1 _24908_ (
    .A(_04698_),
    .ZN(_04699_)
  );
  MUX2_X1 _24909_ (
    .A(_04646_),
    .B(_04699_),
    .S(_08572_),
    .Z(_04700_)
  );
  MUX2_X1 _24910_ (
    .A(_04700_),
    .B(_12986_),
    .S(_02233_),
    .Z(_04701_)
  );
  MUX2_X1 _24911_ (
    .A(ex_reg_rs_msb_1[24]),
    .B(_04701_),
    .S(_02202_),
    .Z(_00173_)
  );
  AND2_X1 _24912_ (
    .A1(_08348_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04702_)
  );
  INV_X1 _24913_ (
    .A(_04702_),
    .ZN(_04703_)
  );
  AND2_X1 _24914_ (
    .A1(_08486_),
    .A2(_08546_),
    .ZN(_04704_)
  );
  INV_X1 _24915_ (
    .A(_04704_),
    .ZN(_04705_)
  );
  AND2_X1 _24916_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04705_),
    .ZN(_04706_)
  );
  AND2_X1 _24917_ (
    .A1(_04703_),
    .A2(_04706_),
    .ZN(_04707_)
  );
  INV_X1 _24918_ (
    .A(_04707_),
    .ZN(_04708_)
  );
  MUX2_X1 _24919_ (
    .A(\rf[15] [27]),
    .B(\rf[11] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04709_)
  );
  AND2_X1 _24920_ (
    .A1(_08544_),
    .A2(_04709_),
    .ZN(_04710_)
  );
  INV_X1 _24921_ (
    .A(_04710_),
    .ZN(_04711_)
  );
  AND2_X1 _24922_ (
    .A1(_08545_),
    .A2(_04711_),
    .ZN(_04712_)
  );
  AND2_X1 _24923_ (
    .A1(_04708_),
    .A2(_04712_),
    .ZN(_04713_)
  );
  INV_X1 _24924_ (
    .A(_04713_),
    .ZN(_04714_)
  );
  AND2_X1 _24925_ (
    .A1(_08369_),
    .A2(_08546_),
    .ZN(_04715_)
  );
  INV_X1 _24926_ (
    .A(_04715_),
    .ZN(_04716_)
  );
  AND2_X1 _24927_ (
    .A1(_08270_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04717_)
  );
  INV_X1 _24928_ (
    .A(_04717_),
    .ZN(_04718_)
  );
  AND2_X1 _24929_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04718_),
    .ZN(_04719_)
  );
  AND2_X1 _24930_ (
    .A1(_04716_),
    .A2(_04719_),
    .ZN(_04720_)
  );
  INV_X1 _24931_ (
    .A(_04720_),
    .ZN(_04721_)
  );
  MUX2_X1 _24932_ (
    .A(\rf[13] [27]),
    .B(\rf[9] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04722_)
  );
  AND2_X1 _24933_ (
    .A1(_08544_),
    .A2(_04722_),
    .ZN(_04723_)
  );
  INV_X1 _24934_ (
    .A(_04723_),
    .ZN(_04724_)
  );
  AND2_X1 _24935_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04724_),
    .ZN(_04725_)
  );
  AND2_X1 _24936_ (
    .A1(_04721_),
    .A2(_04725_),
    .ZN(_04726_)
  );
  INV_X1 _24937_ (
    .A(_04726_),
    .ZN(_04727_)
  );
  AND2_X1 _24938_ (
    .A1(_08547_),
    .A2(_04727_),
    .ZN(_04728_)
  );
  AND2_X1 _24939_ (
    .A1(_04714_),
    .A2(_04728_),
    .ZN(_04729_)
  );
  INV_X1 _24940_ (
    .A(_04729_),
    .ZN(_04730_)
  );
  MUX2_X1 _24941_ (
    .A(\rf[6] [27]),
    .B(\rf[2] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04731_)
  );
  AND2_X1 _24942_ (
    .A1(_08545_),
    .A2(_04731_),
    .ZN(_04732_)
  );
  INV_X1 _24943_ (
    .A(_04732_),
    .ZN(_04733_)
  );
  MUX2_X1 _24944_ (
    .A(\rf[4] [27]),
    .B(\rf[0] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04734_)
  );
  AND2_X1 _24945_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04734_),
    .ZN(_04735_)
  );
  INV_X1 _24946_ (
    .A(_04735_),
    .ZN(_04736_)
  );
  AND2_X1 _24947_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04736_),
    .ZN(_04737_)
  );
  AND2_X1 _24948_ (
    .A1(_04733_),
    .A2(_04737_),
    .ZN(_04738_)
  );
  INV_X1 _24949_ (
    .A(_04738_),
    .ZN(_04739_)
  );
  MUX2_X1 _24950_ (
    .A(\rf[7] [27]),
    .B(\rf[3] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04740_)
  );
  AND2_X1 _24951_ (
    .A1(_08545_),
    .A2(_04740_),
    .ZN(_04741_)
  );
  INV_X1 _24952_ (
    .A(_04741_),
    .ZN(_04742_)
  );
  MUX2_X1 _24953_ (
    .A(\rf[5] [27]),
    .B(\rf[1] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04743_)
  );
  AND2_X1 _24954_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04743_),
    .ZN(_04744_)
  );
  INV_X1 _24955_ (
    .A(_04744_),
    .ZN(_04745_)
  );
  AND2_X1 _24956_ (
    .A1(_08544_),
    .A2(_04745_),
    .ZN(_04746_)
  );
  AND2_X1 _24957_ (
    .A1(_04742_),
    .A2(_04746_),
    .ZN(_04747_)
  );
  INV_X1 _24958_ (
    .A(_04747_),
    .ZN(_04748_)
  );
  AND2_X1 _24959_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_04748_),
    .ZN(_04749_)
  );
  AND2_X1 _24960_ (
    .A1(_04739_),
    .A2(_04749_),
    .ZN(_04750_)
  );
  INV_X1 _24961_ (
    .A(_04750_),
    .ZN(_04751_)
  );
  AND2_X1 _24962_ (
    .A1(_04730_),
    .A2(_04751_),
    .ZN(_04752_)
  );
  AND2_X1 _24963_ (
    .A1(_08331_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04753_)
  );
  INV_X1 _24964_ (
    .A(_04753_),
    .ZN(_04754_)
  );
  AND2_X1 _24965_ (
    .A1(_08430_),
    .A2(_08546_),
    .ZN(_04755_)
  );
  INV_X1 _24966_ (
    .A(_04755_),
    .ZN(_04756_)
  );
  AND2_X1 _24967_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04756_),
    .ZN(_04757_)
  );
  AND2_X1 _24968_ (
    .A1(_04754_),
    .A2(_04757_),
    .ZN(_04758_)
  );
  INV_X1 _24969_ (
    .A(_04758_),
    .ZN(_04759_)
  );
  MUX2_X1 _24970_ (
    .A(\rf[23] [27]),
    .B(\rf[19] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04760_)
  );
  AND2_X1 _24971_ (
    .A1(_08545_),
    .A2(_04760_),
    .ZN(_04761_)
  );
  INV_X1 _24972_ (
    .A(_04761_),
    .ZN(_04762_)
  );
  AND2_X1 _24973_ (
    .A1(_08544_),
    .A2(_04762_),
    .ZN(_04763_)
  );
  AND2_X1 _24974_ (
    .A1(_04759_),
    .A2(_04763_),
    .ZN(_04764_)
  );
  INV_X1 _24975_ (
    .A(_04764_),
    .ZN(_04765_)
  );
  AND2_X1 _24976_ (
    .A1(_08400_),
    .A2(_08546_),
    .ZN(_04766_)
  );
  INV_X1 _24977_ (
    .A(_04766_),
    .ZN(_04767_)
  );
  AND2_X1 _24978_ (
    .A1(_08301_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04768_)
  );
  INV_X1 _24979_ (
    .A(_04768_),
    .ZN(_04769_)
  );
  AND2_X1 _24980_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04769_),
    .ZN(_04770_)
  );
  AND2_X1 _24981_ (
    .A1(_04767_),
    .A2(_04770_),
    .ZN(_04771_)
  );
  INV_X1 _24982_ (
    .A(_04771_),
    .ZN(_04772_)
  );
  MUX2_X1 _24983_ (
    .A(\rf[22] [27]),
    .B(\rf[18] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04773_)
  );
  AND2_X1 _24984_ (
    .A1(_08545_),
    .A2(_04773_),
    .ZN(_04774_)
  );
  INV_X1 _24985_ (
    .A(_04774_),
    .ZN(_04775_)
  );
  AND2_X1 _24986_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04775_),
    .ZN(_04776_)
  );
  AND2_X1 _24987_ (
    .A1(_04772_),
    .A2(_04776_),
    .ZN(_04777_)
  );
  INV_X1 _24988_ (
    .A(_04777_),
    .ZN(_04778_)
  );
  AND2_X1 _24989_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_04765_),
    .ZN(_04779_)
  );
  AND2_X1 _24990_ (
    .A1(_04778_),
    .A2(_04779_),
    .ZN(_04780_)
  );
  INV_X1 _24991_ (
    .A(_04780_),
    .ZN(_04781_)
  );
  AND2_X1 _24992_ (
    .A1(_08455_),
    .A2(_08546_),
    .ZN(_04782_)
  );
  INV_X1 _24993_ (
    .A(_04782_),
    .ZN(_04783_)
  );
  AND2_X1 _24994_ (
    .A1(_08525_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04784_)
  );
  INV_X1 _24995_ (
    .A(_04784_),
    .ZN(_04785_)
  );
  AND2_X1 _24996_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04785_),
    .ZN(_04786_)
  );
  AND2_X1 _24997_ (
    .A1(_04783_),
    .A2(_04786_),
    .ZN(_04787_)
  );
  INV_X1 _24998_ (
    .A(_04787_),
    .ZN(_04788_)
  );
  MUX2_X1 _24999_ (
    .A(\rf[30] [27]),
    .B(\rf[26] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04789_)
  );
  AND2_X1 _25000_ (
    .A1(_08545_),
    .A2(_04789_),
    .ZN(_04790_)
  );
  INV_X1 _25001_ (
    .A(_04790_),
    .ZN(_04791_)
  );
  AND2_X1 _25002_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04791_),
    .ZN(_04792_)
  );
  AND2_X1 _25003_ (
    .A1(_04788_),
    .A2(_04792_),
    .ZN(_04793_)
  );
  INV_X1 _25004_ (
    .A(_04793_),
    .ZN(_04794_)
  );
  MUX2_X1 _25005_ (
    .A(\rf[29] [27]),
    .B(\rf[25] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04795_)
  );
  AND2_X1 _25006_ (
    .A1(\rf[27] [27]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04796_)
  );
  MUX2_X1 _25007_ (
    .A(_04795_),
    .B(_04796_),
    .S(_08545_),
    .Z(_04797_)
  );
  INV_X1 _25008_ (
    .A(_04797_),
    .ZN(_04798_)
  );
  AND2_X1 _25009_ (
    .A1(_08544_),
    .A2(_04798_),
    .ZN(_04799_)
  );
  INV_X1 _25010_ (
    .A(_04799_),
    .ZN(_04800_)
  );
  AND2_X1 _25011_ (
    .A1(_08547_),
    .A2(_04800_),
    .ZN(_04801_)
  );
  AND2_X1 _25012_ (
    .A1(_04794_),
    .A2(_04801_),
    .ZN(_04802_)
  );
  INV_X1 _25013_ (
    .A(_04802_),
    .ZN(_04803_)
  );
  AND2_X1 _25014_ (
    .A1(_04781_),
    .A2(_04803_),
    .ZN(_04804_)
  );
  MUX2_X1 _25015_ (
    .A(_04752_),
    .B(_04804_),
    .S(_08572_),
    .Z(_04805_)
  );
  INV_X1 _25016_ (
    .A(_04805_),
    .ZN(_04806_)
  );
  MUX2_X1 _25017_ (
    .A(_04806_),
    .B(_13102_),
    .S(_02233_),
    .Z(_04807_)
  );
  MUX2_X1 _25018_ (
    .A(ex_reg_rs_msb_1[25]),
    .B(_04807_),
    .S(_02202_),
    .Z(_00174_)
  );
  AND2_X1 _25019_ (
    .A1(_08349_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04808_)
  );
  INV_X1 _25020_ (
    .A(_04808_),
    .ZN(_04809_)
  );
  AND2_X1 _25021_ (
    .A1(_08487_),
    .A2(_08546_),
    .ZN(_04810_)
  );
  INV_X1 _25022_ (
    .A(_04810_),
    .ZN(_04811_)
  );
  AND2_X1 _25023_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04811_),
    .ZN(_04812_)
  );
  AND2_X1 _25024_ (
    .A1(_04809_),
    .A2(_04812_),
    .ZN(_04813_)
  );
  INV_X1 _25025_ (
    .A(_04813_),
    .ZN(_04814_)
  );
  MUX2_X1 _25026_ (
    .A(\rf[15] [28]),
    .B(\rf[11] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04815_)
  );
  AND2_X1 _25027_ (
    .A1(_08544_),
    .A2(_04815_),
    .ZN(_04816_)
  );
  INV_X1 _25028_ (
    .A(_04816_),
    .ZN(_04817_)
  );
  AND2_X1 _25029_ (
    .A1(_08545_),
    .A2(_04817_),
    .ZN(_04818_)
  );
  AND2_X1 _25030_ (
    .A1(_04814_),
    .A2(_04818_),
    .ZN(_04819_)
  );
  INV_X1 _25031_ (
    .A(_04819_),
    .ZN(_04820_)
  );
  AND2_X1 _25032_ (
    .A1(_08370_),
    .A2(_08546_),
    .ZN(_04821_)
  );
  INV_X1 _25033_ (
    .A(_04821_),
    .ZN(_04822_)
  );
  AND2_X1 _25034_ (
    .A1(_08271_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04823_)
  );
  INV_X1 _25035_ (
    .A(_04823_),
    .ZN(_04824_)
  );
  AND2_X1 _25036_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04824_),
    .ZN(_04825_)
  );
  AND2_X1 _25037_ (
    .A1(_04822_),
    .A2(_04825_),
    .ZN(_04826_)
  );
  INV_X1 _25038_ (
    .A(_04826_),
    .ZN(_04827_)
  );
  MUX2_X1 _25039_ (
    .A(\rf[13] [28]),
    .B(\rf[9] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04828_)
  );
  AND2_X1 _25040_ (
    .A1(_08544_),
    .A2(_04828_),
    .ZN(_04829_)
  );
  INV_X1 _25041_ (
    .A(_04829_),
    .ZN(_04830_)
  );
  AND2_X1 _25042_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04830_),
    .ZN(_04831_)
  );
  AND2_X1 _25043_ (
    .A1(_04827_),
    .A2(_04831_),
    .ZN(_04832_)
  );
  INV_X1 _25044_ (
    .A(_04832_),
    .ZN(_04833_)
  );
  AND2_X1 _25045_ (
    .A1(_08547_),
    .A2(_04833_),
    .ZN(_04834_)
  );
  AND2_X1 _25046_ (
    .A1(_04820_),
    .A2(_04834_),
    .ZN(_04835_)
  );
  INV_X1 _25047_ (
    .A(_04835_),
    .ZN(_04836_)
  );
  MUX2_X1 _25048_ (
    .A(\rf[6] [28]),
    .B(\rf[2] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04837_)
  );
  AND2_X1 _25049_ (
    .A1(_08545_),
    .A2(_04837_),
    .ZN(_04838_)
  );
  INV_X1 _25050_ (
    .A(_04838_),
    .ZN(_04839_)
  );
  MUX2_X1 _25051_ (
    .A(\rf[4] [28]),
    .B(\rf[0] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04840_)
  );
  AND2_X1 _25052_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04840_),
    .ZN(_04841_)
  );
  INV_X1 _25053_ (
    .A(_04841_),
    .ZN(_04842_)
  );
  AND2_X1 _25054_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04842_),
    .ZN(_04843_)
  );
  AND2_X1 _25055_ (
    .A1(_04839_),
    .A2(_04843_),
    .ZN(_04844_)
  );
  INV_X1 _25056_ (
    .A(_04844_),
    .ZN(_04845_)
  );
  MUX2_X1 _25057_ (
    .A(\rf[7] [28]),
    .B(\rf[3] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04846_)
  );
  AND2_X1 _25058_ (
    .A1(_08545_),
    .A2(_04846_),
    .ZN(_04847_)
  );
  INV_X1 _25059_ (
    .A(_04847_),
    .ZN(_04848_)
  );
  MUX2_X1 _25060_ (
    .A(\rf[5] [28]),
    .B(\rf[1] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04849_)
  );
  AND2_X1 _25061_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04849_),
    .ZN(_04850_)
  );
  INV_X1 _25062_ (
    .A(_04850_),
    .ZN(_04851_)
  );
  AND2_X1 _25063_ (
    .A1(_08544_),
    .A2(_04851_),
    .ZN(_04852_)
  );
  AND2_X1 _25064_ (
    .A1(_04848_),
    .A2(_04852_),
    .ZN(_04853_)
  );
  INV_X1 _25065_ (
    .A(_04853_),
    .ZN(_04854_)
  );
  AND2_X1 _25066_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_04854_),
    .ZN(_04855_)
  );
  AND2_X1 _25067_ (
    .A1(_04845_),
    .A2(_04855_),
    .ZN(_04856_)
  );
  INV_X1 _25068_ (
    .A(_04856_),
    .ZN(_04857_)
  );
  AND2_X1 _25069_ (
    .A1(_04836_),
    .A2(_04857_),
    .ZN(_04858_)
  );
  AND2_X1 _25070_ (
    .A1(_08332_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04859_)
  );
  INV_X1 _25071_ (
    .A(_04859_),
    .ZN(_04860_)
  );
  AND2_X1 _25072_ (
    .A1(_08431_),
    .A2(_08546_),
    .ZN(_04861_)
  );
  INV_X1 _25073_ (
    .A(_04861_),
    .ZN(_04862_)
  );
  AND2_X1 _25074_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04862_),
    .ZN(_04863_)
  );
  AND2_X1 _25075_ (
    .A1(_04860_),
    .A2(_04863_),
    .ZN(_04864_)
  );
  INV_X1 _25076_ (
    .A(_04864_),
    .ZN(_04865_)
  );
  MUX2_X1 _25077_ (
    .A(\rf[23] [28]),
    .B(\rf[19] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04866_)
  );
  AND2_X1 _25078_ (
    .A1(_08545_),
    .A2(_04866_),
    .ZN(_04867_)
  );
  INV_X1 _25079_ (
    .A(_04867_),
    .ZN(_04868_)
  );
  AND2_X1 _25080_ (
    .A1(_08544_),
    .A2(_04868_),
    .ZN(_04869_)
  );
  AND2_X1 _25081_ (
    .A1(_04865_),
    .A2(_04869_),
    .ZN(_04870_)
  );
  INV_X1 _25082_ (
    .A(_04870_),
    .ZN(_04871_)
  );
  AND2_X1 _25083_ (
    .A1(_08401_),
    .A2(_08546_),
    .ZN(_04872_)
  );
  INV_X1 _25084_ (
    .A(_04872_),
    .ZN(_04873_)
  );
  AND2_X1 _25085_ (
    .A1(_08302_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04874_)
  );
  INV_X1 _25086_ (
    .A(_04874_),
    .ZN(_04875_)
  );
  AND2_X1 _25087_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04875_),
    .ZN(_04876_)
  );
  AND2_X1 _25088_ (
    .A1(_04873_),
    .A2(_04876_),
    .ZN(_04877_)
  );
  INV_X1 _25089_ (
    .A(_04877_),
    .ZN(_04878_)
  );
  MUX2_X1 _25090_ (
    .A(\rf[22] [28]),
    .B(\rf[18] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04879_)
  );
  AND2_X1 _25091_ (
    .A1(_08545_),
    .A2(_04879_),
    .ZN(_04880_)
  );
  INV_X1 _25092_ (
    .A(_04880_),
    .ZN(_04881_)
  );
  AND2_X1 _25093_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04881_),
    .ZN(_04882_)
  );
  AND2_X1 _25094_ (
    .A1(_04878_),
    .A2(_04882_),
    .ZN(_04883_)
  );
  INV_X1 _25095_ (
    .A(_04883_),
    .ZN(_04884_)
  );
  AND2_X1 _25096_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_04871_),
    .ZN(_04885_)
  );
  AND2_X1 _25097_ (
    .A1(_04884_),
    .A2(_04885_),
    .ZN(_04886_)
  );
  INV_X1 _25098_ (
    .A(_04886_),
    .ZN(_04887_)
  );
  AND2_X1 _25099_ (
    .A1(_08456_),
    .A2(_08546_),
    .ZN(_04888_)
  );
  INV_X1 _25100_ (
    .A(_04888_),
    .ZN(_04889_)
  );
  AND2_X1 _25101_ (
    .A1(_08526_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04890_)
  );
  INV_X1 _25102_ (
    .A(_04890_),
    .ZN(_04891_)
  );
  AND2_X1 _25103_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04891_),
    .ZN(_04892_)
  );
  AND2_X1 _25104_ (
    .A1(_04889_),
    .A2(_04892_),
    .ZN(_04893_)
  );
  INV_X1 _25105_ (
    .A(_04893_),
    .ZN(_04894_)
  );
  MUX2_X1 _25106_ (
    .A(\rf[30] [28]),
    .B(\rf[26] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04895_)
  );
  AND2_X1 _25107_ (
    .A1(_08545_),
    .A2(_04895_),
    .ZN(_04896_)
  );
  INV_X1 _25108_ (
    .A(_04896_),
    .ZN(_04897_)
  );
  AND2_X1 _25109_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04897_),
    .ZN(_04898_)
  );
  AND2_X1 _25110_ (
    .A1(_04894_),
    .A2(_04898_),
    .ZN(_04899_)
  );
  INV_X1 _25111_ (
    .A(_04899_),
    .ZN(_04900_)
  );
  MUX2_X1 _25112_ (
    .A(\rf[29] [28]),
    .B(\rf[25] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04901_)
  );
  AND2_X1 _25113_ (
    .A1(\rf[27] [28]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04902_)
  );
  MUX2_X1 _25114_ (
    .A(_04901_),
    .B(_04902_),
    .S(_08545_),
    .Z(_04903_)
  );
  INV_X1 _25115_ (
    .A(_04903_),
    .ZN(_04904_)
  );
  AND2_X1 _25116_ (
    .A1(_08544_),
    .A2(_04904_),
    .ZN(_04905_)
  );
  INV_X1 _25117_ (
    .A(_04905_),
    .ZN(_04906_)
  );
  AND2_X1 _25118_ (
    .A1(_08547_),
    .A2(_04906_),
    .ZN(_04907_)
  );
  AND2_X1 _25119_ (
    .A1(_04900_),
    .A2(_04907_),
    .ZN(_04908_)
  );
  INV_X1 _25120_ (
    .A(_04908_),
    .ZN(_04909_)
  );
  AND2_X1 _25121_ (
    .A1(_04887_),
    .A2(_04909_),
    .ZN(_04910_)
  );
  MUX2_X1 _25122_ (
    .A(_04858_),
    .B(_04910_),
    .S(_08572_),
    .Z(_04911_)
  );
  INV_X1 _25123_ (
    .A(_04911_),
    .ZN(_04912_)
  );
  MUX2_X1 _25124_ (
    .A(_04912_),
    .B(_13218_),
    .S(_02233_),
    .Z(_04913_)
  );
  MUX2_X1 _25125_ (
    .A(ex_reg_rs_msb_1[26]),
    .B(_04913_),
    .S(_02202_),
    .Z(_00175_)
  );
  MUX2_X1 _25126_ (
    .A(\rf[1] [29]),
    .B(\rf[0] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_04914_)
  );
  MUX2_X1 _25127_ (
    .A(\rf[5] [29]),
    .B(\rf[4] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_04915_)
  );
  MUX2_X1 _25128_ (
    .A(_04914_),
    .B(_04915_),
    .S(_08546_),
    .Z(_04916_)
  );
  INV_X1 _25129_ (
    .A(_04916_),
    .ZN(_04917_)
  );
  AND2_X1 _25130_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_04917_),
    .ZN(_04918_)
  );
  INV_X1 _25131_ (
    .A(_04918_),
    .ZN(_04919_)
  );
  MUX2_X1 _25132_ (
    .A(\rf[12] [29]),
    .B(\rf[8] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04920_)
  );
  INV_X1 _25133_ (
    .A(_04920_),
    .ZN(_04921_)
  );
  AND2_X1 _25134_ (
    .A1(_02341_),
    .A2(_04921_),
    .ZN(_04922_)
  );
  INV_X1 _25135_ (
    .A(_04922_),
    .ZN(_04923_)
  );
  MUX2_X1 _25136_ (
    .A(\rf[13] [29]),
    .B(\rf[9] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04924_)
  );
  INV_X1 _25137_ (
    .A(_04924_),
    .ZN(_04925_)
  );
  AND2_X1 _25138_ (
    .A1(_09692_),
    .A2(_04925_),
    .ZN(_04926_)
  );
  INV_X1 _25139_ (
    .A(_04926_),
    .ZN(_04927_)
  );
  AND2_X1 _25140_ (
    .A1(_04923_),
    .A2(_04927_),
    .ZN(_04928_)
  );
  AND2_X1 _25141_ (
    .A1(_04919_),
    .A2(_04928_),
    .ZN(_04929_)
  );
  MUX2_X1 _25142_ (
    .A(\rf[3] [29]),
    .B(\rf[2] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_04930_)
  );
  MUX2_X1 _25143_ (
    .A(\rf[7] [29]),
    .B(\rf[6] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_04931_)
  );
  MUX2_X1 _25144_ (
    .A(_04930_),
    .B(_04931_),
    .S(_08546_),
    .Z(_04932_)
  );
  INV_X1 _25145_ (
    .A(_04932_),
    .ZN(_04933_)
  );
  AND2_X1 _25146_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_04933_),
    .ZN(_04934_)
  );
  INV_X1 _25147_ (
    .A(_04934_),
    .ZN(_04935_)
  );
  MUX2_X1 _25148_ (
    .A(\rf[14] [29]),
    .B(\rf[10] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04936_)
  );
  INV_X1 _25149_ (
    .A(_04936_),
    .ZN(_04937_)
  );
  AND2_X1 _25150_ (
    .A1(_02341_),
    .A2(_04937_),
    .ZN(_04938_)
  );
  INV_X1 _25151_ (
    .A(_04938_),
    .ZN(_04939_)
  );
  MUX2_X1 _25152_ (
    .A(\rf[15] [29]),
    .B(\rf[11] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04940_)
  );
  INV_X1 _25153_ (
    .A(_04940_),
    .ZN(_04941_)
  );
  AND2_X1 _25154_ (
    .A1(_09692_),
    .A2(_04941_),
    .ZN(_04942_)
  );
  INV_X1 _25155_ (
    .A(_04942_),
    .ZN(_04943_)
  );
  AND2_X1 _25156_ (
    .A1(_04939_),
    .A2(_04943_),
    .ZN(_04944_)
  );
  AND2_X1 _25157_ (
    .A1(_04935_),
    .A2(_04944_),
    .ZN(_04945_)
  );
  MUX2_X1 _25158_ (
    .A(_04929_),
    .B(_04945_),
    .S(_08545_),
    .Z(_04946_)
  );
  AND2_X1 _25159_ (
    .A1(_08333_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04947_)
  );
  INV_X1 _25160_ (
    .A(_04947_),
    .ZN(_04948_)
  );
  AND2_X1 _25161_ (
    .A1(_08432_),
    .A2(_08546_),
    .ZN(_04949_)
  );
  INV_X1 _25162_ (
    .A(_04949_),
    .ZN(_04950_)
  );
  AND2_X1 _25163_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04950_),
    .ZN(_04951_)
  );
  AND2_X1 _25164_ (
    .A1(_04948_),
    .A2(_04951_),
    .ZN(_04952_)
  );
  INV_X1 _25165_ (
    .A(_04952_),
    .ZN(_04953_)
  );
  MUX2_X1 _25166_ (
    .A(\rf[23] [29]),
    .B(\rf[19] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04954_)
  );
  AND2_X1 _25167_ (
    .A1(_08545_),
    .A2(_04954_),
    .ZN(_04955_)
  );
  INV_X1 _25168_ (
    .A(_04955_),
    .ZN(_04956_)
  );
  AND2_X1 _25169_ (
    .A1(_08544_),
    .A2(_04956_),
    .ZN(_04957_)
  );
  AND2_X1 _25170_ (
    .A1(_04953_),
    .A2(_04957_),
    .ZN(_04958_)
  );
  INV_X1 _25171_ (
    .A(_04958_),
    .ZN(_04959_)
  );
  AND2_X1 _25172_ (
    .A1(_08402_),
    .A2(_08546_),
    .ZN(_04960_)
  );
  INV_X1 _25173_ (
    .A(_04960_),
    .ZN(_04961_)
  );
  AND2_X1 _25174_ (
    .A1(_08303_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04962_)
  );
  INV_X1 _25175_ (
    .A(_04962_),
    .ZN(_04963_)
  );
  AND2_X1 _25176_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04963_),
    .ZN(_04964_)
  );
  AND2_X1 _25177_ (
    .A1(_04961_),
    .A2(_04964_),
    .ZN(_04965_)
  );
  INV_X1 _25178_ (
    .A(_04965_),
    .ZN(_04966_)
  );
  MUX2_X1 _25179_ (
    .A(\rf[22] [29]),
    .B(\rf[18] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04967_)
  );
  AND2_X1 _25180_ (
    .A1(_08545_),
    .A2(_04967_),
    .ZN(_04968_)
  );
  INV_X1 _25181_ (
    .A(_04968_),
    .ZN(_04969_)
  );
  AND2_X1 _25182_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04969_),
    .ZN(_04970_)
  );
  AND2_X1 _25183_ (
    .A1(_04966_),
    .A2(_04970_),
    .ZN(_04971_)
  );
  INV_X1 _25184_ (
    .A(_04971_),
    .ZN(_04972_)
  );
  AND2_X1 _25185_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_04959_),
    .ZN(_04973_)
  );
  AND2_X1 _25186_ (
    .A1(_04972_),
    .A2(_04973_),
    .ZN(_04974_)
  );
  INV_X1 _25187_ (
    .A(_04974_),
    .ZN(_04975_)
  );
  AND2_X1 _25188_ (
    .A1(_08457_),
    .A2(_08546_),
    .ZN(_04976_)
  );
  INV_X1 _25189_ (
    .A(_04976_),
    .ZN(_04977_)
  );
  AND2_X1 _25190_ (
    .A1(_08527_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04978_)
  );
  INV_X1 _25191_ (
    .A(_04978_),
    .ZN(_04979_)
  );
  AND2_X1 _25192_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_04979_),
    .ZN(_04980_)
  );
  AND2_X1 _25193_ (
    .A1(_04977_),
    .A2(_04980_),
    .ZN(_04981_)
  );
  INV_X1 _25194_ (
    .A(_04981_),
    .ZN(_04982_)
  );
  MUX2_X1 _25195_ (
    .A(\rf[30] [29]),
    .B(\rf[26] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04983_)
  );
  AND2_X1 _25196_ (
    .A1(_08545_),
    .A2(_04983_),
    .ZN(_04984_)
  );
  INV_X1 _25197_ (
    .A(_04984_),
    .ZN(_04985_)
  );
  AND2_X1 _25198_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_04985_),
    .ZN(_04986_)
  );
  AND2_X1 _25199_ (
    .A1(_04982_),
    .A2(_04986_),
    .ZN(_04987_)
  );
  INV_X1 _25200_ (
    .A(_04987_),
    .ZN(_04988_)
  );
  MUX2_X1 _25201_ (
    .A(\rf[29] [29]),
    .B(\rf[25] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_04989_)
  );
  AND2_X1 _25202_ (
    .A1(\rf[27] [29]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_04990_)
  );
  MUX2_X1 _25203_ (
    .A(_04989_),
    .B(_04990_),
    .S(_08545_),
    .Z(_04991_)
  );
  INV_X1 _25204_ (
    .A(_04991_),
    .ZN(_04992_)
  );
  AND2_X1 _25205_ (
    .A1(_08544_),
    .A2(_04992_),
    .ZN(_04993_)
  );
  INV_X1 _25206_ (
    .A(_04993_),
    .ZN(_04994_)
  );
  AND2_X1 _25207_ (
    .A1(_08547_),
    .A2(_04994_),
    .ZN(_04995_)
  );
  AND2_X1 _25208_ (
    .A1(_04988_),
    .A2(_04995_),
    .ZN(_04996_)
  );
  INV_X1 _25209_ (
    .A(_04996_),
    .ZN(_04997_)
  );
  AND2_X1 _25210_ (
    .A1(_04975_),
    .A2(_04997_),
    .ZN(_04998_)
  );
  INV_X1 _25211_ (
    .A(_04998_),
    .ZN(_04999_)
  );
  MUX2_X1 _25212_ (
    .A(_04946_),
    .B(_04999_),
    .S(_08572_),
    .Z(_05000_)
  );
  MUX2_X1 _25213_ (
    .A(_05000_),
    .B(_13338_),
    .S(_02233_),
    .Z(_05001_)
  );
  MUX2_X1 _25214_ (
    .A(ex_reg_rs_msb_1[27]),
    .B(_05001_),
    .S(_02202_),
    .Z(_00176_)
  );
  AND2_X1 _25215_ (
    .A1(_08351_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_05002_)
  );
  INV_X1 _25216_ (
    .A(_05002_),
    .ZN(_05003_)
  );
  AND2_X1 _25217_ (
    .A1(_08489_),
    .A2(_08546_),
    .ZN(_05004_)
  );
  INV_X1 _25218_ (
    .A(_05004_),
    .ZN(_05005_)
  );
  AND2_X1 _25219_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_05005_),
    .ZN(_05006_)
  );
  AND2_X1 _25220_ (
    .A1(_05003_),
    .A2(_05006_),
    .ZN(_05007_)
  );
  INV_X1 _25221_ (
    .A(_05007_),
    .ZN(_05008_)
  );
  MUX2_X1 _25222_ (
    .A(\rf[15] [30]),
    .B(\rf[11] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_05009_)
  );
  AND2_X1 _25223_ (
    .A1(_08544_),
    .A2(_05009_),
    .ZN(_05010_)
  );
  INV_X1 _25224_ (
    .A(_05010_),
    .ZN(_05011_)
  );
  AND2_X1 _25225_ (
    .A1(_08545_),
    .A2(_05011_),
    .ZN(_05012_)
  );
  AND2_X1 _25226_ (
    .A1(_05008_),
    .A2(_05012_),
    .ZN(_05013_)
  );
  INV_X1 _25227_ (
    .A(_05013_),
    .ZN(_05014_)
  );
  AND2_X1 _25228_ (
    .A1(_08372_),
    .A2(_08546_),
    .ZN(_05015_)
  );
  INV_X1 _25229_ (
    .A(_05015_),
    .ZN(_05016_)
  );
  AND2_X1 _25230_ (
    .A1(_08273_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_05017_)
  );
  INV_X1 _25231_ (
    .A(_05017_),
    .ZN(_05018_)
  );
  AND2_X1 _25232_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_05018_),
    .ZN(_05019_)
  );
  AND2_X1 _25233_ (
    .A1(_05016_),
    .A2(_05019_),
    .ZN(_05020_)
  );
  INV_X1 _25234_ (
    .A(_05020_),
    .ZN(_05021_)
  );
  MUX2_X1 _25235_ (
    .A(\rf[13] [30]),
    .B(\rf[9] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_05022_)
  );
  AND2_X1 _25236_ (
    .A1(_08544_),
    .A2(_05022_),
    .ZN(_05023_)
  );
  INV_X1 _25237_ (
    .A(_05023_),
    .ZN(_05024_)
  );
  AND2_X1 _25238_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_05024_),
    .ZN(_05025_)
  );
  AND2_X1 _25239_ (
    .A1(_05021_),
    .A2(_05025_),
    .ZN(_05026_)
  );
  INV_X1 _25240_ (
    .A(_05026_),
    .ZN(_05027_)
  );
  AND2_X1 _25241_ (
    .A1(_08547_),
    .A2(_05027_),
    .ZN(_05028_)
  );
  AND2_X1 _25242_ (
    .A1(_05014_),
    .A2(_05028_),
    .ZN(_05029_)
  );
  INV_X1 _25243_ (
    .A(_05029_),
    .ZN(_05030_)
  );
  MUX2_X1 _25244_ (
    .A(\rf[6] [30]),
    .B(\rf[2] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_05031_)
  );
  AND2_X1 _25245_ (
    .A1(_08545_),
    .A2(_05031_),
    .ZN(_05032_)
  );
  INV_X1 _25246_ (
    .A(_05032_),
    .ZN(_05033_)
  );
  MUX2_X1 _25247_ (
    .A(\rf[4] [30]),
    .B(\rf[0] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_05034_)
  );
  AND2_X1 _25248_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_05034_),
    .ZN(_05035_)
  );
  INV_X1 _25249_ (
    .A(_05035_),
    .ZN(_05036_)
  );
  AND2_X1 _25250_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_05036_),
    .ZN(_05037_)
  );
  AND2_X1 _25251_ (
    .A1(_05033_),
    .A2(_05037_),
    .ZN(_05038_)
  );
  INV_X1 _25252_ (
    .A(_05038_),
    .ZN(_05039_)
  );
  MUX2_X1 _25253_ (
    .A(\rf[7] [30]),
    .B(\rf[3] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_05040_)
  );
  AND2_X1 _25254_ (
    .A1(_08545_),
    .A2(_05040_),
    .ZN(_05041_)
  );
  INV_X1 _25255_ (
    .A(_05041_),
    .ZN(_05042_)
  );
  MUX2_X1 _25256_ (
    .A(\rf[5] [30]),
    .B(\rf[1] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_05043_)
  );
  AND2_X1 _25257_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_05043_),
    .ZN(_05044_)
  );
  INV_X1 _25258_ (
    .A(_05044_),
    .ZN(_05045_)
  );
  AND2_X1 _25259_ (
    .A1(_08544_),
    .A2(_05045_),
    .ZN(_05046_)
  );
  AND2_X1 _25260_ (
    .A1(_05042_),
    .A2(_05046_),
    .ZN(_05047_)
  );
  INV_X1 _25261_ (
    .A(_05047_),
    .ZN(_05048_)
  );
  AND2_X1 _25262_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_05048_),
    .ZN(_05049_)
  );
  AND2_X1 _25263_ (
    .A1(_05039_),
    .A2(_05049_),
    .ZN(_05050_)
  );
  INV_X1 _25264_ (
    .A(_05050_),
    .ZN(_05051_)
  );
  AND2_X1 _25265_ (
    .A1(_05030_),
    .A2(_05051_),
    .ZN(_05052_)
  );
  AND2_X1 _25266_ (
    .A1(_08334_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_05053_)
  );
  INV_X1 _25267_ (
    .A(_05053_),
    .ZN(_05054_)
  );
  AND2_X1 _25268_ (
    .A1(_08433_),
    .A2(_08546_),
    .ZN(_05055_)
  );
  INV_X1 _25269_ (
    .A(_05055_),
    .ZN(_05056_)
  );
  AND2_X1 _25270_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_05056_),
    .ZN(_05057_)
  );
  AND2_X1 _25271_ (
    .A1(_05054_),
    .A2(_05057_),
    .ZN(_05058_)
  );
  INV_X1 _25272_ (
    .A(_05058_),
    .ZN(_05059_)
  );
  MUX2_X1 _25273_ (
    .A(\rf[23] [30]),
    .B(\rf[19] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_05060_)
  );
  AND2_X1 _25274_ (
    .A1(_08545_),
    .A2(_05060_),
    .ZN(_05061_)
  );
  INV_X1 _25275_ (
    .A(_05061_),
    .ZN(_05062_)
  );
  AND2_X1 _25276_ (
    .A1(_08544_),
    .A2(_05062_),
    .ZN(_05063_)
  );
  AND2_X1 _25277_ (
    .A1(_05059_),
    .A2(_05063_),
    .ZN(_05064_)
  );
  INV_X1 _25278_ (
    .A(_05064_),
    .ZN(_05065_)
  );
  AND2_X1 _25279_ (
    .A1(_08403_),
    .A2(_08546_),
    .ZN(_05066_)
  );
  INV_X1 _25280_ (
    .A(_05066_),
    .ZN(_05067_)
  );
  AND2_X1 _25281_ (
    .A1(_08304_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_05068_)
  );
  INV_X1 _25282_ (
    .A(_05068_),
    .ZN(_05069_)
  );
  AND2_X1 _25283_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_05069_),
    .ZN(_05070_)
  );
  AND2_X1 _25284_ (
    .A1(_05067_),
    .A2(_05070_),
    .ZN(_05071_)
  );
  INV_X1 _25285_ (
    .A(_05071_),
    .ZN(_05072_)
  );
  MUX2_X1 _25286_ (
    .A(\rf[22] [30]),
    .B(\rf[18] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_05073_)
  );
  AND2_X1 _25287_ (
    .A1(_08545_),
    .A2(_05073_),
    .ZN(_05074_)
  );
  INV_X1 _25288_ (
    .A(_05074_),
    .ZN(_05075_)
  );
  AND2_X1 _25289_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_05075_),
    .ZN(_05076_)
  );
  AND2_X1 _25290_ (
    .A1(_05072_),
    .A2(_05076_),
    .ZN(_05077_)
  );
  INV_X1 _25291_ (
    .A(_05077_),
    .ZN(_05078_)
  );
  AND2_X1 _25292_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_05065_),
    .ZN(_05079_)
  );
  AND2_X1 _25293_ (
    .A1(_05078_),
    .A2(_05079_),
    .ZN(_05080_)
  );
  INV_X1 _25294_ (
    .A(_05080_),
    .ZN(_05081_)
  );
  AND2_X1 _25295_ (
    .A1(_08458_),
    .A2(_08546_),
    .ZN(_05082_)
  );
  INV_X1 _25296_ (
    .A(_05082_),
    .ZN(_05083_)
  );
  AND2_X1 _25297_ (
    .A1(_08528_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_05084_)
  );
  INV_X1 _25298_ (
    .A(_05084_),
    .ZN(_05085_)
  );
  AND2_X1 _25299_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_05085_),
    .ZN(_05086_)
  );
  AND2_X1 _25300_ (
    .A1(_05083_),
    .A2(_05086_),
    .ZN(_05087_)
  );
  INV_X1 _25301_ (
    .A(_05087_),
    .ZN(_05088_)
  );
  MUX2_X1 _25302_ (
    .A(\rf[30] [30]),
    .B(\rf[26] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_05089_)
  );
  AND2_X1 _25303_ (
    .A1(_08545_),
    .A2(_05089_),
    .ZN(_05090_)
  );
  INV_X1 _25304_ (
    .A(_05090_),
    .ZN(_05091_)
  );
  AND2_X1 _25305_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_05091_),
    .ZN(_05092_)
  );
  AND2_X1 _25306_ (
    .A1(_05088_),
    .A2(_05092_),
    .ZN(_05093_)
  );
  INV_X1 _25307_ (
    .A(_05093_),
    .ZN(_05094_)
  );
  MUX2_X1 _25308_ (
    .A(\rf[29] [30]),
    .B(\rf[25] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_05095_)
  );
  AND2_X1 _25309_ (
    .A1(\rf[27] [30]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_05096_)
  );
  MUX2_X1 _25310_ (
    .A(_05095_),
    .B(_05096_),
    .S(_08545_),
    .Z(_05097_)
  );
  INV_X1 _25311_ (
    .A(_05097_),
    .ZN(_05098_)
  );
  AND2_X1 _25312_ (
    .A1(_08544_),
    .A2(_05098_),
    .ZN(_05099_)
  );
  INV_X1 _25313_ (
    .A(_05099_),
    .ZN(_05100_)
  );
  AND2_X1 _25314_ (
    .A1(_08547_),
    .A2(_05100_),
    .ZN(_05101_)
  );
  AND2_X1 _25315_ (
    .A1(_05094_),
    .A2(_05101_),
    .ZN(_05102_)
  );
  INV_X1 _25316_ (
    .A(_05102_),
    .ZN(_05103_)
  );
  AND2_X1 _25317_ (
    .A1(_05081_),
    .A2(_05103_),
    .ZN(_05104_)
  );
  MUX2_X1 _25318_ (
    .A(_05052_),
    .B(_05104_),
    .S(_08572_),
    .Z(_05105_)
  );
  INV_X1 _25319_ (
    .A(_05105_),
    .ZN(_05106_)
  );
  MUX2_X1 _25320_ (
    .A(_05106_),
    .B(_13349_),
    .S(_02233_),
    .Z(_05107_)
  );
  MUX2_X1 _25321_ (
    .A(ex_reg_rs_msb_1[28]),
    .B(_05107_),
    .S(_02202_),
    .Z(_00177_)
  );
  AND2_X1 _25322_ (
    .A1(_08235_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_05108_)
  );
  INV_X1 _25323_ (
    .A(_05108_),
    .ZN(_05109_)
  );
  AND2_X1 _25324_ (
    .A1(_08233_),
    .A2(_08546_),
    .ZN(_05110_)
  );
  INV_X1 _25325_ (
    .A(_05110_),
    .ZN(_05111_)
  );
  AND2_X1 _25326_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_05111_),
    .ZN(_05112_)
  );
  AND2_X1 _25327_ (
    .A1(_05109_),
    .A2(_05112_),
    .ZN(_05113_)
  );
  INV_X1 _25328_ (
    .A(_05113_),
    .ZN(_05114_)
  );
  MUX2_X1 _25329_ (
    .A(\rf[15] [31]),
    .B(\rf[11] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_05115_)
  );
  AND2_X1 _25330_ (
    .A1(_08544_),
    .A2(_05115_),
    .ZN(_05116_)
  );
  INV_X1 _25331_ (
    .A(_05116_),
    .ZN(_05117_)
  );
  AND2_X1 _25332_ (
    .A1(_08545_),
    .A2(_05117_),
    .ZN(_05118_)
  );
  AND2_X1 _25333_ (
    .A1(_05114_),
    .A2(_05118_),
    .ZN(_05119_)
  );
  INV_X1 _25334_ (
    .A(_05119_),
    .ZN(_05120_)
  );
  AND2_X1 _25335_ (
    .A1(_08234_),
    .A2(_08546_),
    .ZN(_05121_)
  );
  INV_X1 _25336_ (
    .A(_05121_),
    .ZN(_05122_)
  );
  AND2_X1 _25337_ (
    .A1(_08226_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_05123_)
  );
  INV_X1 _25338_ (
    .A(_05123_),
    .ZN(_05124_)
  );
  AND2_X1 _25339_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_05124_),
    .ZN(_05125_)
  );
  AND2_X1 _25340_ (
    .A1(_05122_),
    .A2(_05125_),
    .ZN(_05126_)
  );
  INV_X1 _25341_ (
    .A(_05126_),
    .ZN(_05127_)
  );
  MUX2_X1 _25342_ (
    .A(\rf[13] [31]),
    .B(\rf[9] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_05128_)
  );
  AND2_X1 _25343_ (
    .A1(_08544_),
    .A2(_05128_),
    .ZN(_05129_)
  );
  INV_X1 _25344_ (
    .A(_05129_),
    .ZN(_05130_)
  );
  AND2_X1 _25345_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_05130_),
    .ZN(_05131_)
  );
  AND2_X1 _25346_ (
    .A1(_05127_),
    .A2(_05131_),
    .ZN(_05132_)
  );
  INV_X1 _25347_ (
    .A(_05132_),
    .ZN(_05133_)
  );
  AND2_X1 _25348_ (
    .A1(_08547_),
    .A2(_05133_),
    .ZN(_05134_)
  );
  AND2_X1 _25349_ (
    .A1(_05120_),
    .A2(_05134_),
    .ZN(_05135_)
  );
  INV_X1 _25350_ (
    .A(_05135_),
    .ZN(_05136_)
  );
  MUX2_X1 _25351_ (
    .A(\rf[6] [31]),
    .B(\rf[2] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_05137_)
  );
  AND2_X1 _25352_ (
    .A1(_08545_),
    .A2(_05137_),
    .ZN(_05138_)
  );
  INV_X1 _25353_ (
    .A(_05138_),
    .ZN(_05139_)
  );
  MUX2_X1 _25354_ (
    .A(\rf[4] [31]),
    .B(\rf[0] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_05140_)
  );
  AND2_X1 _25355_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_05140_),
    .ZN(_05141_)
  );
  INV_X1 _25356_ (
    .A(_05141_),
    .ZN(_05142_)
  );
  AND2_X1 _25357_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_05142_),
    .ZN(_05143_)
  );
  AND2_X1 _25358_ (
    .A1(_05139_),
    .A2(_05143_),
    .ZN(_05144_)
  );
  INV_X1 _25359_ (
    .A(_05144_),
    .ZN(_05145_)
  );
  MUX2_X1 _25360_ (
    .A(\rf[7] [31]),
    .B(\rf[3] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_05146_)
  );
  AND2_X1 _25361_ (
    .A1(_08545_),
    .A2(_05146_),
    .ZN(_05147_)
  );
  INV_X1 _25362_ (
    .A(_05147_),
    .ZN(_05148_)
  );
  MUX2_X1 _25363_ (
    .A(\rf[5] [31]),
    .B(\rf[1] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_05149_)
  );
  AND2_X1 _25364_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_05149_),
    .ZN(_05150_)
  );
  INV_X1 _25365_ (
    .A(_05150_),
    .ZN(_05151_)
  );
  AND2_X1 _25366_ (
    .A1(_08544_),
    .A2(_05151_),
    .ZN(_05152_)
  );
  AND2_X1 _25367_ (
    .A1(_05148_),
    .A2(_05152_),
    .ZN(_05153_)
  );
  INV_X1 _25368_ (
    .A(_05153_),
    .ZN(_05154_)
  );
  AND2_X1 _25369_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_05154_),
    .ZN(_05155_)
  );
  AND2_X1 _25370_ (
    .A1(_05145_),
    .A2(_05155_),
    .ZN(_05156_)
  );
  INV_X1 _25371_ (
    .A(_05156_),
    .ZN(_05157_)
  );
  AND2_X1 _25372_ (
    .A1(_05136_),
    .A2(_05157_),
    .ZN(_05158_)
  );
  AND2_X1 _25373_ (
    .A1(_08231_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_05159_)
  );
  INV_X1 _25374_ (
    .A(_05159_),
    .ZN(_05160_)
  );
  AND2_X1 _25375_ (
    .A1(_08229_),
    .A2(_08546_),
    .ZN(_05161_)
  );
  INV_X1 _25376_ (
    .A(_05161_),
    .ZN(_05162_)
  );
  AND2_X1 _25377_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_05162_),
    .ZN(_05163_)
  );
  AND2_X1 _25378_ (
    .A1(_05160_),
    .A2(_05163_),
    .ZN(_05164_)
  );
  INV_X1 _25379_ (
    .A(_05164_),
    .ZN(_05165_)
  );
  MUX2_X1 _25380_ (
    .A(\rf[23] [31]),
    .B(\rf[19] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_05166_)
  );
  AND2_X1 _25381_ (
    .A1(_08545_),
    .A2(_05166_),
    .ZN(_05167_)
  );
  INV_X1 _25382_ (
    .A(_05167_),
    .ZN(_05168_)
  );
  AND2_X1 _25383_ (
    .A1(_08544_),
    .A2(_05168_),
    .ZN(_05169_)
  );
  AND2_X1 _25384_ (
    .A1(_05165_),
    .A2(_05169_),
    .ZN(_05170_)
  );
  INV_X1 _25385_ (
    .A(_05170_),
    .ZN(_05171_)
  );
  AND2_X1 _25386_ (
    .A1(_08230_),
    .A2(_08546_),
    .ZN(_05172_)
  );
  INV_X1 _25387_ (
    .A(_05172_),
    .ZN(_05173_)
  );
  AND2_X1 _25388_ (
    .A1(_08232_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_05174_)
  );
  INV_X1 _25389_ (
    .A(_05174_),
    .ZN(_05175_)
  );
  AND2_X1 _25390_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_05175_),
    .ZN(_05176_)
  );
  AND2_X1 _25391_ (
    .A1(_05173_),
    .A2(_05176_),
    .ZN(_05177_)
  );
  INV_X1 _25392_ (
    .A(_05177_),
    .ZN(_05178_)
  );
  MUX2_X1 _25393_ (
    .A(\rf[22] [31]),
    .B(\rf[18] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_05179_)
  );
  AND2_X1 _25394_ (
    .A1(_08545_),
    .A2(_05179_),
    .ZN(_05180_)
  );
  INV_X1 _25395_ (
    .A(_05180_),
    .ZN(_05181_)
  );
  AND2_X1 _25396_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_05181_),
    .ZN(_05182_)
  );
  AND2_X1 _25397_ (
    .A1(_05178_),
    .A2(_05182_),
    .ZN(_05183_)
  );
  INV_X1 _25398_ (
    .A(_05183_),
    .ZN(_05184_)
  );
  AND2_X1 _25399_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_05171_),
    .ZN(_05185_)
  );
  AND2_X1 _25400_ (
    .A1(_05184_),
    .A2(_05185_),
    .ZN(_05186_)
  );
  INV_X1 _25401_ (
    .A(_05186_),
    .ZN(_05187_)
  );
  AND2_X1 _25402_ (
    .A1(_08227_),
    .A2(_08546_),
    .ZN(_05188_)
  );
  INV_X1 _25403_ (
    .A(_05188_),
    .ZN(_05189_)
  );
  AND2_X1 _25404_ (
    .A1(_08228_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_05190_)
  );
  INV_X1 _25405_ (
    .A(_05190_),
    .ZN(_05191_)
  );
  AND2_X1 _25406_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_05191_),
    .ZN(_05192_)
  );
  AND2_X1 _25407_ (
    .A1(_05189_),
    .A2(_05192_),
    .ZN(_05193_)
  );
  INV_X1 _25408_ (
    .A(_05193_),
    .ZN(_05194_)
  );
  MUX2_X1 _25409_ (
    .A(\rf[30] [31]),
    .B(\rf[26] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_05195_)
  );
  AND2_X1 _25410_ (
    .A1(_08545_),
    .A2(_05195_),
    .ZN(_05196_)
  );
  INV_X1 _25411_ (
    .A(_05196_),
    .ZN(_05197_)
  );
  AND2_X1 _25412_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_05197_),
    .ZN(_05198_)
  );
  AND2_X1 _25413_ (
    .A1(_05194_),
    .A2(_05198_),
    .ZN(_05199_)
  );
  INV_X1 _25414_ (
    .A(_05199_),
    .ZN(_05200_)
  );
  MUX2_X1 _25415_ (
    .A(\rf[29] [31]),
    .B(\rf[25] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_05201_)
  );
  AND2_X1 _25416_ (
    .A1(\rf[27] [31]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_05202_)
  );
  MUX2_X1 _25417_ (
    .A(_05201_),
    .B(_05202_),
    .S(_08545_),
    .Z(_05203_)
  );
  INV_X1 _25418_ (
    .A(_05203_),
    .ZN(_05204_)
  );
  AND2_X1 _25419_ (
    .A1(_08544_),
    .A2(_05204_),
    .ZN(_05205_)
  );
  INV_X1 _25420_ (
    .A(_05205_),
    .ZN(_05206_)
  );
  AND2_X1 _25421_ (
    .A1(_08547_),
    .A2(_05206_),
    .ZN(_05207_)
  );
  AND2_X1 _25422_ (
    .A1(_05200_),
    .A2(_05207_),
    .ZN(_05208_)
  );
  INV_X1 _25423_ (
    .A(_05208_),
    .ZN(_05209_)
  );
  AND2_X1 _25424_ (
    .A1(_05187_),
    .A2(_05209_),
    .ZN(_05210_)
  );
  MUX2_X1 _25425_ (
    .A(_05158_),
    .B(_05210_),
    .S(_08572_),
    .Z(_05211_)
  );
  INV_X1 _25426_ (
    .A(_05211_),
    .ZN(_05212_)
  );
  MUX2_X1 _25427_ (
    .A(_05212_),
    .B(_13465_),
    .S(_02233_),
    .Z(_05213_)
  );
  MUX2_X1 _25428_ (
    .A(ex_reg_rs_msb_1[29]),
    .B(_05213_),
    .S(_02202_),
    .Z(_00178_)
  );
  AND2_X1 _25429_ (
    .A1(_08564_),
    .A2(_08565_),
    .ZN(_05214_)
  );
  AND2_X1 _25430_ (
    .A1(_08566_),
    .A2(_05214_),
    .ZN(_05215_)
  );
  AND2_X1 _25431_ (
    .A1(_08578_),
    .A2(_05215_),
    .ZN(_05216_)
  );
  INV_X1 _25432_ (
    .A(_05216_),
    .ZN(_05217_)
  );
  MUX2_X1 _25433_ (
    .A(ex_reg_rvc),
    .B(_05217_),
    .S(_10244_),
    .Z(_00179_)
  );
  AND2_X1 _25434_ (
    .A1(_08596_),
    .A2(_08624_),
    .ZN(_05218_)
  );
  INV_X1 _25435_ (
    .A(_05218_),
    .ZN(_05219_)
  );
  AND2_X1 _25436_ (
    .A1(mem_reg_cause[4]),
    .A2(_05219_),
    .ZN(_05220_)
  );
  MUX2_X1 _25437_ (
    .A(wb_reg_cause[4]),
    .B(_05220_),
    .S(_13834_),
    .Z(_00180_)
  );
  AND2_X1 _25438_ (
    .A1(mem_reg_cause[5]),
    .A2(_05219_),
    .ZN(_05221_)
  );
  MUX2_X1 _25439_ (
    .A(wb_reg_cause[5]),
    .B(_05221_),
    .S(_13834_),
    .Z(_00181_)
  );
  AND2_X1 _25440_ (
    .A1(mem_reg_cause[6]),
    .A2(_05219_),
    .ZN(_05222_)
  );
  MUX2_X1 _25441_ (
    .A(wb_reg_cause[6]),
    .B(_05222_),
    .S(_13834_),
    .Z(_00182_)
  );
  AND2_X1 _25442_ (
    .A1(mem_reg_cause[7]),
    .A2(_05219_),
    .ZN(_05223_)
  );
  MUX2_X1 _25443_ (
    .A(wb_reg_cause[7]),
    .B(_05223_),
    .S(_13834_),
    .Z(_00183_)
  );
  AND2_X1 _25444_ (
    .A1(mem_reg_cause[8]),
    .A2(_05219_),
    .ZN(_05224_)
  );
  MUX2_X1 _25445_ (
    .A(wb_reg_cause[8]),
    .B(_05224_),
    .S(_13834_),
    .Z(_00184_)
  );
  AND2_X1 _25446_ (
    .A1(mem_reg_cause[9]),
    .A2(_05219_),
    .ZN(_05225_)
  );
  MUX2_X1 _25447_ (
    .A(wb_reg_cause[9]),
    .B(_05225_),
    .S(_13834_),
    .Z(_00185_)
  );
  AND2_X1 _25448_ (
    .A1(mem_reg_cause[10]),
    .A2(_05219_),
    .ZN(_05226_)
  );
  MUX2_X1 _25449_ (
    .A(wb_reg_cause[10]),
    .B(_05226_),
    .S(_13834_),
    .Z(_00186_)
  );
  AND2_X1 _25450_ (
    .A1(mem_reg_cause[11]),
    .A2(_05219_),
    .ZN(_05227_)
  );
  MUX2_X1 _25451_ (
    .A(wb_reg_cause[11]),
    .B(_05227_),
    .S(_13834_),
    .Z(_00187_)
  );
  AND2_X1 _25452_ (
    .A1(mem_reg_cause[12]),
    .A2(_05219_),
    .ZN(_05228_)
  );
  MUX2_X1 _25453_ (
    .A(wb_reg_cause[12]),
    .B(_05228_),
    .S(_13834_),
    .Z(_00188_)
  );
  AND2_X1 _25454_ (
    .A1(mem_reg_cause[13]),
    .A2(_05219_),
    .ZN(_05229_)
  );
  MUX2_X1 _25455_ (
    .A(wb_reg_cause[13]),
    .B(_05229_),
    .S(_13834_),
    .Z(_00189_)
  );
  AND2_X1 _25456_ (
    .A1(mem_reg_cause[14]),
    .A2(_05219_),
    .ZN(_05230_)
  );
  MUX2_X1 _25457_ (
    .A(wb_reg_cause[14]),
    .B(_05230_),
    .S(_13834_),
    .Z(_00190_)
  );
  AND2_X1 _25458_ (
    .A1(mem_reg_cause[15]),
    .A2(_05219_),
    .ZN(_05231_)
  );
  MUX2_X1 _25459_ (
    .A(wb_reg_cause[15]),
    .B(_05231_),
    .S(_13834_),
    .Z(_00191_)
  );
  AND2_X1 _25460_ (
    .A1(mem_reg_cause[16]),
    .A2(_05219_),
    .ZN(_05232_)
  );
  MUX2_X1 _25461_ (
    .A(wb_reg_cause[16]),
    .B(_05232_),
    .S(_13834_),
    .Z(_00192_)
  );
  AND2_X1 _25462_ (
    .A1(mem_reg_cause[17]),
    .A2(_05219_),
    .ZN(_05233_)
  );
  MUX2_X1 _25463_ (
    .A(wb_reg_cause[17]),
    .B(_05233_),
    .S(_13834_),
    .Z(_00193_)
  );
  AND2_X1 _25464_ (
    .A1(mem_reg_cause[18]),
    .A2(_05219_),
    .ZN(_05234_)
  );
  MUX2_X1 _25465_ (
    .A(wb_reg_cause[18]),
    .B(_05234_),
    .S(_13834_),
    .Z(_00194_)
  );
  AND2_X1 _25466_ (
    .A1(mem_reg_cause[19]),
    .A2(_05219_),
    .ZN(_05235_)
  );
  MUX2_X1 _25467_ (
    .A(wb_reg_cause[19]),
    .B(_05235_),
    .S(_13834_),
    .Z(_00195_)
  );
  AND2_X1 _25468_ (
    .A1(mem_reg_cause[20]),
    .A2(_05219_),
    .ZN(_05236_)
  );
  MUX2_X1 _25469_ (
    .A(wb_reg_cause[20]),
    .B(_05236_),
    .S(_13834_),
    .Z(_00196_)
  );
  AND2_X1 _25470_ (
    .A1(mem_reg_cause[21]),
    .A2(_05219_),
    .ZN(_05237_)
  );
  MUX2_X1 _25471_ (
    .A(wb_reg_cause[21]),
    .B(_05237_),
    .S(_13834_),
    .Z(_00197_)
  );
  AND2_X1 _25472_ (
    .A1(mem_reg_cause[22]),
    .A2(_05219_),
    .ZN(_05238_)
  );
  MUX2_X1 _25473_ (
    .A(wb_reg_cause[22]),
    .B(_05238_),
    .S(_13834_),
    .Z(_00198_)
  );
  AND2_X1 _25474_ (
    .A1(mem_reg_cause[23]),
    .A2(_05219_),
    .ZN(_05239_)
  );
  MUX2_X1 _25475_ (
    .A(wb_reg_cause[23]),
    .B(_05239_),
    .S(_13834_),
    .Z(_00199_)
  );
  AND2_X1 _25476_ (
    .A1(mem_reg_cause[24]),
    .A2(_05219_),
    .ZN(_05240_)
  );
  MUX2_X1 _25477_ (
    .A(wb_reg_cause[24]),
    .B(_05240_),
    .S(_13834_),
    .Z(_00200_)
  );
  AND2_X1 _25478_ (
    .A1(mem_reg_cause[25]),
    .A2(_05219_),
    .ZN(_05241_)
  );
  MUX2_X1 _25479_ (
    .A(wb_reg_cause[25]),
    .B(_05241_),
    .S(_13834_),
    .Z(_00201_)
  );
  AND2_X1 _25480_ (
    .A1(mem_reg_cause[26]),
    .A2(_05219_),
    .ZN(_05242_)
  );
  MUX2_X1 _25481_ (
    .A(wb_reg_cause[26]),
    .B(_05242_),
    .S(_13834_),
    .Z(_00202_)
  );
  AND2_X1 _25482_ (
    .A1(mem_reg_cause[27]),
    .A2(_05219_),
    .ZN(_05243_)
  );
  MUX2_X1 _25483_ (
    .A(wb_reg_cause[27]),
    .B(_05243_),
    .S(_13834_),
    .Z(_00203_)
  );
  AND2_X1 _25484_ (
    .A1(mem_reg_cause[28]),
    .A2(_05219_),
    .ZN(_05244_)
  );
  MUX2_X1 _25485_ (
    .A(wb_reg_cause[28]),
    .B(_05244_),
    .S(_13834_),
    .Z(_00204_)
  );
  AND2_X1 _25486_ (
    .A1(mem_reg_cause[29]),
    .A2(_05219_),
    .ZN(_05245_)
  );
  MUX2_X1 _25487_ (
    .A(wb_reg_cause[29]),
    .B(_05245_),
    .S(_13834_),
    .Z(_00205_)
  );
  AND2_X1 _25488_ (
    .A1(mem_reg_cause[30]),
    .A2(_05219_),
    .ZN(_05246_)
  );
  MUX2_X1 _25489_ (
    .A(wb_reg_cause[30]),
    .B(_05246_),
    .S(_13834_),
    .Z(_00206_)
  );
  AND2_X1 _25490_ (
    .A1(mem_reg_cause[31]),
    .A2(_05219_),
    .ZN(_05247_)
  );
  MUX2_X1 _25491_ (
    .A(wb_reg_cause[31]),
    .B(_05247_),
    .S(_13834_),
    .Z(_00207_)
  );
  MUX2_X1 _25492_ (
    .A(mem_reg_pc[0]),
    .B(wb_reg_pc[0]),
    .S(_13833_),
    .Z(_00208_)
  );
  MUX2_X1 _25493_ (
    .A(mem_reg_pc[1]),
    .B(wb_reg_pc[1]),
    .S(_13833_),
    .Z(_00209_)
  );
  MUX2_X1 _25494_ (
    .A(mem_reg_pc[2]),
    .B(wb_reg_pc[2]),
    .S(_13833_),
    .Z(_00210_)
  );
  MUX2_X1 _25495_ (
    .A(mem_reg_pc[3]),
    .B(wb_reg_pc[3]),
    .S(_13833_),
    .Z(_00211_)
  );
  MUX2_X1 _25496_ (
    .A(mem_reg_pc[4]),
    .B(wb_reg_pc[4]),
    .S(_13833_),
    .Z(_00212_)
  );
  MUX2_X1 _25497_ (
    .A(mem_reg_pc[5]),
    .B(wb_reg_pc[5]),
    .S(_13833_),
    .Z(_00213_)
  );
  MUX2_X1 _25498_ (
    .A(mem_reg_pc[6]),
    .B(wb_reg_pc[6]),
    .S(_13833_),
    .Z(_00214_)
  );
  MUX2_X1 _25499_ (
    .A(mem_reg_pc[7]),
    .B(wb_reg_pc[7]),
    .S(_13833_),
    .Z(_00215_)
  );
  MUX2_X1 _25500_ (
    .A(mem_reg_pc[8]),
    .B(wb_reg_pc[8]),
    .S(_13833_),
    .Z(_00216_)
  );
  MUX2_X1 _25501_ (
    .A(mem_reg_pc[9]),
    .B(wb_reg_pc[9]),
    .S(_13833_),
    .Z(_00217_)
  );
  MUX2_X1 _25502_ (
    .A(mem_reg_pc[10]),
    .B(wb_reg_pc[10]),
    .S(_13833_),
    .Z(_00218_)
  );
  MUX2_X1 _25503_ (
    .A(mem_reg_pc[11]),
    .B(wb_reg_pc[11]),
    .S(_13833_),
    .Z(_00219_)
  );
  MUX2_X1 _25504_ (
    .A(mem_reg_pc[12]),
    .B(wb_reg_pc[12]),
    .S(_13833_),
    .Z(_00220_)
  );
  MUX2_X1 _25505_ (
    .A(mem_reg_pc[13]),
    .B(wb_reg_pc[13]),
    .S(_13833_),
    .Z(_00221_)
  );
  MUX2_X1 _25506_ (
    .A(mem_reg_pc[14]),
    .B(wb_reg_pc[14]),
    .S(_13833_),
    .Z(_00222_)
  );
  MUX2_X1 _25507_ (
    .A(mem_reg_pc[15]),
    .B(wb_reg_pc[15]),
    .S(_13833_),
    .Z(_00223_)
  );
  MUX2_X1 _25508_ (
    .A(mem_reg_pc[16]),
    .B(wb_reg_pc[16]),
    .S(_13833_),
    .Z(_00224_)
  );
  MUX2_X1 _25509_ (
    .A(mem_reg_pc[17]),
    .B(wb_reg_pc[17]),
    .S(_13833_),
    .Z(_00225_)
  );
  MUX2_X1 _25510_ (
    .A(mem_reg_pc[18]),
    .B(wb_reg_pc[18]),
    .S(_13833_),
    .Z(_00226_)
  );
  MUX2_X1 _25511_ (
    .A(mem_reg_pc[19]),
    .B(wb_reg_pc[19]),
    .S(_13833_),
    .Z(_00227_)
  );
  MUX2_X1 _25512_ (
    .A(mem_reg_pc[20]),
    .B(wb_reg_pc[20]),
    .S(_13833_),
    .Z(_00228_)
  );
  MUX2_X1 _25513_ (
    .A(mem_reg_pc[21]),
    .B(wb_reg_pc[21]),
    .S(_13833_),
    .Z(_00229_)
  );
  MUX2_X1 _25514_ (
    .A(mem_reg_pc[22]),
    .B(wb_reg_pc[22]),
    .S(_13833_),
    .Z(_00230_)
  );
  MUX2_X1 _25515_ (
    .A(mem_reg_pc[23]),
    .B(wb_reg_pc[23]),
    .S(_13833_),
    .Z(_00231_)
  );
  MUX2_X1 _25516_ (
    .A(mem_reg_pc[24]),
    .B(wb_reg_pc[24]),
    .S(_13833_),
    .Z(_00232_)
  );
  MUX2_X1 _25517_ (
    .A(mem_reg_pc[25]),
    .B(wb_reg_pc[25]),
    .S(_13833_),
    .Z(_00233_)
  );
  MUX2_X1 _25518_ (
    .A(mem_reg_pc[26]),
    .B(wb_reg_pc[26]),
    .S(_13833_),
    .Z(_00234_)
  );
  MUX2_X1 _25519_ (
    .A(mem_reg_pc[27]),
    .B(wb_reg_pc[27]),
    .S(_13833_),
    .Z(_00235_)
  );
  MUX2_X1 _25520_ (
    .A(mem_reg_pc[28]),
    .B(wb_reg_pc[28]),
    .S(_13833_),
    .Z(_00236_)
  );
  MUX2_X1 _25521_ (
    .A(mem_reg_pc[29]),
    .B(wb_reg_pc[29]),
    .S(_13833_),
    .Z(_00237_)
  );
  MUX2_X1 _25522_ (
    .A(mem_reg_pc[30]),
    .B(wb_reg_pc[30]),
    .S(_13833_),
    .Z(_00238_)
  );
  MUX2_X1 _25523_ (
    .A(mem_reg_pc[31]),
    .B(wb_reg_pc[31]),
    .S(_13833_),
    .Z(_00239_)
  );
  AND2_X1 _25524_ (
    .A1(_08606_),
    .A2(_08618_),
    .ZN(_05248_)
  );
  AND2_X1 _25525_ (
    .A1(_08619_),
    .A2(_05248_),
    .ZN(_05249_)
  );
  INV_X1 _25526_ (
    .A(_05249_),
    .ZN(_05250_)
  );
  AND2_X1 _25527_ (
    .A1(mem_reg_flush_pipe),
    .A2(mem_reg_valid),
    .ZN(_05251_)
  );
  INV_X1 _25528_ (
    .A(_05251_),
    .ZN(_05252_)
  );
  AND2_X1 _25529_ (
    .A1(_05250_),
    .A2(_05252_),
    .ZN(_05253_)
  );
  INV_X1 _25530_ (
    .A(_05253_),
    .ZN(_05254_)
  );
  MUX2_X1 _25531_ (
    .A(mem_br_taken),
    .B(alu_io_cmp_out),
    .S(_05253_),
    .Z(_00240_)
  );
  AND2_X1 _25532_ (
    .A1(_08569_),
    .A2(_08570_),
    .ZN(_05255_)
  );
  AND2_X1 _25533_ (
    .A1(_08220_),
    .A2(_08570_),
    .ZN(_05256_)
  );
  INV_X1 _25534_ (
    .A(_05256_),
    .ZN(_05257_)
  );
  AND2_X1 _25535_ (
    .A1(_08221_),
    .A2(_08569_),
    .ZN(_05258_)
  );
  AND2_X1 _25536_ (
    .A1(_05257_),
    .A2(_05258_),
    .ZN(_05259_)
  );
  AND2_X1 _25537_ (
    .A1(mem_reg_wdata[0]),
    .A2(_05259_),
    .ZN(_05260_)
  );
  INV_X1 _25538_ (
    .A(_05260_),
    .ZN(_05261_)
  );
  AND2_X1 _25539_ (
    .A1(wb_reg_wdata[0]),
    .A2(_05256_),
    .ZN(_05262_)
  );
  INV_X1 _25540_ (
    .A(_05262_),
    .ZN(_05263_)
  );
  AND2_X1 _25541_ (
    .A1(_05261_),
    .A2(_05263_),
    .ZN(_05264_)
  );
  INV_X1 _25542_ (
    .A(_05264_),
    .ZN(_05265_)
  );
  MUX2_X1 _25543_ (
    .A(_05265_),
    .B(io_dmem_resp_bits_data_word_bypass[0]),
    .S(_05255_),
    .Z(_05266_)
  );
  MUX2_X1 _25544_ (
    .A(ex_reg_rs_lsb_1[0]),
    .B(_05266_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[0])
  );
  INV_X1 _25545_ (
    .A(_ex_op2_T[0]),
    .ZN(_05267_)
  );
  AND2_X1 _25546_ (
    .A1(ex_ctrl_mem),
    .A2(_05253_),
    .ZN(_05268_)
  );
  AND2_X1 _25547_ (
    .A1(ex_ctrl_rxs2),
    .A2(_05268_),
    .ZN(_05269_)
  );
  INV_X1 _25548_ (
    .A(_05269_),
    .ZN(_05270_)
  );
  AND2_X1 _25549_ (
    .A1(_05267_),
    .A2(_05269_),
    .ZN(_05271_)
  );
  INV_X1 _25550_ (
    .A(_05271_),
    .ZN(_05272_)
  );
  MUX2_X1 _25551_ (
    .A(mem_reg_rs2[0]),
    .B(_ex_op2_T[0]),
    .S(_05269_),
    .Z(_00241_)
  );
  AND2_X1 _25552_ (
    .A1(mem_reg_wdata[1]),
    .A2(_05259_),
    .ZN(_05273_)
  );
  INV_X1 _25553_ (
    .A(_05273_),
    .ZN(_05274_)
  );
  AND2_X1 _25554_ (
    .A1(wb_reg_wdata[1]),
    .A2(_05256_),
    .ZN(_05275_)
  );
  INV_X1 _25555_ (
    .A(_05275_),
    .ZN(_05276_)
  );
  AND2_X1 _25556_ (
    .A1(_05274_),
    .A2(_05276_),
    .ZN(_05277_)
  );
  INV_X1 _25557_ (
    .A(_05277_),
    .ZN(_05278_)
  );
  MUX2_X1 _25558_ (
    .A(_05278_),
    .B(io_dmem_resp_bits_data_word_bypass[1]),
    .S(_05255_),
    .Z(_05279_)
  );
  MUX2_X1 _25559_ (
    .A(ex_reg_rs_lsb_1[1]),
    .B(_05279_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[1])
  );
  INV_X1 _25560_ (
    .A(_ex_op2_T[1]),
    .ZN(_05280_)
  );
  AND2_X1 _25561_ (
    .A1(_05269_),
    .A2(_05280_),
    .ZN(_05281_)
  );
  INV_X1 _25562_ (
    .A(_05281_),
    .ZN(_05282_)
  );
  MUX2_X1 _25563_ (
    .A(mem_reg_rs2[1]),
    .B(_ex_op2_T[1]),
    .S(_05269_),
    .Z(_00242_)
  );
  AND2_X1 _25564_ (
    .A1(mem_reg_wdata[2]),
    .A2(_05259_),
    .ZN(_05283_)
  );
  INV_X1 _25565_ (
    .A(_05283_),
    .ZN(_05284_)
  );
  AND2_X1 _25566_ (
    .A1(wb_reg_wdata[2]),
    .A2(_05256_),
    .ZN(_05285_)
  );
  INV_X1 _25567_ (
    .A(_05285_),
    .ZN(_05286_)
  );
  AND2_X1 _25568_ (
    .A1(_05284_),
    .A2(_05286_),
    .ZN(_05287_)
  );
  INV_X1 _25569_ (
    .A(_05287_),
    .ZN(_05288_)
  );
  MUX2_X1 _25570_ (
    .A(_05288_),
    .B(io_dmem_resp_bits_data_word_bypass[2]),
    .S(_05255_),
    .Z(_05289_)
  );
  MUX2_X1 _25571_ (
    .A(ex_reg_rs_msb_1[0]),
    .B(_05289_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[2])
  );
  INV_X1 _25572_ (
    .A(_ex_op2_T[2]),
    .ZN(_05290_)
  );
  AND2_X1 _25573_ (
    .A1(_05269_),
    .A2(_05290_),
    .ZN(_05291_)
  );
  INV_X1 _25574_ (
    .A(_05291_),
    .ZN(_05292_)
  );
  MUX2_X1 _25575_ (
    .A(mem_reg_rs2[2]),
    .B(_ex_op2_T[2]),
    .S(_05269_),
    .Z(_00243_)
  );
  AND2_X1 _25576_ (
    .A1(mem_reg_wdata[3]),
    .A2(_05259_),
    .ZN(_05293_)
  );
  INV_X1 _25577_ (
    .A(_05293_),
    .ZN(_05294_)
  );
  AND2_X1 _25578_ (
    .A1(wb_reg_wdata[3]),
    .A2(_05256_),
    .ZN(_05295_)
  );
  INV_X1 _25579_ (
    .A(_05295_),
    .ZN(_05296_)
  );
  AND2_X1 _25580_ (
    .A1(_05294_),
    .A2(_05296_),
    .ZN(_05297_)
  );
  INV_X1 _25581_ (
    .A(_05297_),
    .ZN(_05298_)
  );
  MUX2_X1 _25582_ (
    .A(_05298_),
    .B(io_dmem_resp_bits_data_word_bypass[3]),
    .S(_05255_),
    .Z(_05299_)
  );
  MUX2_X1 _25583_ (
    .A(ex_reg_rs_msb_1[1]),
    .B(_05299_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[3])
  );
  INV_X1 _25584_ (
    .A(_ex_op2_T[3]),
    .ZN(_05300_)
  );
  AND2_X1 _25585_ (
    .A1(_05269_),
    .A2(_05300_),
    .ZN(_05301_)
  );
  INV_X1 _25586_ (
    .A(_05301_),
    .ZN(_05302_)
  );
  MUX2_X1 _25587_ (
    .A(mem_reg_rs2[3]),
    .B(_ex_op2_T[3]),
    .S(_05269_),
    .Z(_00244_)
  );
  AND2_X1 _25588_ (
    .A1(mem_reg_wdata[4]),
    .A2(_05259_),
    .ZN(_05303_)
  );
  INV_X1 _25589_ (
    .A(_05303_),
    .ZN(_05304_)
  );
  AND2_X1 _25590_ (
    .A1(wb_reg_wdata[4]),
    .A2(_05256_),
    .ZN(_05305_)
  );
  INV_X1 _25591_ (
    .A(_05305_),
    .ZN(_05306_)
  );
  AND2_X1 _25592_ (
    .A1(_05304_),
    .A2(_05306_),
    .ZN(_05307_)
  );
  INV_X1 _25593_ (
    .A(_05307_),
    .ZN(_05308_)
  );
  MUX2_X1 _25594_ (
    .A(_05308_),
    .B(io_dmem_resp_bits_data_word_bypass[4]),
    .S(_05255_),
    .Z(_05309_)
  );
  MUX2_X1 _25595_ (
    .A(ex_reg_rs_msb_1[2]),
    .B(_05309_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[4])
  );
  INV_X1 _25596_ (
    .A(_ex_op2_T[4]),
    .ZN(_05310_)
  );
  AND2_X1 _25597_ (
    .A1(_05269_),
    .A2(_05310_),
    .ZN(_05311_)
  );
  INV_X1 _25598_ (
    .A(_05311_),
    .ZN(_05312_)
  );
  MUX2_X1 _25599_ (
    .A(mem_reg_rs2[4]),
    .B(_ex_op2_T[4]),
    .S(_05269_),
    .Z(_00245_)
  );
  AND2_X1 _25600_ (
    .A1(mem_reg_wdata[5]),
    .A2(_05259_),
    .ZN(_05313_)
  );
  INV_X1 _25601_ (
    .A(_05313_),
    .ZN(_05314_)
  );
  AND2_X1 _25602_ (
    .A1(wb_reg_wdata[5]),
    .A2(_05256_),
    .ZN(_05315_)
  );
  INV_X1 _25603_ (
    .A(_05315_),
    .ZN(_05316_)
  );
  AND2_X1 _25604_ (
    .A1(_05314_),
    .A2(_05316_),
    .ZN(_05317_)
  );
  INV_X1 _25605_ (
    .A(_05317_),
    .ZN(_05318_)
  );
  MUX2_X1 _25606_ (
    .A(_05318_),
    .B(io_dmem_resp_bits_data_word_bypass[5]),
    .S(_05255_),
    .Z(_05319_)
  );
  MUX2_X1 _25607_ (
    .A(ex_reg_rs_msb_1[3]),
    .B(_05319_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[5])
  );
  INV_X1 _25608_ (
    .A(_ex_op2_T[5]),
    .ZN(_05320_)
  );
  AND2_X1 _25609_ (
    .A1(_05269_),
    .A2(_05320_),
    .ZN(_05321_)
  );
  INV_X1 _25610_ (
    .A(_05321_),
    .ZN(_05322_)
  );
  MUX2_X1 _25611_ (
    .A(mem_reg_rs2[5]),
    .B(_ex_op2_T[5]),
    .S(_05269_),
    .Z(_00246_)
  );
  AND2_X1 _25612_ (
    .A1(mem_reg_wdata[6]),
    .A2(_05259_),
    .ZN(_05323_)
  );
  INV_X1 _25613_ (
    .A(_05323_),
    .ZN(_05324_)
  );
  AND2_X1 _25614_ (
    .A1(wb_reg_wdata[6]),
    .A2(_05256_),
    .ZN(_05325_)
  );
  INV_X1 _25615_ (
    .A(_05325_),
    .ZN(_05326_)
  );
  AND2_X1 _25616_ (
    .A1(_05324_),
    .A2(_05326_),
    .ZN(_05327_)
  );
  INV_X1 _25617_ (
    .A(_05327_),
    .ZN(_05328_)
  );
  MUX2_X1 _25618_ (
    .A(_05328_),
    .B(io_dmem_resp_bits_data_word_bypass[6]),
    .S(_05255_),
    .Z(_05329_)
  );
  MUX2_X1 _25619_ (
    .A(ex_reg_rs_msb_1[4]),
    .B(_05329_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[6])
  );
  MUX2_X1 _25620_ (
    .A(mem_reg_rs2[6]),
    .B(_ex_op2_T[6]),
    .S(_05269_),
    .Z(_00247_)
  );
  AND2_X1 _25621_ (
    .A1(mem_reg_wdata[7]),
    .A2(_05259_),
    .ZN(_05330_)
  );
  INV_X1 _25622_ (
    .A(_05330_),
    .ZN(_05331_)
  );
  AND2_X1 _25623_ (
    .A1(wb_reg_wdata[7]),
    .A2(_05256_),
    .ZN(_05332_)
  );
  INV_X1 _25624_ (
    .A(_05332_),
    .ZN(_05333_)
  );
  AND2_X1 _25625_ (
    .A1(_05331_),
    .A2(_05333_),
    .ZN(_05334_)
  );
  INV_X1 _25626_ (
    .A(_05334_),
    .ZN(_05335_)
  );
  MUX2_X1 _25627_ (
    .A(_05335_),
    .B(io_dmem_resp_bits_data_word_bypass[7]),
    .S(_05255_),
    .Z(_05336_)
  );
  MUX2_X1 _25628_ (
    .A(ex_reg_rs_msb_1[5]),
    .B(_05336_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[7])
  );
  MUX2_X1 _25629_ (
    .A(mem_reg_rs2[7]),
    .B(_ex_op2_T[7]),
    .S(_05269_),
    .Z(_00248_)
  );
  AND2_X1 _25630_ (
    .A1(_08153_),
    .A2(_08154_),
    .ZN(_05337_)
  );
  INV_X1 _25631_ (
    .A(_05337_),
    .ZN(_05338_)
  );
  AND2_X1 _25632_ (
    .A1(mem_reg_wdata[8]),
    .A2(_05259_),
    .ZN(_05339_)
  );
  INV_X1 _25633_ (
    .A(_05339_),
    .ZN(_05340_)
  );
  AND2_X1 _25634_ (
    .A1(wb_reg_wdata[8]),
    .A2(_05256_),
    .ZN(_05341_)
  );
  INV_X1 _25635_ (
    .A(_05341_),
    .ZN(_05342_)
  );
  AND2_X1 _25636_ (
    .A1(_05340_),
    .A2(_05342_),
    .ZN(_05343_)
  );
  INV_X1 _25637_ (
    .A(_05343_),
    .ZN(_05344_)
  );
  MUX2_X1 _25638_ (
    .A(_05344_),
    .B(io_dmem_resp_bits_data_word_bypass[8]),
    .S(_05255_),
    .Z(_05345_)
  );
  MUX2_X1 _25639_ (
    .A(ex_reg_rs_msb_1[6]),
    .B(_05345_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[8])
  );
  AND2_X1 _25640_ (
    .A1(_05338_),
    .A2(_ex_op2_T[8]),
    .ZN(_05346_)
  );
  INV_X1 _25641_ (
    .A(_05346_),
    .ZN(_05347_)
  );
  AND2_X1 _25642_ (
    .A1(_05269_),
    .A2(_05338_),
    .ZN(_05348_)
  );
  INV_X1 _25643_ (
    .A(_05348_),
    .ZN(_05349_)
  );
  AND2_X1 _25644_ (
    .A1(_05272_),
    .A2(_05349_),
    .ZN(_05350_)
  );
  INV_X1 _25645_ (
    .A(_05350_),
    .ZN(_05351_)
  );
  AND2_X1 _25646_ (
    .A1(_05347_),
    .A2(_05351_),
    .ZN(_05352_)
  );
  INV_X1 _25647_ (
    .A(_05352_),
    .ZN(_05353_)
  );
  AND2_X1 _25648_ (
    .A1(_08043_),
    .A2(_05270_),
    .ZN(_05354_)
  );
  INV_X1 _25649_ (
    .A(_05354_),
    .ZN(_05355_)
  );
  AND2_X1 _25650_ (
    .A1(_05353_),
    .A2(_05355_),
    .ZN(_00249_)
  );
  AND2_X1 _25651_ (
    .A1(mem_reg_wdata[9]),
    .A2(_05259_),
    .ZN(_05356_)
  );
  INV_X1 _25652_ (
    .A(_05356_),
    .ZN(_05357_)
  );
  AND2_X1 _25653_ (
    .A1(wb_reg_wdata[9]),
    .A2(_05256_),
    .ZN(_05358_)
  );
  INV_X1 _25654_ (
    .A(_05358_),
    .ZN(_05359_)
  );
  AND2_X1 _25655_ (
    .A1(_05357_),
    .A2(_05359_),
    .ZN(_05360_)
  );
  INV_X1 _25656_ (
    .A(_05360_),
    .ZN(_05361_)
  );
  MUX2_X1 _25657_ (
    .A(_05361_),
    .B(io_dmem_resp_bits_data_word_bypass[9]),
    .S(_05255_),
    .Z(_05362_)
  );
  MUX2_X1 _25658_ (
    .A(ex_reg_rs_msb_1[7]),
    .B(_05362_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[9])
  );
  AND2_X1 _25659_ (
    .A1(_05338_),
    .A2(_ex_op2_T[9]),
    .ZN(_05363_)
  );
  INV_X1 _25660_ (
    .A(_05363_),
    .ZN(_05364_)
  );
  AND2_X1 _25661_ (
    .A1(_05282_),
    .A2(_05349_),
    .ZN(_05365_)
  );
  INV_X1 _25662_ (
    .A(_05365_),
    .ZN(_05366_)
  );
  AND2_X1 _25663_ (
    .A1(_05364_),
    .A2(_05366_),
    .ZN(_05367_)
  );
  INV_X1 _25664_ (
    .A(_05367_),
    .ZN(_05368_)
  );
  AND2_X1 _25665_ (
    .A1(_08044_),
    .A2(_05270_),
    .ZN(_05369_)
  );
  INV_X1 _25666_ (
    .A(_05369_),
    .ZN(_05370_)
  );
  AND2_X1 _25667_ (
    .A1(_05368_),
    .A2(_05370_),
    .ZN(_00250_)
  );
  AND2_X1 _25668_ (
    .A1(mem_reg_wdata[10]),
    .A2(_05259_),
    .ZN(_05371_)
  );
  INV_X1 _25669_ (
    .A(_05371_),
    .ZN(_05372_)
  );
  AND2_X1 _25670_ (
    .A1(wb_reg_wdata[10]),
    .A2(_05256_),
    .ZN(_05373_)
  );
  INV_X1 _25671_ (
    .A(_05373_),
    .ZN(_05374_)
  );
  AND2_X1 _25672_ (
    .A1(_05372_),
    .A2(_05374_),
    .ZN(_05375_)
  );
  INV_X1 _25673_ (
    .A(_05375_),
    .ZN(_05376_)
  );
  MUX2_X1 _25674_ (
    .A(_05376_),
    .B(io_dmem_resp_bits_data_word_bypass[10]),
    .S(_05255_),
    .Z(_05377_)
  );
  MUX2_X1 _25675_ (
    .A(ex_reg_rs_msb_1[8]),
    .B(_05377_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[10])
  );
  AND2_X1 _25676_ (
    .A1(_05338_),
    .A2(_ex_op2_T[10]),
    .ZN(_05378_)
  );
  INV_X1 _25677_ (
    .A(_05378_),
    .ZN(_05379_)
  );
  AND2_X1 _25678_ (
    .A1(_05292_),
    .A2(_05349_),
    .ZN(_05380_)
  );
  INV_X1 _25679_ (
    .A(_05380_),
    .ZN(_05381_)
  );
  AND2_X1 _25680_ (
    .A1(_05379_),
    .A2(_05381_),
    .ZN(_05382_)
  );
  INV_X1 _25681_ (
    .A(_05382_),
    .ZN(_05383_)
  );
  AND2_X1 _25682_ (
    .A1(_08045_),
    .A2(_05270_),
    .ZN(_05384_)
  );
  INV_X1 _25683_ (
    .A(_05384_),
    .ZN(_05385_)
  );
  AND2_X1 _25684_ (
    .A1(_05383_),
    .A2(_05385_),
    .ZN(_00251_)
  );
  AND2_X1 _25685_ (
    .A1(mem_reg_wdata[11]),
    .A2(_05259_),
    .ZN(_05386_)
  );
  INV_X1 _25686_ (
    .A(_05386_),
    .ZN(_05387_)
  );
  AND2_X1 _25687_ (
    .A1(wb_reg_wdata[11]),
    .A2(_05256_),
    .ZN(_05388_)
  );
  INV_X1 _25688_ (
    .A(_05388_),
    .ZN(_05389_)
  );
  AND2_X1 _25689_ (
    .A1(_05387_),
    .A2(_05389_),
    .ZN(_05390_)
  );
  INV_X1 _25690_ (
    .A(_05390_),
    .ZN(_05391_)
  );
  MUX2_X1 _25691_ (
    .A(_05391_),
    .B(io_dmem_resp_bits_data_word_bypass[11]),
    .S(_05255_),
    .Z(_05392_)
  );
  MUX2_X1 _25692_ (
    .A(ex_reg_rs_msb_1[9]),
    .B(_05392_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[11])
  );
  AND2_X1 _25693_ (
    .A1(_05338_),
    .A2(_ex_op2_T[11]),
    .ZN(_05393_)
  );
  INV_X1 _25694_ (
    .A(_05393_),
    .ZN(_05394_)
  );
  AND2_X1 _25695_ (
    .A1(_05302_),
    .A2(_05349_),
    .ZN(_05395_)
  );
  INV_X1 _25696_ (
    .A(_05395_),
    .ZN(_05396_)
  );
  AND2_X1 _25697_ (
    .A1(_05394_),
    .A2(_05396_),
    .ZN(_05397_)
  );
  INV_X1 _25698_ (
    .A(_05397_),
    .ZN(_05398_)
  );
  AND2_X1 _25699_ (
    .A1(_08046_),
    .A2(_05270_),
    .ZN(_05399_)
  );
  INV_X1 _25700_ (
    .A(_05399_),
    .ZN(_05400_)
  );
  AND2_X1 _25701_ (
    .A1(_05398_),
    .A2(_05400_),
    .ZN(_00252_)
  );
  AND2_X1 _25702_ (
    .A1(mem_reg_wdata[12]),
    .A2(_05259_),
    .ZN(_05401_)
  );
  INV_X1 _25703_ (
    .A(_05401_),
    .ZN(_05402_)
  );
  AND2_X1 _25704_ (
    .A1(wb_reg_wdata[12]),
    .A2(_05256_),
    .ZN(_05403_)
  );
  INV_X1 _25705_ (
    .A(_05403_),
    .ZN(_05404_)
  );
  AND2_X1 _25706_ (
    .A1(_05402_),
    .A2(_05404_),
    .ZN(_05405_)
  );
  INV_X1 _25707_ (
    .A(_05405_),
    .ZN(_05406_)
  );
  MUX2_X1 _25708_ (
    .A(_05406_),
    .B(io_dmem_resp_bits_data_word_bypass[12]),
    .S(_05255_),
    .Z(_05407_)
  );
  MUX2_X1 _25709_ (
    .A(ex_reg_rs_msb_1[10]),
    .B(_05407_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[12])
  );
  AND2_X1 _25710_ (
    .A1(_05338_),
    .A2(_ex_op2_T[12]),
    .ZN(_05408_)
  );
  INV_X1 _25711_ (
    .A(_05408_),
    .ZN(_05409_)
  );
  AND2_X1 _25712_ (
    .A1(_05312_),
    .A2(_05349_),
    .ZN(_05410_)
  );
  INV_X1 _25713_ (
    .A(_05410_),
    .ZN(_05411_)
  );
  AND2_X1 _25714_ (
    .A1(_05409_),
    .A2(_05411_),
    .ZN(_05412_)
  );
  INV_X1 _25715_ (
    .A(_05412_),
    .ZN(_05413_)
  );
  AND2_X1 _25716_ (
    .A1(_08047_),
    .A2(_05270_),
    .ZN(_05414_)
  );
  INV_X1 _25717_ (
    .A(_05414_),
    .ZN(_05415_)
  );
  AND2_X1 _25718_ (
    .A1(_05413_),
    .A2(_05415_),
    .ZN(_00253_)
  );
  AND2_X1 _25719_ (
    .A1(mem_reg_wdata[13]),
    .A2(_05259_),
    .ZN(_05416_)
  );
  INV_X1 _25720_ (
    .A(_05416_),
    .ZN(_05417_)
  );
  AND2_X1 _25721_ (
    .A1(wb_reg_wdata[13]),
    .A2(_05256_),
    .ZN(_05418_)
  );
  INV_X1 _25722_ (
    .A(_05418_),
    .ZN(_05419_)
  );
  AND2_X1 _25723_ (
    .A1(_05417_),
    .A2(_05419_),
    .ZN(_05420_)
  );
  INV_X1 _25724_ (
    .A(_05420_),
    .ZN(_05421_)
  );
  MUX2_X1 _25725_ (
    .A(_05421_),
    .B(io_dmem_resp_bits_data_word_bypass[13]),
    .S(_05255_),
    .Z(_05422_)
  );
  MUX2_X1 _25726_ (
    .A(ex_reg_rs_msb_1[11]),
    .B(_05422_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[13])
  );
  AND2_X1 _25727_ (
    .A1(_05338_),
    .A2(_ex_op2_T[13]),
    .ZN(_05423_)
  );
  INV_X1 _25728_ (
    .A(_05423_),
    .ZN(_05424_)
  );
  AND2_X1 _25729_ (
    .A1(_05322_),
    .A2(_05349_),
    .ZN(_05425_)
  );
  INV_X1 _25730_ (
    .A(_05425_),
    .ZN(_05426_)
  );
  AND2_X1 _25731_ (
    .A1(_05424_),
    .A2(_05426_),
    .ZN(_05427_)
  );
  INV_X1 _25732_ (
    .A(_05427_),
    .ZN(_05428_)
  );
  AND2_X1 _25733_ (
    .A1(_08048_),
    .A2(_05270_),
    .ZN(_05429_)
  );
  INV_X1 _25734_ (
    .A(_05429_),
    .ZN(_05430_)
  );
  AND2_X1 _25735_ (
    .A1(_05428_),
    .A2(_05430_),
    .ZN(_00254_)
  );
  AND2_X1 _25736_ (
    .A1(mem_reg_wdata[14]),
    .A2(_05259_),
    .ZN(_05431_)
  );
  INV_X1 _25737_ (
    .A(_05431_),
    .ZN(_05432_)
  );
  AND2_X1 _25738_ (
    .A1(wb_reg_wdata[14]),
    .A2(_05256_),
    .ZN(_05433_)
  );
  INV_X1 _25739_ (
    .A(_05433_),
    .ZN(_05434_)
  );
  AND2_X1 _25740_ (
    .A1(_05432_),
    .A2(_05434_),
    .ZN(_05435_)
  );
  INV_X1 _25741_ (
    .A(_05435_),
    .ZN(_05436_)
  );
  MUX2_X1 _25742_ (
    .A(_05436_),
    .B(io_dmem_resp_bits_data_word_bypass[14]),
    .S(_05255_),
    .Z(_05437_)
  );
  MUX2_X1 _25743_ (
    .A(ex_reg_rs_msb_1[12]),
    .B(_05437_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[14])
  );
  AND2_X1 _25744_ (
    .A1(_05338_),
    .A2(_ex_op2_T[14]),
    .ZN(_05438_)
  );
  INV_X1 _25745_ (
    .A(_05438_),
    .ZN(_05439_)
  );
  AND2_X1 _25746_ (
    .A1(_ex_op2_T[6]),
    .A2(_05337_),
    .ZN(_05440_)
  );
  INV_X1 _25747_ (
    .A(_05440_),
    .ZN(_05441_)
  );
  MUX2_X1 _25748_ (
    .A(_ex_op2_T[6]),
    .B(_ex_op2_T[14]),
    .S(_05338_),
    .Z(_05442_)
  );
  MUX2_X1 _25749_ (
    .A(mem_reg_rs2[14]),
    .B(_05442_),
    .S(_05269_),
    .Z(_00255_)
  );
  AND2_X1 _25750_ (
    .A1(mem_reg_wdata[15]),
    .A2(_05259_),
    .ZN(_05443_)
  );
  INV_X1 _25751_ (
    .A(_05443_),
    .ZN(_05444_)
  );
  AND2_X1 _25752_ (
    .A1(wb_reg_wdata[15]),
    .A2(_05256_),
    .ZN(_05445_)
  );
  INV_X1 _25753_ (
    .A(_05445_),
    .ZN(_05446_)
  );
  AND2_X1 _25754_ (
    .A1(_05444_),
    .A2(_05446_),
    .ZN(_05447_)
  );
  INV_X1 _25755_ (
    .A(_05447_),
    .ZN(_05448_)
  );
  MUX2_X1 _25756_ (
    .A(_05448_),
    .B(io_dmem_resp_bits_data_word_bypass[15]),
    .S(_05255_),
    .Z(_05449_)
  );
  MUX2_X1 _25757_ (
    .A(ex_reg_rs_msb_1[13]),
    .B(_05449_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[15])
  );
  AND2_X1 _25758_ (
    .A1(_05338_),
    .A2(_ex_op2_T[15]),
    .ZN(_05450_)
  );
  INV_X1 _25759_ (
    .A(_05450_),
    .ZN(_05451_)
  );
  AND2_X1 _25760_ (
    .A1(_ex_op2_T[7]),
    .A2(_05337_),
    .ZN(_05452_)
  );
  INV_X1 _25761_ (
    .A(_05452_),
    .ZN(_05453_)
  );
  MUX2_X1 _25762_ (
    .A(_ex_op2_T[7]),
    .B(_ex_op2_T[15]),
    .S(_05338_),
    .Z(_05454_)
  );
  MUX2_X1 _25763_ (
    .A(mem_reg_rs2[15]),
    .B(_05454_),
    .S(_05269_),
    .Z(_00256_)
  );
  AND2_X1 _25764_ (
    .A1(_08154_),
    .A2(_08557_),
    .ZN(_05455_)
  );
  INV_X1 _25765_ (
    .A(_05455_),
    .ZN(_05456_)
  );
  AND2_X1 _25766_ (
    .A1(_05338_),
    .A2(_05456_),
    .ZN(_05457_)
  );
  INV_X1 _25767_ (
    .A(_05457_),
    .ZN(_05458_)
  );
  AND2_X1 _25768_ (
    .A1(mem_reg_wdata[16]),
    .A2(_05259_),
    .ZN(_05459_)
  );
  INV_X1 _25769_ (
    .A(_05459_),
    .ZN(_05460_)
  );
  AND2_X1 _25770_ (
    .A1(wb_reg_wdata[16]),
    .A2(_05256_),
    .ZN(_05461_)
  );
  INV_X1 _25771_ (
    .A(_05461_),
    .ZN(_05462_)
  );
  AND2_X1 _25772_ (
    .A1(_05460_),
    .A2(_05462_),
    .ZN(_05463_)
  );
  INV_X1 _25773_ (
    .A(_05463_),
    .ZN(_05464_)
  );
  MUX2_X1 _25774_ (
    .A(_05464_),
    .B(io_dmem_resp_bits_data_word_bypass[16]),
    .S(_05255_),
    .Z(_05465_)
  );
  MUX2_X1 _25775_ (
    .A(ex_reg_rs_msb_1[14]),
    .B(_05465_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[16])
  );
  MUX2_X1 _25776_ (
    .A(_ex_op2_T[0]),
    .B(_ex_op2_T[16]),
    .S(_05457_),
    .Z(_05466_)
  );
  MUX2_X1 _25777_ (
    .A(mem_reg_rs2[16]),
    .B(_05466_),
    .S(_05269_),
    .Z(_00257_)
  );
  AND2_X1 _25778_ (
    .A1(mem_reg_wdata[17]),
    .A2(_05259_),
    .ZN(_05467_)
  );
  INV_X1 _25779_ (
    .A(_05467_),
    .ZN(_05468_)
  );
  AND2_X1 _25780_ (
    .A1(wb_reg_wdata[17]),
    .A2(_05256_),
    .ZN(_05469_)
  );
  INV_X1 _25781_ (
    .A(_05469_),
    .ZN(_05470_)
  );
  AND2_X1 _25782_ (
    .A1(_05468_),
    .A2(_05470_),
    .ZN(_05471_)
  );
  INV_X1 _25783_ (
    .A(_05471_),
    .ZN(_05472_)
  );
  MUX2_X1 _25784_ (
    .A(_05472_),
    .B(io_dmem_resp_bits_data_word_bypass[17]),
    .S(_05255_),
    .Z(_05473_)
  );
  MUX2_X1 _25785_ (
    .A(ex_reg_rs_msb_1[15]),
    .B(_05473_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[17])
  );
  MUX2_X1 _25786_ (
    .A(_ex_op2_T[1]),
    .B(_ex_op2_T[17]),
    .S(_05457_),
    .Z(_05474_)
  );
  MUX2_X1 _25787_ (
    .A(mem_reg_rs2[17]),
    .B(_05474_),
    .S(_05269_),
    .Z(_00258_)
  );
  AND2_X1 _25788_ (
    .A1(mem_reg_wdata[18]),
    .A2(_05259_),
    .ZN(_05475_)
  );
  INV_X1 _25789_ (
    .A(_05475_),
    .ZN(_05476_)
  );
  AND2_X1 _25790_ (
    .A1(wb_reg_wdata[18]),
    .A2(_05256_),
    .ZN(_05477_)
  );
  INV_X1 _25791_ (
    .A(_05477_),
    .ZN(_05478_)
  );
  AND2_X1 _25792_ (
    .A1(_05476_),
    .A2(_05478_),
    .ZN(_05479_)
  );
  INV_X1 _25793_ (
    .A(_05479_),
    .ZN(_05480_)
  );
  MUX2_X1 _25794_ (
    .A(_05480_),
    .B(io_dmem_resp_bits_data_word_bypass[18]),
    .S(_05255_),
    .Z(_05481_)
  );
  MUX2_X1 _25795_ (
    .A(ex_reg_rs_msb_1[16]),
    .B(_05481_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[18])
  );
  MUX2_X1 _25796_ (
    .A(_ex_op2_T[2]),
    .B(_ex_op2_T[18]),
    .S(_05457_),
    .Z(_05482_)
  );
  MUX2_X1 _25797_ (
    .A(mem_reg_rs2[18]),
    .B(_05482_),
    .S(_05269_),
    .Z(_00259_)
  );
  AND2_X1 _25798_ (
    .A1(mem_reg_wdata[19]),
    .A2(_05259_),
    .ZN(_05483_)
  );
  INV_X1 _25799_ (
    .A(_05483_),
    .ZN(_05484_)
  );
  AND2_X1 _25800_ (
    .A1(wb_reg_wdata[19]),
    .A2(_05256_),
    .ZN(_05485_)
  );
  INV_X1 _25801_ (
    .A(_05485_),
    .ZN(_05486_)
  );
  AND2_X1 _25802_ (
    .A1(_05484_),
    .A2(_05486_),
    .ZN(_05487_)
  );
  INV_X1 _25803_ (
    .A(_05487_),
    .ZN(_05488_)
  );
  MUX2_X1 _25804_ (
    .A(_05488_),
    .B(io_dmem_resp_bits_data_word_bypass[19]),
    .S(_05255_),
    .Z(_05489_)
  );
  MUX2_X1 _25805_ (
    .A(ex_reg_rs_msb_1[17]),
    .B(_05489_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[19])
  );
  MUX2_X1 _25806_ (
    .A(_ex_op2_T[3]),
    .B(_ex_op2_T[19]),
    .S(_05457_),
    .Z(_05490_)
  );
  MUX2_X1 _25807_ (
    .A(mem_reg_rs2[19]),
    .B(_05490_),
    .S(_05269_),
    .Z(_00260_)
  );
  AND2_X1 _25808_ (
    .A1(mem_reg_wdata[20]),
    .A2(_05259_),
    .ZN(_05491_)
  );
  INV_X1 _25809_ (
    .A(_05491_),
    .ZN(_05492_)
  );
  AND2_X1 _25810_ (
    .A1(wb_reg_wdata[20]),
    .A2(_05256_),
    .ZN(_05493_)
  );
  INV_X1 _25811_ (
    .A(_05493_),
    .ZN(_05494_)
  );
  AND2_X1 _25812_ (
    .A1(_05492_),
    .A2(_05494_),
    .ZN(_05495_)
  );
  INV_X1 _25813_ (
    .A(_05495_),
    .ZN(_05496_)
  );
  MUX2_X1 _25814_ (
    .A(_05496_),
    .B(io_dmem_resp_bits_data_word_bypass[20]),
    .S(_05255_),
    .Z(_05497_)
  );
  MUX2_X1 _25815_ (
    .A(ex_reg_rs_msb_1[18]),
    .B(_05497_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[20])
  );
  MUX2_X1 _25816_ (
    .A(_ex_op2_T[4]),
    .B(_ex_op2_T[20]),
    .S(_05457_),
    .Z(_05498_)
  );
  MUX2_X1 _25817_ (
    .A(mem_reg_rs2[20]),
    .B(_05498_),
    .S(_05269_),
    .Z(_00261_)
  );
  AND2_X1 _25818_ (
    .A1(mem_reg_wdata[21]),
    .A2(_05259_),
    .ZN(_05499_)
  );
  INV_X1 _25819_ (
    .A(_05499_),
    .ZN(_05500_)
  );
  AND2_X1 _25820_ (
    .A1(wb_reg_wdata[21]),
    .A2(_05256_),
    .ZN(_05501_)
  );
  INV_X1 _25821_ (
    .A(_05501_),
    .ZN(_05502_)
  );
  AND2_X1 _25822_ (
    .A1(_05500_),
    .A2(_05502_),
    .ZN(_05503_)
  );
  INV_X1 _25823_ (
    .A(_05503_),
    .ZN(_05504_)
  );
  MUX2_X1 _25824_ (
    .A(_05504_),
    .B(io_dmem_resp_bits_data_word_bypass[21]),
    .S(_05255_),
    .Z(_05505_)
  );
  MUX2_X1 _25825_ (
    .A(ex_reg_rs_msb_1[19]),
    .B(_05505_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[21])
  );
  MUX2_X1 _25826_ (
    .A(_ex_op2_T[5]),
    .B(_ex_op2_T[21]),
    .S(_05457_),
    .Z(_05506_)
  );
  MUX2_X1 _25827_ (
    .A(mem_reg_rs2[21]),
    .B(_05506_),
    .S(_05269_),
    .Z(_00262_)
  );
  AND2_X1 _25828_ (
    .A1(mem_reg_wdata[22]),
    .A2(_05259_),
    .ZN(_05507_)
  );
  INV_X1 _25829_ (
    .A(_05507_),
    .ZN(_05508_)
  );
  AND2_X1 _25830_ (
    .A1(wb_reg_wdata[22]),
    .A2(_05256_),
    .ZN(_05509_)
  );
  INV_X1 _25831_ (
    .A(_05509_),
    .ZN(_05510_)
  );
  AND2_X1 _25832_ (
    .A1(_05508_),
    .A2(_05510_),
    .ZN(_05511_)
  );
  INV_X1 _25833_ (
    .A(_05511_),
    .ZN(_05512_)
  );
  MUX2_X1 _25834_ (
    .A(_05512_),
    .B(io_dmem_resp_bits_data_word_bypass[22]),
    .S(_05255_),
    .Z(_05513_)
  );
  MUX2_X1 _25835_ (
    .A(ex_reg_rs_msb_1[20]),
    .B(_05513_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[22])
  );
  MUX2_X1 _25836_ (
    .A(_ex_op2_T[6]),
    .B(_ex_op2_T[22]),
    .S(_05457_),
    .Z(_05514_)
  );
  MUX2_X1 _25837_ (
    .A(mem_reg_rs2[22]),
    .B(_05514_),
    .S(_05269_),
    .Z(_00263_)
  );
  AND2_X1 _25838_ (
    .A1(mem_reg_wdata[23]),
    .A2(_05259_),
    .ZN(_05515_)
  );
  INV_X1 _25839_ (
    .A(_05515_),
    .ZN(_05516_)
  );
  AND2_X1 _25840_ (
    .A1(wb_reg_wdata[23]),
    .A2(_05256_),
    .ZN(_05517_)
  );
  INV_X1 _25841_ (
    .A(_05517_),
    .ZN(_05518_)
  );
  AND2_X1 _25842_ (
    .A1(_05516_),
    .A2(_05518_),
    .ZN(_05519_)
  );
  INV_X1 _25843_ (
    .A(_05519_),
    .ZN(_05520_)
  );
  MUX2_X1 _25844_ (
    .A(_05520_),
    .B(io_dmem_resp_bits_data_word_bypass[23]),
    .S(_05255_),
    .Z(_05521_)
  );
  MUX2_X1 _25845_ (
    .A(ex_reg_rs_msb_1[21]),
    .B(_05521_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[23])
  );
  MUX2_X1 _25846_ (
    .A(_ex_op2_T[7]),
    .B(_ex_op2_T[23]),
    .S(_05457_),
    .Z(_05522_)
  );
  MUX2_X1 _25847_ (
    .A(mem_reg_rs2[23]),
    .B(_05522_),
    .S(_05269_),
    .Z(_00264_)
  );
  AND2_X1 _25848_ (
    .A1(_05352_),
    .A2(_05458_),
    .ZN(_05523_)
  );
  INV_X1 _25849_ (
    .A(_05523_),
    .ZN(_05524_)
  );
  AND2_X1 _25850_ (
    .A1(mem_reg_wdata[24]),
    .A2(_05259_),
    .ZN(_05525_)
  );
  INV_X1 _25851_ (
    .A(_05525_),
    .ZN(_05526_)
  );
  AND2_X1 _25852_ (
    .A1(wb_reg_wdata[24]),
    .A2(_05256_),
    .ZN(_05527_)
  );
  INV_X1 _25853_ (
    .A(_05527_),
    .ZN(_05528_)
  );
  AND2_X1 _25854_ (
    .A1(_05526_),
    .A2(_05528_),
    .ZN(_05529_)
  );
  INV_X1 _25855_ (
    .A(_05529_),
    .ZN(_05530_)
  );
  MUX2_X1 _25856_ (
    .A(_05530_),
    .B(io_dmem_resp_bits_data_word_bypass[24]),
    .S(_05255_),
    .Z(_05531_)
  );
  MUX2_X1 _25857_ (
    .A(ex_reg_rs_msb_1[22]),
    .B(_05531_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[24])
  );
  INV_X1 _25858_ (
    .A(_ex_op2_T[24]),
    .ZN(_05532_)
  );
  AND2_X1 _25859_ (
    .A1(_05456_),
    .A2(_05532_),
    .ZN(_05533_)
  );
  AND2_X1 _25860_ (
    .A1(_05351_),
    .A2(_05533_),
    .ZN(_05534_)
  );
  INV_X1 _25861_ (
    .A(_05534_),
    .ZN(_05535_)
  );
  AND2_X1 _25862_ (
    .A1(_08049_),
    .A2(_05270_),
    .ZN(_05536_)
  );
  INV_X1 _25863_ (
    .A(_05536_),
    .ZN(_05537_)
  );
  AND2_X1 _25864_ (
    .A1(_05535_),
    .A2(_05537_),
    .ZN(_05538_)
  );
  AND2_X1 _25865_ (
    .A1(_05524_),
    .A2(_05538_),
    .ZN(_00265_)
  );
  AND2_X1 _25866_ (
    .A1(_05367_),
    .A2(_05458_),
    .ZN(_05539_)
  );
  INV_X1 _25867_ (
    .A(_05539_),
    .ZN(_05540_)
  );
  AND2_X1 _25868_ (
    .A1(_08050_),
    .A2(_05270_),
    .ZN(_05541_)
  );
  INV_X1 _25869_ (
    .A(_05541_),
    .ZN(_05542_)
  );
  AND2_X1 _25870_ (
    .A1(mem_reg_wdata[25]),
    .A2(_05259_),
    .ZN(_05543_)
  );
  INV_X1 _25871_ (
    .A(_05543_),
    .ZN(_05544_)
  );
  AND2_X1 _25872_ (
    .A1(wb_reg_wdata[25]),
    .A2(_05256_),
    .ZN(_05545_)
  );
  INV_X1 _25873_ (
    .A(_05545_),
    .ZN(_05546_)
  );
  AND2_X1 _25874_ (
    .A1(_05544_),
    .A2(_05546_),
    .ZN(_05547_)
  );
  INV_X1 _25875_ (
    .A(_05547_),
    .ZN(_05548_)
  );
  MUX2_X1 _25876_ (
    .A(_05548_),
    .B(io_dmem_resp_bits_data_word_bypass[25]),
    .S(_05255_),
    .Z(_05549_)
  );
  MUX2_X1 _25877_ (
    .A(ex_reg_rs_msb_1[23]),
    .B(_05549_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[25])
  );
  INV_X1 _25878_ (
    .A(_ex_op2_T[25]),
    .ZN(_05550_)
  );
  AND2_X1 _25879_ (
    .A1(_05456_),
    .A2(_05550_),
    .ZN(_05551_)
  );
  AND2_X1 _25880_ (
    .A1(_05366_),
    .A2(_05551_),
    .ZN(_05552_)
  );
  INV_X1 _25881_ (
    .A(_05552_),
    .ZN(_05553_)
  );
  AND2_X1 _25882_ (
    .A1(_05542_),
    .A2(_05553_),
    .ZN(_05554_)
  );
  AND2_X1 _25883_ (
    .A1(_05540_),
    .A2(_05554_),
    .ZN(_00266_)
  );
  AND2_X1 _25884_ (
    .A1(_05382_),
    .A2(_05458_),
    .ZN(_05555_)
  );
  INV_X1 _25885_ (
    .A(_05555_),
    .ZN(_05556_)
  );
  AND2_X1 _25886_ (
    .A1(mem_reg_wdata[26]),
    .A2(_05259_),
    .ZN(_05557_)
  );
  INV_X1 _25887_ (
    .A(_05557_),
    .ZN(_05558_)
  );
  AND2_X1 _25888_ (
    .A1(wb_reg_wdata[26]),
    .A2(_05256_),
    .ZN(_05559_)
  );
  INV_X1 _25889_ (
    .A(_05559_),
    .ZN(_05560_)
  );
  AND2_X1 _25890_ (
    .A1(_05558_),
    .A2(_05560_),
    .ZN(_05561_)
  );
  INV_X1 _25891_ (
    .A(_05561_),
    .ZN(_05562_)
  );
  MUX2_X1 _25892_ (
    .A(_05562_),
    .B(io_dmem_resp_bits_data_word_bypass[26]),
    .S(_05255_),
    .Z(_05563_)
  );
  MUX2_X1 _25893_ (
    .A(ex_reg_rs_msb_1[24]),
    .B(_05563_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[26])
  );
  INV_X1 _25894_ (
    .A(_ex_op2_T[26]),
    .ZN(_05564_)
  );
  AND2_X1 _25895_ (
    .A1(_05456_),
    .A2(_05564_),
    .ZN(_05565_)
  );
  AND2_X1 _25896_ (
    .A1(_05381_),
    .A2(_05565_),
    .ZN(_05566_)
  );
  INV_X1 _25897_ (
    .A(_05566_),
    .ZN(_05567_)
  );
  AND2_X1 _25898_ (
    .A1(_08051_),
    .A2(_05270_),
    .ZN(_05568_)
  );
  INV_X1 _25899_ (
    .A(_05568_),
    .ZN(_05569_)
  );
  AND2_X1 _25900_ (
    .A1(_05567_),
    .A2(_05569_),
    .ZN(_05570_)
  );
  AND2_X1 _25901_ (
    .A1(_05556_),
    .A2(_05570_),
    .ZN(_00267_)
  );
  AND2_X1 _25902_ (
    .A1(_05397_),
    .A2(_05458_),
    .ZN(_05571_)
  );
  INV_X1 _25903_ (
    .A(_05571_),
    .ZN(_05572_)
  );
  AND2_X1 _25904_ (
    .A1(mem_reg_wdata[27]),
    .A2(_05259_),
    .ZN(_05573_)
  );
  INV_X1 _25905_ (
    .A(_05573_),
    .ZN(_05574_)
  );
  AND2_X1 _25906_ (
    .A1(wb_reg_wdata[27]),
    .A2(_05256_),
    .ZN(_05575_)
  );
  INV_X1 _25907_ (
    .A(_05575_),
    .ZN(_05576_)
  );
  AND2_X1 _25908_ (
    .A1(_05574_),
    .A2(_05576_),
    .ZN(_05577_)
  );
  INV_X1 _25909_ (
    .A(_05577_),
    .ZN(_05578_)
  );
  MUX2_X1 _25910_ (
    .A(_05578_),
    .B(io_dmem_resp_bits_data_word_bypass[27]),
    .S(_05255_),
    .Z(_05579_)
  );
  MUX2_X1 _25911_ (
    .A(ex_reg_rs_msb_1[25]),
    .B(_05579_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[27])
  );
  INV_X1 _25912_ (
    .A(_ex_op2_T[27]),
    .ZN(_05580_)
  );
  AND2_X1 _25913_ (
    .A1(_05456_),
    .A2(_05580_),
    .ZN(_05581_)
  );
  AND2_X1 _25914_ (
    .A1(_05396_),
    .A2(_05581_),
    .ZN(_05582_)
  );
  INV_X1 _25915_ (
    .A(_05582_),
    .ZN(_05583_)
  );
  AND2_X1 _25916_ (
    .A1(_08052_),
    .A2(_05270_),
    .ZN(_05584_)
  );
  INV_X1 _25917_ (
    .A(_05584_),
    .ZN(_05585_)
  );
  AND2_X1 _25918_ (
    .A1(_05583_),
    .A2(_05585_),
    .ZN(_05586_)
  );
  AND2_X1 _25919_ (
    .A1(_05572_),
    .A2(_05586_),
    .ZN(_00268_)
  );
  AND2_X1 _25920_ (
    .A1(_05412_),
    .A2(_05458_),
    .ZN(_05587_)
  );
  INV_X1 _25921_ (
    .A(_05587_),
    .ZN(_05588_)
  );
  AND2_X1 _25922_ (
    .A1(mem_reg_wdata[28]),
    .A2(_05259_),
    .ZN(_05589_)
  );
  INV_X1 _25923_ (
    .A(_05589_),
    .ZN(_05590_)
  );
  AND2_X1 _25924_ (
    .A1(wb_reg_wdata[28]),
    .A2(_05256_),
    .ZN(_05591_)
  );
  INV_X1 _25925_ (
    .A(_05591_),
    .ZN(_05592_)
  );
  AND2_X1 _25926_ (
    .A1(_05590_),
    .A2(_05592_),
    .ZN(_05593_)
  );
  INV_X1 _25927_ (
    .A(_05593_),
    .ZN(_05594_)
  );
  MUX2_X1 _25928_ (
    .A(_05594_),
    .B(io_dmem_resp_bits_data_word_bypass[28]),
    .S(_05255_),
    .Z(_05595_)
  );
  MUX2_X1 _25929_ (
    .A(ex_reg_rs_msb_1[26]),
    .B(_05595_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[28])
  );
  INV_X1 _25930_ (
    .A(_ex_op2_T[28]),
    .ZN(_05596_)
  );
  AND2_X1 _25931_ (
    .A1(_05456_),
    .A2(_05596_),
    .ZN(_05597_)
  );
  AND2_X1 _25932_ (
    .A1(_05411_),
    .A2(_05597_),
    .ZN(_05598_)
  );
  INV_X1 _25933_ (
    .A(_05598_),
    .ZN(_05599_)
  );
  AND2_X1 _25934_ (
    .A1(_08053_),
    .A2(_05270_),
    .ZN(_05600_)
  );
  INV_X1 _25935_ (
    .A(_05600_),
    .ZN(_05601_)
  );
  AND2_X1 _25936_ (
    .A1(_05599_),
    .A2(_05601_),
    .ZN(_05602_)
  );
  AND2_X1 _25937_ (
    .A1(_05588_),
    .A2(_05602_),
    .ZN(_00269_)
  );
  AND2_X1 _25938_ (
    .A1(_05427_),
    .A2(_05458_),
    .ZN(_05603_)
  );
  INV_X1 _25939_ (
    .A(_05603_),
    .ZN(_05604_)
  );
  AND2_X1 _25940_ (
    .A1(mem_reg_wdata[29]),
    .A2(_05259_),
    .ZN(_05605_)
  );
  INV_X1 _25941_ (
    .A(_05605_),
    .ZN(_05606_)
  );
  AND2_X1 _25942_ (
    .A1(wb_reg_wdata[29]),
    .A2(_05256_),
    .ZN(_05607_)
  );
  INV_X1 _25943_ (
    .A(_05607_),
    .ZN(_05608_)
  );
  AND2_X1 _25944_ (
    .A1(_05606_),
    .A2(_05608_),
    .ZN(_05609_)
  );
  INV_X1 _25945_ (
    .A(_05609_),
    .ZN(_05610_)
  );
  MUX2_X1 _25946_ (
    .A(_05610_),
    .B(io_dmem_resp_bits_data_word_bypass[29]),
    .S(_05255_),
    .Z(_05611_)
  );
  MUX2_X1 _25947_ (
    .A(ex_reg_rs_msb_1[27]),
    .B(_05611_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[29])
  );
  INV_X1 _25948_ (
    .A(_ex_op2_T[29]),
    .ZN(_05612_)
  );
  AND2_X1 _25949_ (
    .A1(_05456_),
    .A2(_05612_),
    .ZN(_05613_)
  );
  AND2_X1 _25950_ (
    .A1(_05426_),
    .A2(_05613_),
    .ZN(_05614_)
  );
  INV_X1 _25951_ (
    .A(_05614_),
    .ZN(_05615_)
  );
  AND2_X1 _25952_ (
    .A1(_08054_),
    .A2(_05270_),
    .ZN(_05616_)
  );
  INV_X1 _25953_ (
    .A(_05616_),
    .ZN(_05617_)
  );
  AND2_X1 _25954_ (
    .A1(_05615_),
    .A2(_05617_),
    .ZN(_05618_)
  );
  AND2_X1 _25955_ (
    .A1(_05604_),
    .A2(_05618_),
    .ZN(_00270_)
  );
  AND2_X1 _25956_ (
    .A1(_08055_),
    .A2(_05270_),
    .ZN(_05619_)
  );
  INV_X1 _25957_ (
    .A(_05619_),
    .ZN(_05620_)
  );
  AND2_X1 _25958_ (
    .A1(mem_reg_wdata[30]),
    .A2(_05259_),
    .ZN(_05621_)
  );
  INV_X1 _25959_ (
    .A(_05621_),
    .ZN(_05622_)
  );
  AND2_X1 _25960_ (
    .A1(wb_reg_wdata[30]),
    .A2(_05256_),
    .ZN(_05623_)
  );
  INV_X1 _25961_ (
    .A(_05623_),
    .ZN(_05624_)
  );
  AND2_X1 _25962_ (
    .A1(_05622_),
    .A2(_05624_),
    .ZN(_05625_)
  );
  INV_X1 _25963_ (
    .A(_05625_),
    .ZN(_05626_)
  );
  MUX2_X1 _25964_ (
    .A(_05626_),
    .B(io_dmem_resp_bits_data_word_bypass[30]),
    .S(_05255_),
    .Z(_05627_)
  );
  MUX2_X1 _25965_ (
    .A(ex_reg_rs_msb_1[28]),
    .B(_05627_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[30])
  );
  INV_X1 _25966_ (
    .A(_ex_op2_T[30]),
    .ZN(_05628_)
  );
  AND2_X1 _25967_ (
    .A1(_05456_),
    .A2(_05628_),
    .ZN(_05629_)
  );
  INV_X1 _25968_ (
    .A(_05629_),
    .ZN(_05630_)
  );
  AND2_X1 _25969_ (
    .A1(_05439_),
    .A2(_05458_),
    .ZN(_05631_)
  );
  INV_X1 _25970_ (
    .A(_05631_),
    .ZN(_05632_)
  );
  AND2_X1 _25971_ (
    .A1(_05630_),
    .A2(_05632_),
    .ZN(_05633_)
  );
  INV_X1 _25972_ (
    .A(_05633_),
    .ZN(_05634_)
  );
  AND2_X1 _25973_ (
    .A1(_05269_),
    .A2(_05634_),
    .ZN(_05635_)
  );
  AND2_X1 _25974_ (
    .A1(_05441_),
    .A2(_05635_),
    .ZN(_05636_)
  );
  INV_X1 _25975_ (
    .A(_05636_),
    .ZN(_05637_)
  );
  AND2_X1 _25976_ (
    .A1(_05620_),
    .A2(_05637_),
    .ZN(_00271_)
  );
  AND2_X1 _25977_ (
    .A1(_08056_),
    .A2(_05270_),
    .ZN(_05638_)
  );
  INV_X1 _25978_ (
    .A(_05638_),
    .ZN(_05639_)
  );
  AND2_X1 _25979_ (
    .A1(mem_reg_wdata[31]),
    .A2(_05259_),
    .ZN(_05640_)
  );
  INV_X1 _25980_ (
    .A(_05640_),
    .ZN(_05641_)
  );
  AND2_X1 _25981_ (
    .A1(wb_reg_wdata[31]),
    .A2(_05256_),
    .ZN(_05642_)
  );
  INV_X1 _25982_ (
    .A(_05642_),
    .ZN(_05643_)
  );
  AND2_X1 _25983_ (
    .A1(_05641_),
    .A2(_05643_),
    .ZN(_05644_)
  );
  INV_X1 _25984_ (
    .A(_05644_),
    .ZN(_05645_)
  );
  MUX2_X1 _25985_ (
    .A(_05645_),
    .B(io_dmem_resp_bits_data_word_bypass[31]),
    .S(_05255_),
    .Z(_05646_)
  );
  MUX2_X1 _25986_ (
    .A(ex_reg_rs_msb_1[29]),
    .B(_05646_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[31])
  );
  INV_X1 _25987_ (
    .A(_ex_op2_T[31]),
    .ZN(_05647_)
  );
  AND2_X1 _25988_ (
    .A1(_05456_),
    .A2(_05647_),
    .ZN(_05648_)
  );
  INV_X1 _25989_ (
    .A(_05648_),
    .ZN(_05649_)
  );
  AND2_X1 _25990_ (
    .A1(_05451_),
    .A2(_05458_),
    .ZN(_05650_)
  );
  INV_X1 _25991_ (
    .A(_05650_),
    .ZN(_05651_)
  );
  AND2_X1 _25992_ (
    .A1(_05649_),
    .A2(_05651_),
    .ZN(_05652_)
  );
  INV_X1 _25993_ (
    .A(_05652_),
    .ZN(_05653_)
  );
  AND2_X1 _25994_ (
    .A1(_05269_),
    .A2(_05653_),
    .ZN(_05654_)
  );
  AND2_X1 _25995_ (
    .A1(_05453_),
    .A2(_05654_),
    .ZN(_05655_)
  );
  INV_X1 _25996_ (
    .A(_05655_),
    .ZN(_05656_)
  );
  AND2_X1 _25997_ (
    .A1(_05639_),
    .A2(_05656_),
    .ZN(_00272_)
  );
  MUX2_X1 _25998_ (
    .A(mem_reg_wdata[0]),
    .B(alu_io_out[0]),
    .S(_05253_),
    .Z(_00273_)
  );
  MUX2_X1 _25999_ (
    .A(mem_reg_wdata[1]),
    .B(alu_io_out[1]),
    .S(_05253_),
    .Z(_00274_)
  );
  MUX2_X1 _26000_ (
    .A(mem_reg_wdata[2]),
    .B(alu_io_out[2]),
    .S(_05253_),
    .Z(_00275_)
  );
  MUX2_X1 _26001_ (
    .A(mem_reg_wdata[3]),
    .B(alu_io_out[3]),
    .S(_05253_),
    .Z(_00276_)
  );
  MUX2_X1 _26002_ (
    .A(mem_reg_wdata[4]),
    .B(alu_io_out[4]),
    .S(_05253_),
    .Z(_00277_)
  );
  MUX2_X1 _26003_ (
    .A(mem_reg_wdata[5]),
    .B(alu_io_out[5]),
    .S(_05253_),
    .Z(_00278_)
  );
  MUX2_X1 _26004_ (
    .A(mem_reg_wdata[6]),
    .B(alu_io_out[6]),
    .S(_05253_),
    .Z(_00279_)
  );
  MUX2_X1 _26005_ (
    .A(mem_reg_wdata[7]),
    .B(alu_io_out[7]),
    .S(_05253_),
    .Z(_00280_)
  );
  MUX2_X1 _26006_ (
    .A(mem_reg_wdata[8]),
    .B(alu_io_out[8]),
    .S(_05253_),
    .Z(_00281_)
  );
  MUX2_X1 _26007_ (
    .A(mem_reg_wdata[9]),
    .B(alu_io_out[9]),
    .S(_05253_),
    .Z(_00282_)
  );
  MUX2_X1 _26008_ (
    .A(mem_reg_wdata[10]),
    .B(alu_io_out[10]),
    .S(_05253_),
    .Z(_00283_)
  );
  MUX2_X1 _26009_ (
    .A(mem_reg_wdata[11]),
    .B(alu_io_out[11]),
    .S(_05253_),
    .Z(_00284_)
  );
  MUX2_X1 _26010_ (
    .A(mem_reg_wdata[12]),
    .B(alu_io_out[12]),
    .S(_05253_),
    .Z(_00285_)
  );
  MUX2_X1 _26011_ (
    .A(mem_reg_wdata[13]),
    .B(alu_io_out[13]),
    .S(_05253_),
    .Z(_00286_)
  );
  MUX2_X1 _26012_ (
    .A(mem_reg_wdata[14]),
    .B(alu_io_out[14]),
    .S(_05253_),
    .Z(_00287_)
  );
  MUX2_X1 _26013_ (
    .A(mem_reg_wdata[15]),
    .B(alu_io_out[15]),
    .S(_05253_),
    .Z(_00288_)
  );
  MUX2_X1 _26014_ (
    .A(mem_reg_wdata[16]),
    .B(alu_io_out[16]),
    .S(_05253_),
    .Z(_00289_)
  );
  MUX2_X1 _26015_ (
    .A(mem_reg_wdata[17]),
    .B(alu_io_out[17]),
    .S(_05253_),
    .Z(_00290_)
  );
  MUX2_X1 _26016_ (
    .A(mem_reg_wdata[18]),
    .B(alu_io_out[18]),
    .S(_05253_),
    .Z(_00291_)
  );
  MUX2_X1 _26017_ (
    .A(mem_reg_wdata[19]),
    .B(alu_io_out[19]),
    .S(_05253_),
    .Z(_00292_)
  );
  MUX2_X1 _26018_ (
    .A(mem_reg_wdata[20]),
    .B(alu_io_out[20]),
    .S(_05253_),
    .Z(_00293_)
  );
  MUX2_X1 _26019_ (
    .A(mem_reg_wdata[21]),
    .B(alu_io_out[21]),
    .S(_05253_),
    .Z(_00294_)
  );
  MUX2_X1 _26020_ (
    .A(mem_reg_wdata[22]),
    .B(alu_io_out[22]),
    .S(_05253_),
    .Z(_00295_)
  );
  MUX2_X1 _26021_ (
    .A(mem_reg_wdata[23]),
    .B(alu_io_out[23]),
    .S(_05253_),
    .Z(_00296_)
  );
  MUX2_X1 _26022_ (
    .A(mem_reg_wdata[24]),
    .B(alu_io_out[24]),
    .S(_05253_),
    .Z(_00297_)
  );
  MUX2_X1 _26023_ (
    .A(mem_reg_wdata[25]),
    .B(alu_io_out[25]),
    .S(_05253_),
    .Z(_00298_)
  );
  MUX2_X1 _26024_ (
    .A(mem_reg_wdata[26]),
    .B(alu_io_out[26]),
    .S(_05253_),
    .Z(_00299_)
  );
  MUX2_X1 _26025_ (
    .A(mem_reg_wdata[27]),
    .B(alu_io_out[27]),
    .S(_05253_),
    .Z(_00300_)
  );
  MUX2_X1 _26026_ (
    .A(mem_reg_wdata[28]),
    .B(alu_io_out[28]),
    .S(_05253_),
    .Z(_00301_)
  );
  MUX2_X1 _26027_ (
    .A(mem_reg_wdata[29]),
    .B(alu_io_out[29]),
    .S(_05253_),
    .Z(_00302_)
  );
  MUX2_X1 _26028_ (
    .A(mem_reg_wdata[30]),
    .B(alu_io_out[30]),
    .S(_05253_),
    .Z(_00303_)
  );
  MUX2_X1 _26029_ (
    .A(mem_reg_wdata[31]),
    .B(alu_io_out[31]),
    .S(_05253_),
    .Z(_00304_)
  );
  MUX2_X1 _26030_ (
    .A(mem_reg_raw_inst[0]),
    .B(ex_reg_raw_inst[0]),
    .S(_05253_),
    .Z(_00305_)
  );
  MUX2_X1 _26031_ (
    .A(mem_reg_raw_inst[1]),
    .B(ex_reg_raw_inst[1]),
    .S(_05253_),
    .Z(_00306_)
  );
  MUX2_X1 _26032_ (
    .A(mem_reg_raw_inst[2]),
    .B(ex_reg_raw_inst[2]),
    .S(_05253_),
    .Z(_00307_)
  );
  MUX2_X1 _26033_ (
    .A(mem_reg_raw_inst[3]),
    .B(ex_reg_raw_inst[3]),
    .S(_05253_),
    .Z(_00308_)
  );
  MUX2_X1 _26034_ (
    .A(mem_reg_raw_inst[4]),
    .B(ex_reg_raw_inst[4]),
    .S(_05253_),
    .Z(_00309_)
  );
  MUX2_X1 _26035_ (
    .A(mem_reg_raw_inst[5]),
    .B(ex_reg_raw_inst[5]),
    .S(_05253_),
    .Z(_00310_)
  );
  MUX2_X1 _26036_ (
    .A(mem_reg_raw_inst[6]),
    .B(ex_reg_raw_inst[6]),
    .S(_05253_),
    .Z(_00311_)
  );
  MUX2_X1 _26037_ (
    .A(mem_reg_raw_inst[7]),
    .B(ex_reg_raw_inst[7]),
    .S(_05253_),
    .Z(_00312_)
  );
  MUX2_X1 _26038_ (
    .A(mem_reg_raw_inst[8]),
    .B(ex_reg_raw_inst[8]),
    .S(_05253_),
    .Z(_00313_)
  );
  MUX2_X1 _26039_ (
    .A(mem_reg_raw_inst[9]),
    .B(ex_reg_raw_inst[9]),
    .S(_05253_),
    .Z(_00314_)
  );
  MUX2_X1 _26040_ (
    .A(mem_reg_raw_inst[10]),
    .B(ex_reg_raw_inst[10]),
    .S(_05253_),
    .Z(_00315_)
  );
  MUX2_X1 _26041_ (
    .A(mem_reg_raw_inst[11]),
    .B(ex_reg_raw_inst[11]),
    .S(_05253_),
    .Z(_00316_)
  );
  MUX2_X1 _26042_ (
    .A(mem_reg_raw_inst[12]),
    .B(ex_reg_raw_inst[12]),
    .S(_05253_),
    .Z(_00317_)
  );
  MUX2_X1 _26043_ (
    .A(mem_reg_raw_inst[13]),
    .B(ex_reg_raw_inst[13]),
    .S(_05253_),
    .Z(_00318_)
  );
  MUX2_X1 _26044_ (
    .A(mem_reg_raw_inst[14]),
    .B(ex_reg_raw_inst[14]),
    .S(_05253_),
    .Z(_00319_)
  );
  MUX2_X1 _26045_ (
    .A(mem_reg_raw_inst[15]),
    .B(ex_reg_raw_inst[15]),
    .S(_05253_),
    .Z(_00320_)
  );
  MUX2_X1 _26046_ (
    .A(mem_reg_inst[7]),
    .B(ex_reg_inst[7]),
    .S(_05253_),
    .Z(_00321_)
  );
  MUX2_X1 _26047_ (
    .A(mem_reg_inst[8]),
    .B(ex_reg_inst[8]),
    .S(_05253_),
    .Z(_00322_)
  );
  MUX2_X1 _26048_ (
    .A(mem_reg_inst[9]),
    .B(ex_reg_inst[9]),
    .S(_05253_),
    .Z(_00323_)
  );
  MUX2_X1 _26049_ (
    .A(mem_reg_inst[10]),
    .B(ex_reg_inst[10]),
    .S(_05253_),
    .Z(_00324_)
  );
  MUX2_X1 _26050_ (
    .A(mem_reg_inst[11]),
    .B(ex_reg_inst[11]),
    .S(_05253_),
    .Z(_00325_)
  );
  MUX2_X1 _26051_ (
    .A(mem_reg_inst[12]),
    .B(ex_reg_inst[12]),
    .S(_05253_),
    .Z(_00326_)
  );
  MUX2_X1 _26052_ (
    .A(mem_reg_inst[13]),
    .B(ex_reg_inst[13]),
    .S(_05253_),
    .Z(_00327_)
  );
  MUX2_X1 _26053_ (
    .A(mem_reg_inst[14]),
    .B(ex_reg_inst[14]),
    .S(_05253_),
    .Z(_00328_)
  );
  MUX2_X1 _26054_ (
    .A(mem_reg_inst[15]),
    .B(ex_reg_inst[15]),
    .S(_05253_),
    .Z(_00329_)
  );
  MUX2_X1 _26055_ (
    .A(mem_reg_inst[16]),
    .B(ex_reg_inst[16]),
    .S(_05253_),
    .Z(_00330_)
  );
  MUX2_X1 _26056_ (
    .A(mem_reg_inst[17]),
    .B(ex_reg_inst[17]),
    .S(_05253_),
    .Z(_00331_)
  );
  MUX2_X1 _26057_ (
    .A(mem_reg_inst[18]),
    .B(ex_reg_inst[18]),
    .S(_05253_),
    .Z(_00332_)
  );
  MUX2_X1 _26058_ (
    .A(mem_reg_inst[19]),
    .B(ex_reg_inst[19]),
    .S(_05253_),
    .Z(_00333_)
  );
  MUX2_X1 _26059_ (
    .A(mem_reg_inst[20]),
    .B(ex_reg_inst[20]),
    .S(_05253_),
    .Z(_00334_)
  );
  MUX2_X1 _26060_ (
    .A(mem_reg_inst[21]),
    .B(ex_reg_inst[21]),
    .S(_05253_),
    .Z(_00335_)
  );
  MUX2_X1 _26061_ (
    .A(mem_reg_inst[22]),
    .B(ex_reg_inst[22]),
    .S(_05253_),
    .Z(_00336_)
  );
  MUX2_X1 _26062_ (
    .A(mem_reg_inst[23]),
    .B(ex_reg_inst[23]),
    .S(_05253_),
    .Z(_00337_)
  );
  MUX2_X1 _26063_ (
    .A(mem_reg_inst[24]),
    .B(ex_reg_inst[24]),
    .S(_05253_),
    .Z(_00338_)
  );
  MUX2_X1 _26064_ (
    .A(mem_reg_inst[25]),
    .B(ex_reg_inst[25]),
    .S(_05253_),
    .Z(_00339_)
  );
  MUX2_X1 _26065_ (
    .A(mem_reg_inst[26]),
    .B(ex_reg_inst[26]),
    .S(_05253_),
    .Z(_00340_)
  );
  MUX2_X1 _26066_ (
    .A(mem_reg_inst[27]),
    .B(ex_reg_inst[27]),
    .S(_05253_),
    .Z(_00341_)
  );
  MUX2_X1 _26067_ (
    .A(mem_reg_inst[28]),
    .B(ex_reg_inst[28]),
    .S(_05253_),
    .Z(_00342_)
  );
  MUX2_X1 _26068_ (
    .A(mem_reg_inst[29]),
    .B(ex_reg_inst[29]),
    .S(_05253_),
    .Z(_00343_)
  );
  MUX2_X1 _26069_ (
    .A(mem_reg_inst[30]),
    .B(ex_reg_inst[30]),
    .S(_05253_),
    .Z(_00344_)
  );
  MUX2_X1 _26070_ (
    .A(mem_reg_inst[31]),
    .B(ex_reg_inst[31]),
    .S(_05253_),
    .Z(_00345_)
  );
  MUX2_X1 _26071_ (
    .A(mem_reg_pc[0]),
    .B(ex_reg_pc[0]),
    .S(_05253_),
    .Z(_00346_)
  );
  MUX2_X1 _26072_ (
    .A(mem_reg_pc[1]),
    .B(ex_reg_pc[1]),
    .S(_05253_),
    .Z(_00347_)
  );
  MUX2_X1 _26073_ (
    .A(mem_reg_pc[2]),
    .B(ex_reg_pc[2]),
    .S(_05253_),
    .Z(_00348_)
  );
  MUX2_X1 _26074_ (
    .A(mem_reg_pc[3]),
    .B(ex_reg_pc[3]),
    .S(_05253_),
    .Z(_00349_)
  );
  MUX2_X1 _26075_ (
    .A(mem_reg_pc[4]),
    .B(ex_reg_pc[4]),
    .S(_05253_),
    .Z(_00350_)
  );
  MUX2_X1 _26076_ (
    .A(mem_reg_pc[5]),
    .B(ex_reg_pc[5]),
    .S(_05253_),
    .Z(_00351_)
  );
  MUX2_X1 _26077_ (
    .A(mem_reg_pc[6]),
    .B(ex_reg_pc[6]),
    .S(_05253_),
    .Z(_00352_)
  );
  MUX2_X1 _26078_ (
    .A(mem_reg_pc[7]),
    .B(ex_reg_pc[7]),
    .S(_05253_),
    .Z(_00353_)
  );
  MUX2_X1 _26079_ (
    .A(mem_reg_pc[8]),
    .B(ex_reg_pc[8]),
    .S(_05253_),
    .Z(_00354_)
  );
  MUX2_X1 _26080_ (
    .A(mem_reg_pc[9]),
    .B(ex_reg_pc[9]),
    .S(_05253_),
    .Z(_00355_)
  );
  MUX2_X1 _26081_ (
    .A(mem_reg_pc[10]),
    .B(ex_reg_pc[10]),
    .S(_05253_),
    .Z(_00356_)
  );
  MUX2_X1 _26082_ (
    .A(mem_reg_pc[11]),
    .B(ex_reg_pc[11]),
    .S(_05253_),
    .Z(_00357_)
  );
  MUX2_X1 _26083_ (
    .A(mem_reg_pc[12]),
    .B(ex_reg_pc[12]),
    .S(_05253_),
    .Z(_00358_)
  );
  MUX2_X1 _26084_ (
    .A(mem_reg_pc[13]),
    .B(ex_reg_pc[13]),
    .S(_05253_),
    .Z(_00359_)
  );
  MUX2_X1 _26085_ (
    .A(mem_reg_pc[14]),
    .B(ex_reg_pc[14]),
    .S(_05253_),
    .Z(_00360_)
  );
  MUX2_X1 _26086_ (
    .A(mem_reg_pc[15]),
    .B(ex_reg_pc[15]),
    .S(_05253_),
    .Z(_00361_)
  );
  MUX2_X1 _26087_ (
    .A(mem_reg_pc[16]),
    .B(ex_reg_pc[16]),
    .S(_05253_),
    .Z(_00362_)
  );
  MUX2_X1 _26088_ (
    .A(mem_reg_pc[17]),
    .B(ex_reg_pc[17]),
    .S(_05253_),
    .Z(_00363_)
  );
  MUX2_X1 _26089_ (
    .A(mem_reg_pc[18]),
    .B(ex_reg_pc[18]),
    .S(_05253_),
    .Z(_00364_)
  );
  MUX2_X1 _26090_ (
    .A(mem_reg_pc[19]),
    .B(ex_reg_pc[19]),
    .S(_05253_),
    .Z(_00365_)
  );
  MUX2_X1 _26091_ (
    .A(mem_reg_pc[20]),
    .B(ex_reg_pc[20]),
    .S(_05253_),
    .Z(_00366_)
  );
  MUX2_X1 _26092_ (
    .A(mem_reg_pc[21]),
    .B(ex_reg_pc[21]),
    .S(_05253_),
    .Z(_00367_)
  );
  MUX2_X1 _26093_ (
    .A(mem_reg_pc[22]),
    .B(ex_reg_pc[22]),
    .S(_05253_),
    .Z(_00368_)
  );
  MUX2_X1 _26094_ (
    .A(mem_reg_pc[23]),
    .B(ex_reg_pc[23]),
    .S(_05253_),
    .Z(_00369_)
  );
  MUX2_X1 _26095_ (
    .A(mem_reg_pc[24]),
    .B(ex_reg_pc[24]),
    .S(_05253_),
    .Z(_00370_)
  );
  MUX2_X1 _26096_ (
    .A(mem_reg_pc[25]),
    .B(ex_reg_pc[25]),
    .S(_05253_),
    .Z(_00371_)
  );
  MUX2_X1 _26097_ (
    .A(mem_reg_pc[26]),
    .B(ex_reg_pc[26]),
    .S(_05253_),
    .Z(_00372_)
  );
  MUX2_X1 _26098_ (
    .A(mem_reg_pc[27]),
    .B(ex_reg_pc[27]),
    .S(_05253_),
    .Z(_00373_)
  );
  MUX2_X1 _26099_ (
    .A(mem_reg_pc[28]),
    .B(ex_reg_pc[28]),
    .S(_05253_),
    .Z(_00374_)
  );
  MUX2_X1 _26100_ (
    .A(mem_reg_pc[29]),
    .B(ex_reg_pc[29]),
    .S(_05253_),
    .Z(_00375_)
  );
  MUX2_X1 _26101_ (
    .A(mem_reg_pc[30]),
    .B(ex_reg_pc[30]),
    .S(_05253_),
    .Z(_00376_)
  );
  MUX2_X1 _26102_ (
    .A(mem_reg_pc[31]),
    .B(ex_reg_pc[31]),
    .S(_05253_),
    .Z(_00377_)
  );
  AND2_X1 _26103_ (
    .A1(mem_reg_store),
    .A2(_05254_),
    .ZN(_05657_)
  );
  INV_X1 _26104_ (
    .A(_05657_),
    .ZN(_05658_)
  );
  AND2_X1 _26105_ (
    .A1(ex_ctrl_mem_cmd[2]),
    .A2(_00025_),
    .ZN(_05659_)
  );
  INV_X1 _26106_ (
    .A(_05659_),
    .ZN(_05660_)
  );
  AND2_X1 _26107_ (
    .A1(_08556_),
    .A2(_05660_),
    .ZN(_05661_)
  );
  INV_X1 _26108_ (
    .A(_05661_),
    .ZN(_05662_)
  );
  AND2_X1 _26109_ (
    .A1(_08213_),
    .A2(_08555_),
    .ZN(_05663_)
  );
  AND2_X1 _26110_ (
    .A1(_08210_),
    .A2(_08211_),
    .ZN(_05664_)
  );
  AND2_X1 _26111_ (
    .A1(_05663_),
    .A2(_05664_),
    .ZN(_05665_)
  );
  INV_X1 _26112_ (
    .A(_05665_),
    .ZN(_05666_)
  );
  AND2_X1 _26113_ (
    .A1(_05662_),
    .A2(_05666_),
    .ZN(_05667_)
  );
  INV_X1 _26114_ (
    .A(_05667_),
    .ZN(_05668_)
  );
  AND2_X1 _26115_ (
    .A1(ex_ctrl_mem_cmd[0]),
    .A2(_00027_),
    .ZN(_05669_)
  );
  INV_X1 _26116_ (
    .A(_05669_),
    .ZN(_05670_)
  );
  AND2_X1 _26117_ (
    .A1(ex_ctrl_mem_cmd[1]),
    .A2(_00026_),
    .ZN(_05671_)
  );
  INV_X1 _26118_ (
    .A(_05671_),
    .ZN(_05672_)
  );
  AND2_X1 _26119_ (
    .A1(_05670_),
    .A2(_05672_),
    .ZN(_05673_)
  );
  AND2_X1 _26120_ (
    .A1(_05668_),
    .A2(_05673_),
    .ZN(_05674_)
  );
  INV_X1 _26121_ (
    .A(_05674_),
    .ZN(_05675_)
  );
  AND2_X1 _26122_ (
    .A1(_08554_),
    .A2(_05663_),
    .ZN(_05676_)
  );
  INV_X1 _26123_ (
    .A(_05676_),
    .ZN(_05677_)
  );
  AND2_X1 _26124_ (
    .A1(_08212_),
    .A2(_08213_),
    .ZN(_05678_)
  );
  AND2_X1 _26125_ (
    .A1(_08211_),
    .A2(_05678_),
    .ZN(_05679_)
  );
  INV_X1 _26126_ (
    .A(_05679_),
    .ZN(_05680_)
  );
  AND2_X1 _26127_ (
    .A1(_05677_),
    .A2(_05680_),
    .ZN(_05681_)
  );
  INV_X1 _26128_ (
    .A(_05681_),
    .ZN(_05682_)
  );
  AND2_X1 _26129_ (
    .A1(_08553_),
    .A2(_05682_),
    .ZN(_05683_)
  );
  INV_X1 _26130_ (
    .A(_05683_),
    .ZN(_05684_)
  );
  AND2_X1 _26131_ (
    .A1(_05675_),
    .A2(_05684_),
    .ZN(_05685_)
  );
  INV_X1 _26132_ (
    .A(_05685_),
    .ZN(_05686_)
  );
  AND2_X1 _26133_ (
    .A1(_05268_),
    .A2(_05686_),
    .ZN(_05687_)
  );
  INV_X1 _26134_ (
    .A(_05687_),
    .ZN(_05688_)
  );
  AND2_X1 _26135_ (
    .A1(_05658_),
    .A2(_05688_),
    .ZN(_05689_)
  );
  INV_X1 _26136_ (
    .A(_05689_),
    .ZN(_00378_)
  );
  AND2_X1 _26137_ (
    .A1(mem_reg_load),
    .A2(_05254_),
    .ZN(_05690_)
  );
  INV_X1 _26138_ (
    .A(_05690_),
    .ZN(_05691_)
  );
  AND2_X1 _26139_ (
    .A1(_08210_),
    .A2(_05682_),
    .ZN(_05692_)
  );
  INV_X1 _26140_ (
    .A(_05692_),
    .ZN(_05693_)
  );
  AND2_X1 _26141_ (
    .A1(_08553_),
    .A2(_05676_),
    .ZN(_05694_)
  );
  INV_X1 _26142_ (
    .A(_05694_),
    .ZN(_05695_)
  );
  AND2_X1 _26143_ (
    .A1(_05675_),
    .A2(_05695_),
    .ZN(_05696_)
  );
  AND2_X1 _26144_ (
    .A1(_05693_),
    .A2(_05696_),
    .ZN(_05697_)
  );
  INV_X1 _26145_ (
    .A(_05697_),
    .ZN(_05698_)
  );
  AND2_X1 _26146_ (
    .A1(_05268_),
    .A2(_05698_),
    .ZN(_05699_)
  );
  INV_X1 _26147_ (
    .A(_05699_),
    .ZN(_05700_)
  );
  AND2_X1 _26148_ (
    .A1(_05691_),
    .A2(_05700_),
    .ZN(_05701_)
  );
  INV_X1 _26149_ (
    .A(_05701_),
    .ZN(_00379_)
  );
  AND2_X1 _26150_ (
    .A1(_08621_),
    .A2(_05695_),
    .ZN(_05702_)
  );
  INV_X1 _26151_ (
    .A(_05702_),
    .ZN(_05703_)
  );
  MUX2_X1 _26152_ (
    .A(mem_reg_slow_bypass),
    .B(_05703_),
    .S(_05253_),
    .Z(_00380_)
  );
  MUX2_X1 _26153_ (
    .A(mem_reg_cause[0]),
    .B(ex_reg_cause[0]),
    .S(_05253_),
    .Z(_00381_)
  );
  MUX2_X1 _26154_ (
    .A(mem_reg_cause[1]),
    .B(ex_reg_cause[1]),
    .S(_05253_),
    .Z(_00382_)
  );
  MUX2_X1 _26155_ (
    .A(mem_reg_cause[2]),
    .B(ex_reg_cause[2]),
    .S(_05253_),
    .Z(_00383_)
  );
  MUX2_X1 _26156_ (
    .A(mem_reg_cause[3]),
    .B(ex_reg_cause[3]),
    .S(_05253_),
    .Z(_00384_)
  );
  MUX2_X1 _26157_ (
    .A(mem_reg_cause[4]),
    .B(ex_reg_cause[4]),
    .S(_05253_),
    .Z(_00385_)
  );
  MUX2_X1 _26158_ (
    .A(mem_reg_cause[5]),
    .B(ex_reg_cause[5]),
    .S(_05253_),
    .Z(_00386_)
  );
  MUX2_X1 _26159_ (
    .A(mem_reg_cause[6]),
    .B(ex_reg_cause[6]),
    .S(_05253_),
    .Z(_00387_)
  );
  MUX2_X1 _26160_ (
    .A(mem_reg_cause[7]),
    .B(ex_reg_cause[7]),
    .S(_05253_),
    .Z(_00388_)
  );
  MUX2_X1 _26161_ (
    .A(mem_reg_cause[8]),
    .B(ex_reg_cause[8]),
    .S(_05253_),
    .Z(_00389_)
  );
  MUX2_X1 _26162_ (
    .A(mem_reg_cause[9]),
    .B(ex_reg_cause[9]),
    .S(_05253_),
    .Z(_00390_)
  );
  MUX2_X1 _26163_ (
    .A(mem_reg_cause[10]),
    .B(ex_reg_cause[10]),
    .S(_05253_),
    .Z(_00391_)
  );
  MUX2_X1 _26164_ (
    .A(mem_reg_cause[11]),
    .B(ex_reg_cause[11]),
    .S(_05253_),
    .Z(_00392_)
  );
  MUX2_X1 _26165_ (
    .A(mem_reg_cause[12]),
    .B(ex_reg_cause[12]),
    .S(_05253_),
    .Z(_00393_)
  );
  MUX2_X1 _26166_ (
    .A(mem_reg_cause[13]),
    .B(ex_reg_cause[13]),
    .S(_05253_),
    .Z(_00394_)
  );
  MUX2_X1 _26167_ (
    .A(mem_reg_cause[14]),
    .B(ex_reg_cause[14]),
    .S(_05253_),
    .Z(_00395_)
  );
  MUX2_X1 _26168_ (
    .A(mem_reg_cause[15]),
    .B(ex_reg_cause[15]),
    .S(_05253_),
    .Z(_00396_)
  );
  MUX2_X1 _26169_ (
    .A(mem_reg_cause[16]),
    .B(ex_reg_cause[16]),
    .S(_05253_),
    .Z(_00397_)
  );
  MUX2_X1 _26170_ (
    .A(mem_reg_cause[17]),
    .B(ex_reg_cause[17]),
    .S(_05253_),
    .Z(_00398_)
  );
  MUX2_X1 _26171_ (
    .A(mem_reg_cause[18]),
    .B(ex_reg_cause[18]),
    .S(_05253_),
    .Z(_00399_)
  );
  MUX2_X1 _26172_ (
    .A(mem_reg_cause[19]),
    .B(ex_reg_cause[19]),
    .S(_05253_),
    .Z(_00400_)
  );
  MUX2_X1 _26173_ (
    .A(mem_reg_cause[20]),
    .B(ex_reg_cause[20]),
    .S(_05253_),
    .Z(_00401_)
  );
  MUX2_X1 _26174_ (
    .A(mem_reg_cause[21]),
    .B(ex_reg_cause[21]),
    .S(_05253_),
    .Z(_00402_)
  );
  MUX2_X1 _26175_ (
    .A(mem_reg_cause[22]),
    .B(ex_reg_cause[22]),
    .S(_05253_),
    .Z(_00403_)
  );
  MUX2_X1 _26176_ (
    .A(mem_reg_cause[23]),
    .B(ex_reg_cause[23]),
    .S(_05253_),
    .Z(_00404_)
  );
  MUX2_X1 _26177_ (
    .A(mem_reg_cause[24]),
    .B(ex_reg_cause[24]),
    .S(_05253_),
    .Z(_00405_)
  );
  MUX2_X1 _26178_ (
    .A(mem_reg_cause[25]),
    .B(ex_reg_cause[25]),
    .S(_05253_),
    .Z(_00406_)
  );
  MUX2_X1 _26179_ (
    .A(mem_reg_cause[26]),
    .B(ex_reg_cause[26]),
    .S(_05253_),
    .Z(_00407_)
  );
  MUX2_X1 _26180_ (
    .A(mem_reg_cause[27]),
    .B(ex_reg_cause[27]),
    .S(_05253_),
    .Z(_00408_)
  );
  MUX2_X1 _26181_ (
    .A(mem_reg_cause[28]),
    .B(ex_reg_cause[28]),
    .S(_05253_),
    .Z(_00409_)
  );
  MUX2_X1 _26182_ (
    .A(mem_reg_cause[29]),
    .B(ex_reg_cause[29]),
    .S(_05253_),
    .Z(_00410_)
  );
  MUX2_X1 _26183_ (
    .A(mem_reg_cause[30]),
    .B(ex_reg_cause[30]),
    .S(_05253_),
    .Z(_00411_)
  );
  MUX2_X1 _26184_ (
    .A(mem_reg_cause[31]),
    .B(ex_reg_cause[31]),
    .S(_05253_),
    .Z(_00412_)
  );
  AND2_X1 _26185_ (
    .A1(ex_ctrl_jalr),
    .A2(bpu_io_status_debug),
    .ZN(_05704_)
  );
  INV_X1 _26186_ (
    .A(_05704_),
    .ZN(_05705_)
  );
  AND2_X1 _26187_ (
    .A1(_08187_),
    .A2(_05705_),
    .ZN(_05706_)
  );
  INV_X1 _26188_ (
    .A(_05706_),
    .ZN(_05707_)
  );
  MUX2_X1 _26189_ (
    .A(mem_reg_flush_pipe),
    .B(_05707_),
    .S(_05253_),
    .Z(_00413_)
  );
  MUX2_X1 _26190_ (
    .A(mem_reg_rvc),
    .B(ex_reg_rvc),
    .S(_05253_),
    .Z(_00414_)
  );
  AND2_X1 _26191_ (
    .A1(_09298_),
    .A2(_10245_),
    .ZN(_05708_)
  );
  MUX2_X1 _26192_ (
    .A(ibuf_io_inst_0_bits_raw[0]),
    .B(ex_reg_raw_inst[0]),
    .S(_05708_),
    .Z(_00415_)
  );
  MUX2_X1 _26193_ (
    .A(ibuf_io_inst_0_bits_raw[1]),
    .B(ex_reg_raw_inst[1]),
    .S(_05708_),
    .Z(_00416_)
  );
  MUX2_X1 _26194_ (
    .A(ibuf_io_inst_0_bits_raw[2]),
    .B(ex_reg_raw_inst[2]),
    .S(_05708_),
    .Z(_00417_)
  );
  MUX2_X1 _26195_ (
    .A(ibuf_io_inst_0_bits_raw[3]),
    .B(ex_reg_raw_inst[3]),
    .S(_05708_),
    .Z(_00418_)
  );
  MUX2_X1 _26196_ (
    .A(ibuf_io_inst_0_bits_raw[4]),
    .B(ex_reg_raw_inst[4]),
    .S(_05708_),
    .Z(_00419_)
  );
  MUX2_X1 _26197_ (
    .A(ibuf_io_inst_0_bits_raw[5]),
    .B(ex_reg_raw_inst[5]),
    .S(_05708_),
    .Z(_00420_)
  );
  MUX2_X1 _26198_ (
    .A(ibuf_io_inst_0_bits_raw[6]),
    .B(ex_reg_raw_inst[6]),
    .S(_05708_),
    .Z(_00421_)
  );
  MUX2_X1 _26199_ (
    .A(ibuf_io_inst_0_bits_raw[7]),
    .B(ex_reg_raw_inst[7]),
    .S(_05708_),
    .Z(_00422_)
  );
  MUX2_X1 _26200_ (
    .A(ibuf_io_inst_0_bits_raw[8]),
    .B(ex_reg_raw_inst[8]),
    .S(_05708_),
    .Z(_00423_)
  );
  MUX2_X1 _26201_ (
    .A(ibuf_io_inst_0_bits_raw[9]),
    .B(ex_reg_raw_inst[9]),
    .S(_05708_),
    .Z(_00424_)
  );
  MUX2_X1 _26202_ (
    .A(ibuf_io_inst_0_bits_raw[10]),
    .B(ex_reg_raw_inst[10]),
    .S(_05708_),
    .Z(_00425_)
  );
  MUX2_X1 _26203_ (
    .A(ibuf_io_inst_0_bits_raw[11]),
    .B(ex_reg_raw_inst[11]),
    .S(_05708_),
    .Z(_00426_)
  );
  MUX2_X1 _26204_ (
    .A(ibuf_io_inst_0_bits_raw[12]),
    .B(ex_reg_raw_inst[12]),
    .S(_05708_),
    .Z(_00427_)
  );
  MUX2_X1 _26205_ (
    .A(ibuf_io_inst_0_bits_raw[13]),
    .B(ex_reg_raw_inst[13]),
    .S(_05708_),
    .Z(_00428_)
  );
  MUX2_X1 _26206_ (
    .A(ibuf_io_inst_0_bits_raw[14]),
    .B(ex_reg_raw_inst[14]),
    .S(_05708_),
    .Z(_00429_)
  );
  MUX2_X1 _26207_ (
    .A(ibuf_io_inst_0_bits_raw[15]),
    .B(ex_reg_raw_inst[15]),
    .S(_05708_),
    .Z(_00430_)
  );
  MUX2_X1 _26208_ (
    .A(csr_io_decode_0_inst[7]),
    .B(ex_reg_inst[7]),
    .S(_05708_),
    .Z(_00431_)
  );
  MUX2_X1 _26209_ (
    .A(csr_io_decode_0_inst[8]),
    .B(ex_reg_inst[8]),
    .S(_05708_),
    .Z(_00432_)
  );
  MUX2_X1 _26210_ (
    .A(csr_io_decode_0_inst[9]),
    .B(ex_reg_inst[9]),
    .S(_05708_),
    .Z(_00433_)
  );
  MUX2_X1 _26211_ (
    .A(csr_io_decode_0_inst[10]),
    .B(ex_reg_inst[10]),
    .S(_05708_),
    .Z(_00434_)
  );
  MUX2_X1 _26212_ (
    .A(csr_io_decode_0_inst[11]),
    .B(ex_reg_inst[11]),
    .S(_05708_),
    .Z(_00435_)
  );
  MUX2_X1 _26213_ (
    .A(csr_io_decode_0_inst[12]),
    .B(ex_reg_inst[12]),
    .S(_05708_),
    .Z(_00436_)
  );
  MUX2_X1 _26214_ (
    .A(csr_io_decode_0_inst[13]),
    .B(ex_reg_inst[13]),
    .S(_05708_),
    .Z(_00437_)
  );
  MUX2_X1 _26215_ (
    .A(csr_io_decode_0_inst[14]),
    .B(ex_reg_inst[14]),
    .S(_05708_),
    .Z(_00438_)
  );
  MUX2_X1 _26216_ (
    .A(csr_io_decode_0_inst[15]),
    .B(ex_reg_inst[15]),
    .S(_05708_),
    .Z(_00439_)
  );
  MUX2_X1 _26217_ (
    .A(csr_io_decode_0_inst[16]),
    .B(ex_reg_inst[16]),
    .S(_05708_),
    .Z(_00440_)
  );
  MUX2_X1 _26218_ (
    .A(csr_io_decode_0_inst[17]),
    .B(ex_reg_inst[17]),
    .S(_05708_),
    .Z(_00441_)
  );
  MUX2_X1 _26219_ (
    .A(csr_io_decode_0_inst[18]),
    .B(ex_reg_inst[18]),
    .S(_05708_),
    .Z(_00442_)
  );
  MUX2_X1 _26220_ (
    .A(csr_io_decode_0_inst[19]),
    .B(ex_reg_inst[19]),
    .S(_05708_),
    .Z(_00443_)
  );
  MUX2_X1 _26221_ (
    .A(csr_io_decode_0_inst[20]),
    .B(ex_reg_inst[20]),
    .S(_05708_),
    .Z(_00444_)
  );
  MUX2_X1 _26222_ (
    .A(csr_io_decode_0_inst[21]),
    .B(ex_reg_inst[21]),
    .S(_05708_),
    .Z(_00445_)
  );
  MUX2_X1 _26223_ (
    .A(csr_io_decode_0_inst[22]),
    .B(ex_reg_inst[22]),
    .S(_05708_),
    .Z(_00446_)
  );
  MUX2_X1 _26224_ (
    .A(csr_io_decode_0_inst[23]),
    .B(ex_reg_inst[23]),
    .S(_05708_),
    .Z(_00447_)
  );
  MUX2_X1 _26225_ (
    .A(csr_io_decode_0_inst[24]),
    .B(ex_reg_inst[24]),
    .S(_05708_),
    .Z(_00448_)
  );
  MUX2_X1 _26226_ (
    .A(csr_io_decode_0_inst[25]),
    .B(ex_reg_inst[25]),
    .S(_05708_),
    .Z(_00449_)
  );
  MUX2_X1 _26227_ (
    .A(csr_io_decode_0_inst[26]),
    .B(ex_reg_inst[26]),
    .S(_05708_),
    .Z(_00450_)
  );
  MUX2_X1 _26228_ (
    .A(csr_io_decode_0_inst[27]),
    .B(ex_reg_inst[27]),
    .S(_05708_),
    .Z(_00451_)
  );
  MUX2_X1 _26229_ (
    .A(csr_io_decode_0_inst[28]),
    .B(ex_reg_inst[28]),
    .S(_05708_),
    .Z(_00452_)
  );
  MUX2_X1 _26230_ (
    .A(csr_io_decode_0_inst[29]),
    .B(ex_reg_inst[29]),
    .S(_05708_),
    .Z(_00453_)
  );
  MUX2_X1 _26231_ (
    .A(csr_io_decode_0_inst[30]),
    .B(ex_reg_inst[30]),
    .S(_05708_),
    .Z(_00454_)
  );
  MUX2_X1 _26232_ (
    .A(csr_io_decode_0_inst[31]),
    .B(ex_reg_inst[31]),
    .S(_05708_),
    .Z(_00455_)
  );
  MUX2_X1 _26233_ (
    .A(ex_reg_mem_size[0]),
    .B(csr_io_decode_0_inst[12]),
    .S(_10244_),
    .Z(_00456_)
  );
  MUX2_X1 _26234_ (
    .A(ex_reg_mem_size[1]),
    .B(csr_io_decode_0_inst[13]),
    .S(_10244_),
    .Z(_00457_)
  );
  AND2_X1 _26235_ (
    .A1(ex_reg_cause[5]),
    .A2(_05708_),
    .ZN(_05709_)
  );
  INV_X1 _26236_ (
    .A(_05709_),
    .ZN(_05710_)
  );
  AND2_X1 _26237_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[5]),
    .ZN(_05711_)
  );
  INV_X1 _26238_ (
    .A(_05711_),
    .ZN(_05712_)
  );
  AND2_X1 _26239_ (
    .A1(_05710_),
    .A2(_05712_),
    .ZN(_05713_)
  );
  INV_X1 _26240_ (
    .A(_05713_),
    .ZN(_00458_)
  );
  AND2_X1 _26241_ (
    .A1(ex_reg_cause[6]),
    .A2(_05708_),
    .ZN(_05714_)
  );
  INV_X1 _26242_ (
    .A(_05714_),
    .ZN(_05715_)
  );
  AND2_X1 _26243_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[6]),
    .ZN(_05716_)
  );
  INV_X1 _26244_ (
    .A(_05716_),
    .ZN(_05717_)
  );
  AND2_X1 _26245_ (
    .A1(_05715_),
    .A2(_05717_),
    .ZN(_05718_)
  );
  INV_X1 _26246_ (
    .A(_05718_),
    .ZN(_00459_)
  );
  AND2_X1 _26247_ (
    .A1(ex_reg_cause[7]),
    .A2(_05708_),
    .ZN(_05719_)
  );
  INV_X1 _26248_ (
    .A(_05719_),
    .ZN(_05720_)
  );
  AND2_X1 _26249_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[7]),
    .ZN(_05721_)
  );
  INV_X1 _26250_ (
    .A(_05721_),
    .ZN(_05722_)
  );
  AND2_X1 _26251_ (
    .A1(_05720_),
    .A2(_05722_),
    .ZN(_05723_)
  );
  INV_X1 _26252_ (
    .A(_05723_),
    .ZN(_00460_)
  );
  AND2_X1 _26253_ (
    .A1(ex_reg_cause[8]),
    .A2(_05708_),
    .ZN(_05724_)
  );
  INV_X1 _26254_ (
    .A(_05724_),
    .ZN(_05725_)
  );
  AND2_X1 _26255_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[8]),
    .ZN(_05726_)
  );
  INV_X1 _26256_ (
    .A(_05726_),
    .ZN(_05727_)
  );
  AND2_X1 _26257_ (
    .A1(_05725_),
    .A2(_05727_),
    .ZN(_05728_)
  );
  INV_X1 _26258_ (
    .A(_05728_),
    .ZN(_00461_)
  );
  AND2_X1 _26259_ (
    .A1(ex_reg_cause[9]),
    .A2(_05708_),
    .ZN(_05729_)
  );
  INV_X1 _26260_ (
    .A(_05729_),
    .ZN(_05730_)
  );
  AND2_X1 _26261_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[9]),
    .ZN(_05731_)
  );
  INV_X1 _26262_ (
    .A(_05731_),
    .ZN(_05732_)
  );
  AND2_X1 _26263_ (
    .A1(_05730_),
    .A2(_05732_),
    .ZN(_05733_)
  );
  INV_X1 _26264_ (
    .A(_05733_),
    .ZN(_00462_)
  );
  AND2_X1 _26265_ (
    .A1(ex_reg_cause[10]),
    .A2(_05708_),
    .ZN(_05734_)
  );
  INV_X1 _26266_ (
    .A(_05734_),
    .ZN(_05735_)
  );
  AND2_X1 _26267_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[10]),
    .ZN(_05736_)
  );
  INV_X1 _26268_ (
    .A(_05736_),
    .ZN(_05737_)
  );
  AND2_X1 _26269_ (
    .A1(_05735_),
    .A2(_05737_),
    .ZN(_05738_)
  );
  INV_X1 _26270_ (
    .A(_05738_),
    .ZN(_00463_)
  );
  AND2_X1 _26271_ (
    .A1(ex_reg_cause[11]),
    .A2(_05708_),
    .ZN(_05739_)
  );
  INV_X1 _26272_ (
    .A(_05739_),
    .ZN(_05740_)
  );
  AND2_X1 _26273_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[11]),
    .ZN(_05741_)
  );
  INV_X1 _26274_ (
    .A(_05741_),
    .ZN(_05742_)
  );
  AND2_X1 _26275_ (
    .A1(_05740_),
    .A2(_05742_),
    .ZN(_05743_)
  );
  INV_X1 _26276_ (
    .A(_05743_),
    .ZN(_00464_)
  );
  AND2_X1 _26277_ (
    .A1(ex_reg_cause[12]),
    .A2(_05708_),
    .ZN(_05744_)
  );
  INV_X1 _26278_ (
    .A(_05744_),
    .ZN(_05745_)
  );
  AND2_X1 _26279_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[12]),
    .ZN(_05746_)
  );
  INV_X1 _26280_ (
    .A(_05746_),
    .ZN(_05747_)
  );
  AND2_X1 _26281_ (
    .A1(_05745_),
    .A2(_05747_),
    .ZN(_05748_)
  );
  INV_X1 _26282_ (
    .A(_05748_),
    .ZN(_00465_)
  );
  AND2_X1 _26283_ (
    .A1(ex_reg_cause[13]),
    .A2(_05708_),
    .ZN(_05749_)
  );
  INV_X1 _26284_ (
    .A(_05749_),
    .ZN(_05750_)
  );
  AND2_X1 _26285_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[13]),
    .ZN(_05751_)
  );
  INV_X1 _26286_ (
    .A(_05751_),
    .ZN(_05752_)
  );
  AND2_X1 _26287_ (
    .A1(_05750_),
    .A2(_05752_),
    .ZN(_05753_)
  );
  INV_X1 _26288_ (
    .A(_05753_),
    .ZN(_00466_)
  );
  AND2_X1 _26289_ (
    .A1(ex_reg_cause[14]),
    .A2(_05708_),
    .ZN(_05754_)
  );
  INV_X1 _26290_ (
    .A(_05754_),
    .ZN(_05755_)
  );
  AND2_X1 _26291_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[14]),
    .ZN(_05756_)
  );
  INV_X1 _26292_ (
    .A(_05756_),
    .ZN(_05757_)
  );
  AND2_X1 _26293_ (
    .A1(_05755_),
    .A2(_05757_),
    .ZN(_05758_)
  );
  INV_X1 _26294_ (
    .A(_05758_),
    .ZN(_00467_)
  );
  AND2_X1 _26295_ (
    .A1(ex_reg_cause[15]),
    .A2(_05708_),
    .ZN(_05759_)
  );
  INV_X1 _26296_ (
    .A(_05759_),
    .ZN(_05760_)
  );
  AND2_X1 _26297_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[15]),
    .ZN(_05761_)
  );
  INV_X1 _26298_ (
    .A(_05761_),
    .ZN(_05762_)
  );
  AND2_X1 _26299_ (
    .A1(_05760_),
    .A2(_05762_),
    .ZN(_05763_)
  );
  INV_X1 _26300_ (
    .A(_05763_),
    .ZN(_00468_)
  );
  AND2_X1 _26301_ (
    .A1(ex_reg_cause[16]),
    .A2(_05708_),
    .ZN(_05764_)
  );
  INV_X1 _26302_ (
    .A(_05764_),
    .ZN(_05765_)
  );
  AND2_X1 _26303_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[16]),
    .ZN(_05766_)
  );
  INV_X1 _26304_ (
    .A(_05766_),
    .ZN(_05767_)
  );
  AND2_X1 _26305_ (
    .A1(_05765_),
    .A2(_05767_),
    .ZN(_05768_)
  );
  INV_X1 _26306_ (
    .A(_05768_),
    .ZN(_00469_)
  );
  AND2_X1 _26307_ (
    .A1(ex_reg_cause[17]),
    .A2(_05708_),
    .ZN(_05769_)
  );
  INV_X1 _26308_ (
    .A(_05769_),
    .ZN(_05770_)
  );
  AND2_X1 _26309_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[17]),
    .ZN(_05771_)
  );
  INV_X1 _26310_ (
    .A(_05771_),
    .ZN(_05772_)
  );
  AND2_X1 _26311_ (
    .A1(_05770_),
    .A2(_05772_),
    .ZN(_05773_)
  );
  INV_X1 _26312_ (
    .A(_05773_),
    .ZN(_00470_)
  );
  AND2_X1 _26313_ (
    .A1(ex_reg_cause[18]),
    .A2(_05708_),
    .ZN(_05774_)
  );
  INV_X1 _26314_ (
    .A(_05774_),
    .ZN(_05775_)
  );
  AND2_X1 _26315_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[18]),
    .ZN(_05776_)
  );
  INV_X1 _26316_ (
    .A(_05776_),
    .ZN(_05777_)
  );
  AND2_X1 _26317_ (
    .A1(_05775_),
    .A2(_05777_),
    .ZN(_05778_)
  );
  INV_X1 _26318_ (
    .A(_05778_),
    .ZN(_00471_)
  );
  AND2_X1 _26319_ (
    .A1(ex_reg_cause[19]),
    .A2(_05708_),
    .ZN(_05779_)
  );
  INV_X1 _26320_ (
    .A(_05779_),
    .ZN(_05780_)
  );
  AND2_X1 _26321_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[19]),
    .ZN(_05781_)
  );
  INV_X1 _26322_ (
    .A(_05781_),
    .ZN(_05782_)
  );
  AND2_X1 _26323_ (
    .A1(_05780_),
    .A2(_05782_),
    .ZN(_05783_)
  );
  INV_X1 _26324_ (
    .A(_05783_),
    .ZN(_00472_)
  );
  AND2_X1 _26325_ (
    .A1(ex_reg_cause[20]),
    .A2(_05708_),
    .ZN(_05784_)
  );
  INV_X1 _26326_ (
    .A(_05784_),
    .ZN(_05785_)
  );
  AND2_X1 _26327_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[20]),
    .ZN(_05786_)
  );
  INV_X1 _26328_ (
    .A(_05786_),
    .ZN(_05787_)
  );
  AND2_X1 _26329_ (
    .A1(_05785_),
    .A2(_05787_),
    .ZN(_05788_)
  );
  INV_X1 _26330_ (
    .A(_05788_),
    .ZN(_00473_)
  );
  AND2_X1 _26331_ (
    .A1(ex_reg_cause[21]),
    .A2(_05708_),
    .ZN(_05789_)
  );
  INV_X1 _26332_ (
    .A(_05789_),
    .ZN(_05790_)
  );
  AND2_X1 _26333_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[21]),
    .ZN(_05791_)
  );
  INV_X1 _26334_ (
    .A(_05791_),
    .ZN(_05792_)
  );
  AND2_X1 _26335_ (
    .A1(_05790_),
    .A2(_05792_),
    .ZN(_05793_)
  );
  INV_X1 _26336_ (
    .A(_05793_),
    .ZN(_00474_)
  );
  AND2_X1 _26337_ (
    .A1(ex_reg_cause[22]),
    .A2(_05708_),
    .ZN(_05794_)
  );
  INV_X1 _26338_ (
    .A(_05794_),
    .ZN(_05795_)
  );
  AND2_X1 _26339_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[22]),
    .ZN(_05796_)
  );
  INV_X1 _26340_ (
    .A(_05796_),
    .ZN(_05797_)
  );
  AND2_X1 _26341_ (
    .A1(_05795_),
    .A2(_05797_),
    .ZN(_05798_)
  );
  INV_X1 _26342_ (
    .A(_05798_),
    .ZN(_00475_)
  );
  AND2_X1 _26343_ (
    .A1(ex_reg_cause[23]),
    .A2(_05708_),
    .ZN(_05799_)
  );
  INV_X1 _26344_ (
    .A(_05799_),
    .ZN(_05800_)
  );
  AND2_X1 _26345_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[23]),
    .ZN(_05801_)
  );
  INV_X1 _26346_ (
    .A(_05801_),
    .ZN(_05802_)
  );
  AND2_X1 _26347_ (
    .A1(_05800_),
    .A2(_05802_),
    .ZN(_05803_)
  );
  INV_X1 _26348_ (
    .A(_05803_),
    .ZN(_00476_)
  );
  AND2_X1 _26349_ (
    .A1(ex_reg_cause[24]),
    .A2(_05708_),
    .ZN(_05804_)
  );
  INV_X1 _26350_ (
    .A(_05804_),
    .ZN(_05805_)
  );
  AND2_X1 _26351_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[24]),
    .ZN(_05806_)
  );
  INV_X1 _26352_ (
    .A(_05806_),
    .ZN(_05807_)
  );
  AND2_X1 _26353_ (
    .A1(_05805_),
    .A2(_05807_),
    .ZN(_05808_)
  );
  INV_X1 _26354_ (
    .A(_05808_),
    .ZN(_00477_)
  );
  AND2_X1 _26355_ (
    .A1(ex_reg_cause[25]),
    .A2(_05708_),
    .ZN(_05809_)
  );
  INV_X1 _26356_ (
    .A(_05809_),
    .ZN(_05810_)
  );
  AND2_X1 _26357_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[25]),
    .ZN(_05811_)
  );
  INV_X1 _26358_ (
    .A(_05811_),
    .ZN(_05812_)
  );
  AND2_X1 _26359_ (
    .A1(_05810_),
    .A2(_05812_),
    .ZN(_05813_)
  );
  INV_X1 _26360_ (
    .A(_05813_),
    .ZN(_00478_)
  );
  AND2_X1 _26361_ (
    .A1(ex_reg_cause[26]),
    .A2(_05708_),
    .ZN(_05814_)
  );
  INV_X1 _26362_ (
    .A(_05814_),
    .ZN(_05815_)
  );
  AND2_X1 _26363_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[26]),
    .ZN(_05816_)
  );
  INV_X1 _26364_ (
    .A(_05816_),
    .ZN(_05817_)
  );
  AND2_X1 _26365_ (
    .A1(_05815_),
    .A2(_05817_),
    .ZN(_05818_)
  );
  INV_X1 _26366_ (
    .A(_05818_),
    .ZN(_00479_)
  );
  AND2_X1 _26367_ (
    .A1(ex_reg_cause[27]),
    .A2(_05708_),
    .ZN(_05819_)
  );
  INV_X1 _26368_ (
    .A(_05819_),
    .ZN(_05820_)
  );
  AND2_X1 _26369_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[27]),
    .ZN(_05821_)
  );
  INV_X1 _26370_ (
    .A(_05821_),
    .ZN(_05822_)
  );
  AND2_X1 _26371_ (
    .A1(_05820_),
    .A2(_05822_),
    .ZN(_05823_)
  );
  INV_X1 _26372_ (
    .A(_05823_),
    .ZN(_00480_)
  );
  AND2_X1 _26373_ (
    .A1(ex_reg_cause[28]),
    .A2(_05708_),
    .ZN(_05824_)
  );
  INV_X1 _26374_ (
    .A(_05824_),
    .ZN(_05825_)
  );
  AND2_X1 _26375_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[28]),
    .ZN(_05826_)
  );
  INV_X1 _26376_ (
    .A(_05826_),
    .ZN(_05827_)
  );
  AND2_X1 _26377_ (
    .A1(_05825_),
    .A2(_05827_),
    .ZN(_05828_)
  );
  INV_X1 _26378_ (
    .A(_05828_),
    .ZN(_00481_)
  );
  AND2_X1 _26379_ (
    .A1(ex_reg_cause[29]),
    .A2(_05708_),
    .ZN(_05829_)
  );
  INV_X1 _26380_ (
    .A(_05829_),
    .ZN(_05830_)
  );
  AND2_X1 _26381_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[29]),
    .ZN(_05831_)
  );
  INV_X1 _26382_ (
    .A(_05831_),
    .ZN(_05832_)
  );
  AND2_X1 _26383_ (
    .A1(_05830_),
    .A2(_05832_),
    .ZN(_05833_)
  );
  INV_X1 _26384_ (
    .A(_05833_),
    .ZN(_00482_)
  );
  AND2_X1 _26385_ (
    .A1(ex_reg_cause[30]),
    .A2(_05708_),
    .ZN(_05834_)
  );
  INV_X1 _26386_ (
    .A(_05834_),
    .ZN(_05835_)
  );
  AND2_X1 _26387_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[30]),
    .ZN(_05836_)
  );
  INV_X1 _26388_ (
    .A(_05836_),
    .ZN(_05837_)
  );
  AND2_X1 _26389_ (
    .A1(_05835_),
    .A2(_05837_),
    .ZN(_05838_)
  );
  INV_X1 _26390_ (
    .A(_05838_),
    .ZN(_00483_)
  );
  AND2_X1 _26391_ (
    .A1(ex_reg_cause[31]),
    .A2(_05708_),
    .ZN(_05839_)
  );
  INV_X1 _26392_ (
    .A(_05839_),
    .ZN(_05840_)
  );
  AND2_X1 _26393_ (
    .A1(csr_io_interrupt_cause[31]),
    .A2(csr_io_interrupt),
    .ZN(_05841_)
  );
  INV_X1 _26394_ (
    .A(_05841_),
    .ZN(_05842_)
  );
  AND2_X1 _26395_ (
    .A1(_05840_),
    .A2(_05842_),
    .ZN(_05843_)
  );
  INV_X1 _26396_ (
    .A(_05843_),
    .ZN(_00484_)
  );
  MUX2_X1 _26397_ (
    .A(bpu_io_pc[0]),
    .B(ex_reg_pc[0]),
    .S(_05708_),
    .Z(_00485_)
  );
  MUX2_X1 _26398_ (
    .A(bpu_io_pc[1]),
    .B(ex_reg_pc[1]),
    .S(_05708_),
    .Z(_00486_)
  );
  MUX2_X1 _26399_ (
    .A(bpu_io_pc[2]),
    .B(ex_reg_pc[2]),
    .S(_05708_),
    .Z(_00487_)
  );
  MUX2_X1 _26400_ (
    .A(bpu_io_pc[3]),
    .B(ex_reg_pc[3]),
    .S(_05708_),
    .Z(_00488_)
  );
  MUX2_X1 _26401_ (
    .A(bpu_io_pc[4]),
    .B(ex_reg_pc[4]),
    .S(_05708_),
    .Z(_00489_)
  );
  MUX2_X1 _26402_ (
    .A(bpu_io_pc[5]),
    .B(ex_reg_pc[5]),
    .S(_05708_),
    .Z(_00490_)
  );
  MUX2_X1 _26403_ (
    .A(bpu_io_pc[6]),
    .B(ex_reg_pc[6]),
    .S(_05708_),
    .Z(_00491_)
  );
  MUX2_X1 _26404_ (
    .A(bpu_io_pc[7]),
    .B(ex_reg_pc[7]),
    .S(_05708_),
    .Z(_00492_)
  );
  MUX2_X1 _26405_ (
    .A(bpu_io_pc[8]),
    .B(ex_reg_pc[8]),
    .S(_05708_),
    .Z(_00493_)
  );
  MUX2_X1 _26406_ (
    .A(bpu_io_pc[9]),
    .B(ex_reg_pc[9]),
    .S(_05708_),
    .Z(_00494_)
  );
  MUX2_X1 _26407_ (
    .A(bpu_io_pc[10]),
    .B(ex_reg_pc[10]),
    .S(_05708_),
    .Z(_00495_)
  );
  MUX2_X1 _26408_ (
    .A(bpu_io_pc[11]),
    .B(ex_reg_pc[11]),
    .S(_05708_),
    .Z(_00496_)
  );
  MUX2_X1 _26409_ (
    .A(bpu_io_pc[12]),
    .B(ex_reg_pc[12]),
    .S(_05708_),
    .Z(_00497_)
  );
  MUX2_X1 _26410_ (
    .A(bpu_io_pc[13]),
    .B(ex_reg_pc[13]),
    .S(_05708_),
    .Z(_00498_)
  );
  MUX2_X1 _26411_ (
    .A(bpu_io_pc[14]),
    .B(ex_reg_pc[14]),
    .S(_05708_),
    .Z(_00499_)
  );
  MUX2_X1 _26412_ (
    .A(bpu_io_pc[15]),
    .B(ex_reg_pc[15]),
    .S(_05708_),
    .Z(_00500_)
  );
  MUX2_X1 _26413_ (
    .A(bpu_io_pc[16]),
    .B(ex_reg_pc[16]),
    .S(_05708_),
    .Z(_00501_)
  );
  MUX2_X1 _26414_ (
    .A(bpu_io_pc[17]),
    .B(ex_reg_pc[17]),
    .S(_05708_),
    .Z(_00502_)
  );
  MUX2_X1 _26415_ (
    .A(bpu_io_pc[18]),
    .B(ex_reg_pc[18]),
    .S(_05708_),
    .Z(_00503_)
  );
  MUX2_X1 _26416_ (
    .A(bpu_io_pc[19]),
    .B(ex_reg_pc[19]),
    .S(_05708_),
    .Z(_00504_)
  );
  MUX2_X1 _26417_ (
    .A(bpu_io_pc[20]),
    .B(ex_reg_pc[20]),
    .S(_05708_),
    .Z(_00505_)
  );
  MUX2_X1 _26418_ (
    .A(bpu_io_pc[21]),
    .B(ex_reg_pc[21]),
    .S(_05708_),
    .Z(_00506_)
  );
  MUX2_X1 _26419_ (
    .A(bpu_io_pc[22]),
    .B(ex_reg_pc[22]),
    .S(_05708_),
    .Z(_00507_)
  );
  MUX2_X1 _26420_ (
    .A(bpu_io_pc[23]),
    .B(ex_reg_pc[23]),
    .S(_05708_),
    .Z(_00508_)
  );
  MUX2_X1 _26421_ (
    .A(bpu_io_pc[24]),
    .B(ex_reg_pc[24]),
    .S(_05708_),
    .Z(_00509_)
  );
  MUX2_X1 _26422_ (
    .A(bpu_io_pc[25]),
    .B(ex_reg_pc[25]),
    .S(_05708_),
    .Z(_00510_)
  );
  MUX2_X1 _26423_ (
    .A(bpu_io_pc[26]),
    .B(ex_reg_pc[26]),
    .S(_05708_),
    .Z(_00511_)
  );
  MUX2_X1 _26424_ (
    .A(bpu_io_pc[27]),
    .B(ex_reg_pc[27]),
    .S(_05708_),
    .Z(_00512_)
  );
  MUX2_X1 _26425_ (
    .A(bpu_io_pc[28]),
    .B(ex_reg_pc[28]),
    .S(_05708_),
    .Z(_00513_)
  );
  MUX2_X1 _26426_ (
    .A(bpu_io_pc[29]),
    .B(ex_reg_pc[29]),
    .S(_05708_),
    .Z(_00514_)
  );
  MUX2_X1 _26427_ (
    .A(bpu_io_pc[30]),
    .B(ex_reg_pc[30]),
    .S(_05708_),
    .Z(_00515_)
  );
  MUX2_X1 _26428_ (
    .A(bpu_io_pc[31]),
    .B(ex_reg_pc[31]),
    .S(_05708_),
    .Z(_00516_)
  );
  AND2_X1 _26429_ (
    .A1(mem_ctrl_mem),
    .A2(_09881_),
    .ZN(_05844_)
  );
  MUX2_X1 _26430_ (
    .A(ex_reg_load_use),
    .B(_05844_),
    .S(_ex_reg_valid_T),
    .Z(_00517_)
  );
  AND2_X1 _26431_ (
    .A1(_08187_),
    .A2(_10078_),
    .ZN(_05845_)
  );
  INV_X1 _26432_ (
    .A(_05845_),
    .ZN(_05846_)
  );
  AND2_X1 _26433_ (
    .A1(csr_io_decode_0_write_flush),
    .A2(_09263_),
    .ZN(_05847_)
  );
  AND2_X1 _26434_ (
    .A1(_09274_),
    .A2(_05847_),
    .ZN(_05848_)
  );
  INV_X1 _26435_ (
    .A(_05848_),
    .ZN(_05849_)
  );
  AND2_X1 _26436_ (
    .A1(_09269_),
    .A2(_05849_),
    .ZN(_05850_)
  );
  AND2_X1 _26437_ (
    .A1(_09472_),
    .A2(_ex_reg_valid_T),
    .ZN(_05851_)
  );
  AND2_X1 _26438_ (
    .A1(_05850_),
    .A2(_05851_),
    .ZN(_05852_)
  );
  INV_X1 _26439_ (
    .A(_05852_),
    .ZN(_05853_)
  );
  AND2_X1 _26440_ (
    .A1(_05846_),
    .A2(_05853_),
    .ZN(_00518_)
  );
  MUX2_X1 _26441_ (
    .A(mem_ctrl_fence_i),
    .B(wb_ctrl_fence_i),
    .S(_13833_),
    .Z(_00519_)
  );
  MUX2_X1 _26442_ (
    .A(mem_ctrl_csr[0]),
    .B(wb_ctrl_csr[0]),
    .S(_13833_),
    .Z(_00520_)
  );
  MUX2_X1 _26443_ (
    .A(mem_ctrl_csr[1]),
    .B(wb_ctrl_csr[1]),
    .S(_13833_),
    .Z(_00521_)
  );
  MUX2_X1 _26444_ (
    .A(mem_ctrl_csr[2]),
    .B(wb_ctrl_csr[2]),
    .S(_13833_),
    .Z(_00522_)
  );
  MUX2_X1 _26445_ (
    .A(mem_ctrl_wxd),
    .B(wb_ctrl_wxd),
    .S(_13833_),
    .Z(_00523_)
  );
  MUX2_X1 _26446_ (
    .A(mem_ctrl_div),
    .B(wb_ctrl_div),
    .S(_13833_),
    .Z(_00524_)
  );
  MUX2_X1 _26447_ (
    .A(mem_ctrl_mem),
    .B(wb_ctrl_mem),
    .S(_13833_),
    .Z(_00525_)
  );
  MUX2_X1 _26448_ (
    .A(mem_reg_inst[7]),
    .B(wb_reg_inst[7]),
    .S(_13833_),
    .Z(_00526_)
  );
  MUX2_X1 _26449_ (
    .A(mem_reg_inst[8]),
    .B(wb_reg_inst[8]),
    .S(_13833_),
    .Z(_00527_)
  );
  MUX2_X1 _26450_ (
    .A(mem_reg_inst[9]),
    .B(wb_reg_inst[9]),
    .S(_13833_),
    .Z(_00528_)
  );
  MUX2_X1 _26451_ (
    .A(mem_reg_inst[10]),
    .B(wb_reg_inst[10]),
    .S(_13833_),
    .Z(_00529_)
  );
  MUX2_X1 _26452_ (
    .A(mem_reg_inst[11]),
    .B(wb_reg_inst[11]),
    .S(_13833_),
    .Z(_00530_)
  );
  MUX2_X1 _26453_ (
    .A(mem_reg_inst[16]),
    .B(wb_reg_inst[16]),
    .S(_13833_),
    .Z(_00531_)
  );
  MUX2_X1 _26454_ (
    .A(mem_reg_inst[17]),
    .B(wb_reg_inst[17]),
    .S(_13833_),
    .Z(_00532_)
  );
  MUX2_X1 _26455_ (
    .A(mem_reg_inst[18]),
    .B(wb_reg_inst[18]),
    .S(_13833_),
    .Z(_00533_)
  );
  MUX2_X1 _26456_ (
    .A(mem_reg_inst[19]),
    .B(wb_reg_inst[19]),
    .S(_13833_),
    .Z(_00534_)
  );
  MUX2_X1 _26457_ (
    .A(mem_reg_inst[20]),
    .B(wb_reg_inst[20]),
    .S(_13833_),
    .Z(_00535_)
  );
  MUX2_X1 _26458_ (
    .A(mem_reg_inst[21]),
    .B(wb_reg_inst[21]),
    .S(_13833_),
    .Z(_00536_)
  );
  MUX2_X1 _26459_ (
    .A(mem_reg_inst[22]),
    .B(wb_reg_inst[22]),
    .S(_13833_),
    .Z(_00537_)
  );
  MUX2_X1 _26460_ (
    .A(mem_reg_inst[23]),
    .B(wb_reg_inst[23]),
    .S(_13833_),
    .Z(_00538_)
  );
  MUX2_X1 _26461_ (
    .A(mem_reg_inst[24]),
    .B(wb_reg_inst[24]),
    .S(_13833_),
    .Z(_00539_)
  );
  MUX2_X1 _26462_ (
    .A(mem_reg_inst[25]),
    .B(wb_reg_inst[25]),
    .S(_13833_),
    .Z(_00540_)
  );
  MUX2_X1 _26463_ (
    .A(mem_reg_inst[26]),
    .B(wb_reg_inst[26]),
    .S(_13833_),
    .Z(_00541_)
  );
  MUX2_X1 _26464_ (
    .A(mem_reg_inst[27]),
    .B(wb_reg_inst[27]),
    .S(_13833_),
    .Z(_00542_)
  );
  MUX2_X1 _26465_ (
    .A(mem_reg_inst[28]),
    .B(wb_reg_inst[28]),
    .S(_13833_),
    .Z(_00543_)
  );
  MUX2_X1 _26466_ (
    .A(mem_reg_inst[29]),
    .B(wb_reg_inst[29]),
    .S(_13833_),
    .Z(_00544_)
  );
  MUX2_X1 _26467_ (
    .A(mem_reg_inst[30]),
    .B(wb_reg_inst[30]),
    .S(_13833_),
    .Z(_00545_)
  );
  MUX2_X1 _26468_ (
    .A(mem_reg_inst[31]),
    .B(wb_reg_inst[31]),
    .S(_13833_),
    .Z(_00546_)
  );
  AND2_X1 _26469_ (
    .A1(_08209_),
    .A2(_05705_),
    .ZN(_05854_)
  );
  INV_X1 _26470_ (
    .A(_05854_),
    .ZN(_05855_)
  );
  MUX2_X1 _26471_ (
    .A(mem_ctrl_fence_i),
    .B(_05855_),
    .S(_05253_),
    .Z(_00547_)
  );
  MUX2_X1 _26472_ (
    .A(mem_ctrl_csr[0]),
    .B(ex_ctrl_csr[0]),
    .S(_05253_),
    .Z(_00548_)
  );
  MUX2_X1 _26473_ (
    .A(mem_ctrl_csr[1]),
    .B(ex_ctrl_csr[1]),
    .S(_05253_),
    .Z(_00549_)
  );
  MUX2_X1 _26474_ (
    .A(mem_ctrl_csr[2]),
    .B(ex_ctrl_csr[2]),
    .S(_05253_),
    .Z(_00550_)
  );
  MUX2_X1 _26475_ (
    .A(mem_ctrl_wxd),
    .B(ex_ctrl_wxd),
    .S(_05253_),
    .Z(_00551_)
  );
  MUX2_X1 _26476_ (
    .A(mem_ctrl_div),
    .B(ex_ctrl_div),
    .S(_05253_),
    .Z(_00552_)
  );
  MUX2_X1 _26477_ (
    .A(mem_ctrl_mem),
    .B(ex_ctrl_mem),
    .S(_05253_),
    .Z(_00553_)
  );
  MUX2_X1 _26478_ (
    .A(mem_ctrl_jalr),
    .B(ex_ctrl_jalr),
    .S(_05253_),
    .Z(_00554_)
  );
  MUX2_X1 _26479_ (
    .A(mem_ctrl_jal),
    .B(ex_ctrl_jal),
    .S(_05253_),
    .Z(_00555_)
  );
  MUX2_X1 _26480_ (
    .A(mem_ctrl_branch),
    .B(ex_ctrl_branch),
    .S(_05253_),
    .Z(_00556_)
  );
  MUX2_X1 _26481_ (
    .A(ex_ctrl_csr[1]),
    .B(_09241_),
    .S(_10244_),
    .Z(_00557_)
  );
  MUX2_X1 _26482_ (
    .A(ex_ctrl_fence_i),
    .B(_09471_),
    .S(_ex_reg_valid_T),
    .Z(_00558_)
  );
  MUX2_X1 _26483_ (
    .A(ex_ctrl_wxd),
    .B(_09317_),
    .S(_10244_),
    .Z(_00559_)
  );
  MUX2_X1 _26484_ (
    .A(ex_ctrl_div),
    .B(_09283_),
    .S(_10244_),
    .Z(_00560_)
  );
  AND2_X1 _26485_ (
    .A1(_09079_),
    .A2(_09089_),
    .ZN(_05856_)
  );
  INV_X1 _26486_ (
    .A(_05856_),
    .ZN(_05857_)
  );
  AND2_X1 _26487_ (
    .A1(csr_io_decode_0_inst[29]),
    .A2(_09057_),
    .ZN(_05858_)
  );
  INV_X1 _26488_ (
    .A(_05858_),
    .ZN(_05859_)
  );
  AND2_X1 _26489_ (
    .A1(_08529_),
    .A2(_09683_),
    .ZN(_05860_)
  );
  INV_X1 _26490_ (
    .A(_05860_),
    .ZN(_05861_)
  );
  AND2_X1 _26491_ (
    .A1(_05859_),
    .A2(_05861_),
    .ZN(_05862_)
  );
  AND2_X1 _26492_ (
    .A1(_05857_),
    .A2(_05862_),
    .ZN(_05863_)
  );
  INV_X1 _26493_ (
    .A(_05863_),
    .ZN(_05864_)
  );
  MUX2_X1 _26494_ (
    .A(ex_ctrl_mem_cmd[0]),
    .B(_05864_),
    .S(_ex_reg_valid_T),
    .Z(_00561_)
  );
  AND2_X1 _26495_ (
    .A1(csr_io_decode_0_inst[30]),
    .A2(_09057_),
    .ZN(_05865_)
  );
  INV_X1 _26496_ (
    .A(_05865_),
    .ZN(_05866_)
  );
  AND2_X1 _26497_ (
    .A1(_09088_),
    .A2(_05857_),
    .ZN(_05867_)
  );
  AND2_X1 _26498_ (
    .A1(_05866_),
    .A2(_05867_),
    .ZN(_05868_)
  );
  INV_X1 _26499_ (
    .A(_05868_),
    .ZN(_05869_)
  );
  MUX2_X1 _26500_ (
    .A(ex_ctrl_mem_cmd[1]),
    .B(_05869_),
    .S(_ex_reg_valid_T),
    .Z(_00562_)
  );
  AND2_X1 _26501_ (
    .A1(csr_io_decode_0_inst[31]),
    .A2(_09057_),
    .ZN(_05870_)
  );
  INV_X1 _26502_ (
    .A(_05870_),
    .ZN(_05871_)
  );
  AND2_X1 _26503_ (
    .A1(_09092_),
    .A2(_05871_),
    .ZN(_05872_)
  );
  INV_X1 _26504_ (
    .A(_05872_),
    .ZN(_05873_)
  );
  MUX2_X1 _26505_ (
    .A(ex_ctrl_mem_cmd[2]),
    .B(_05873_),
    .S(_ex_reg_valid_T),
    .Z(_00563_)
  );
  MUX2_X1 _26506_ (
    .A(ex_ctrl_mem_cmd[3]),
    .B(_09057_),
    .S(_ex_reg_valid_T),
    .Z(_00564_)
  );
  AND2_X1 _26507_ (
    .A1(_08135_),
    .A2(_08146_),
    .ZN(_05874_)
  );
  INV_X1 _26508_ (
    .A(_05874_),
    .ZN(_05875_)
  );
  AND2_X1 _26509_ (
    .A1(_09096_),
    .A2(_05875_),
    .ZN(_05876_)
  );
  INV_X1 _26510_ (
    .A(_05876_),
    .ZN(_05877_)
  );
  AND2_X1 _26511_ (
    .A1(_09040_),
    .A2(_05877_),
    .ZN(_05878_)
  );
  AND2_X1 _26512_ (
    .A1(_08987_),
    .A2(_09014_),
    .ZN(_05879_)
  );
  INV_X1 _26513_ (
    .A(_05879_),
    .ZN(_05880_)
  );
  AND2_X1 _26514_ (
    .A1(_05878_),
    .A2(_05880_),
    .ZN(_05881_)
  );
  INV_X1 _26515_ (
    .A(_05881_),
    .ZN(_05882_)
  );
  AND2_X1 _26516_ (
    .A1(csr_io_decode_0_inst[12]),
    .A2(_05882_),
    .ZN(_05883_)
  );
  INV_X1 _26517_ (
    .A(_05883_),
    .ZN(_05884_)
  );
  AND2_X1 _26518_ (
    .A1(_09020_),
    .A2(_09305_),
    .ZN(_05885_)
  );
  AND2_X1 _26519_ (
    .A1(_09048_),
    .A2(_05885_),
    .ZN(_05886_)
  );
  INV_X1 _26520_ (
    .A(_05886_),
    .ZN(_05887_)
  );
  AND2_X1 _26521_ (
    .A1(_09299_),
    .A2(_05887_),
    .ZN(_05888_)
  );
  AND2_X1 _26522_ (
    .A1(_05884_),
    .A2(_05888_),
    .ZN(_05889_)
  );
  INV_X1 _26523_ (
    .A(_05889_),
    .ZN(_05890_)
  );
  AND2_X1 _26524_ (
    .A1(_08581_),
    .A2(_08582_),
    .ZN(_05891_)
  );
  AND2_X1 _26525_ (
    .A1(_05215_),
    .A2(_05891_),
    .ZN(_05892_)
  );
  INV_X1 _26526_ (
    .A(_05892_),
    .ZN(_05893_)
  );
  AND2_X1 _26527_ (
    .A1(_07941_),
    .A2(_08583_),
    .ZN(_05894_)
  );
  AND2_X1 _26528_ (
    .A1(_09294_),
    .A2(_05894_),
    .ZN(_05895_)
  );
  AND2_X1 _26529_ (
    .A1(_05892_),
    .A2(_05895_),
    .ZN(_05896_)
  );
  INV_X1 _26530_ (
    .A(_05896_),
    .ZN(_05897_)
  );
  AND2_X1 _26531_ (
    .A1(_05890_),
    .A2(_05896_),
    .ZN(_05898_)
  );
  MUX2_X1 _26532_ (
    .A(ex_ctrl_alu_fn[0]),
    .B(_05898_),
    .S(_ex_reg_valid_T),
    .Z(_00565_)
  );
  AND2_X1 _26533_ (
    .A1(_08146_),
    .A2(_09000_),
    .ZN(_05899_)
  );
  INV_X1 _26534_ (
    .A(_05899_),
    .ZN(_05900_)
  );
  AND2_X1 _26535_ (
    .A1(csr_io_decode_0_inst[13]),
    .A2(_05900_),
    .ZN(_05901_)
  );
  AND2_X1 _26536_ (
    .A1(csr_io_decode_0_inst[4]),
    .A2(_08989_),
    .ZN(_05902_)
  );
  AND2_X1 _26537_ (
    .A1(_09307_),
    .A2(_05902_),
    .ZN(_05903_)
  );
  INV_X1 _26538_ (
    .A(_05903_),
    .ZN(_05904_)
  );
  AND2_X1 _26539_ (
    .A1(_09097_),
    .A2(_05904_),
    .ZN(_05905_)
  );
  INV_X1 _26540_ (
    .A(_05905_),
    .ZN(_05906_)
  );
  AND2_X1 _26541_ (
    .A1(_05901_),
    .A2(_05906_),
    .ZN(_05907_)
  );
  INV_X1 _26542_ (
    .A(_05907_),
    .ZN(_05908_)
  );
  AND2_X1 _26543_ (
    .A1(_08997_),
    .A2(_09306_),
    .ZN(_05909_)
  );
  INV_X1 _26544_ (
    .A(_05909_),
    .ZN(_05910_)
  );
  AND2_X1 _26545_ (
    .A1(_09037_),
    .A2(_05910_),
    .ZN(_05911_)
  );
  INV_X1 _26546_ (
    .A(_05911_),
    .ZN(_05912_)
  );
  AND2_X1 _26547_ (
    .A1(_09023_),
    .A2(_05874_),
    .ZN(_05913_)
  );
  AND2_X1 _26548_ (
    .A1(_08990_),
    .A2(_05913_),
    .ZN(_05914_)
  );
  AND2_X1 _26549_ (
    .A1(_09095_),
    .A2(_05914_),
    .ZN(_05915_)
  );
  INV_X1 _26550_ (
    .A(_05915_),
    .ZN(_05916_)
  );
  AND2_X1 _26551_ (
    .A1(_09043_),
    .A2(_05916_),
    .ZN(_05917_)
  );
  INV_X1 _26552_ (
    .A(_05917_),
    .ZN(_05918_)
  );
  AND2_X1 _26553_ (
    .A1(csr_io_decode_0_inst[30]),
    .A2(_09029_),
    .ZN(_05919_)
  );
  AND2_X1 _26554_ (
    .A1(_05918_),
    .A2(_05919_),
    .ZN(_05920_)
  );
  INV_X1 _26555_ (
    .A(_05920_),
    .ZN(_05921_)
  );
  AND2_X1 _26556_ (
    .A1(_05912_),
    .A2(_05921_),
    .ZN(_05922_)
  );
  AND2_X1 _26557_ (
    .A1(_05908_),
    .A2(_05922_),
    .ZN(_05923_)
  );
  INV_X1 _26558_ (
    .A(_05923_),
    .ZN(_05924_)
  );
  AND2_X1 _26559_ (
    .A1(_05896_),
    .A2(_05924_),
    .ZN(_05925_)
  );
  MUX2_X1 _26560_ (
    .A(ex_ctrl_alu_fn[1]),
    .B(_05925_),
    .S(_ex_reg_valid_T),
    .Z(_00566_)
  );
  AND2_X1 _26561_ (
    .A1(_09048_),
    .A2(_09075_),
    .ZN(_05926_)
  );
  INV_X1 _26562_ (
    .A(_05926_),
    .ZN(_05927_)
  );
  AND2_X1 _26563_ (
    .A1(_09033_),
    .A2(_05927_),
    .ZN(_05928_)
  );
  INV_X1 _26564_ (
    .A(_05928_),
    .ZN(_05929_)
  );
  AND2_X1 _26565_ (
    .A1(csr_io_decode_0_inst[14]),
    .A2(_05929_),
    .ZN(_05930_)
  );
  INV_X1 _26566_ (
    .A(_05930_),
    .ZN(_05931_)
  );
  AND2_X1 _26567_ (
    .A1(csr_io_decode_0_inst[13]),
    .A2(_08146_),
    .ZN(_05932_)
  );
  INV_X1 _26568_ (
    .A(_05932_),
    .ZN(_05933_)
  );
  AND2_X1 _26569_ (
    .A1(_08135_),
    .A2(_05933_),
    .ZN(_05934_)
  );
  INV_X1 _26570_ (
    .A(_05934_),
    .ZN(_05935_)
  );
  AND2_X1 _26571_ (
    .A1(_09096_),
    .A2(_05935_),
    .ZN(_05936_)
  );
  INV_X1 _26572_ (
    .A(_05936_),
    .ZN(_05937_)
  );
  AND2_X1 _26573_ (
    .A1(_09040_),
    .A2(_09050_),
    .ZN(_05938_)
  );
  AND2_X1 _26574_ (
    .A1(_05937_),
    .A2(_05938_),
    .ZN(_05939_)
  );
  AND2_X1 _26575_ (
    .A1(_05931_),
    .A2(_05939_),
    .ZN(_05940_)
  );
  INV_X1 _26576_ (
    .A(_05940_),
    .ZN(_05941_)
  );
  AND2_X1 _26577_ (
    .A1(_05896_),
    .A2(_05941_),
    .ZN(_05942_)
  );
  MUX2_X1 _26578_ (
    .A(ex_ctrl_alu_fn[2]),
    .B(_05942_),
    .S(_ex_reg_valid_T),
    .Z(_00567_)
  );
  AND2_X1 _26579_ (
    .A1(_09060_),
    .A2(_05902_),
    .ZN(_05943_)
  );
  INV_X1 _26580_ (
    .A(_05943_),
    .ZN(_05944_)
  );
  AND2_X1 _26581_ (
    .A1(_09047_),
    .A2(_05913_),
    .ZN(_05945_)
  );
  AND2_X1 _26582_ (
    .A1(_09094_),
    .A2(_05945_),
    .ZN(_05946_)
  );
  AND2_X1 _26583_ (
    .A1(_09030_),
    .A2(_05946_),
    .ZN(_05947_)
  );
  INV_X1 _26584_ (
    .A(_05947_),
    .ZN(_05948_)
  );
  AND2_X1 _26585_ (
    .A1(_09040_),
    .A2(_05948_),
    .ZN(_05949_)
  );
  AND2_X1 _26586_ (
    .A1(_05944_),
    .A2(_05949_),
    .ZN(_05950_)
  );
  AND2_X1 _26587_ (
    .A1(_05921_),
    .A2(_05950_),
    .ZN(_05951_)
  );
  INV_X1 _26588_ (
    .A(_05951_),
    .ZN(_05952_)
  );
  AND2_X1 _26589_ (
    .A1(_05896_),
    .A2(_05952_),
    .ZN(_05953_)
  );
  MUX2_X1 _26590_ (
    .A(ex_ctrl_alu_fn[3]),
    .B(_05953_),
    .S(_ex_reg_valid_T),
    .Z(_00568_)
  );
  MUX2_X1 _26591_ (
    .A(ex_ctrl_mem),
    .B(_09501_),
    .S(_ex_reg_valid_T),
    .Z(_00569_)
  );
  AND2_X1 _26592_ (
    .A1(_08991_),
    .A2(_09038_),
    .ZN(_05954_)
  );
  AND2_X1 _26593_ (
    .A1(_08987_),
    .A2(_05954_),
    .ZN(_05955_)
  );
  INV_X1 _26594_ (
    .A(_05955_),
    .ZN(_05956_)
  );
  AND2_X1 _26595_ (
    .A1(_05880_),
    .A2(_05956_),
    .ZN(_05957_)
  );
  AND2_X1 _26596_ (
    .A1(_09246_),
    .A2(_05957_),
    .ZN(_05958_)
  );
  INV_X1 _26597_ (
    .A(_05958_),
    .ZN(_05959_)
  );
  MUX2_X1 _26598_ (
    .A(ex_ctrl_sel_imm[0]),
    .B(_05959_),
    .S(_10244_),
    .Z(_00570_)
  );
  AND2_X1 _26599_ (
    .A1(_09187_),
    .A2(_09246_),
    .ZN(_05960_)
  );
  INV_X1 _26600_ (
    .A(_05960_),
    .ZN(_05961_)
  );
  MUX2_X1 _26601_ (
    .A(ex_ctrl_sel_imm[1]),
    .B(_05961_),
    .S(_10244_),
    .Z(_00571_)
  );
  AND2_X1 _26602_ (
    .A1(_08531_),
    .A2(_09300_),
    .ZN(_05962_)
  );
  INV_X1 _26603_ (
    .A(_05962_),
    .ZN(_05963_)
  );
  AND2_X1 _26604_ (
    .A1(_09019_),
    .A2(_05954_),
    .ZN(_05964_)
  );
  INV_X1 _26605_ (
    .A(_05964_),
    .ZN(_05965_)
  );
  AND2_X1 _26606_ (
    .A1(_09050_),
    .A2(_09304_),
    .ZN(_05966_)
  );
  AND2_X1 _26607_ (
    .A1(_05965_),
    .A2(_05966_),
    .ZN(_05967_)
  );
  AND2_X1 _26608_ (
    .A1(_05963_),
    .A2(_05967_),
    .ZN(_05968_)
  );
  AND2_X1 _26609_ (
    .A1(_09311_),
    .A2(_05968_),
    .ZN(_05969_)
  );
  INV_X1 _26610_ (
    .A(_05969_),
    .ZN(_05970_)
  );
  MUX2_X1 _26611_ (
    .A(ex_ctrl_sel_imm[2]),
    .B(_05970_),
    .S(_10244_),
    .Z(_00572_)
  );
  AND2_X1 _26612_ (
    .A1(_09108_),
    .A2(_05895_),
    .ZN(_05971_)
  );
  INV_X1 _26613_ (
    .A(_05971_),
    .ZN(_05972_)
  );
  AND2_X1 _26614_ (
    .A1(_05892_),
    .A2(_05972_),
    .ZN(_05973_)
  );
  MUX2_X1 _26615_ (
    .A(ex_ctrl_sel_alu1[0]),
    .B(_05973_),
    .S(_10244_),
    .Z(_00573_)
  );
  AND2_X1 _26616_ (
    .A1(_08531_),
    .A2(_09186_),
    .ZN(_05974_)
  );
  INV_X1 _26617_ (
    .A(_05974_),
    .ZN(_05975_)
  );
  AND2_X1 _26618_ (
    .A1(_09244_),
    .A2(_05975_),
    .ZN(_05976_)
  );
  INV_X1 _26619_ (
    .A(_05976_),
    .ZN(_05977_)
  );
  AND2_X1 _26620_ (
    .A1(_05895_),
    .A2(_05977_),
    .ZN(_05978_)
  );
  INV_X1 _26621_ (
    .A(_05978_),
    .ZN(_05979_)
  );
  AND2_X1 _26622_ (
    .A1(_05892_),
    .A2(_05979_),
    .ZN(_05980_)
  );
  INV_X1 _26623_ (
    .A(_05980_),
    .ZN(_05981_)
  );
  MUX2_X1 _26624_ (
    .A(ex_ctrl_sel_alu1[1]),
    .B(_05981_),
    .S(_10244_),
    .Z(_00574_)
  );
  AND2_X1 _26625_ (
    .A1(_09011_),
    .A2(_05960_),
    .ZN(_05982_)
  );
  AND2_X1 _26626_ (
    .A1(_05968_),
    .A2(_05982_),
    .ZN(_05983_)
  );
  INV_X1 _26627_ (
    .A(_05983_),
    .ZN(_05984_)
  );
  AND2_X1 _26628_ (
    .A1(_05895_),
    .A2(_05984_),
    .ZN(_05985_)
  );
  INV_X1 _26629_ (
    .A(_05985_),
    .ZN(_05986_)
  );
  AND2_X1 _26630_ (
    .A1(_05215_),
    .A2(_05986_),
    .ZN(_05987_)
  );
  INV_X1 _26631_ (
    .A(_05987_),
    .ZN(_05988_)
  );
  AND2_X1 _26632_ (
    .A1(_05891_),
    .A2(_05988_),
    .ZN(_05989_)
  );
  MUX2_X1 _26633_ (
    .A(ex_ctrl_sel_alu2[0]),
    .B(_05989_),
    .S(_10244_),
    .Z(_00575_)
  );
  MUX2_X1 _26634_ (
    .A(ex_ctrl_rxs2),
    .B(_09691_),
    .S(_10244_),
    .Z(_00576_)
  );
  MUX2_X1 _26635_ (
    .A(ex_ctrl_jalr),
    .B(_09303_),
    .S(_10244_),
    .Z(_00577_)
  );
  MUX2_X1 _26636_ (
    .A(ex_ctrl_jal),
    .B(_09245_),
    .S(_10244_),
    .Z(_00578_)
  );
  AND2_X1 _26637_ (
    .A1(_09037_),
    .A2(_09061_),
    .ZN(_05990_)
  );
  MUX2_X1 _26638_ (
    .A(ex_ctrl_branch),
    .B(_05990_),
    .S(_10244_),
    .Z(_00579_)
  );
  AND2_X1 _26639_ (
    .A1(_09840_),
    .A2(_13693_),
    .ZN(_05991_)
  );
  AND2_X1 _26640_ (
    .A1(_13827_),
    .A2(_05991_),
    .ZN(_05992_)
  );
  INV_X1 _26641_ (
    .A(_05992_),
    .ZN(_05993_)
  );
  AND2_X1 _26642_ (
    .A1(_09696_),
    .A2(_05993_),
    .ZN(_05994_)
  );
  AND2_X1 _26643_ (
    .A1(_08494_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_05995_)
  );
  INV_X1 _26644_ (
    .A(_05995_),
    .ZN(_05996_)
  );
  AND2_X1 _26645_ (
    .A1(_08467_),
    .A2(_08546_),
    .ZN(_05997_)
  );
  INV_X1 _26646_ (
    .A(_05997_),
    .ZN(_05998_)
  );
  AND2_X1 _26647_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_05998_),
    .ZN(_05999_)
  );
  AND2_X1 _26648_ (
    .A1(_05996_),
    .A2(_05999_),
    .ZN(_06000_)
  );
  INV_X1 _26649_ (
    .A(_06000_),
    .ZN(_06001_)
  );
  AND2_X1 _26650_ (
    .A1(\rf[27] [0]),
    .A2(_09705_),
    .ZN(_06002_)
  );
  INV_X1 _26651_ (
    .A(_06002_),
    .ZN(_06003_)
  );
  MUX2_X1 _26652_ (
    .A(\rf[13] [0]),
    .B(\rf[9] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06004_)
  );
  AND2_X1 _26653_ (
    .A1(_08257_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_06005_)
  );
  INV_X1 _26654_ (
    .A(_06005_),
    .ZN(_06006_)
  );
  AND2_X1 _26655_ (
    .A1(_08356_),
    .A2(_08546_),
    .ZN(_06007_)
  );
  INV_X1 _26656_ (
    .A(_06007_),
    .ZN(_06008_)
  );
  MUX2_X1 _26657_ (
    .A(\rf[15] [0]),
    .B(\rf[11] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06009_)
  );
  AND2_X1 _26658_ (
    .A1(_08473_),
    .A2(_08546_),
    .ZN(_06010_)
  );
  INV_X1 _26659_ (
    .A(_06010_),
    .ZN(_06011_)
  );
  AND2_X1 _26660_ (
    .A1(_08335_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_06012_)
  );
  INV_X1 _26661_ (
    .A(_06012_),
    .ZN(_06013_)
  );
  MUX2_X1 _26662_ (
    .A(\rf[29] [0]),
    .B(\rf[25] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06014_)
  );
  AND2_X1 _26663_ (
    .A1(_08544_),
    .A2(_06014_),
    .ZN(_06015_)
  );
  INV_X1 _26664_ (
    .A(_06015_),
    .ZN(_06016_)
  );
  AND2_X1 _26665_ (
    .A1(_08434_),
    .A2(_08546_),
    .ZN(_06017_)
  );
  INV_X1 _26666_ (
    .A(_06017_),
    .ZN(_06018_)
  );
  AND2_X1 _26667_ (
    .A1(_08504_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_06019_)
  );
  INV_X1 _26668_ (
    .A(_06019_),
    .ZN(_06020_)
  );
  AND2_X1 _26669_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_06020_),
    .ZN(_06021_)
  );
  AND2_X1 _26670_ (
    .A1(_06018_),
    .A2(_06021_),
    .ZN(_06022_)
  );
  INV_X1 _26671_ (
    .A(_06022_),
    .ZN(_06023_)
  );
  AND2_X1 _26672_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_06023_),
    .ZN(_06024_)
  );
  AND2_X1 _26673_ (
    .A1(_06016_),
    .A2(_06024_),
    .ZN(_06025_)
  );
  INV_X1 _26674_ (
    .A(_06025_),
    .ZN(_06026_)
  );
  AND2_X1 _26675_ (
    .A1(_08545_),
    .A2(_06003_),
    .ZN(_06027_)
  );
  AND2_X1 _26676_ (
    .A1(_06001_),
    .A2(_06027_),
    .ZN(_06028_)
  );
  INV_X1 _26677_ (
    .A(_06028_),
    .ZN(_06029_)
  );
  AND2_X1 _26678_ (
    .A1(_08547_),
    .A2(_06029_),
    .ZN(_06030_)
  );
  AND2_X1 _26679_ (
    .A1(_06026_),
    .A2(_06030_),
    .ZN(_06031_)
  );
  INV_X1 _26680_ (
    .A(_06031_),
    .ZN(_06032_)
  );
  MUX2_X1 _26681_ (
    .A(\rf[21] [0]),
    .B(\rf[17] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06033_)
  );
  AND2_X1 _26682_ (
    .A1(_08544_),
    .A2(_06033_),
    .ZN(_06034_)
  );
  INV_X1 _26683_ (
    .A(_06034_),
    .ZN(_06035_)
  );
  AND2_X1 _26684_ (
    .A1(_08373_),
    .A2(_08546_),
    .ZN(_06036_)
  );
  INV_X1 _26685_ (
    .A(_06036_),
    .ZN(_06037_)
  );
  AND2_X1 _26686_ (
    .A1(_08274_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_06038_)
  );
  INV_X1 _26687_ (
    .A(_06038_),
    .ZN(_06039_)
  );
  AND2_X1 _26688_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_06039_),
    .ZN(_06040_)
  );
  AND2_X1 _26689_ (
    .A1(_06037_),
    .A2(_06040_),
    .ZN(_06041_)
  );
  INV_X1 _26690_ (
    .A(_06041_),
    .ZN(_06042_)
  );
  AND2_X1 _26691_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_06035_),
    .ZN(_06043_)
  );
  AND2_X1 _26692_ (
    .A1(_06042_),
    .A2(_06043_),
    .ZN(_06044_)
  );
  INV_X1 _26693_ (
    .A(_06044_),
    .ZN(_06045_)
  );
  AND2_X1 _26694_ (
    .A1(_08352_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_06046_)
  );
  INV_X1 _26695_ (
    .A(_06046_),
    .ZN(_06047_)
  );
  AND2_X1 _26696_ (
    .A1(_08490_),
    .A2(_08546_),
    .ZN(_06048_)
  );
  INV_X1 _26697_ (
    .A(_06048_),
    .ZN(_06049_)
  );
  AND2_X1 _26698_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_06049_),
    .ZN(_06050_)
  );
  AND2_X1 _26699_ (
    .A1(_06047_),
    .A2(_06050_),
    .ZN(_06051_)
  );
  INV_X1 _26700_ (
    .A(_06051_),
    .ZN(_06052_)
  );
  MUX2_X1 _26701_ (
    .A(\rf[23] [0]),
    .B(\rf[19] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06053_)
  );
  AND2_X1 _26702_ (
    .A1(_08544_),
    .A2(_06053_),
    .ZN(_06054_)
  );
  INV_X1 _26703_ (
    .A(_06054_),
    .ZN(_06055_)
  );
  AND2_X1 _26704_ (
    .A1(_08545_),
    .A2(_06055_),
    .ZN(_06056_)
  );
  AND2_X1 _26705_ (
    .A1(_06052_),
    .A2(_06056_),
    .ZN(_06057_)
  );
  INV_X1 _26706_ (
    .A(_06057_),
    .ZN(_06058_)
  );
  AND2_X1 _26707_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_06058_),
    .ZN(_06059_)
  );
  AND2_X1 _26708_ (
    .A1(_06045_),
    .A2(_06059_),
    .ZN(_06060_)
  );
  INV_X1 _26709_ (
    .A(_06060_),
    .ZN(_06061_)
  );
  AND2_X1 _26710_ (
    .A1(_08572_),
    .A2(_06061_),
    .ZN(_06062_)
  );
  AND2_X1 _26711_ (
    .A1(_06032_),
    .A2(_06062_),
    .ZN(_06063_)
  );
  INV_X1 _26712_ (
    .A(_06063_),
    .ZN(_06064_)
  );
  AND2_X1 _26713_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_06011_),
    .ZN(_06065_)
  );
  AND2_X1 _26714_ (
    .A1(_06013_),
    .A2(_06065_),
    .ZN(_06066_)
  );
  INV_X1 _26715_ (
    .A(_06066_),
    .ZN(_06067_)
  );
  AND2_X1 _26716_ (
    .A1(_08544_),
    .A2(_06009_),
    .ZN(_06068_)
  );
  INV_X1 _26717_ (
    .A(_06068_),
    .ZN(_06069_)
  );
  AND2_X1 _26718_ (
    .A1(_08545_),
    .A2(_06069_),
    .ZN(_06070_)
  );
  AND2_X1 _26719_ (
    .A1(_06067_),
    .A2(_06070_),
    .ZN(_06071_)
  );
  INV_X1 _26720_ (
    .A(_06071_),
    .ZN(_06072_)
  );
  AND2_X1 _26721_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_06006_),
    .ZN(_06073_)
  );
  AND2_X1 _26722_ (
    .A1(_06008_),
    .A2(_06073_),
    .ZN(_06074_)
  );
  INV_X1 _26723_ (
    .A(_06074_),
    .ZN(_06075_)
  );
  AND2_X1 _26724_ (
    .A1(_08544_),
    .A2(_06004_),
    .ZN(_06076_)
  );
  INV_X1 _26725_ (
    .A(_06076_),
    .ZN(_06077_)
  );
  AND2_X1 _26726_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_06077_),
    .ZN(_06078_)
  );
  AND2_X1 _26727_ (
    .A1(_06075_),
    .A2(_06078_),
    .ZN(_06079_)
  );
  INV_X1 _26728_ (
    .A(_06079_),
    .ZN(_06080_)
  );
  AND2_X1 _26729_ (
    .A1(_08547_),
    .A2(_06080_),
    .ZN(_06081_)
  );
  AND2_X1 _26730_ (
    .A1(_06072_),
    .A2(_06081_),
    .ZN(_06082_)
  );
  INV_X1 _26731_ (
    .A(_06082_),
    .ZN(_06083_)
  );
  AND2_X1 _26732_ (
    .A1(_08253_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_06084_)
  );
  INV_X1 _26733_ (
    .A(_06084_),
    .ZN(_06085_)
  );
  AND2_X1 _26734_ (
    .A1(_08248_),
    .A2(_08546_),
    .ZN(_06086_)
  );
  INV_X1 _26735_ (
    .A(_06086_),
    .ZN(_06087_)
  );
  AND2_X1 _26736_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_06087_),
    .ZN(_06088_)
  );
  AND2_X1 _26737_ (
    .A1(_06085_),
    .A2(_06088_),
    .ZN(_06089_)
  );
  INV_X1 _26738_ (
    .A(_06089_),
    .ZN(_06090_)
  );
  MUX2_X1 _26739_ (
    .A(\rf[5] [0]),
    .B(\rf[1] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06091_)
  );
  AND2_X1 _26740_ (
    .A1(_08544_),
    .A2(_06091_),
    .ZN(_06092_)
  );
  INV_X1 _26741_ (
    .A(_06092_),
    .ZN(_06093_)
  );
  AND2_X1 _26742_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_06093_),
    .ZN(_06094_)
  );
  AND2_X1 _26743_ (
    .A1(_06090_),
    .A2(_06094_),
    .ZN(_06095_)
  );
  INV_X1 _26744_ (
    .A(_06095_),
    .ZN(_06096_)
  );
  MUX2_X1 _26745_ (
    .A(\rf[7] [0]),
    .B(\rf[3] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06097_)
  );
  AND2_X1 _26746_ (
    .A1(_08544_),
    .A2(_06097_),
    .ZN(_06098_)
  );
  INV_X1 _26747_ (
    .A(_06098_),
    .ZN(_06099_)
  );
  AND2_X1 _26748_ (
    .A1(_08500_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_06100_)
  );
  INV_X1 _26749_ (
    .A(_06100_),
    .ZN(_06101_)
  );
  AND2_X1 _26750_ (
    .A1(_08244_),
    .A2(_08546_),
    .ZN(_06102_)
  );
  INV_X1 _26751_ (
    .A(_06102_),
    .ZN(_06103_)
  );
  AND2_X1 _26752_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_06103_),
    .ZN(_06104_)
  );
  AND2_X1 _26753_ (
    .A1(_06101_),
    .A2(_06104_),
    .ZN(_06105_)
  );
  INV_X1 _26754_ (
    .A(_06105_),
    .ZN(_06106_)
  );
  AND2_X1 _26755_ (
    .A1(_06099_),
    .A2(_06106_),
    .ZN(_06107_)
  );
  AND2_X1 _26756_ (
    .A1(_08545_),
    .A2(_06107_),
    .ZN(_06108_)
  );
  INV_X1 _26757_ (
    .A(_06108_),
    .ZN(_06109_)
  );
  AND2_X1 _26758_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_06096_),
    .ZN(_06110_)
  );
  AND2_X1 _26759_ (
    .A1(_06109_),
    .A2(_06110_),
    .ZN(_06111_)
  );
  INV_X1 _26760_ (
    .A(_06111_),
    .ZN(_06112_)
  );
  AND2_X1 _26761_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[4]),
    .A2(_06083_),
    .ZN(_06113_)
  );
  AND2_X1 _26762_ (
    .A1(_06112_),
    .A2(_06113_),
    .ZN(_06114_)
  );
  INV_X1 _26763_ (
    .A(_06114_),
    .ZN(_06115_)
  );
  AND2_X1 _26764_ (
    .A1(_06064_),
    .A2(_06115_),
    .ZN(_06116_)
  );
  AND2_X1 _26765_ (
    .A1(_13580_),
    .A2(_02233_),
    .ZN(_06117_)
  );
  INV_X1 _26766_ (
    .A(_06117_),
    .ZN(_06118_)
  );
  AND2_X1 _26767_ (
    .A1(_02234_),
    .A2(_06116_),
    .ZN(_06119_)
  );
  INV_X1 _26768_ (
    .A(_06119_),
    .ZN(_06120_)
  );
  AND2_X1 _26769_ (
    .A1(_02201_),
    .A2(_06118_),
    .ZN(_06121_)
  );
  AND2_X1 _26770_ (
    .A1(_06120_),
    .A2(_06121_),
    .ZN(_06122_)
  );
  INV_X1 _26771_ (
    .A(_06122_),
    .ZN(_06123_)
  );
  AND2_X1 _26772_ (
    .A1(_05994_),
    .A2(_06123_),
    .ZN(_06124_)
  );
  MUX2_X1 _26773_ (
    .A(ex_reg_rs_lsb_1[0]),
    .B(_06124_),
    .S(_10244_),
    .Z(_00580_)
  );
  AND2_X1 _26774_ (
    .A1(_08495_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_06125_)
  );
  INV_X1 _26775_ (
    .A(_06125_),
    .ZN(_06126_)
  );
  AND2_X1 _26776_ (
    .A1(_08468_),
    .A2(_08546_),
    .ZN(_06127_)
  );
  INV_X1 _26777_ (
    .A(_06127_),
    .ZN(_06128_)
  );
  AND2_X1 _26778_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_06128_),
    .ZN(_06129_)
  );
  AND2_X1 _26779_ (
    .A1(_06126_),
    .A2(_06129_),
    .ZN(_06130_)
  );
  INV_X1 _26780_ (
    .A(_06130_),
    .ZN(_06131_)
  );
  AND2_X1 _26781_ (
    .A1(\rf[27] [1]),
    .A2(_09705_),
    .ZN(_06132_)
  );
  INV_X1 _26782_ (
    .A(_06132_),
    .ZN(_06133_)
  );
  MUX2_X1 _26783_ (
    .A(\rf[13] [1]),
    .B(\rf[9] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06134_)
  );
  AND2_X1 _26784_ (
    .A1(_08258_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_06135_)
  );
  INV_X1 _26785_ (
    .A(_06135_),
    .ZN(_06136_)
  );
  AND2_X1 _26786_ (
    .A1(_08357_),
    .A2(_08546_),
    .ZN(_06137_)
  );
  INV_X1 _26787_ (
    .A(_06137_),
    .ZN(_06138_)
  );
  MUX2_X1 _26788_ (
    .A(\rf[15] [1]),
    .B(\rf[11] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06139_)
  );
  AND2_X1 _26789_ (
    .A1(_08474_),
    .A2(_08546_),
    .ZN(_06140_)
  );
  INV_X1 _26790_ (
    .A(_06140_),
    .ZN(_06141_)
  );
  AND2_X1 _26791_ (
    .A1(_08336_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_06142_)
  );
  INV_X1 _26792_ (
    .A(_06142_),
    .ZN(_06143_)
  );
  MUX2_X1 _26793_ (
    .A(\rf[29] [1]),
    .B(\rf[25] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06144_)
  );
  AND2_X1 _26794_ (
    .A1(_08544_),
    .A2(_06144_),
    .ZN(_06145_)
  );
  INV_X1 _26795_ (
    .A(_06145_),
    .ZN(_06146_)
  );
  AND2_X1 _26796_ (
    .A1(_08435_),
    .A2(_08546_),
    .ZN(_06147_)
  );
  INV_X1 _26797_ (
    .A(_06147_),
    .ZN(_06148_)
  );
  AND2_X1 _26798_ (
    .A1(_08505_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_06149_)
  );
  INV_X1 _26799_ (
    .A(_06149_),
    .ZN(_06150_)
  );
  AND2_X1 _26800_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_06150_),
    .ZN(_06151_)
  );
  AND2_X1 _26801_ (
    .A1(_06148_),
    .A2(_06151_),
    .ZN(_06152_)
  );
  INV_X1 _26802_ (
    .A(_06152_),
    .ZN(_06153_)
  );
  AND2_X1 _26803_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_06153_),
    .ZN(_06154_)
  );
  AND2_X1 _26804_ (
    .A1(_06146_),
    .A2(_06154_),
    .ZN(_06155_)
  );
  INV_X1 _26805_ (
    .A(_06155_),
    .ZN(_06156_)
  );
  AND2_X1 _26806_ (
    .A1(_08545_),
    .A2(_06133_),
    .ZN(_06157_)
  );
  AND2_X1 _26807_ (
    .A1(_06131_),
    .A2(_06157_),
    .ZN(_06158_)
  );
  INV_X1 _26808_ (
    .A(_06158_),
    .ZN(_06159_)
  );
  AND2_X1 _26809_ (
    .A1(_08547_),
    .A2(_06159_),
    .ZN(_06160_)
  );
  AND2_X1 _26810_ (
    .A1(_06156_),
    .A2(_06160_),
    .ZN(_06161_)
  );
  INV_X1 _26811_ (
    .A(_06161_),
    .ZN(_06162_)
  );
  MUX2_X1 _26812_ (
    .A(\rf[21] [1]),
    .B(\rf[17] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06163_)
  );
  AND2_X1 _26813_ (
    .A1(_08544_),
    .A2(_06163_),
    .ZN(_06164_)
  );
  INV_X1 _26814_ (
    .A(_06164_),
    .ZN(_06165_)
  );
  AND2_X1 _26815_ (
    .A1(_08374_),
    .A2(_08546_),
    .ZN(_06166_)
  );
  INV_X1 _26816_ (
    .A(_06166_),
    .ZN(_06167_)
  );
  AND2_X1 _26817_ (
    .A1(_08275_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_06168_)
  );
  INV_X1 _26818_ (
    .A(_06168_),
    .ZN(_06169_)
  );
  AND2_X1 _26819_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_06169_),
    .ZN(_06170_)
  );
  AND2_X1 _26820_ (
    .A1(_06167_),
    .A2(_06170_),
    .ZN(_06171_)
  );
  INV_X1 _26821_ (
    .A(_06171_),
    .ZN(_06172_)
  );
  AND2_X1 _26822_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_06165_),
    .ZN(_06173_)
  );
  AND2_X1 _26823_ (
    .A1(_06172_),
    .A2(_06173_),
    .ZN(_06174_)
  );
  INV_X1 _26824_ (
    .A(_06174_),
    .ZN(_06175_)
  );
  AND2_X1 _26825_ (
    .A1(_08353_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_06176_)
  );
  INV_X1 _26826_ (
    .A(_06176_),
    .ZN(_06177_)
  );
  AND2_X1 _26827_ (
    .A1(_08491_),
    .A2(_08546_),
    .ZN(_06178_)
  );
  INV_X1 _26828_ (
    .A(_06178_),
    .ZN(_06179_)
  );
  AND2_X1 _26829_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_06179_),
    .ZN(_06180_)
  );
  AND2_X1 _26830_ (
    .A1(_06177_),
    .A2(_06180_),
    .ZN(_06181_)
  );
  INV_X1 _26831_ (
    .A(_06181_),
    .ZN(_06182_)
  );
  MUX2_X1 _26832_ (
    .A(\rf[23] [1]),
    .B(\rf[19] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06183_)
  );
  AND2_X1 _26833_ (
    .A1(_08544_),
    .A2(_06183_),
    .ZN(_06184_)
  );
  INV_X1 _26834_ (
    .A(_06184_),
    .ZN(_06185_)
  );
  AND2_X1 _26835_ (
    .A1(_08545_),
    .A2(_06185_),
    .ZN(_06186_)
  );
  AND2_X1 _26836_ (
    .A1(_06182_),
    .A2(_06186_),
    .ZN(_06187_)
  );
  INV_X1 _26837_ (
    .A(_06187_),
    .ZN(_06188_)
  );
  AND2_X1 _26838_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_06188_),
    .ZN(_06189_)
  );
  AND2_X1 _26839_ (
    .A1(_06175_),
    .A2(_06189_),
    .ZN(_06190_)
  );
  INV_X1 _26840_ (
    .A(_06190_),
    .ZN(_06191_)
  );
  AND2_X1 _26841_ (
    .A1(_08572_),
    .A2(_06191_),
    .ZN(_06192_)
  );
  AND2_X1 _26842_ (
    .A1(_06162_),
    .A2(_06192_),
    .ZN(_06193_)
  );
  INV_X1 _26843_ (
    .A(_06193_),
    .ZN(_06194_)
  );
  AND2_X1 _26844_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_06141_),
    .ZN(_06195_)
  );
  AND2_X1 _26845_ (
    .A1(_06143_),
    .A2(_06195_),
    .ZN(_06196_)
  );
  INV_X1 _26846_ (
    .A(_06196_),
    .ZN(_06197_)
  );
  AND2_X1 _26847_ (
    .A1(_08544_),
    .A2(_06139_),
    .ZN(_06198_)
  );
  INV_X1 _26848_ (
    .A(_06198_),
    .ZN(_06199_)
  );
  AND2_X1 _26849_ (
    .A1(_08545_),
    .A2(_06199_),
    .ZN(_06200_)
  );
  AND2_X1 _26850_ (
    .A1(_06197_),
    .A2(_06200_),
    .ZN(_06201_)
  );
  INV_X1 _26851_ (
    .A(_06201_),
    .ZN(_06202_)
  );
  AND2_X1 _26852_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_06136_),
    .ZN(_06203_)
  );
  AND2_X1 _26853_ (
    .A1(_06138_),
    .A2(_06203_),
    .ZN(_06204_)
  );
  INV_X1 _26854_ (
    .A(_06204_),
    .ZN(_06205_)
  );
  AND2_X1 _26855_ (
    .A1(_08544_),
    .A2(_06134_),
    .ZN(_06206_)
  );
  INV_X1 _26856_ (
    .A(_06206_),
    .ZN(_06207_)
  );
  AND2_X1 _26857_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_06207_),
    .ZN(_06208_)
  );
  AND2_X1 _26858_ (
    .A1(_06205_),
    .A2(_06208_),
    .ZN(_06209_)
  );
  INV_X1 _26859_ (
    .A(_06209_),
    .ZN(_06210_)
  );
  AND2_X1 _26860_ (
    .A1(_08547_),
    .A2(_06210_),
    .ZN(_06211_)
  );
  AND2_X1 _26861_ (
    .A1(_06202_),
    .A2(_06211_),
    .ZN(_06212_)
  );
  INV_X1 _26862_ (
    .A(_06212_),
    .ZN(_06213_)
  );
  AND2_X1 _26863_ (
    .A1(_08254_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_06214_)
  );
  INV_X1 _26864_ (
    .A(_06214_),
    .ZN(_06215_)
  );
  AND2_X1 _26865_ (
    .A1(_08249_),
    .A2(_08546_),
    .ZN(_06216_)
  );
  INV_X1 _26866_ (
    .A(_06216_),
    .ZN(_06217_)
  );
  AND2_X1 _26867_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_06217_),
    .ZN(_06218_)
  );
  AND2_X1 _26868_ (
    .A1(_06215_),
    .A2(_06218_),
    .ZN(_06219_)
  );
  INV_X1 _26869_ (
    .A(_06219_),
    .ZN(_06220_)
  );
  MUX2_X1 _26870_ (
    .A(\rf[5] [1]),
    .B(\rf[1] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06221_)
  );
  AND2_X1 _26871_ (
    .A1(_08544_),
    .A2(_06221_),
    .ZN(_06222_)
  );
  INV_X1 _26872_ (
    .A(_06222_),
    .ZN(_06223_)
  );
  AND2_X1 _26873_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_06223_),
    .ZN(_06224_)
  );
  AND2_X1 _26874_ (
    .A1(_06220_),
    .A2(_06224_),
    .ZN(_06225_)
  );
  INV_X1 _26875_ (
    .A(_06225_),
    .ZN(_06226_)
  );
  MUX2_X1 _26876_ (
    .A(\rf[7] [1]),
    .B(\rf[3] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06227_)
  );
  AND2_X1 _26877_ (
    .A1(_08544_),
    .A2(_06227_),
    .ZN(_06228_)
  );
  INV_X1 _26878_ (
    .A(_06228_),
    .ZN(_06229_)
  );
  AND2_X1 _26879_ (
    .A1(_08501_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_06230_)
  );
  INV_X1 _26880_ (
    .A(_06230_),
    .ZN(_06231_)
  );
  AND2_X1 _26881_ (
    .A1(_08245_),
    .A2(_08546_),
    .ZN(_06232_)
  );
  INV_X1 _26882_ (
    .A(_06232_),
    .ZN(_06233_)
  );
  AND2_X1 _26883_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_06233_),
    .ZN(_06234_)
  );
  AND2_X1 _26884_ (
    .A1(_06231_),
    .A2(_06234_),
    .ZN(_06235_)
  );
  INV_X1 _26885_ (
    .A(_06235_),
    .ZN(_06236_)
  );
  AND2_X1 _26886_ (
    .A1(_06229_),
    .A2(_06236_),
    .ZN(_06237_)
  );
  AND2_X1 _26887_ (
    .A1(_08545_),
    .A2(_06237_),
    .ZN(_06238_)
  );
  INV_X1 _26888_ (
    .A(_06238_),
    .ZN(_06239_)
  );
  AND2_X1 _26889_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_06226_),
    .ZN(_06240_)
  );
  AND2_X1 _26890_ (
    .A1(_06239_),
    .A2(_06240_),
    .ZN(_06241_)
  );
  INV_X1 _26891_ (
    .A(_06241_),
    .ZN(_06242_)
  );
  AND2_X1 _26892_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[4]),
    .A2(_06213_),
    .ZN(_06243_)
  );
  AND2_X1 _26893_ (
    .A1(_06242_),
    .A2(_06243_),
    .ZN(_06244_)
  );
  INV_X1 _26894_ (
    .A(_06244_),
    .ZN(_06245_)
  );
  AND2_X1 _26895_ (
    .A1(_06194_),
    .A2(_06245_),
    .ZN(_06246_)
  );
  MUX2_X1 _26896_ (
    .A(_13820_),
    .B(_06246_),
    .S(_02234_),
    .Z(_06247_)
  );
  INV_X1 _26897_ (
    .A(_06247_),
    .ZN(_06248_)
  );
  AND2_X1 _26898_ (
    .A1(_02201_),
    .A2(_06248_),
    .ZN(_06249_)
  );
  INV_X1 _26899_ (
    .A(_06249_),
    .ZN(_06250_)
  );
  AND2_X1 _26900_ (
    .A1(_13828_),
    .A2(_06250_),
    .ZN(_06251_)
  );
  MUX2_X1 _26901_ (
    .A(ex_reg_rs_lsb_1[1]),
    .B(_06251_),
    .S(_10244_),
    .Z(_00581_)
  );
  AND2_X1 _26902_ (
    .A1(_09083_),
    .A2(_09258_),
    .ZN(_06252_)
  );
  AND2_X1 _26903_ (
    .A1(_ex_reg_valid_T),
    .A2(_06252_),
    .ZN(_06253_)
  );
  INV_X1 _26904_ (
    .A(_06253_),
    .ZN(_06254_)
  );
  AND2_X1 _26905_ (
    .A1(_07940_),
    .A2(_06254_),
    .ZN(_06255_)
  );
  INV_X1 _26906_ (
    .A(_06255_),
    .ZN(_06256_)
  );
  AND2_X1 _26907_ (
    .A1(_08573_),
    .A2(_08574_),
    .ZN(_06257_)
  );
  AND2_X1 _26908_ (
    .A1(_08575_),
    .A2(_08577_),
    .ZN(_06258_)
  );
  AND2_X1 _26909_ (
    .A1(_06257_),
    .A2(_06258_),
    .ZN(_06259_)
  );
  AND2_X1 _26910_ (
    .A1(_08576_),
    .A2(_06259_),
    .ZN(_06260_)
  );
  INV_X1 _26911_ (
    .A(_06260_),
    .ZN(_06261_)
  );
  AND2_X1 _26912_ (
    .A1(_08628_),
    .A2(_06261_),
    .ZN(_06262_)
  );
  AND2_X1 _26913_ (
    .A1(_10075_),
    .A2(_06262_),
    .ZN(_06263_)
  );
  AND2_X1 _26914_ (
    .A1(_06256_),
    .A2(_06263_),
    .ZN(_00582_)
  );
  AND2_X1 _26915_ (
    .A1(csr_io_decode_0_inst[26]),
    .A2(_09289_),
    .ZN(_06264_)
  );
  INV_X1 _26916_ (
    .A(_06264_),
    .ZN(_06265_)
  );
  AND2_X1 _26917_ (
    .A1(_09251_),
    .A2(_06265_),
    .ZN(_06266_)
  );
  INV_X1 _26918_ (
    .A(_06266_),
    .ZN(_06267_)
  );
  AND2_X1 _26919_ (
    .A1(_ex_reg_valid_T),
    .A2(_06267_),
    .ZN(_06268_)
  );
  INV_X1 _26920_ (
    .A(_06268_),
    .ZN(_06269_)
  );
  AND2_X1 _26921_ (
    .A1(_09495_),
    .A2(_06269_),
    .ZN(_06270_)
  );
  INV_X1 _26922_ (
    .A(_06270_),
    .ZN(_06271_)
  );
  AND2_X1 _26923_ (
    .A1(_07954_),
    .A2(_06271_),
    .ZN(_00583_)
  );
  AND2_X1 _26924_ (
    .A1(ibuf_io_inst_0_bits_xcpt1_pf_inst),
    .A2(_05891_),
    .ZN(_06272_)
  );
  INV_X1 _26925_ (
    .A(_06272_),
    .ZN(_06273_)
  );
  AND2_X1 _26926_ (
    .A1(_08583_),
    .A2(_06273_),
    .ZN(_06274_)
  );
  INV_X1 _26927_ (
    .A(_06274_),
    .ZN(_06275_)
  );
  AND2_X1 _26928_ (
    .A1(_07941_),
    .A2(_06275_),
    .ZN(_06276_)
  );
  INV_X1 _26929_ (
    .A(_06276_),
    .ZN(_06277_)
  );
  AND2_X1 _26930_ (
    .A1(ibuf_io_inst_0_bits_xcpt1_ae_inst),
    .A2(_08565_),
    .ZN(_06278_)
  );
  INV_X1 _26931_ (
    .A(_06278_),
    .ZN(_06279_)
  );
  AND2_X1 _26932_ (
    .A1(_05891_),
    .A2(_06279_),
    .ZN(_06280_)
  );
  INV_X1 _26933_ (
    .A(_06280_),
    .ZN(_06281_)
  );
  MUX2_X1 _26934_ (
    .A(csr_io_interrupt_cause[0]),
    .B(_06281_),
    .S(_07941_),
    .Z(_06282_)
  );
  AND2_X1 _26935_ (
    .A1(_06277_),
    .A2(_06282_),
    .ZN(_06283_)
  );
  MUX2_X1 _26936_ (
    .A(_06283_),
    .B(ex_reg_cause[0]),
    .S(_05708_),
    .Z(_00584_)
  );
  AND2_X1 _26937_ (
    .A1(csr_io_interrupt),
    .A2(_08579_),
    .ZN(_06284_)
  );
  INV_X1 _26938_ (
    .A(_06284_),
    .ZN(_06285_)
  );
  AND2_X1 _26939_ (
    .A1(_08582_),
    .A2(_05894_),
    .ZN(_06286_)
  );
  AND2_X1 _26940_ (
    .A1(_05893_),
    .A2(_06286_),
    .ZN(_06287_)
  );
  INV_X1 _26941_ (
    .A(_06287_),
    .ZN(_06288_)
  );
  AND2_X1 _26942_ (
    .A1(_06285_),
    .A2(_06288_),
    .ZN(_06289_)
  );
  MUX2_X1 _26943_ (
    .A(_06289_),
    .B(ex_reg_cause[1]),
    .S(_05708_),
    .Z(_00585_)
  );
  AND2_X1 _26944_ (
    .A1(ibuf_io_inst_0_bits_xcpt1_gf_inst),
    .A2(_08566_),
    .ZN(_06290_)
  );
  AND2_X1 _26945_ (
    .A1(_05891_),
    .A2(_06290_),
    .ZN(_06291_)
  );
  AND2_X1 _26946_ (
    .A1(_05894_),
    .A2(_06291_),
    .ZN(_06292_)
  );
  INV_X1 _26947_ (
    .A(_06292_),
    .ZN(_06293_)
  );
  MUX2_X1 _26948_ (
    .A(_08580_),
    .B(_06274_),
    .S(_07941_),
    .Z(_06294_)
  );
  AND2_X1 _26949_ (
    .A1(_06293_),
    .A2(_06294_),
    .ZN(_06295_)
  );
  INV_X1 _26950_ (
    .A(_06295_),
    .ZN(_06296_)
  );
  MUX2_X1 _26951_ (
    .A(_06296_),
    .B(ex_reg_cause[2]),
    .S(_05708_),
    .Z(_00586_)
  );
  MUX2_X1 _26952_ (
    .A(csr_io_interrupt_cause[3]),
    .B(_06275_),
    .S(_07941_),
    .Z(_06297_)
  );
  MUX2_X1 _26953_ (
    .A(_06297_),
    .B(ex_reg_cause[3]),
    .S(_05708_),
    .Z(_00587_)
  );
  AND2_X1 _26954_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[4]),
    .ZN(_06298_)
  );
  INV_X1 _26955_ (
    .A(_06298_),
    .ZN(_06299_)
  );
  AND2_X1 _26956_ (
    .A1(_06293_),
    .A2(_06299_),
    .ZN(_06300_)
  );
  INV_X1 _26957_ (
    .A(_06300_),
    .ZN(_06301_)
  );
  MUX2_X1 _26958_ (
    .A(_06301_),
    .B(ex_reg_cause[4]),
    .S(_05708_),
    .Z(_00588_)
  );
  AND2_X1 _26959_ (
    .A1(_09261_),
    .A2(_09274_),
    .ZN(_06302_)
  );
  MUX2_X1 _26960_ (
    .A(ex_ctrl_csr[0]),
    .B(_06302_),
    .S(_10244_),
    .Z(_00589_)
  );
  AND2_X1 _26961_ (
    .A1(_09267_),
    .A2(_09274_),
    .ZN(_06303_)
  );
  MUX2_X1 _26962_ (
    .A(ex_ctrl_csr[2]),
    .B(_06303_),
    .S(_10244_),
    .Z(_00590_)
  );
  AND2_X1 _26963_ (
    .A1(_08222_),
    .A2(_13833_),
    .ZN(_06304_)
  );
  INV_X1 _26964_ (
    .A(_06304_),
    .ZN(_06305_)
  );
  AND2_X1 _26965_ (
    .A1(mem_reg_load),
    .A2(bpu_io_debug_ld),
    .ZN(_06306_)
  );
  INV_X1 _26966_ (
    .A(_06306_),
    .ZN(_06307_)
  );
  AND2_X1 _26967_ (
    .A1(mem_reg_store),
    .A2(bpu_io_debug_st),
    .ZN(_06308_)
  );
  INV_X1 _26968_ (
    .A(_06308_),
    .ZN(_06309_)
  );
  AND2_X1 _26969_ (
    .A1(_06307_),
    .A2(_06309_),
    .ZN(_06310_)
  );
  INV_X1 _26970_ (
    .A(_06310_),
    .ZN(_06311_)
  );
  AND2_X1 _26971_ (
    .A1(mem_reg_valid),
    .A2(_13845_),
    .ZN(_06312_)
  );
  INV_X1 _26972_ (
    .A(_06312_),
    .ZN(_06313_)
  );
  AND2_X1 _26973_ (
    .A1(_05218_),
    .A2(_06313_),
    .ZN(_06314_)
  );
  INV_X1 _26974_ (
    .A(_06314_),
    .ZN(_06315_)
  );
  AND2_X1 _26975_ (
    .A1(_06310_),
    .A2(_06314_),
    .ZN(_06316_)
  );
  INV_X1 _26976_ (
    .A(_06316_),
    .ZN(_06317_)
  );
  AND2_X1 _26977_ (
    .A1(mem_reg_cause[0]),
    .A2(_05219_),
    .ZN(_06318_)
  );
  INV_X1 _26978_ (
    .A(_06318_),
    .ZN(_06319_)
  );
  AND2_X1 _26979_ (
    .A1(_13834_),
    .A2(_06319_),
    .ZN(_06320_)
  );
  AND2_X1 _26980_ (
    .A1(_06317_),
    .A2(_06320_),
    .ZN(_06321_)
  );
  INV_X1 _26981_ (
    .A(_06321_),
    .ZN(_06322_)
  );
  AND2_X1 _26982_ (
    .A1(_06305_),
    .A2(_06322_),
    .ZN(_00591_)
  );
  AND2_X1 _26983_ (
    .A1(_08223_),
    .A2(_13833_),
    .ZN(_06323_)
  );
  INV_X1 _26984_ (
    .A(_06323_),
    .ZN(_06324_)
  );
  AND2_X1 _26985_ (
    .A1(mem_reg_cause[1]),
    .A2(_05219_),
    .ZN(_06325_)
  );
  INV_X1 _26986_ (
    .A(_06325_),
    .ZN(_06326_)
  );
  AND2_X1 _26987_ (
    .A1(_13834_),
    .A2(_06326_),
    .ZN(_06327_)
  );
  AND2_X1 _26988_ (
    .A1(_06315_),
    .A2(_06327_),
    .ZN(_06328_)
  );
  INV_X1 _26989_ (
    .A(_06328_),
    .ZN(_06329_)
  );
  AND2_X1 _26990_ (
    .A1(_06324_),
    .A2(_06329_),
    .ZN(_00592_)
  );
  AND2_X1 _26991_ (
    .A1(_08224_),
    .A2(_13833_),
    .ZN(_06330_)
  );
  INV_X1 _26992_ (
    .A(_06330_),
    .ZN(_06331_)
  );
  AND2_X1 _26993_ (
    .A1(_06311_),
    .A2(_06314_),
    .ZN(_06332_)
  );
  INV_X1 _26994_ (
    .A(_06332_),
    .ZN(_06333_)
  );
  AND2_X1 _26995_ (
    .A1(mem_reg_cause[2]),
    .A2(_05219_),
    .ZN(_06334_)
  );
  INV_X1 _26996_ (
    .A(_06334_),
    .ZN(_06335_)
  );
  AND2_X1 _26997_ (
    .A1(_13834_),
    .A2(_06335_),
    .ZN(_06336_)
  );
  AND2_X1 _26998_ (
    .A1(_06333_),
    .A2(_06336_),
    .ZN(_06337_)
  );
  INV_X1 _26999_ (
    .A(_06337_),
    .ZN(_06338_)
  );
  AND2_X1 _27000_ (
    .A1(_06331_),
    .A2(_06338_),
    .ZN(_00593_)
  );
  AND2_X1 _27001_ (
    .A1(_08225_),
    .A2(_13833_),
    .ZN(_06339_)
  );
  INV_X1 _27002_ (
    .A(_06339_),
    .ZN(_06340_)
  );
  AND2_X1 _27003_ (
    .A1(mem_reg_cause[3]),
    .A2(_05219_),
    .ZN(_06341_)
  );
  INV_X1 _27004_ (
    .A(_06341_),
    .ZN(_06342_)
  );
  AND2_X1 _27005_ (
    .A1(_13834_),
    .A2(_06342_),
    .ZN(_06343_)
  );
  AND2_X1 _27006_ (
    .A1(_06333_),
    .A2(_06343_),
    .ZN(_06344_)
  );
  INV_X1 _27007_ (
    .A(_06344_),
    .ZN(_06345_)
  );
  AND2_X1 _27008_ (
    .A1(_06340_),
    .A2(_06345_),
    .ZN(_00594_)
  );
  AND2_X1 _27009_ (
    .A1(_10088_),
    .A2(_10100_),
    .ZN(_06346_)
  );
  INV_X1 _27010_ (
    .A(_06346_),
    .ZN(_06347_)
  );
  AND2_X1 _27011_ (
    .A1(_10086_),
    .A2(_06346_),
    .ZN(_06348_)
  );
  AND2_X1 _27012_ (
    .A1(_10095_),
    .A2(_10100_),
    .ZN(_06349_)
  );
  INV_X1 _27013_ (
    .A(_06349_),
    .ZN(_06350_)
  );
  AND2_X1 _27014_ (
    .A1(_10093_),
    .A2(_06349_),
    .ZN(_06351_)
  );
  AND2_X1 _27015_ (
    .A1(_10091_),
    .A2(_06351_),
    .ZN(_06352_)
  );
  AND2_X1 _27016_ (
    .A1(_06348_),
    .A2(_06352_),
    .ZN(_06353_)
  );
  AND2_X1 _27017_ (
    .A1(_10100_),
    .A2(_13465_),
    .ZN(_06354_)
  );
  MUX2_X1 _27018_ (
    .A(\rf[9] [31]),
    .B(_06354_),
    .S(_06353_),
    .Z(_00595_)
  );
  AND2_X1 _27019_ (
    .A1(_10085_),
    .A2(_10100_),
    .ZN(_06355_)
  );
  INV_X1 _27020_ (
    .A(_06355_),
    .ZN(_06356_)
  );
  AND2_X1 _27021_ (
    .A1(_06347_),
    .A2(_06356_),
    .ZN(_06357_)
  );
  AND2_X1 _27022_ (
    .A1(_06352_),
    .A2(_06357_),
    .ZN(_06358_)
  );
  MUX2_X1 _27023_ (
    .A(\rf[8] [31]),
    .B(_06354_),
    .S(_06358_),
    .Z(_00596_)
  );
  AND2_X1 _27024_ (
    .A1(_10085_),
    .A2(_06346_),
    .ZN(_06359_)
  );
  AND2_X1 _27025_ (
    .A1(_10090_),
    .A2(_10100_),
    .ZN(_06360_)
  );
  INV_X1 _27026_ (
    .A(_06360_),
    .ZN(_06361_)
  );
  AND2_X1 _27027_ (
    .A1(_10092_),
    .A2(_10100_),
    .ZN(_06362_)
  );
  INV_X1 _27028_ (
    .A(_06362_),
    .ZN(_06363_)
  );
  AND2_X1 _27029_ (
    .A1(_06350_),
    .A2(_06363_),
    .ZN(_06364_)
  );
  AND2_X1 _27030_ (
    .A1(_06360_),
    .A2(_06364_),
    .ZN(_06365_)
  );
  AND2_X1 _27031_ (
    .A1(_06359_),
    .A2(_06365_),
    .ZN(_06366_)
  );
  MUX2_X1 _27032_ (
    .A(\rf[7] [31]),
    .B(_13465_),
    .S(_06366_),
    .Z(_00597_)
  );
  AND2_X1 _27033_ (
    .A1(_10087_),
    .A2(_06355_),
    .ZN(_06367_)
  );
  AND2_X1 _27034_ (
    .A1(_06365_),
    .A2(_06367_),
    .ZN(_06368_)
  );
  MUX2_X1 _27035_ (
    .A(\rf[6] [31]),
    .B(_06354_),
    .S(_06368_),
    .Z(_00598_)
  );
  AND2_X1 _27036_ (
    .A1(_06348_),
    .A2(_06365_),
    .ZN(_06369_)
  );
  MUX2_X1 _27037_ (
    .A(\rf[5] [31]),
    .B(_06354_),
    .S(_06369_),
    .Z(_00599_)
  );
  AND2_X1 _27038_ (
    .A1(_06357_),
    .A2(_06365_),
    .ZN(_06370_)
  );
  MUX2_X1 _27039_ (
    .A(\rf[4] [31]),
    .B(_06354_),
    .S(_06370_),
    .Z(_00600_)
  );
  AND2_X1 _27040_ (
    .A1(_06361_),
    .A2(_06364_),
    .ZN(_06371_)
  );
  AND2_X1 _27041_ (
    .A1(_06359_),
    .A2(_06371_),
    .ZN(_06372_)
  );
  MUX2_X1 _27042_ (
    .A(\rf[3] [31]),
    .B(_06354_),
    .S(_06372_),
    .Z(_00601_)
  );
  AND2_X1 _27043_ (
    .A1(_10097_),
    .A2(_06367_),
    .ZN(_06373_)
  );
  MUX2_X1 _27044_ (
    .A(\rf[30] [31]),
    .B(_06354_),
    .S(_06373_),
    .Z(_00602_)
  );
  AND2_X1 _27045_ (
    .A1(_06367_),
    .A2(_06371_),
    .ZN(_06374_)
  );
  MUX2_X1 _27046_ (
    .A(\rf[2] [31]),
    .B(_06354_),
    .S(_06374_),
    .Z(_00603_)
  );
  AND2_X1 _27047_ (
    .A1(_10097_),
    .A2(_06348_),
    .ZN(_06375_)
  );
  MUX2_X1 _27048_ (
    .A(\rf[29] [31]),
    .B(_06354_),
    .S(_06375_),
    .Z(_00604_)
  );
  AND2_X1 _27049_ (
    .A1(_10100_),
    .A2(_06357_),
    .ZN(_06376_)
  );
  AND2_X1 _27050_ (
    .A1(_10097_),
    .A2(_06376_),
    .ZN(_06377_)
  );
  MUX2_X1 _27051_ (
    .A(\rf[28] [31]),
    .B(_06354_),
    .S(_06377_),
    .Z(_00605_)
  );
  AND2_X1 _27052_ (
    .A1(_10091_),
    .A2(_10096_),
    .ZN(_06378_)
  );
  AND2_X1 _27053_ (
    .A1(_06359_),
    .A2(_06378_),
    .ZN(_06379_)
  );
  MUX2_X1 _27054_ (
    .A(\rf[27] [31]),
    .B(_06354_),
    .S(_06379_),
    .Z(_00606_)
  );
  AND2_X1 _27055_ (
    .A1(_06367_),
    .A2(_06378_),
    .ZN(_06380_)
  );
  MUX2_X1 _27056_ (
    .A(\rf[26] [31]),
    .B(_06354_),
    .S(_06380_),
    .Z(_00607_)
  );
  AND2_X1 _27057_ (
    .A1(_06348_),
    .A2(_06378_),
    .ZN(_06381_)
  );
  MUX2_X1 _27058_ (
    .A(\rf[25] [31]),
    .B(_06354_),
    .S(_06381_),
    .Z(_00608_)
  );
  AND2_X1 _27059_ (
    .A1(_06376_),
    .A2(_06378_),
    .ZN(_06382_)
  );
  MUX2_X1 _27060_ (
    .A(\rf[24] [31]),
    .B(_13465_),
    .S(_06382_),
    .Z(_00609_)
  );
  AND2_X1 _27061_ (
    .A1(_10094_),
    .A2(_06362_),
    .ZN(_06383_)
  );
  AND2_X1 _27062_ (
    .A1(_10090_),
    .A2(_06383_),
    .ZN(_06384_)
  );
  AND2_X1 _27063_ (
    .A1(_06359_),
    .A2(_06384_),
    .ZN(_06385_)
  );
  MUX2_X1 _27064_ (
    .A(\rf[23] [31]),
    .B(_06354_),
    .S(_06385_),
    .Z(_00610_)
  );
  AND2_X1 _27065_ (
    .A1(_06367_),
    .A2(_06384_),
    .ZN(_06386_)
  );
  MUX2_X1 _27066_ (
    .A(\rf[22] [31]),
    .B(_06354_),
    .S(_06386_),
    .Z(_00611_)
  );
  AND2_X1 _27067_ (
    .A1(_06348_),
    .A2(_06384_),
    .ZN(_06387_)
  );
  MUX2_X1 _27068_ (
    .A(\rf[21] [31]),
    .B(_06354_),
    .S(_06387_),
    .Z(_00612_)
  );
  AND2_X1 _27069_ (
    .A1(_06357_),
    .A2(_06384_),
    .ZN(_06388_)
  );
  MUX2_X1 _27070_ (
    .A(\rf[20] [31]),
    .B(_06354_),
    .S(_06388_),
    .Z(_00613_)
  );
  AND2_X1 _27071_ (
    .A1(_06348_),
    .A2(_06371_),
    .ZN(_06389_)
  );
  MUX2_X1 _27072_ (
    .A(\rf[1] [31]),
    .B(_06354_),
    .S(_06389_),
    .Z(_00614_)
  );
  AND2_X1 _27073_ (
    .A1(_10091_),
    .A2(_06383_),
    .ZN(_06390_)
  );
  AND2_X1 _27074_ (
    .A1(_06359_),
    .A2(_06390_),
    .ZN(_06391_)
  );
  MUX2_X1 _27075_ (
    .A(\rf[19] [31]),
    .B(_13465_),
    .S(_06391_),
    .Z(_00615_)
  );
  AND2_X1 _27076_ (
    .A1(_06367_),
    .A2(_06390_),
    .ZN(_06392_)
  );
  MUX2_X1 _27077_ (
    .A(\rf[18] [31]),
    .B(_06354_),
    .S(_06392_),
    .Z(_00616_)
  );
  AND2_X1 _27078_ (
    .A1(_06348_),
    .A2(_06390_),
    .ZN(_06393_)
  );
  MUX2_X1 _27079_ (
    .A(\rf[17] [31]),
    .B(_06354_),
    .S(_06393_),
    .Z(_00617_)
  );
  AND2_X1 _27080_ (
    .A1(_06357_),
    .A2(_06390_),
    .ZN(_06394_)
  );
  MUX2_X1 _27081_ (
    .A(\rf[16] [31]),
    .B(_06354_),
    .S(_06394_),
    .Z(_00618_)
  );
  AND2_X1 _27082_ (
    .A1(_10090_),
    .A2(_06351_),
    .ZN(_06395_)
  );
  AND2_X1 _27083_ (
    .A1(_06359_),
    .A2(_06395_),
    .ZN(_06396_)
  );
  MUX2_X1 _27084_ (
    .A(\rf[15] [31]),
    .B(_06354_),
    .S(_06396_),
    .Z(_00619_)
  );
  AND2_X1 _27085_ (
    .A1(_06367_),
    .A2(_06395_),
    .ZN(_06397_)
  );
  MUX2_X1 _27086_ (
    .A(\rf[14] [31]),
    .B(_06354_),
    .S(_06397_),
    .Z(_00620_)
  );
  AND2_X1 _27087_ (
    .A1(_06348_),
    .A2(_06395_),
    .ZN(_06398_)
  );
  MUX2_X1 _27088_ (
    .A(\rf[13] [31]),
    .B(_06354_),
    .S(_06398_),
    .Z(_00621_)
  );
  AND2_X1 _27089_ (
    .A1(_06357_),
    .A2(_06395_),
    .ZN(_06399_)
  );
  MUX2_X1 _27090_ (
    .A(\rf[12] [31]),
    .B(_06354_),
    .S(_06399_),
    .Z(_00622_)
  );
  AND2_X1 _27091_ (
    .A1(_06352_),
    .A2(_06359_),
    .ZN(_06400_)
  );
  MUX2_X1 _27092_ (
    .A(\rf[11] [31]),
    .B(_13465_),
    .S(_06400_),
    .Z(_00623_)
  );
  AND2_X1 _27093_ (
    .A1(_06352_),
    .A2(_06367_),
    .ZN(_06401_)
  );
  MUX2_X1 _27094_ (
    .A(\rf[10] [31]),
    .B(_06354_),
    .S(_06401_),
    .Z(_00624_)
  );
  AND2_X1 _27095_ (
    .A1(_06371_),
    .A2(_06376_),
    .ZN(_06402_)
  );
  MUX2_X1 _27096_ (
    .A(\rf[0] [31]),
    .B(_13465_),
    .S(_06402_),
    .Z(_00625_)
  );
  AND2_X1 _27097_ (
    .A1(_10100_),
    .A2(_13580_),
    .ZN(_06403_)
  );
  MUX2_X1 _27098_ (
    .A(\rf[25] [0]),
    .B(_06403_),
    .S(_06381_),
    .Z(_00626_)
  );
  AND2_X1 _27099_ (
    .A1(_10100_),
    .A2(_13820_),
    .ZN(_06404_)
  );
  MUX2_X1 _27100_ (
    .A(\rf[25] [1]),
    .B(_06404_),
    .S(_06381_),
    .Z(_00627_)
  );
  AND2_X1 _27101_ (
    .A1(_10100_),
    .A2(_10137_),
    .ZN(_06405_)
  );
  MUX2_X1 _27102_ (
    .A(\rf[25] [2]),
    .B(_06405_),
    .S(_06381_),
    .Z(_00628_)
  );
  AND2_X1 _27103_ (
    .A1(_10100_),
    .A2(_10250_),
    .ZN(_06406_)
  );
  MUX2_X1 _27104_ (
    .A(\rf[25] [3]),
    .B(_06406_),
    .S(_06381_),
    .Z(_00629_)
  );
  AND2_X1 _27105_ (
    .A1(_10100_),
    .A2(_10389_),
    .ZN(_06407_)
  );
  MUX2_X1 _27106_ (
    .A(\rf[25] [4]),
    .B(_06407_),
    .S(_06381_),
    .Z(_00630_)
  );
  AND2_X1 _27107_ (
    .A1(_10100_),
    .A2(_10505_),
    .ZN(_06408_)
  );
  MUX2_X1 _27108_ (
    .A(\rf[25] [5]),
    .B(_06408_),
    .S(_06381_),
    .Z(_00631_)
  );
  AND2_X1 _27109_ (
    .A1(_10100_),
    .A2(_10620_),
    .ZN(_06409_)
  );
  MUX2_X1 _27110_ (
    .A(\rf[25] [6]),
    .B(_06409_),
    .S(_06381_),
    .Z(_00632_)
  );
  AND2_X1 _27111_ (
    .A1(_10100_),
    .A2(_10733_),
    .ZN(_06410_)
  );
  MUX2_X1 _27112_ (
    .A(\rf[25] [7]),
    .B(_06410_),
    .S(_06381_),
    .Z(_00633_)
  );
  AND2_X1 _27113_ (
    .A1(_10100_),
    .A2(_10846_),
    .ZN(_06411_)
  );
  MUX2_X1 _27114_ (
    .A(\rf[25] [8]),
    .B(_06411_),
    .S(_06381_),
    .Z(_00634_)
  );
  AND2_X1 _27115_ (
    .A1(_10100_),
    .A2(_10956_),
    .ZN(_06412_)
  );
  MUX2_X1 _27116_ (
    .A(\rf[25] [9]),
    .B(_06412_),
    .S(_06381_),
    .Z(_00635_)
  );
  AND2_X1 _27117_ (
    .A1(_10100_),
    .A2(_11066_),
    .ZN(_06413_)
  );
  MUX2_X1 _27118_ (
    .A(\rf[25] [10]),
    .B(_06413_),
    .S(_06381_),
    .Z(_00636_)
  );
  AND2_X1 _27119_ (
    .A1(_10100_),
    .A2(_11205_),
    .ZN(_06414_)
  );
  MUX2_X1 _27120_ (
    .A(\rf[25] [11]),
    .B(_06414_),
    .S(_06381_),
    .Z(_00637_)
  );
  AND2_X1 _27121_ (
    .A1(_10100_),
    .A2(_11315_),
    .ZN(_06415_)
  );
  MUX2_X1 _27122_ (
    .A(\rf[25] [12]),
    .B(_06415_),
    .S(_06381_),
    .Z(_00638_)
  );
  AND2_X1 _27123_ (
    .A1(_10100_),
    .A2(_11428_),
    .ZN(_06416_)
  );
  MUX2_X1 _27124_ (
    .A(\rf[25] [13]),
    .B(_06416_),
    .S(_06381_),
    .Z(_00639_)
  );
  AND2_X1 _27125_ (
    .A1(_10100_),
    .A2(_11541_),
    .ZN(_06417_)
  );
  MUX2_X1 _27126_ (
    .A(\rf[25] [14]),
    .B(_06417_),
    .S(_06381_),
    .Z(_00640_)
  );
  AND2_X1 _27127_ (
    .A1(_10100_),
    .A2(_11656_),
    .ZN(_06418_)
  );
  MUX2_X1 _27128_ (
    .A(\rf[25] [15]),
    .B(_06418_),
    .S(_06381_),
    .Z(_00641_)
  );
  AND2_X1 _27129_ (
    .A1(_10100_),
    .A2(_11766_),
    .ZN(_06419_)
  );
  MUX2_X1 _27130_ (
    .A(\rf[25] [16]),
    .B(_06419_),
    .S(_06381_),
    .Z(_00642_)
  );
  AND2_X1 _27131_ (
    .A1(_10100_),
    .A2(_11882_),
    .ZN(_06420_)
  );
  MUX2_X1 _27132_ (
    .A(\rf[25] [17]),
    .B(_06420_),
    .S(_06381_),
    .Z(_00643_)
  );
  AND2_X1 _27133_ (
    .A1(_10100_),
    .A2(_12088_),
    .ZN(_06421_)
  );
  MUX2_X1 _27134_ (
    .A(\rf[25] [18]),
    .B(_06421_),
    .S(_06381_),
    .Z(_00644_)
  );
  AND2_X1 _27135_ (
    .A1(_10100_),
    .A2(_12099_),
    .ZN(_06422_)
  );
  MUX2_X1 _27136_ (
    .A(\rf[25] [19]),
    .B(_06422_),
    .S(_06381_),
    .Z(_00645_)
  );
  AND2_X1 _27137_ (
    .A1(_10100_),
    .A2(_12305_),
    .ZN(_06423_)
  );
  MUX2_X1 _27138_ (
    .A(\rf[25] [20]),
    .B(_06423_),
    .S(_06381_),
    .Z(_00646_)
  );
  AND2_X1 _27139_ (
    .A1(_10100_),
    .A2(_12316_),
    .ZN(_06424_)
  );
  MUX2_X1 _27140_ (
    .A(\rf[25] [21]),
    .B(_06424_),
    .S(_06381_),
    .Z(_00647_)
  );
  AND2_X1 _27141_ (
    .A1(_10100_),
    .A2(_12537_),
    .ZN(_06425_)
  );
  MUX2_X1 _27142_ (
    .A(\rf[25] [22]),
    .B(_06425_),
    .S(_06381_),
    .Z(_00648_)
  );
  AND2_X1 _27143_ (
    .A1(_10100_),
    .A2(_12638_),
    .ZN(_06426_)
  );
  MUX2_X1 _27144_ (
    .A(\rf[25] [23]),
    .B(_06426_),
    .S(_06381_),
    .Z(_00649_)
  );
  AND2_X1 _27145_ (
    .A1(_10100_),
    .A2(_12649_),
    .ZN(_06427_)
  );
  MUX2_X1 _27146_ (
    .A(\rf[25] [24]),
    .B(_06427_),
    .S(_06381_),
    .Z(_00650_)
  );
  AND2_X1 _27147_ (
    .A1(_10100_),
    .A2(_12765_),
    .ZN(_06428_)
  );
  MUX2_X1 _27148_ (
    .A(\rf[25] [25]),
    .B(_06428_),
    .S(_06381_),
    .Z(_00651_)
  );
  AND2_X1 _27149_ (
    .A1(_10100_),
    .A2(_12986_),
    .ZN(_06429_)
  );
  MUX2_X1 _27150_ (
    .A(\rf[25] [26]),
    .B(_06429_),
    .S(_06381_),
    .Z(_00652_)
  );
  AND2_X1 _27151_ (
    .A1(_10100_),
    .A2(_13102_),
    .ZN(_06430_)
  );
  MUX2_X1 _27152_ (
    .A(\rf[25] [27]),
    .B(_06430_),
    .S(_06381_),
    .Z(_00653_)
  );
  AND2_X1 _27153_ (
    .A1(_10100_),
    .A2(_13218_),
    .ZN(_06431_)
  );
  MUX2_X1 _27154_ (
    .A(\rf[25] [28]),
    .B(_06431_),
    .S(_06381_),
    .Z(_00654_)
  );
  AND2_X1 _27155_ (
    .A1(_10100_),
    .A2(_13338_),
    .ZN(_06432_)
  );
  MUX2_X1 _27156_ (
    .A(\rf[25] [29]),
    .B(_06432_),
    .S(_06381_),
    .Z(_00655_)
  );
  AND2_X1 _27157_ (
    .A1(_10100_),
    .A2(_13349_),
    .ZN(_06433_)
  );
  MUX2_X1 _27158_ (
    .A(\rf[25] [30]),
    .B(_06433_),
    .S(_06381_),
    .Z(_00656_)
  );
  MUX2_X1 _27159_ (
    .A(\rf[23] [0]),
    .B(_13580_),
    .S(_06385_),
    .Z(_00657_)
  );
  MUX2_X1 _27160_ (
    .A(\rf[23] [1]),
    .B(_06404_),
    .S(_06385_),
    .Z(_00658_)
  );
  MUX2_X1 _27161_ (
    .A(\rf[23] [2]),
    .B(_10137_),
    .S(_06385_),
    .Z(_00659_)
  );
  MUX2_X1 _27162_ (
    .A(\rf[23] [3]),
    .B(_10250_),
    .S(_06385_),
    .Z(_00660_)
  );
  MUX2_X1 _27163_ (
    .A(\rf[23] [4]),
    .B(_10389_),
    .S(_06385_),
    .Z(_00661_)
  );
  MUX2_X1 _27164_ (
    .A(\rf[23] [5]),
    .B(_10505_),
    .S(_06385_),
    .Z(_00662_)
  );
  MUX2_X1 _27165_ (
    .A(\rf[23] [6]),
    .B(_10620_),
    .S(_06385_),
    .Z(_00663_)
  );
  MUX2_X1 _27166_ (
    .A(\rf[23] [7]),
    .B(_06410_),
    .S(_06385_),
    .Z(_00664_)
  );
  MUX2_X1 _27167_ (
    .A(\rf[23] [8]),
    .B(_10846_),
    .S(_06385_),
    .Z(_00665_)
  );
  MUX2_X1 _27168_ (
    .A(\rf[23] [9]),
    .B(_10956_),
    .S(_06385_),
    .Z(_00666_)
  );
  MUX2_X1 _27169_ (
    .A(\rf[23] [10]),
    .B(_06413_),
    .S(_06385_),
    .Z(_00667_)
  );
  MUX2_X1 _27170_ (
    .A(\rf[23] [11]),
    .B(_11205_),
    .S(_06385_),
    .Z(_00668_)
  );
  MUX2_X1 _27171_ (
    .A(\rf[23] [12]),
    .B(_11315_),
    .S(_06385_),
    .Z(_00669_)
  );
  MUX2_X1 _27172_ (
    .A(\rf[23] [13]),
    .B(_11428_),
    .S(_06385_),
    .Z(_00670_)
  );
  MUX2_X1 _27173_ (
    .A(\rf[23] [14]),
    .B(_11541_),
    .S(_06385_),
    .Z(_00671_)
  );
  MUX2_X1 _27174_ (
    .A(\rf[23] [15]),
    .B(_11656_),
    .S(_06385_),
    .Z(_00672_)
  );
  MUX2_X1 _27175_ (
    .A(\rf[23] [16]),
    .B(_06419_),
    .S(_06385_),
    .Z(_00673_)
  );
  MUX2_X1 _27176_ (
    .A(\rf[23] [17]),
    .B(_11882_),
    .S(_06385_),
    .Z(_00674_)
  );
  MUX2_X1 _27177_ (
    .A(\rf[23] [18]),
    .B(_12088_),
    .S(_06385_),
    .Z(_00675_)
  );
  MUX2_X1 _27178_ (
    .A(\rf[23] [19]),
    .B(_06422_),
    .S(_06385_),
    .Z(_00676_)
  );
  MUX2_X1 _27179_ (
    .A(\rf[23] [20]),
    .B(_12305_),
    .S(_06385_),
    .Z(_00677_)
  );
  MUX2_X1 _27180_ (
    .A(\rf[23] [21]),
    .B(_06424_),
    .S(_06385_),
    .Z(_00678_)
  );
  MUX2_X1 _27181_ (
    .A(\rf[23] [22]),
    .B(_12537_),
    .S(_06385_),
    .Z(_00679_)
  );
  MUX2_X1 _27182_ (
    .A(\rf[23] [23]),
    .B(_12638_),
    .S(_06385_),
    .Z(_00680_)
  );
  MUX2_X1 _27183_ (
    .A(\rf[23] [24]),
    .B(_12649_),
    .S(_06385_),
    .Z(_00681_)
  );
  MUX2_X1 _27184_ (
    .A(\rf[23] [25]),
    .B(_12765_),
    .S(_06385_),
    .Z(_00682_)
  );
  MUX2_X1 _27185_ (
    .A(\rf[23] [26]),
    .B(_12986_),
    .S(_06385_),
    .Z(_00683_)
  );
  MUX2_X1 _27186_ (
    .A(\rf[23] [27]),
    .B(_13102_),
    .S(_06385_),
    .Z(_00684_)
  );
  MUX2_X1 _27187_ (
    .A(\rf[23] [28]),
    .B(_13218_),
    .S(_06385_),
    .Z(_00685_)
  );
  MUX2_X1 _27188_ (
    .A(\rf[23] [29]),
    .B(_13338_),
    .S(_06385_),
    .Z(_00686_)
  );
  MUX2_X1 _27189_ (
    .A(\rf[23] [30]),
    .B(_13349_),
    .S(_06385_),
    .Z(_00687_)
  );
  MUX2_X1 _27190_ (
    .A(\rf[4] [26]),
    .B(_06429_),
    .S(_06370_),
    .Z(_00688_)
  );
  MUX2_X1 _27191_ (
    .A(\rf[4] [28]),
    .B(_06431_),
    .S(_06370_),
    .Z(_00689_)
  );
  MUX2_X1 _27192_ (
    .A(\rf[4] [30]),
    .B(_06433_),
    .S(_06370_),
    .Z(_00690_)
  );
  MUX2_X1 _27193_ (
    .A(\rf[6] [0]),
    .B(_06403_),
    .S(_06368_),
    .Z(_00691_)
  );
  MUX2_X1 _27194_ (
    .A(\rf[6] [1]),
    .B(_06404_),
    .S(_06368_),
    .Z(_00692_)
  );
  MUX2_X1 _27195_ (
    .A(\rf[6] [2]),
    .B(_06405_),
    .S(_06368_),
    .Z(_00693_)
  );
  MUX2_X1 _27196_ (
    .A(\rf[6] [3]),
    .B(_06406_),
    .S(_06368_),
    .Z(_00694_)
  );
  MUX2_X1 _27197_ (
    .A(\rf[6] [4]),
    .B(_06407_),
    .S(_06368_),
    .Z(_00695_)
  );
  MUX2_X1 _27198_ (
    .A(\rf[6] [5]),
    .B(_06408_),
    .S(_06368_),
    .Z(_00696_)
  );
  MUX2_X1 _27199_ (
    .A(\rf[6] [6]),
    .B(_06409_),
    .S(_06368_),
    .Z(_00697_)
  );
  MUX2_X1 _27200_ (
    .A(\rf[6] [7]),
    .B(_06410_),
    .S(_06368_),
    .Z(_00698_)
  );
  MUX2_X1 _27201_ (
    .A(\rf[6] [8]),
    .B(_06411_),
    .S(_06368_),
    .Z(_00699_)
  );
  MUX2_X1 _27202_ (
    .A(\rf[6] [9]),
    .B(_06412_),
    .S(_06368_),
    .Z(_00700_)
  );
  MUX2_X1 _27203_ (
    .A(\rf[6] [10]),
    .B(_06413_),
    .S(_06368_),
    .Z(_00701_)
  );
  MUX2_X1 _27204_ (
    .A(\rf[6] [11]),
    .B(_06414_),
    .S(_06368_),
    .Z(_00702_)
  );
  MUX2_X1 _27205_ (
    .A(\rf[6] [12]),
    .B(_06415_),
    .S(_06368_),
    .Z(_00703_)
  );
  MUX2_X1 _27206_ (
    .A(\rf[6] [13]),
    .B(_06416_),
    .S(_06368_),
    .Z(_00704_)
  );
  MUX2_X1 _27207_ (
    .A(\rf[6] [14]),
    .B(_06417_),
    .S(_06368_),
    .Z(_00705_)
  );
  MUX2_X1 _27208_ (
    .A(\rf[6] [15]),
    .B(_06418_),
    .S(_06368_),
    .Z(_00706_)
  );
  MUX2_X1 _27209_ (
    .A(\rf[6] [16]),
    .B(_06419_),
    .S(_06368_),
    .Z(_00707_)
  );
  MUX2_X1 _27210_ (
    .A(\rf[6] [17]),
    .B(_06420_),
    .S(_06368_),
    .Z(_00708_)
  );
  MUX2_X1 _27211_ (
    .A(\rf[6] [18]),
    .B(_06421_),
    .S(_06368_),
    .Z(_00709_)
  );
  MUX2_X1 _27212_ (
    .A(\rf[6] [19]),
    .B(_06422_),
    .S(_06368_),
    .Z(_00710_)
  );
  MUX2_X1 _27213_ (
    .A(\rf[6] [20]),
    .B(_06423_),
    .S(_06368_),
    .Z(_00711_)
  );
  MUX2_X1 _27214_ (
    .A(\rf[6] [21]),
    .B(_06424_),
    .S(_06368_),
    .Z(_00712_)
  );
  MUX2_X1 _27215_ (
    .A(\rf[6] [22]),
    .B(_06425_),
    .S(_06368_),
    .Z(_00713_)
  );
  MUX2_X1 _27216_ (
    .A(\rf[6] [23]),
    .B(_06426_),
    .S(_06368_),
    .Z(_00714_)
  );
  MUX2_X1 _27217_ (
    .A(\rf[6] [24]),
    .B(_06427_),
    .S(_06368_),
    .Z(_00715_)
  );
  MUX2_X1 _27218_ (
    .A(\rf[6] [25]),
    .B(_06428_),
    .S(_06368_),
    .Z(_00716_)
  );
  MUX2_X1 _27219_ (
    .A(\rf[6] [26]),
    .B(_06429_),
    .S(_06368_),
    .Z(_00717_)
  );
  MUX2_X1 _27220_ (
    .A(\rf[6] [27]),
    .B(_06430_),
    .S(_06368_),
    .Z(_00718_)
  );
  MUX2_X1 _27221_ (
    .A(\rf[6] [28]),
    .B(_06431_),
    .S(_06368_),
    .Z(_00719_)
  );
  MUX2_X1 _27222_ (
    .A(\rf[6] [29]),
    .B(_06432_),
    .S(_06368_),
    .Z(_00720_)
  );
  MUX2_X1 _27223_ (
    .A(\rf[6] [30]),
    .B(_06433_),
    .S(_06368_),
    .Z(_00721_)
  );
  MUX2_X1 _27224_ (
    .A(\rf[4] [0]),
    .B(_06403_),
    .S(_06370_),
    .Z(_00722_)
  );
  MUX2_X1 _27225_ (
    .A(\rf[4] [1]),
    .B(_06404_),
    .S(_06370_),
    .Z(_00723_)
  );
  MUX2_X1 _27226_ (
    .A(\rf[4] [2]),
    .B(_06405_),
    .S(_06370_),
    .Z(_00724_)
  );
  MUX2_X1 _27227_ (
    .A(\rf[4] [3]),
    .B(_06406_),
    .S(_06370_),
    .Z(_00725_)
  );
  MUX2_X1 _27228_ (
    .A(\rf[4] [4]),
    .B(_06407_),
    .S(_06370_),
    .Z(_00726_)
  );
  MUX2_X1 _27229_ (
    .A(\rf[4] [5]),
    .B(_06408_),
    .S(_06370_),
    .Z(_00727_)
  );
  MUX2_X1 _27230_ (
    .A(\rf[4] [6]),
    .B(_06409_),
    .S(_06370_),
    .Z(_00728_)
  );
  MUX2_X1 _27231_ (
    .A(\rf[4] [7]),
    .B(_06410_),
    .S(_06370_),
    .Z(_00729_)
  );
  MUX2_X1 _27232_ (
    .A(\rf[4] [8]),
    .B(_06411_),
    .S(_06370_),
    .Z(_00730_)
  );
  MUX2_X1 _27233_ (
    .A(\rf[4] [9]),
    .B(_06412_),
    .S(_06370_),
    .Z(_00731_)
  );
  MUX2_X1 _27234_ (
    .A(\rf[4] [10]),
    .B(_06413_),
    .S(_06370_),
    .Z(_00732_)
  );
  MUX2_X1 _27235_ (
    .A(\rf[4] [11]),
    .B(_06414_),
    .S(_06370_),
    .Z(_00733_)
  );
  MUX2_X1 _27236_ (
    .A(\rf[4] [12]),
    .B(_06415_),
    .S(_06370_),
    .Z(_00734_)
  );
  MUX2_X1 _27237_ (
    .A(\rf[4] [13]),
    .B(_06416_),
    .S(_06370_),
    .Z(_00735_)
  );
  MUX2_X1 _27238_ (
    .A(\rf[4] [14]),
    .B(_06417_),
    .S(_06370_),
    .Z(_00736_)
  );
  MUX2_X1 _27239_ (
    .A(\rf[4] [15]),
    .B(_06418_),
    .S(_06370_),
    .Z(_00737_)
  );
  MUX2_X1 _27240_ (
    .A(\rf[4] [16]),
    .B(_06419_),
    .S(_06370_),
    .Z(_00738_)
  );
  MUX2_X1 _27241_ (
    .A(\rf[4] [17]),
    .B(_06420_),
    .S(_06370_),
    .Z(_00739_)
  );
  MUX2_X1 _27242_ (
    .A(\rf[4] [18]),
    .B(_06421_),
    .S(_06370_),
    .Z(_00740_)
  );
  MUX2_X1 _27243_ (
    .A(\rf[4] [19]),
    .B(_06422_),
    .S(_06370_),
    .Z(_00741_)
  );
  MUX2_X1 _27244_ (
    .A(\rf[4] [20]),
    .B(_06423_),
    .S(_06370_),
    .Z(_00742_)
  );
  MUX2_X1 _27245_ (
    .A(\rf[4] [21]),
    .B(_06424_),
    .S(_06370_),
    .Z(_00743_)
  );
  MUX2_X1 _27246_ (
    .A(\rf[4] [23]),
    .B(_06426_),
    .S(_06370_),
    .Z(_00744_)
  );
  MUX2_X1 _27247_ (
    .A(\rf[4] [24]),
    .B(_06427_),
    .S(_06370_),
    .Z(_00745_)
  );
  MUX2_X1 _27248_ (
    .A(\rf[4] [22]),
    .B(_06425_),
    .S(_06370_),
    .Z(_00746_)
  );
  AND2_X1 _27249_ (
    .A1(_09050_),
    .A2(_05957_),
    .ZN(_06434_)
  );
  AND2_X1 _27250_ (
    .A1(_09045_),
    .A2(_06434_),
    .ZN(_06435_)
  );
  AND2_X1 _27251_ (
    .A1(_09035_),
    .A2(_06435_),
    .ZN(_06436_)
  );
  AND2_X1 _27252_ (
    .A1(_09188_),
    .A2(_06436_),
    .ZN(_06437_)
  );
  INV_X1 _27253_ (
    .A(_06437_),
    .ZN(_06438_)
  );
  AND2_X1 _27254_ (
    .A1(_05896_),
    .A2(_06438_),
    .ZN(_06439_)
  );
  MUX2_X1 _27255_ (
    .A(ex_ctrl_sel_alu2[1]),
    .B(_06439_),
    .S(_ex_reg_valid_T),
    .Z(_00747_)
  );
  MUX2_X1 _27256_ (
    .A(\rf[4] [25]),
    .B(_06428_),
    .S(_06370_),
    .Z(_00748_)
  );
  MUX2_X1 _27257_ (
    .A(\rf[4] [27]),
    .B(_06430_),
    .S(_06370_),
    .Z(_00749_)
  );
  MUX2_X1 _27258_ (
    .A(\rf[4] [29]),
    .B(_06432_),
    .S(_06370_),
    .Z(_00750_)
  );
  MUX2_X1 _27259_ (
    .A(\rf[0] [0]),
    .B(_13580_),
    .S(_06402_),
    .Z(_00751_)
  );
  MUX2_X1 _27260_ (
    .A(\rf[0] [1]),
    .B(_13820_),
    .S(_06402_),
    .Z(_00752_)
  );
  MUX2_X1 _27261_ (
    .A(\rf[0] [2]),
    .B(_10137_),
    .S(_06402_),
    .Z(_00753_)
  );
  MUX2_X1 _27262_ (
    .A(\rf[0] [3]),
    .B(_10250_),
    .S(_06402_),
    .Z(_00754_)
  );
  MUX2_X1 _27263_ (
    .A(\rf[0] [4]),
    .B(_10389_),
    .S(_06402_),
    .Z(_00755_)
  );
  MUX2_X1 _27264_ (
    .A(\rf[0] [5]),
    .B(_10505_),
    .S(_06402_),
    .Z(_00756_)
  );
  MUX2_X1 _27265_ (
    .A(\rf[0] [6]),
    .B(_10620_),
    .S(_06402_),
    .Z(_00757_)
  );
  MUX2_X1 _27266_ (
    .A(\rf[0] [7]),
    .B(_10733_),
    .S(_06402_),
    .Z(_00758_)
  );
  MUX2_X1 _27267_ (
    .A(\rf[0] [8]),
    .B(_10846_),
    .S(_06402_),
    .Z(_00759_)
  );
  MUX2_X1 _27268_ (
    .A(\rf[0] [9]),
    .B(_10956_),
    .S(_06402_),
    .Z(_00760_)
  );
  MUX2_X1 _27269_ (
    .A(\rf[0] [10]),
    .B(_11066_),
    .S(_06402_),
    .Z(_00761_)
  );
  MUX2_X1 _27270_ (
    .A(\rf[0] [11]),
    .B(_11205_),
    .S(_06402_),
    .Z(_00762_)
  );
  MUX2_X1 _27271_ (
    .A(\rf[0] [12]),
    .B(_11315_),
    .S(_06402_),
    .Z(_00763_)
  );
  MUX2_X1 _27272_ (
    .A(\rf[0] [13]),
    .B(_11428_),
    .S(_06402_),
    .Z(_00764_)
  );
  MUX2_X1 _27273_ (
    .A(\rf[0] [14]),
    .B(_11541_),
    .S(_06402_),
    .Z(_00765_)
  );
  MUX2_X1 _27274_ (
    .A(\rf[0] [15]),
    .B(_11656_),
    .S(_06402_),
    .Z(_00766_)
  );
  MUX2_X1 _27275_ (
    .A(\rf[0] [16]),
    .B(_11766_),
    .S(_06402_),
    .Z(_00767_)
  );
  MUX2_X1 _27276_ (
    .A(\rf[0] [17]),
    .B(_11882_),
    .S(_06402_),
    .Z(_00768_)
  );
  MUX2_X1 _27277_ (
    .A(\rf[0] [18]),
    .B(_12088_),
    .S(_06402_),
    .Z(_00769_)
  );
  MUX2_X1 _27278_ (
    .A(\rf[0] [19]),
    .B(_12099_),
    .S(_06402_),
    .Z(_00770_)
  );
  MUX2_X1 _27279_ (
    .A(\rf[0] [20]),
    .B(_12305_),
    .S(_06402_),
    .Z(_00771_)
  );
  MUX2_X1 _27280_ (
    .A(\rf[0] [21]),
    .B(_12316_),
    .S(_06402_),
    .Z(_00772_)
  );
  MUX2_X1 _27281_ (
    .A(\rf[0] [22]),
    .B(_12537_),
    .S(_06402_),
    .Z(_00773_)
  );
  MUX2_X1 _27282_ (
    .A(\rf[0] [23]),
    .B(_12638_),
    .S(_06402_),
    .Z(_00774_)
  );
  MUX2_X1 _27283_ (
    .A(\rf[0] [24]),
    .B(_12649_),
    .S(_06402_),
    .Z(_00775_)
  );
  MUX2_X1 _27284_ (
    .A(\rf[0] [25]),
    .B(_12765_),
    .S(_06402_),
    .Z(_00776_)
  );
  MUX2_X1 _27285_ (
    .A(\rf[0] [26]),
    .B(_12986_),
    .S(_06402_),
    .Z(_00777_)
  );
  MUX2_X1 _27286_ (
    .A(\rf[0] [27]),
    .B(_13102_),
    .S(_06402_),
    .Z(_00778_)
  );
  MUX2_X1 _27287_ (
    .A(\rf[0] [28]),
    .B(_13218_),
    .S(_06402_),
    .Z(_00779_)
  );
  MUX2_X1 _27288_ (
    .A(\rf[0] [29]),
    .B(_13338_),
    .S(_06402_),
    .Z(_00780_)
  );
  MUX2_X1 _27289_ (
    .A(\rf[0] [30]),
    .B(_13349_),
    .S(_06402_),
    .Z(_00781_)
  );
  MUX2_X1 _27290_ (
    .A(\rf[15] [0]),
    .B(_06403_),
    .S(_06396_),
    .Z(_00782_)
  );
  MUX2_X1 _27291_ (
    .A(\rf[15] [1]),
    .B(_06404_),
    .S(_06396_),
    .Z(_00783_)
  );
  MUX2_X1 _27292_ (
    .A(\rf[15] [2]),
    .B(_10137_),
    .S(_06396_),
    .Z(_00784_)
  );
  MUX2_X1 _27293_ (
    .A(\rf[15] [3]),
    .B(_10250_),
    .S(_06396_),
    .Z(_00785_)
  );
  MUX2_X1 _27294_ (
    .A(\rf[15] [4]),
    .B(_10389_),
    .S(_06396_),
    .Z(_00786_)
  );
  MUX2_X1 _27295_ (
    .A(\rf[15] [5]),
    .B(_10505_),
    .S(_06396_),
    .Z(_00787_)
  );
  MUX2_X1 _27296_ (
    .A(\rf[15] [6]),
    .B(_06409_),
    .S(_06396_),
    .Z(_00788_)
  );
  MUX2_X1 _27297_ (
    .A(\rf[15] [7]),
    .B(_06410_),
    .S(_06396_),
    .Z(_00789_)
  );
  MUX2_X1 _27298_ (
    .A(\rf[15] [8]),
    .B(_10846_),
    .S(_06396_),
    .Z(_00790_)
  );
  MUX2_X1 _27299_ (
    .A(\rf[15] [9]),
    .B(_10956_),
    .S(_06396_),
    .Z(_00791_)
  );
  MUX2_X1 _27300_ (
    .A(\rf[15] [10]),
    .B(_11066_),
    .S(_06396_),
    .Z(_00792_)
  );
  MUX2_X1 _27301_ (
    .A(\rf[15] [11]),
    .B(_11205_),
    .S(_06396_),
    .Z(_00793_)
  );
  MUX2_X1 _27302_ (
    .A(\rf[15] [12]),
    .B(_11315_),
    .S(_06396_),
    .Z(_00794_)
  );
  MUX2_X1 _27303_ (
    .A(\rf[15] [13]),
    .B(_11428_),
    .S(_06396_),
    .Z(_00795_)
  );
  MUX2_X1 _27304_ (
    .A(\rf[15] [14]),
    .B(_11541_),
    .S(_06396_),
    .Z(_00796_)
  );
  MUX2_X1 _27305_ (
    .A(\rf[15] [15]),
    .B(_11656_),
    .S(_06396_),
    .Z(_00797_)
  );
  MUX2_X1 _27306_ (
    .A(\rf[15] [16]),
    .B(_06419_),
    .S(_06396_),
    .Z(_00798_)
  );
  MUX2_X1 _27307_ (
    .A(\rf[15] [17]),
    .B(_11882_),
    .S(_06396_),
    .Z(_00799_)
  );
  MUX2_X1 _27308_ (
    .A(\rf[15] [18]),
    .B(_06421_),
    .S(_06396_),
    .Z(_00800_)
  );
  MUX2_X1 _27309_ (
    .A(\rf[15] [19]),
    .B(_06422_),
    .S(_06396_),
    .Z(_00801_)
  );
  MUX2_X1 _27310_ (
    .A(\rf[15] [20]),
    .B(_12305_),
    .S(_06396_),
    .Z(_00802_)
  );
  MUX2_X1 _27311_ (
    .A(\rf[15] [21]),
    .B(_12316_),
    .S(_06396_),
    .Z(_00803_)
  );
  MUX2_X1 _27312_ (
    .A(\rf[15] [22]),
    .B(_12537_),
    .S(_06396_),
    .Z(_00804_)
  );
  MUX2_X1 _27313_ (
    .A(\rf[15] [23]),
    .B(_12638_),
    .S(_06396_),
    .Z(_00805_)
  );
  MUX2_X1 _27314_ (
    .A(\rf[15] [24]),
    .B(_12649_),
    .S(_06396_),
    .Z(_00806_)
  );
  MUX2_X1 _27315_ (
    .A(\rf[15] [25]),
    .B(_12765_),
    .S(_06396_),
    .Z(_00807_)
  );
  MUX2_X1 _27316_ (
    .A(\rf[15] [26]),
    .B(_12986_),
    .S(_06396_),
    .Z(_00808_)
  );
  MUX2_X1 _27317_ (
    .A(\rf[15] [27]),
    .B(_13102_),
    .S(_06396_),
    .Z(_00809_)
  );
  MUX2_X1 _27318_ (
    .A(\rf[15] [28]),
    .B(_06431_),
    .S(_06396_),
    .Z(_00810_)
  );
  MUX2_X1 _27319_ (
    .A(\rf[15] [29]),
    .B(_13338_),
    .S(_06396_),
    .Z(_00811_)
  );
  MUX2_X1 _27320_ (
    .A(\rf[15] [30]),
    .B(_13349_),
    .S(_06396_),
    .Z(_00812_)
  );
  MUX2_X1 _27321_ (
    .A(\rf[8] [0]),
    .B(_06403_),
    .S(_06358_),
    .Z(_00813_)
  );
  MUX2_X1 _27322_ (
    .A(\rf[8] [1]),
    .B(_06404_),
    .S(_06358_),
    .Z(_00814_)
  );
  MUX2_X1 _27323_ (
    .A(\rf[8] [2]),
    .B(_06405_),
    .S(_06358_),
    .Z(_00815_)
  );
  MUX2_X1 _27324_ (
    .A(\rf[8] [3]),
    .B(_06406_),
    .S(_06358_),
    .Z(_00816_)
  );
  MUX2_X1 _27325_ (
    .A(\rf[8] [4]),
    .B(_06407_),
    .S(_06358_),
    .Z(_00817_)
  );
  MUX2_X1 _27326_ (
    .A(\rf[8] [5]),
    .B(_06408_),
    .S(_06358_),
    .Z(_00818_)
  );
  MUX2_X1 _27327_ (
    .A(\rf[8] [6]),
    .B(_06409_),
    .S(_06358_),
    .Z(_00819_)
  );
  MUX2_X1 _27328_ (
    .A(\rf[8] [7]),
    .B(_06410_),
    .S(_06358_),
    .Z(_00820_)
  );
  MUX2_X1 _27329_ (
    .A(\rf[8] [8]),
    .B(_06411_),
    .S(_06358_),
    .Z(_00821_)
  );
  MUX2_X1 _27330_ (
    .A(\rf[8] [9]),
    .B(_06412_),
    .S(_06358_),
    .Z(_00822_)
  );
  MUX2_X1 _27331_ (
    .A(\rf[8] [10]),
    .B(_06413_),
    .S(_06358_),
    .Z(_00823_)
  );
  MUX2_X1 _27332_ (
    .A(\rf[8] [11]),
    .B(_06414_),
    .S(_06358_),
    .Z(_00824_)
  );
  MUX2_X1 _27333_ (
    .A(\rf[8] [12]),
    .B(_06415_),
    .S(_06358_),
    .Z(_00825_)
  );
  MUX2_X1 _27334_ (
    .A(\rf[8] [13]),
    .B(_06416_),
    .S(_06358_),
    .Z(_00826_)
  );
  MUX2_X1 _27335_ (
    .A(\rf[8] [14]),
    .B(_06417_),
    .S(_06358_),
    .Z(_00827_)
  );
  MUX2_X1 _27336_ (
    .A(\rf[8] [15]),
    .B(_06418_),
    .S(_06358_),
    .Z(_00828_)
  );
  MUX2_X1 _27337_ (
    .A(\rf[8] [16]),
    .B(_06419_),
    .S(_06358_),
    .Z(_00829_)
  );
  MUX2_X1 _27338_ (
    .A(\rf[8] [17]),
    .B(_06420_),
    .S(_06358_),
    .Z(_00830_)
  );
  MUX2_X1 _27339_ (
    .A(\rf[8] [18]),
    .B(_06421_),
    .S(_06358_),
    .Z(_00831_)
  );
  MUX2_X1 _27340_ (
    .A(\rf[8] [19]),
    .B(_06422_),
    .S(_06358_),
    .Z(_00832_)
  );
  MUX2_X1 _27341_ (
    .A(\rf[8] [20]),
    .B(_06423_),
    .S(_06358_),
    .Z(_00833_)
  );
  MUX2_X1 _27342_ (
    .A(\rf[8] [21]),
    .B(_06424_),
    .S(_06358_),
    .Z(_00834_)
  );
  MUX2_X1 _27343_ (
    .A(\rf[8] [22]),
    .B(_06425_),
    .S(_06358_),
    .Z(_00835_)
  );
  MUX2_X1 _27344_ (
    .A(\rf[8] [23]),
    .B(_06426_),
    .S(_06358_),
    .Z(_00836_)
  );
  MUX2_X1 _27345_ (
    .A(\rf[8] [24]),
    .B(_06427_),
    .S(_06358_),
    .Z(_00837_)
  );
  MUX2_X1 _27346_ (
    .A(\rf[8] [25]),
    .B(_06428_),
    .S(_06358_),
    .Z(_00838_)
  );
  MUX2_X1 _27347_ (
    .A(\rf[8] [26]),
    .B(_06429_),
    .S(_06358_),
    .Z(_00839_)
  );
  MUX2_X1 _27348_ (
    .A(\rf[8] [27]),
    .B(_06430_),
    .S(_06358_),
    .Z(_00840_)
  );
  MUX2_X1 _27349_ (
    .A(\rf[8] [28]),
    .B(_06431_),
    .S(_06358_),
    .Z(_00841_)
  );
  MUX2_X1 _27350_ (
    .A(\rf[8] [29]),
    .B(_06432_),
    .S(_06358_),
    .Z(_00842_)
  );
  MUX2_X1 _27351_ (
    .A(\rf[8] [30]),
    .B(_06433_),
    .S(_06358_),
    .Z(_00843_)
  );
  MUX2_X1 _27352_ (
    .A(\rf[16] [0]),
    .B(_06403_),
    .S(_06394_),
    .Z(_00844_)
  );
  MUX2_X1 _27353_ (
    .A(\rf[16] [1]),
    .B(_06404_),
    .S(_06394_),
    .Z(_00845_)
  );
  MUX2_X1 _27354_ (
    .A(\rf[16] [2]),
    .B(_06405_),
    .S(_06394_),
    .Z(_00846_)
  );
  MUX2_X1 _27355_ (
    .A(\rf[16] [3]),
    .B(_06406_),
    .S(_06394_),
    .Z(_00847_)
  );
  MUX2_X1 _27356_ (
    .A(\rf[16] [4]),
    .B(_06407_),
    .S(_06394_),
    .Z(_00848_)
  );
  MUX2_X1 _27357_ (
    .A(\rf[16] [5]),
    .B(_06408_),
    .S(_06394_),
    .Z(_00849_)
  );
  MUX2_X1 _27358_ (
    .A(\rf[16] [6]),
    .B(_06409_),
    .S(_06394_),
    .Z(_00850_)
  );
  MUX2_X1 _27359_ (
    .A(\rf[16] [7]),
    .B(_06410_),
    .S(_06394_),
    .Z(_00851_)
  );
  MUX2_X1 _27360_ (
    .A(\rf[16] [8]),
    .B(_06411_),
    .S(_06394_),
    .Z(_00852_)
  );
  MUX2_X1 _27361_ (
    .A(\rf[16] [9]),
    .B(_06412_),
    .S(_06394_),
    .Z(_00853_)
  );
  MUX2_X1 _27362_ (
    .A(\rf[16] [10]),
    .B(_06413_),
    .S(_06394_),
    .Z(_00854_)
  );
  MUX2_X1 _27363_ (
    .A(\rf[16] [11]),
    .B(_06414_),
    .S(_06394_),
    .Z(_00855_)
  );
  MUX2_X1 _27364_ (
    .A(\rf[16] [12]),
    .B(_06415_),
    .S(_06394_),
    .Z(_00856_)
  );
  MUX2_X1 _27365_ (
    .A(\rf[16] [13]),
    .B(_06416_),
    .S(_06394_),
    .Z(_00857_)
  );
  MUX2_X1 _27366_ (
    .A(\rf[16] [14]),
    .B(_06417_),
    .S(_06394_),
    .Z(_00858_)
  );
  MUX2_X1 _27367_ (
    .A(\rf[16] [15]),
    .B(_06418_),
    .S(_06394_),
    .Z(_00859_)
  );
  MUX2_X1 _27368_ (
    .A(\rf[16] [16]),
    .B(_06419_),
    .S(_06394_),
    .Z(_00860_)
  );
  MUX2_X1 _27369_ (
    .A(\rf[16] [17]),
    .B(_06420_),
    .S(_06394_),
    .Z(_00861_)
  );
  MUX2_X1 _27370_ (
    .A(\rf[16] [18]),
    .B(_06421_),
    .S(_06394_),
    .Z(_00862_)
  );
  MUX2_X1 _27371_ (
    .A(\rf[16] [19]),
    .B(_06422_),
    .S(_06394_),
    .Z(_00863_)
  );
  MUX2_X1 _27372_ (
    .A(\rf[16] [20]),
    .B(_06423_),
    .S(_06394_),
    .Z(_00864_)
  );
  MUX2_X1 _27373_ (
    .A(\rf[16] [21]),
    .B(_06424_),
    .S(_06394_),
    .Z(_00865_)
  );
  MUX2_X1 _27374_ (
    .A(\rf[16] [22]),
    .B(_06425_),
    .S(_06394_),
    .Z(_00866_)
  );
  MUX2_X1 _27375_ (
    .A(\rf[16] [23]),
    .B(_06426_),
    .S(_06394_),
    .Z(_00867_)
  );
  MUX2_X1 _27376_ (
    .A(\rf[16] [24]),
    .B(_06427_),
    .S(_06394_),
    .Z(_00868_)
  );
  MUX2_X1 _27377_ (
    .A(\rf[16] [25]),
    .B(_06428_),
    .S(_06394_),
    .Z(_00869_)
  );
  MUX2_X1 _27378_ (
    .A(\rf[16] [26]),
    .B(_06429_),
    .S(_06394_),
    .Z(_00870_)
  );
  MUX2_X1 _27379_ (
    .A(\rf[16] [27]),
    .B(_06430_),
    .S(_06394_),
    .Z(_00871_)
  );
  MUX2_X1 _27380_ (
    .A(\rf[16] [28]),
    .B(_06431_),
    .S(_06394_),
    .Z(_00872_)
  );
  MUX2_X1 _27381_ (
    .A(\rf[16] [29]),
    .B(_06432_),
    .S(_06394_),
    .Z(_00873_)
  );
  MUX2_X1 _27382_ (
    .A(\rf[16] [30]),
    .B(_06433_),
    .S(_06394_),
    .Z(_00874_)
  );
  MUX2_X1 _27383_ (
    .A(\rf[17] [0]),
    .B(_06403_),
    .S(_06393_),
    .Z(_00875_)
  );
  MUX2_X1 _27384_ (
    .A(\rf[17] [1]),
    .B(_06404_),
    .S(_06393_),
    .Z(_00876_)
  );
  MUX2_X1 _27385_ (
    .A(\rf[17] [2]),
    .B(_06405_),
    .S(_06393_),
    .Z(_00877_)
  );
  MUX2_X1 _27386_ (
    .A(\rf[17] [3]),
    .B(_06406_),
    .S(_06393_),
    .Z(_00878_)
  );
  MUX2_X1 _27387_ (
    .A(\rf[17] [4]),
    .B(_06407_),
    .S(_06393_),
    .Z(_00879_)
  );
  MUX2_X1 _27388_ (
    .A(\rf[17] [5]),
    .B(_06408_),
    .S(_06393_),
    .Z(_00880_)
  );
  MUX2_X1 _27389_ (
    .A(\rf[17] [6]),
    .B(_06409_),
    .S(_06393_),
    .Z(_00881_)
  );
  MUX2_X1 _27390_ (
    .A(\rf[17] [7]),
    .B(_06410_),
    .S(_06393_),
    .Z(_00882_)
  );
  MUX2_X1 _27391_ (
    .A(\rf[17] [8]),
    .B(_06411_),
    .S(_06393_),
    .Z(_00883_)
  );
  MUX2_X1 _27392_ (
    .A(\rf[17] [9]),
    .B(_06412_),
    .S(_06393_),
    .Z(_00884_)
  );
  MUX2_X1 _27393_ (
    .A(\rf[17] [10]),
    .B(_06413_),
    .S(_06393_),
    .Z(_00885_)
  );
  MUX2_X1 _27394_ (
    .A(\rf[17] [11]),
    .B(_06414_),
    .S(_06393_),
    .Z(_00886_)
  );
  MUX2_X1 _27395_ (
    .A(\rf[17] [12]),
    .B(_06415_),
    .S(_06393_),
    .Z(_00887_)
  );
  MUX2_X1 _27396_ (
    .A(\rf[17] [13]),
    .B(_06416_),
    .S(_06393_),
    .Z(_00888_)
  );
  MUX2_X1 _27397_ (
    .A(\rf[17] [14]),
    .B(_06417_),
    .S(_06393_),
    .Z(_00889_)
  );
  MUX2_X1 _27398_ (
    .A(\rf[17] [15]),
    .B(_06418_),
    .S(_06393_),
    .Z(_00890_)
  );
  MUX2_X1 _27399_ (
    .A(\rf[17] [16]),
    .B(_06419_),
    .S(_06393_),
    .Z(_00891_)
  );
  MUX2_X1 _27400_ (
    .A(\rf[17] [17]),
    .B(_06420_),
    .S(_06393_),
    .Z(_00892_)
  );
  MUX2_X1 _27401_ (
    .A(\rf[17] [18]),
    .B(_06421_),
    .S(_06393_),
    .Z(_00893_)
  );
  MUX2_X1 _27402_ (
    .A(\rf[17] [19]),
    .B(_06422_),
    .S(_06393_),
    .Z(_00894_)
  );
  MUX2_X1 _27403_ (
    .A(\rf[17] [20]),
    .B(_06423_),
    .S(_06393_),
    .Z(_00895_)
  );
  MUX2_X1 _27404_ (
    .A(\rf[17] [21]),
    .B(_06424_),
    .S(_06393_),
    .Z(_00896_)
  );
  MUX2_X1 _27405_ (
    .A(\rf[17] [22]),
    .B(_06425_),
    .S(_06393_),
    .Z(_00897_)
  );
  MUX2_X1 _27406_ (
    .A(\rf[17] [23]),
    .B(_06426_),
    .S(_06393_),
    .Z(_00898_)
  );
  MUX2_X1 _27407_ (
    .A(\rf[17] [24]),
    .B(_06427_),
    .S(_06393_),
    .Z(_00899_)
  );
  MUX2_X1 _27408_ (
    .A(\rf[17] [25]),
    .B(_06428_),
    .S(_06393_),
    .Z(_00900_)
  );
  MUX2_X1 _27409_ (
    .A(\rf[17] [26]),
    .B(_06429_),
    .S(_06393_),
    .Z(_00901_)
  );
  MUX2_X1 _27410_ (
    .A(\rf[17] [27]),
    .B(_06430_),
    .S(_06393_),
    .Z(_00902_)
  );
  MUX2_X1 _27411_ (
    .A(\rf[17] [28]),
    .B(_06431_),
    .S(_06393_),
    .Z(_00903_)
  );
  MUX2_X1 _27412_ (
    .A(\rf[17] [29]),
    .B(_06432_),
    .S(_06393_),
    .Z(_00904_)
  );
  MUX2_X1 _27413_ (
    .A(\rf[17] [30]),
    .B(_06433_),
    .S(_06393_),
    .Z(_00905_)
  );
  MUX2_X1 _27414_ (
    .A(\rf[10] [0]),
    .B(_06403_),
    .S(_06401_),
    .Z(_00906_)
  );
  MUX2_X1 _27415_ (
    .A(\rf[10] [1]),
    .B(_06404_),
    .S(_06401_),
    .Z(_00907_)
  );
  MUX2_X1 _27416_ (
    .A(\rf[10] [2]),
    .B(_06405_),
    .S(_06401_),
    .Z(_00908_)
  );
  MUX2_X1 _27417_ (
    .A(\rf[10] [3]),
    .B(_06406_),
    .S(_06401_),
    .Z(_00909_)
  );
  MUX2_X1 _27418_ (
    .A(\rf[10] [4]),
    .B(_06407_),
    .S(_06401_),
    .Z(_00910_)
  );
  MUX2_X1 _27419_ (
    .A(\rf[10] [5]),
    .B(_06408_),
    .S(_06401_),
    .Z(_00911_)
  );
  MUX2_X1 _27420_ (
    .A(\rf[10] [6]),
    .B(_06409_),
    .S(_06401_),
    .Z(_00912_)
  );
  MUX2_X1 _27421_ (
    .A(\rf[10] [7]),
    .B(_06410_),
    .S(_06401_),
    .Z(_00913_)
  );
  MUX2_X1 _27422_ (
    .A(\rf[10] [8]),
    .B(_06411_),
    .S(_06401_),
    .Z(_00914_)
  );
  MUX2_X1 _27423_ (
    .A(\rf[10] [9]),
    .B(_06412_),
    .S(_06401_),
    .Z(_00915_)
  );
  MUX2_X1 _27424_ (
    .A(\rf[10] [10]),
    .B(_06413_),
    .S(_06401_),
    .Z(_00916_)
  );
  MUX2_X1 _27425_ (
    .A(\rf[10] [11]),
    .B(_06414_),
    .S(_06401_),
    .Z(_00917_)
  );
  MUX2_X1 _27426_ (
    .A(\rf[10] [12]),
    .B(_06415_),
    .S(_06401_),
    .Z(_00918_)
  );
  MUX2_X1 _27427_ (
    .A(\rf[10] [13]),
    .B(_06416_),
    .S(_06401_),
    .Z(_00919_)
  );
  MUX2_X1 _27428_ (
    .A(\rf[10] [14]),
    .B(_06417_),
    .S(_06401_),
    .Z(_00920_)
  );
  MUX2_X1 _27429_ (
    .A(\rf[10] [15]),
    .B(_06418_),
    .S(_06401_),
    .Z(_00921_)
  );
  MUX2_X1 _27430_ (
    .A(\rf[10] [16]),
    .B(_06419_),
    .S(_06401_),
    .Z(_00922_)
  );
  MUX2_X1 _27431_ (
    .A(\rf[10] [17]),
    .B(_06420_),
    .S(_06401_),
    .Z(_00923_)
  );
  MUX2_X1 _27432_ (
    .A(\rf[10] [18]),
    .B(_06421_),
    .S(_06401_),
    .Z(_00924_)
  );
  MUX2_X1 _27433_ (
    .A(\rf[10] [19]),
    .B(_06422_),
    .S(_06401_),
    .Z(_00925_)
  );
  MUX2_X1 _27434_ (
    .A(\rf[10] [20]),
    .B(_06423_),
    .S(_06401_),
    .Z(_00926_)
  );
  MUX2_X1 _27435_ (
    .A(\rf[10] [21]),
    .B(_06424_),
    .S(_06401_),
    .Z(_00927_)
  );
  MUX2_X1 _27436_ (
    .A(\rf[10] [22]),
    .B(_06425_),
    .S(_06401_),
    .Z(_00928_)
  );
  MUX2_X1 _27437_ (
    .A(\rf[10] [23]),
    .B(_06426_),
    .S(_06401_),
    .Z(_00929_)
  );
  MUX2_X1 _27438_ (
    .A(\rf[10] [24]),
    .B(_06427_),
    .S(_06401_),
    .Z(_00930_)
  );
  MUX2_X1 _27439_ (
    .A(\rf[10] [25]),
    .B(_06428_),
    .S(_06401_),
    .Z(_00931_)
  );
  MUX2_X1 _27440_ (
    .A(\rf[10] [26]),
    .B(_06429_),
    .S(_06401_),
    .Z(_00932_)
  );
  MUX2_X1 _27441_ (
    .A(\rf[10] [27]),
    .B(_06430_),
    .S(_06401_),
    .Z(_00933_)
  );
  MUX2_X1 _27442_ (
    .A(\rf[10] [28]),
    .B(_06431_),
    .S(_06401_),
    .Z(_00934_)
  );
  MUX2_X1 _27443_ (
    .A(\rf[10] [29]),
    .B(_06432_),
    .S(_06401_),
    .Z(_00935_)
  );
  MUX2_X1 _27444_ (
    .A(\rf[10] [30]),
    .B(_06433_),
    .S(_06401_),
    .Z(_00936_)
  );
  MUX2_X1 _27445_ (
    .A(\rf[18] [0]),
    .B(_06403_),
    .S(_06392_),
    .Z(_00937_)
  );
  MUX2_X1 _27446_ (
    .A(\rf[18] [1]),
    .B(_06404_),
    .S(_06392_),
    .Z(_00938_)
  );
  MUX2_X1 _27447_ (
    .A(\rf[18] [2]),
    .B(_06405_),
    .S(_06392_),
    .Z(_00939_)
  );
  MUX2_X1 _27448_ (
    .A(\rf[18] [3]),
    .B(_06406_),
    .S(_06392_),
    .Z(_00940_)
  );
  MUX2_X1 _27449_ (
    .A(\rf[18] [4]),
    .B(_06407_),
    .S(_06392_),
    .Z(_00941_)
  );
  MUX2_X1 _27450_ (
    .A(\rf[18] [5]),
    .B(_06408_),
    .S(_06392_),
    .Z(_00942_)
  );
  MUX2_X1 _27451_ (
    .A(\rf[18] [6]),
    .B(_06409_),
    .S(_06392_),
    .Z(_00943_)
  );
  MUX2_X1 _27452_ (
    .A(\rf[18] [7]),
    .B(_06410_),
    .S(_06392_),
    .Z(_00944_)
  );
  MUX2_X1 _27453_ (
    .A(\rf[18] [8]),
    .B(_06411_),
    .S(_06392_),
    .Z(_00945_)
  );
  MUX2_X1 _27454_ (
    .A(\rf[18] [9]),
    .B(_06412_),
    .S(_06392_),
    .Z(_00946_)
  );
  MUX2_X1 _27455_ (
    .A(\rf[18] [10]),
    .B(_06413_),
    .S(_06392_),
    .Z(_00947_)
  );
  MUX2_X1 _27456_ (
    .A(\rf[18] [11]),
    .B(_06414_),
    .S(_06392_),
    .Z(_00948_)
  );
  MUX2_X1 _27457_ (
    .A(\rf[18] [12]),
    .B(_06415_),
    .S(_06392_),
    .Z(_00949_)
  );
  MUX2_X1 _27458_ (
    .A(\rf[18] [13]),
    .B(_06416_),
    .S(_06392_),
    .Z(_00950_)
  );
  MUX2_X1 _27459_ (
    .A(\rf[18] [14]),
    .B(_06417_),
    .S(_06392_),
    .Z(_00951_)
  );
  MUX2_X1 _27460_ (
    .A(\rf[18] [15]),
    .B(_06418_),
    .S(_06392_),
    .Z(_00952_)
  );
  MUX2_X1 _27461_ (
    .A(\rf[18] [16]),
    .B(_06419_),
    .S(_06392_),
    .Z(_00953_)
  );
  MUX2_X1 _27462_ (
    .A(\rf[18] [17]),
    .B(_06420_),
    .S(_06392_),
    .Z(_00954_)
  );
  MUX2_X1 _27463_ (
    .A(\rf[18] [18]),
    .B(_06421_),
    .S(_06392_),
    .Z(_00955_)
  );
  MUX2_X1 _27464_ (
    .A(\rf[18] [19]),
    .B(_06422_),
    .S(_06392_),
    .Z(_00956_)
  );
  MUX2_X1 _27465_ (
    .A(\rf[18] [20]),
    .B(_06423_),
    .S(_06392_),
    .Z(_00957_)
  );
  MUX2_X1 _27466_ (
    .A(\rf[18] [21]),
    .B(_06424_),
    .S(_06392_),
    .Z(_00958_)
  );
  MUX2_X1 _27467_ (
    .A(\rf[18] [22]),
    .B(_06425_),
    .S(_06392_),
    .Z(_00959_)
  );
  MUX2_X1 _27468_ (
    .A(\rf[18] [23]),
    .B(_06426_),
    .S(_06392_),
    .Z(_00960_)
  );
  MUX2_X1 _27469_ (
    .A(\rf[18] [24]),
    .B(_06427_),
    .S(_06392_),
    .Z(_00961_)
  );
  MUX2_X1 _27470_ (
    .A(\rf[18] [25]),
    .B(_06428_),
    .S(_06392_),
    .Z(_00962_)
  );
  MUX2_X1 _27471_ (
    .A(\rf[18] [26]),
    .B(_06429_),
    .S(_06392_),
    .Z(_00963_)
  );
  MUX2_X1 _27472_ (
    .A(\rf[18] [27]),
    .B(_06430_),
    .S(_06392_),
    .Z(_00964_)
  );
  MUX2_X1 _27473_ (
    .A(\rf[18] [28]),
    .B(_06431_),
    .S(_06392_),
    .Z(_00965_)
  );
  MUX2_X1 _27474_ (
    .A(\rf[18] [29]),
    .B(_06432_),
    .S(_06392_),
    .Z(_00966_)
  );
  MUX2_X1 _27475_ (
    .A(\rf[18] [30]),
    .B(_06433_),
    .S(_06392_),
    .Z(_00967_)
  );
  MUX2_X1 _27476_ (
    .A(\rf[11] [0]),
    .B(_06403_),
    .S(_06400_),
    .Z(_00968_)
  );
  MUX2_X1 _27477_ (
    .A(\rf[11] [1]),
    .B(_06404_),
    .S(_06400_),
    .Z(_00969_)
  );
  MUX2_X1 _27478_ (
    .A(\rf[11] [2]),
    .B(_10137_),
    .S(_06400_),
    .Z(_00970_)
  );
  MUX2_X1 _27479_ (
    .A(\rf[11] [3]),
    .B(_10250_),
    .S(_06400_),
    .Z(_00971_)
  );
  MUX2_X1 _27480_ (
    .A(\rf[11] [4]),
    .B(_10389_),
    .S(_06400_),
    .Z(_00972_)
  );
  MUX2_X1 _27481_ (
    .A(\rf[11] [5]),
    .B(_10505_),
    .S(_06400_),
    .Z(_00973_)
  );
  MUX2_X1 _27482_ (
    .A(\rf[11] [6]),
    .B(_06409_),
    .S(_06400_),
    .Z(_00974_)
  );
  MUX2_X1 _27483_ (
    .A(\rf[11] [7]),
    .B(_06410_),
    .S(_06400_),
    .Z(_00975_)
  );
  MUX2_X1 _27484_ (
    .A(\rf[11] [8]),
    .B(_06411_),
    .S(_06400_),
    .Z(_00976_)
  );
  MUX2_X1 _27485_ (
    .A(\rf[11] [9]),
    .B(_06412_),
    .S(_06400_),
    .Z(_00977_)
  );
  MUX2_X1 _27486_ (
    .A(\rf[11] [10]),
    .B(_06413_),
    .S(_06400_),
    .Z(_00978_)
  );
  MUX2_X1 _27487_ (
    .A(\rf[11] [11]),
    .B(_11205_),
    .S(_06400_),
    .Z(_00979_)
  );
  MUX2_X1 _27488_ (
    .A(\rf[11] [12]),
    .B(_11315_),
    .S(_06400_),
    .Z(_00980_)
  );
  MUX2_X1 _27489_ (
    .A(\rf[11] [13]),
    .B(_11428_),
    .S(_06400_),
    .Z(_00981_)
  );
  MUX2_X1 _27490_ (
    .A(\rf[11] [14]),
    .B(_06417_),
    .S(_06400_),
    .Z(_00982_)
  );
  MUX2_X1 _27491_ (
    .A(\rf[11] [15]),
    .B(_11656_),
    .S(_06400_),
    .Z(_00983_)
  );
  MUX2_X1 _27492_ (
    .A(\rf[11] [16]),
    .B(_06419_),
    .S(_06400_),
    .Z(_00984_)
  );
  MUX2_X1 _27493_ (
    .A(\rf[11] [17]),
    .B(_11882_),
    .S(_06400_),
    .Z(_00985_)
  );
  MUX2_X1 _27494_ (
    .A(\rf[11] [18]),
    .B(_06421_),
    .S(_06400_),
    .Z(_00986_)
  );
  MUX2_X1 _27495_ (
    .A(\rf[11] [19]),
    .B(_06422_),
    .S(_06400_),
    .Z(_00987_)
  );
  MUX2_X1 _27496_ (
    .A(\rf[11] [20]),
    .B(_12305_),
    .S(_06400_),
    .Z(_00988_)
  );
  MUX2_X1 _27497_ (
    .A(\rf[11] [21]),
    .B(_06424_),
    .S(_06400_),
    .Z(_00989_)
  );
  MUX2_X1 _27498_ (
    .A(\rf[11] [22]),
    .B(_12537_),
    .S(_06400_),
    .Z(_00990_)
  );
  MUX2_X1 _27499_ (
    .A(\rf[11] [23]),
    .B(_12638_),
    .S(_06400_),
    .Z(_00991_)
  );
  MUX2_X1 _27500_ (
    .A(\rf[11] [24]),
    .B(_12649_),
    .S(_06400_),
    .Z(_00992_)
  );
  MUX2_X1 _27501_ (
    .A(\rf[11] [25]),
    .B(_06428_),
    .S(_06400_),
    .Z(_00993_)
  );
  MUX2_X1 _27502_ (
    .A(\rf[11] [26]),
    .B(_12986_),
    .S(_06400_),
    .Z(_00994_)
  );
  MUX2_X1 _27503_ (
    .A(\rf[11] [27]),
    .B(_06430_),
    .S(_06400_),
    .Z(_00995_)
  );
  MUX2_X1 _27504_ (
    .A(\rf[11] [28]),
    .B(_06431_),
    .S(_06400_),
    .Z(_00996_)
  );
  MUX2_X1 _27505_ (
    .A(\rf[11] [29]),
    .B(_06432_),
    .S(_06400_),
    .Z(_00997_)
  );
  MUX2_X1 _27506_ (
    .A(\rf[11] [30]),
    .B(_13349_),
    .S(_06400_),
    .Z(_00998_)
  );
  MUX2_X1 _27507_ (
    .A(\rf[19] [0]),
    .B(_13580_),
    .S(_06391_),
    .Z(_00999_)
  );
  MUX2_X1 _27508_ (
    .A(\rf[19] [1]),
    .B(_06404_),
    .S(_06391_),
    .Z(_01000_)
  );
  MUX2_X1 _27509_ (
    .A(\rf[19] [2]),
    .B(_10137_),
    .S(_06391_),
    .Z(_01001_)
  );
  MUX2_X1 _27510_ (
    .A(\rf[19] [3]),
    .B(_10250_),
    .S(_06391_),
    .Z(_01002_)
  );
  MUX2_X1 _27511_ (
    .A(\rf[19] [4]),
    .B(_10389_),
    .S(_06391_),
    .Z(_01003_)
  );
  MUX2_X1 _27512_ (
    .A(\rf[19] [5]),
    .B(_10505_),
    .S(_06391_),
    .Z(_01004_)
  );
  MUX2_X1 _27513_ (
    .A(\rf[19] [6]),
    .B(_10620_),
    .S(_06391_),
    .Z(_01005_)
  );
  MUX2_X1 _27514_ (
    .A(\rf[19] [7]),
    .B(_06410_),
    .S(_06391_),
    .Z(_01006_)
  );
  MUX2_X1 _27515_ (
    .A(\rf[19] [8]),
    .B(_10846_),
    .S(_06391_),
    .Z(_01007_)
  );
  MUX2_X1 _27516_ (
    .A(\rf[19] [9]),
    .B(_10956_),
    .S(_06391_),
    .Z(_01008_)
  );
  MUX2_X1 _27517_ (
    .A(\rf[19] [10]),
    .B(_11066_),
    .S(_06391_),
    .Z(_01009_)
  );
  MUX2_X1 _27518_ (
    .A(\rf[19] [11]),
    .B(_11205_),
    .S(_06391_),
    .Z(_01010_)
  );
  MUX2_X1 _27519_ (
    .A(\rf[19] [12]),
    .B(_11315_),
    .S(_06391_),
    .Z(_01011_)
  );
  MUX2_X1 _27520_ (
    .A(\rf[19] [13]),
    .B(_11428_),
    .S(_06391_),
    .Z(_01012_)
  );
  MUX2_X1 _27521_ (
    .A(\rf[19] [14]),
    .B(_11541_),
    .S(_06391_),
    .Z(_01013_)
  );
  MUX2_X1 _27522_ (
    .A(\rf[19] [15]),
    .B(_11656_),
    .S(_06391_),
    .Z(_01014_)
  );
  MUX2_X1 _27523_ (
    .A(\rf[19] [16]),
    .B(_06419_),
    .S(_06391_),
    .Z(_01015_)
  );
  MUX2_X1 _27524_ (
    .A(\rf[19] [17]),
    .B(_11882_),
    .S(_06391_),
    .Z(_01016_)
  );
  MUX2_X1 _27525_ (
    .A(\rf[19] [18]),
    .B(_12088_),
    .S(_06391_),
    .Z(_01017_)
  );
  MUX2_X1 _27526_ (
    .A(\rf[19] [19]),
    .B(_06422_),
    .S(_06391_),
    .Z(_01018_)
  );
  MUX2_X1 _27527_ (
    .A(\rf[19] [20]),
    .B(_12305_),
    .S(_06391_),
    .Z(_01019_)
  );
  MUX2_X1 _27528_ (
    .A(\rf[19] [21]),
    .B(_06424_),
    .S(_06391_),
    .Z(_01020_)
  );
  MUX2_X1 _27529_ (
    .A(\rf[19] [22]),
    .B(_12537_),
    .S(_06391_),
    .Z(_01021_)
  );
  MUX2_X1 _27530_ (
    .A(\rf[19] [23]),
    .B(_12638_),
    .S(_06391_),
    .Z(_01022_)
  );
  MUX2_X1 _27531_ (
    .A(\rf[19] [24]),
    .B(_12649_),
    .S(_06391_),
    .Z(_01023_)
  );
  MUX2_X1 _27532_ (
    .A(\rf[19] [25]),
    .B(_06428_),
    .S(_06391_),
    .Z(_01024_)
  );
  MUX2_X1 _27533_ (
    .A(\rf[19] [26]),
    .B(_12986_),
    .S(_06391_),
    .Z(_01025_)
  );
  MUX2_X1 _27534_ (
    .A(\rf[19] [27]),
    .B(_13102_),
    .S(_06391_),
    .Z(_01026_)
  );
  MUX2_X1 _27535_ (
    .A(\rf[19] [28]),
    .B(_13218_),
    .S(_06391_),
    .Z(_01027_)
  );
  MUX2_X1 _27536_ (
    .A(\rf[19] [29]),
    .B(_13338_),
    .S(_06391_),
    .Z(_01028_)
  );
  MUX2_X1 _27537_ (
    .A(\rf[19] [30]),
    .B(_13349_),
    .S(_06391_),
    .Z(_01029_)
  );
  MUX2_X1 _27538_ (
    .A(\rf[12] [0]),
    .B(_06403_),
    .S(_06399_),
    .Z(_01030_)
  );
  MUX2_X1 _27539_ (
    .A(\rf[12] [1]),
    .B(_06404_),
    .S(_06399_),
    .Z(_01031_)
  );
  MUX2_X1 _27540_ (
    .A(\rf[12] [2]),
    .B(_06405_),
    .S(_06399_),
    .Z(_01032_)
  );
  MUX2_X1 _27541_ (
    .A(\rf[12] [3]),
    .B(_06406_),
    .S(_06399_),
    .Z(_01033_)
  );
  MUX2_X1 _27542_ (
    .A(\rf[12] [4]),
    .B(_06407_),
    .S(_06399_),
    .Z(_01034_)
  );
  MUX2_X1 _27543_ (
    .A(\rf[12] [5]),
    .B(_06408_),
    .S(_06399_),
    .Z(_01035_)
  );
  MUX2_X1 _27544_ (
    .A(\rf[12] [6]),
    .B(_06409_),
    .S(_06399_),
    .Z(_01036_)
  );
  MUX2_X1 _27545_ (
    .A(\rf[12] [7]),
    .B(_06410_),
    .S(_06399_),
    .Z(_01037_)
  );
  MUX2_X1 _27546_ (
    .A(\rf[12] [8]),
    .B(_06411_),
    .S(_06399_),
    .Z(_01038_)
  );
  MUX2_X1 _27547_ (
    .A(\rf[12] [9]),
    .B(_06412_),
    .S(_06399_),
    .Z(_01039_)
  );
  MUX2_X1 _27548_ (
    .A(\rf[12] [10]),
    .B(_06413_),
    .S(_06399_),
    .Z(_01040_)
  );
  MUX2_X1 _27549_ (
    .A(\rf[12] [11]),
    .B(_06414_),
    .S(_06399_),
    .Z(_01041_)
  );
  MUX2_X1 _27550_ (
    .A(\rf[12] [12]),
    .B(_06415_),
    .S(_06399_),
    .Z(_01042_)
  );
  MUX2_X1 _27551_ (
    .A(\rf[12] [13]),
    .B(_06416_),
    .S(_06399_),
    .Z(_01043_)
  );
  MUX2_X1 _27552_ (
    .A(\rf[12] [14]),
    .B(_06417_),
    .S(_06399_),
    .Z(_01044_)
  );
  MUX2_X1 _27553_ (
    .A(\rf[12] [15]),
    .B(_06418_),
    .S(_06399_),
    .Z(_01045_)
  );
  MUX2_X1 _27554_ (
    .A(\rf[12] [16]),
    .B(_06419_),
    .S(_06399_),
    .Z(_01046_)
  );
  MUX2_X1 _27555_ (
    .A(\rf[12] [17]),
    .B(_06420_),
    .S(_06399_),
    .Z(_01047_)
  );
  MUX2_X1 _27556_ (
    .A(\rf[12] [18]),
    .B(_06421_),
    .S(_06399_),
    .Z(_01048_)
  );
  MUX2_X1 _27557_ (
    .A(\rf[12] [19]),
    .B(_06422_),
    .S(_06399_),
    .Z(_01049_)
  );
  MUX2_X1 _27558_ (
    .A(\rf[12] [20]),
    .B(_06423_),
    .S(_06399_),
    .Z(_01050_)
  );
  MUX2_X1 _27559_ (
    .A(\rf[12] [21]),
    .B(_06424_),
    .S(_06399_),
    .Z(_01051_)
  );
  MUX2_X1 _27560_ (
    .A(\rf[12] [22]),
    .B(_06425_),
    .S(_06399_),
    .Z(_01052_)
  );
  MUX2_X1 _27561_ (
    .A(\rf[12] [23]),
    .B(_06426_),
    .S(_06399_),
    .Z(_01053_)
  );
  MUX2_X1 _27562_ (
    .A(\rf[12] [24]),
    .B(_06427_),
    .S(_06399_),
    .Z(_01054_)
  );
  MUX2_X1 _27563_ (
    .A(\rf[12] [25]),
    .B(_06428_),
    .S(_06399_),
    .Z(_01055_)
  );
  MUX2_X1 _27564_ (
    .A(\rf[12] [26]),
    .B(_06429_),
    .S(_06399_),
    .Z(_01056_)
  );
  MUX2_X1 _27565_ (
    .A(\rf[12] [27]),
    .B(_06430_),
    .S(_06399_),
    .Z(_01057_)
  );
  MUX2_X1 _27566_ (
    .A(\rf[12] [28]),
    .B(_06431_),
    .S(_06399_),
    .Z(_01058_)
  );
  MUX2_X1 _27567_ (
    .A(\rf[12] [29]),
    .B(_06432_),
    .S(_06399_),
    .Z(_01059_)
  );
  MUX2_X1 _27568_ (
    .A(\rf[12] [30]),
    .B(_06433_),
    .S(_06399_),
    .Z(_01060_)
  );
  MUX2_X1 _27569_ (
    .A(\rf[20] [0]),
    .B(_06403_),
    .S(_06388_),
    .Z(_01061_)
  );
  MUX2_X1 _27570_ (
    .A(\rf[20] [1]),
    .B(_06404_),
    .S(_06388_),
    .Z(_01062_)
  );
  MUX2_X1 _27571_ (
    .A(\rf[20] [2]),
    .B(_06405_),
    .S(_06388_),
    .Z(_01063_)
  );
  MUX2_X1 _27572_ (
    .A(\rf[20] [3]),
    .B(_06406_),
    .S(_06388_),
    .Z(_01064_)
  );
  MUX2_X1 _27573_ (
    .A(\rf[20] [4]),
    .B(_06407_),
    .S(_06388_),
    .Z(_01065_)
  );
  MUX2_X1 _27574_ (
    .A(\rf[20] [5]),
    .B(_06408_),
    .S(_06388_),
    .Z(_01066_)
  );
  MUX2_X1 _27575_ (
    .A(\rf[20] [6]),
    .B(_06409_),
    .S(_06388_),
    .Z(_01067_)
  );
  MUX2_X1 _27576_ (
    .A(\rf[20] [7]),
    .B(_06410_),
    .S(_06388_),
    .Z(_01068_)
  );
  MUX2_X1 _27577_ (
    .A(\rf[20] [8]),
    .B(_06411_),
    .S(_06388_),
    .Z(_01069_)
  );
  MUX2_X1 _27578_ (
    .A(\rf[20] [9]),
    .B(_06412_),
    .S(_06388_),
    .Z(_01070_)
  );
  MUX2_X1 _27579_ (
    .A(\rf[20] [10]),
    .B(_06413_),
    .S(_06388_),
    .Z(_01071_)
  );
  MUX2_X1 _27580_ (
    .A(\rf[20] [11]),
    .B(_06414_),
    .S(_06388_),
    .Z(_01072_)
  );
  MUX2_X1 _27581_ (
    .A(\rf[20] [12]),
    .B(_06415_),
    .S(_06388_),
    .Z(_01073_)
  );
  MUX2_X1 _27582_ (
    .A(\rf[20] [13]),
    .B(_06416_),
    .S(_06388_),
    .Z(_01074_)
  );
  MUX2_X1 _27583_ (
    .A(\rf[20] [14]),
    .B(_06417_),
    .S(_06388_),
    .Z(_01075_)
  );
  MUX2_X1 _27584_ (
    .A(\rf[20] [15]),
    .B(_06418_),
    .S(_06388_),
    .Z(_01076_)
  );
  MUX2_X1 _27585_ (
    .A(\rf[20] [16]),
    .B(_06419_),
    .S(_06388_),
    .Z(_01077_)
  );
  MUX2_X1 _27586_ (
    .A(\rf[20] [17]),
    .B(_06420_),
    .S(_06388_),
    .Z(_01078_)
  );
  MUX2_X1 _27587_ (
    .A(\rf[20] [18]),
    .B(_06421_),
    .S(_06388_),
    .Z(_01079_)
  );
  MUX2_X1 _27588_ (
    .A(\rf[20] [19]),
    .B(_06422_),
    .S(_06388_),
    .Z(_01080_)
  );
  MUX2_X1 _27589_ (
    .A(\rf[20] [20]),
    .B(_06423_),
    .S(_06388_),
    .Z(_01081_)
  );
  MUX2_X1 _27590_ (
    .A(\rf[20] [21]),
    .B(_06424_),
    .S(_06388_),
    .Z(_01082_)
  );
  MUX2_X1 _27591_ (
    .A(\rf[20] [22]),
    .B(_06425_),
    .S(_06388_),
    .Z(_01083_)
  );
  MUX2_X1 _27592_ (
    .A(\rf[20] [23]),
    .B(_06426_),
    .S(_06388_),
    .Z(_01084_)
  );
  MUX2_X1 _27593_ (
    .A(\rf[20] [24]),
    .B(_06427_),
    .S(_06388_),
    .Z(_01085_)
  );
  MUX2_X1 _27594_ (
    .A(\rf[20] [25]),
    .B(_06428_),
    .S(_06388_),
    .Z(_01086_)
  );
  MUX2_X1 _27595_ (
    .A(\rf[20] [26]),
    .B(_06429_),
    .S(_06388_),
    .Z(_01087_)
  );
  MUX2_X1 _27596_ (
    .A(\rf[20] [27]),
    .B(_06430_),
    .S(_06388_),
    .Z(_01088_)
  );
  MUX2_X1 _27597_ (
    .A(\rf[20] [28]),
    .B(_06431_),
    .S(_06388_),
    .Z(_01089_)
  );
  MUX2_X1 _27598_ (
    .A(\rf[20] [29]),
    .B(_06432_),
    .S(_06388_),
    .Z(_01090_)
  );
  MUX2_X1 _27599_ (
    .A(\rf[20] [30]),
    .B(_06433_),
    .S(_06388_),
    .Z(_01091_)
  );
  MUX2_X1 _27600_ (
    .A(\rf[9] [0]),
    .B(_06403_),
    .S(_06353_),
    .Z(_01092_)
  );
  MUX2_X1 _27601_ (
    .A(\rf[9] [1]),
    .B(_06404_),
    .S(_06353_),
    .Z(_01093_)
  );
  MUX2_X1 _27602_ (
    .A(\rf[9] [2]),
    .B(_06405_),
    .S(_06353_),
    .Z(_01094_)
  );
  MUX2_X1 _27603_ (
    .A(\rf[9] [3]),
    .B(_06406_),
    .S(_06353_),
    .Z(_01095_)
  );
  MUX2_X1 _27604_ (
    .A(\rf[9] [4]),
    .B(_06407_),
    .S(_06353_),
    .Z(_01096_)
  );
  MUX2_X1 _27605_ (
    .A(\rf[9] [5]),
    .B(_06408_),
    .S(_06353_),
    .Z(_01097_)
  );
  MUX2_X1 _27606_ (
    .A(\rf[9] [6]),
    .B(_06409_),
    .S(_06353_),
    .Z(_01098_)
  );
  MUX2_X1 _27607_ (
    .A(\rf[9] [7]),
    .B(_06410_),
    .S(_06353_),
    .Z(_01099_)
  );
  MUX2_X1 _27608_ (
    .A(\rf[9] [8]),
    .B(_06411_),
    .S(_06353_),
    .Z(_01100_)
  );
  MUX2_X1 _27609_ (
    .A(\rf[9] [9]),
    .B(_06412_),
    .S(_06353_),
    .Z(_01101_)
  );
  MUX2_X1 _27610_ (
    .A(\rf[9] [10]),
    .B(_06413_),
    .S(_06353_),
    .Z(_01102_)
  );
  MUX2_X1 _27611_ (
    .A(\rf[9] [11]),
    .B(_06414_),
    .S(_06353_),
    .Z(_01103_)
  );
  MUX2_X1 _27612_ (
    .A(\rf[9] [12]),
    .B(_06415_),
    .S(_06353_),
    .Z(_01104_)
  );
  MUX2_X1 _27613_ (
    .A(\rf[9] [13]),
    .B(_06416_),
    .S(_06353_),
    .Z(_01105_)
  );
  MUX2_X1 _27614_ (
    .A(\rf[9] [14]),
    .B(_06417_),
    .S(_06353_),
    .Z(_01106_)
  );
  MUX2_X1 _27615_ (
    .A(\rf[9] [15]),
    .B(_06418_),
    .S(_06353_),
    .Z(_01107_)
  );
  MUX2_X1 _27616_ (
    .A(\rf[9] [16]),
    .B(_06419_),
    .S(_06353_),
    .Z(_01108_)
  );
  MUX2_X1 _27617_ (
    .A(\rf[9] [17]),
    .B(_06420_),
    .S(_06353_),
    .Z(_01109_)
  );
  MUX2_X1 _27618_ (
    .A(\rf[9] [18]),
    .B(_06421_),
    .S(_06353_),
    .Z(_01110_)
  );
  MUX2_X1 _27619_ (
    .A(\rf[9] [19]),
    .B(_06422_),
    .S(_06353_),
    .Z(_01111_)
  );
  MUX2_X1 _27620_ (
    .A(\rf[9] [20]),
    .B(_06423_),
    .S(_06353_),
    .Z(_01112_)
  );
  MUX2_X1 _27621_ (
    .A(\rf[9] [21]),
    .B(_06424_),
    .S(_06353_),
    .Z(_01113_)
  );
  MUX2_X1 _27622_ (
    .A(\rf[9] [22]),
    .B(_06425_),
    .S(_06353_),
    .Z(_01114_)
  );
  MUX2_X1 _27623_ (
    .A(\rf[9] [23]),
    .B(_06426_),
    .S(_06353_),
    .Z(_01115_)
  );
  MUX2_X1 _27624_ (
    .A(\rf[9] [24]),
    .B(_06427_),
    .S(_06353_),
    .Z(_01116_)
  );
  MUX2_X1 _27625_ (
    .A(\rf[9] [25]),
    .B(_06428_),
    .S(_06353_),
    .Z(_01117_)
  );
  MUX2_X1 _27626_ (
    .A(\rf[9] [26]),
    .B(_06429_),
    .S(_06353_),
    .Z(_01118_)
  );
  MUX2_X1 _27627_ (
    .A(\rf[9] [27]),
    .B(_06430_),
    .S(_06353_),
    .Z(_01119_)
  );
  MUX2_X1 _27628_ (
    .A(\rf[9] [28]),
    .B(_06431_),
    .S(_06353_),
    .Z(_01120_)
  );
  MUX2_X1 _27629_ (
    .A(\rf[9] [29]),
    .B(_06432_),
    .S(_06353_),
    .Z(_01121_)
  );
  MUX2_X1 _27630_ (
    .A(\rf[9] [30]),
    .B(_06433_),
    .S(_06353_),
    .Z(_01122_)
  );
  MUX2_X1 _27631_ (
    .A(\rf[21] [0]),
    .B(_06403_),
    .S(_06387_),
    .Z(_01123_)
  );
  MUX2_X1 _27632_ (
    .A(\rf[21] [1]),
    .B(_06404_),
    .S(_06387_),
    .Z(_01124_)
  );
  MUX2_X1 _27633_ (
    .A(\rf[21] [2]),
    .B(_06405_),
    .S(_06387_),
    .Z(_01125_)
  );
  MUX2_X1 _27634_ (
    .A(\rf[21] [3]),
    .B(_06406_),
    .S(_06387_),
    .Z(_01126_)
  );
  MUX2_X1 _27635_ (
    .A(\rf[21] [4]),
    .B(_06407_),
    .S(_06387_),
    .Z(_01127_)
  );
  MUX2_X1 _27636_ (
    .A(\rf[21] [5]),
    .B(_06408_),
    .S(_06387_),
    .Z(_01128_)
  );
  MUX2_X1 _27637_ (
    .A(\rf[21] [6]),
    .B(_06409_),
    .S(_06387_),
    .Z(_01129_)
  );
  MUX2_X1 _27638_ (
    .A(\rf[21] [7]),
    .B(_06410_),
    .S(_06387_),
    .Z(_01130_)
  );
  MUX2_X1 _27639_ (
    .A(\rf[21] [8]),
    .B(_06411_),
    .S(_06387_),
    .Z(_01131_)
  );
  MUX2_X1 _27640_ (
    .A(\rf[21] [9]),
    .B(_06412_),
    .S(_06387_),
    .Z(_01132_)
  );
  MUX2_X1 _27641_ (
    .A(\rf[21] [10]),
    .B(_06413_),
    .S(_06387_),
    .Z(_01133_)
  );
  MUX2_X1 _27642_ (
    .A(\rf[21] [11]),
    .B(_06414_),
    .S(_06387_),
    .Z(_01134_)
  );
  MUX2_X1 _27643_ (
    .A(\rf[21] [12]),
    .B(_06415_),
    .S(_06387_),
    .Z(_01135_)
  );
  MUX2_X1 _27644_ (
    .A(\rf[21] [13]),
    .B(_06416_),
    .S(_06387_),
    .Z(_01136_)
  );
  MUX2_X1 _27645_ (
    .A(\rf[21] [14]),
    .B(_06417_),
    .S(_06387_),
    .Z(_01137_)
  );
  MUX2_X1 _27646_ (
    .A(\rf[21] [15]),
    .B(_06418_),
    .S(_06387_),
    .Z(_01138_)
  );
  MUX2_X1 _27647_ (
    .A(\rf[21] [16]),
    .B(_06419_),
    .S(_06387_),
    .Z(_01139_)
  );
  MUX2_X1 _27648_ (
    .A(\rf[21] [17]),
    .B(_06420_),
    .S(_06387_),
    .Z(_01140_)
  );
  MUX2_X1 _27649_ (
    .A(\rf[21] [18]),
    .B(_06421_),
    .S(_06387_),
    .Z(_01141_)
  );
  MUX2_X1 _27650_ (
    .A(\rf[21] [19]),
    .B(_06422_),
    .S(_06387_),
    .Z(_01142_)
  );
  MUX2_X1 _27651_ (
    .A(\rf[21] [20]),
    .B(_06423_),
    .S(_06387_),
    .Z(_01143_)
  );
  MUX2_X1 _27652_ (
    .A(\rf[21] [21]),
    .B(_06424_),
    .S(_06387_),
    .Z(_01144_)
  );
  MUX2_X1 _27653_ (
    .A(\rf[21] [22]),
    .B(_06425_),
    .S(_06387_),
    .Z(_01145_)
  );
  MUX2_X1 _27654_ (
    .A(\rf[21] [23]),
    .B(_06426_),
    .S(_06387_),
    .Z(_01146_)
  );
  MUX2_X1 _27655_ (
    .A(\rf[21] [24]),
    .B(_06427_),
    .S(_06387_),
    .Z(_01147_)
  );
  MUX2_X1 _27656_ (
    .A(\rf[21] [25]),
    .B(_06428_),
    .S(_06387_),
    .Z(_01148_)
  );
  MUX2_X1 _27657_ (
    .A(\rf[21] [26]),
    .B(_06429_),
    .S(_06387_),
    .Z(_01149_)
  );
  MUX2_X1 _27658_ (
    .A(\rf[21] [27]),
    .B(_06430_),
    .S(_06387_),
    .Z(_01150_)
  );
  MUX2_X1 _27659_ (
    .A(\rf[21] [28]),
    .B(_06431_),
    .S(_06387_),
    .Z(_01151_)
  );
  MUX2_X1 _27660_ (
    .A(\rf[21] [29]),
    .B(_06432_),
    .S(_06387_),
    .Z(_01152_)
  );
  MUX2_X1 _27661_ (
    .A(\rf[21] [30]),
    .B(_06433_),
    .S(_06387_),
    .Z(_01153_)
  );
  MUX2_X1 _27662_ (
    .A(\rf[13] [0]),
    .B(_06403_),
    .S(_06398_),
    .Z(_01154_)
  );
  MUX2_X1 _27663_ (
    .A(\rf[13] [1]),
    .B(_06404_),
    .S(_06398_),
    .Z(_01155_)
  );
  MUX2_X1 _27664_ (
    .A(\rf[13] [2]),
    .B(_06405_),
    .S(_06398_),
    .Z(_01156_)
  );
  MUX2_X1 _27665_ (
    .A(\rf[13] [3]),
    .B(_06406_),
    .S(_06398_),
    .Z(_01157_)
  );
  MUX2_X1 _27666_ (
    .A(\rf[13] [4]),
    .B(_06407_),
    .S(_06398_),
    .Z(_01158_)
  );
  MUX2_X1 _27667_ (
    .A(\rf[13] [5]),
    .B(_06408_),
    .S(_06398_),
    .Z(_01159_)
  );
  MUX2_X1 _27668_ (
    .A(\rf[13] [6]),
    .B(_06409_),
    .S(_06398_),
    .Z(_01160_)
  );
  MUX2_X1 _27669_ (
    .A(\rf[13] [7]),
    .B(_06410_),
    .S(_06398_),
    .Z(_01161_)
  );
  MUX2_X1 _27670_ (
    .A(\rf[13] [8]),
    .B(_06411_),
    .S(_06398_),
    .Z(_01162_)
  );
  MUX2_X1 _27671_ (
    .A(\rf[13] [9]),
    .B(_06412_),
    .S(_06398_),
    .Z(_01163_)
  );
  MUX2_X1 _27672_ (
    .A(\rf[13] [10]),
    .B(_06413_),
    .S(_06398_),
    .Z(_01164_)
  );
  MUX2_X1 _27673_ (
    .A(\rf[13] [11]),
    .B(_06414_),
    .S(_06398_),
    .Z(_01165_)
  );
  MUX2_X1 _27674_ (
    .A(\rf[13] [12]),
    .B(_06415_),
    .S(_06398_),
    .Z(_01166_)
  );
  MUX2_X1 _27675_ (
    .A(\rf[13] [13]),
    .B(_06416_),
    .S(_06398_),
    .Z(_01167_)
  );
  MUX2_X1 _27676_ (
    .A(\rf[13] [14]),
    .B(_06417_),
    .S(_06398_),
    .Z(_01168_)
  );
  MUX2_X1 _27677_ (
    .A(\rf[13] [15]),
    .B(_06418_),
    .S(_06398_),
    .Z(_01169_)
  );
  MUX2_X1 _27678_ (
    .A(\rf[13] [16]),
    .B(_06419_),
    .S(_06398_),
    .Z(_01170_)
  );
  MUX2_X1 _27679_ (
    .A(\rf[13] [17]),
    .B(_06420_),
    .S(_06398_),
    .Z(_01171_)
  );
  MUX2_X1 _27680_ (
    .A(\rf[13] [18]),
    .B(_06421_),
    .S(_06398_),
    .Z(_01172_)
  );
  MUX2_X1 _27681_ (
    .A(\rf[13] [19]),
    .B(_06422_),
    .S(_06398_),
    .Z(_01173_)
  );
  MUX2_X1 _27682_ (
    .A(\rf[13] [20]),
    .B(_06423_),
    .S(_06398_),
    .Z(_01174_)
  );
  MUX2_X1 _27683_ (
    .A(\rf[13] [21]),
    .B(_06424_),
    .S(_06398_),
    .Z(_01175_)
  );
  MUX2_X1 _27684_ (
    .A(\rf[13] [22]),
    .B(_06425_),
    .S(_06398_),
    .Z(_01176_)
  );
  MUX2_X1 _27685_ (
    .A(\rf[13] [23]),
    .B(_06426_),
    .S(_06398_),
    .Z(_01177_)
  );
  MUX2_X1 _27686_ (
    .A(\rf[13] [24]),
    .B(_06427_),
    .S(_06398_),
    .Z(_01178_)
  );
  MUX2_X1 _27687_ (
    .A(\rf[13] [25]),
    .B(_06428_),
    .S(_06398_),
    .Z(_01179_)
  );
  MUX2_X1 _27688_ (
    .A(\rf[13] [26]),
    .B(_06429_),
    .S(_06398_),
    .Z(_01180_)
  );
  MUX2_X1 _27689_ (
    .A(\rf[13] [27]),
    .B(_06430_),
    .S(_06398_),
    .Z(_01181_)
  );
  MUX2_X1 _27690_ (
    .A(\rf[13] [28]),
    .B(_06431_),
    .S(_06398_),
    .Z(_01182_)
  );
  MUX2_X1 _27691_ (
    .A(\rf[13] [29]),
    .B(_06432_),
    .S(_06398_),
    .Z(_01183_)
  );
  MUX2_X1 _27692_ (
    .A(\rf[13] [30]),
    .B(_06433_),
    .S(_06398_),
    .Z(_01184_)
  );
  MUX2_X1 _27693_ (
    .A(\rf[28] [0]),
    .B(_06403_),
    .S(_06377_),
    .Z(_01185_)
  );
  MUX2_X1 _27694_ (
    .A(\rf[28] [1]),
    .B(_06404_),
    .S(_06377_),
    .Z(_01186_)
  );
  MUX2_X1 _27695_ (
    .A(\rf[28] [2]),
    .B(_06405_),
    .S(_06377_),
    .Z(_01187_)
  );
  MUX2_X1 _27696_ (
    .A(\rf[28] [3]),
    .B(_06406_),
    .S(_06377_),
    .Z(_01188_)
  );
  MUX2_X1 _27697_ (
    .A(\rf[28] [4]),
    .B(_06407_),
    .S(_06377_),
    .Z(_01189_)
  );
  MUX2_X1 _27698_ (
    .A(\rf[28] [5]),
    .B(_06408_),
    .S(_06377_),
    .Z(_01190_)
  );
  MUX2_X1 _27699_ (
    .A(\rf[28] [6]),
    .B(_06409_),
    .S(_06377_),
    .Z(_01191_)
  );
  MUX2_X1 _27700_ (
    .A(\rf[28] [7]),
    .B(_06410_),
    .S(_06377_),
    .Z(_01192_)
  );
  MUX2_X1 _27701_ (
    .A(\rf[28] [8]),
    .B(_06411_),
    .S(_06377_),
    .Z(_01193_)
  );
  MUX2_X1 _27702_ (
    .A(\rf[28] [9]),
    .B(_06412_),
    .S(_06377_),
    .Z(_01194_)
  );
  MUX2_X1 _27703_ (
    .A(\rf[28] [10]),
    .B(_06413_),
    .S(_06377_),
    .Z(_01195_)
  );
  MUX2_X1 _27704_ (
    .A(\rf[28] [11]),
    .B(_06414_),
    .S(_06377_),
    .Z(_01196_)
  );
  MUX2_X1 _27705_ (
    .A(\rf[28] [12]),
    .B(_06415_),
    .S(_06377_),
    .Z(_01197_)
  );
  MUX2_X1 _27706_ (
    .A(\rf[28] [13]),
    .B(_06416_),
    .S(_06377_),
    .Z(_01198_)
  );
  MUX2_X1 _27707_ (
    .A(\rf[28] [14]),
    .B(_06417_),
    .S(_06377_),
    .Z(_01199_)
  );
  MUX2_X1 _27708_ (
    .A(\rf[28] [15]),
    .B(_06418_),
    .S(_06377_),
    .Z(_01200_)
  );
  MUX2_X1 _27709_ (
    .A(\rf[28] [16]),
    .B(_06419_),
    .S(_06377_),
    .Z(_01201_)
  );
  MUX2_X1 _27710_ (
    .A(\rf[28] [17]),
    .B(_06420_),
    .S(_06377_),
    .Z(_01202_)
  );
  MUX2_X1 _27711_ (
    .A(\rf[28] [18]),
    .B(_06421_),
    .S(_06377_),
    .Z(_01203_)
  );
  MUX2_X1 _27712_ (
    .A(\rf[28] [19]),
    .B(_06422_),
    .S(_06377_),
    .Z(_01204_)
  );
  MUX2_X1 _27713_ (
    .A(\rf[28] [20]),
    .B(_06423_),
    .S(_06377_),
    .Z(_01205_)
  );
  MUX2_X1 _27714_ (
    .A(\rf[28] [21]),
    .B(_06424_),
    .S(_06377_),
    .Z(_01206_)
  );
  MUX2_X1 _27715_ (
    .A(\rf[28] [22]),
    .B(_06425_),
    .S(_06377_),
    .Z(_01207_)
  );
  MUX2_X1 _27716_ (
    .A(\rf[28] [23]),
    .B(_06426_),
    .S(_06377_),
    .Z(_01208_)
  );
  MUX2_X1 _27717_ (
    .A(\rf[28] [24]),
    .B(_06427_),
    .S(_06377_),
    .Z(_01209_)
  );
  MUX2_X1 _27718_ (
    .A(\rf[28] [25]),
    .B(_06428_),
    .S(_06377_),
    .Z(_01210_)
  );
  MUX2_X1 _27719_ (
    .A(\rf[28] [26]),
    .B(_06429_),
    .S(_06377_),
    .Z(_01211_)
  );
  MUX2_X1 _27720_ (
    .A(\rf[28] [27]),
    .B(_06430_),
    .S(_06377_),
    .Z(_01212_)
  );
  MUX2_X1 _27721_ (
    .A(\rf[28] [28]),
    .B(_06431_),
    .S(_06377_),
    .Z(_01213_)
  );
  MUX2_X1 _27722_ (
    .A(\rf[28] [29]),
    .B(_06432_),
    .S(_06377_),
    .Z(_01214_)
  );
  MUX2_X1 _27723_ (
    .A(\rf[28] [30]),
    .B(_06433_),
    .S(_06377_),
    .Z(_01215_)
  );
  MUX2_X1 _27724_ (
    .A(\rf[29] [0]),
    .B(_06403_),
    .S(_06375_),
    .Z(_01216_)
  );
  MUX2_X1 _27725_ (
    .A(\rf[29] [1]),
    .B(_06404_),
    .S(_06375_),
    .Z(_01217_)
  );
  MUX2_X1 _27726_ (
    .A(\rf[29] [2]),
    .B(_06405_),
    .S(_06375_),
    .Z(_01218_)
  );
  MUX2_X1 _27727_ (
    .A(\rf[29] [3]),
    .B(_06406_),
    .S(_06375_),
    .Z(_01219_)
  );
  MUX2_X1 _27728_ (
    .A(\rf[29] [4]),
    .B(_06407_),
    .S(_06375_),
    .Z(_01220_)
  );
  MUX2_X1 _27729_ (
    .A(\rf[29] [5]),
    .B(_06408_),
    .S(_06375_),
    .Z(_01221_)
  );
  MUX2_X1 _27730_ (
    .A(\rf[29] [6]),
    .B(_06409_),
    .S(_06375_),
    .Z(_01222_)
  );
  MUX2_X1 _27731_ (
    .A(\rf[29] [7]),
    .B(_06410_),
    .S(_06375_),
    .Z(_01223_)
  );
  MUX2_X1 _27732_ (
    .A(\rf[29] [8]),
    .B(_06411_),
    .S(_06375_),
    .Z(_01224_)
  );
  MUX2_X1 _27733_ (
    .A(\rf[29] [9]),
    .B(_06412_),
    .S(_06375_),
    .Z(_01225_)
  );
  MUX2_X1 _27734_ (
    .A(\rf[29] [10]),
    .B(_06413_),
    .S(_06375_),
    .Z(_01226_)
  );
  MUX2_X1 _27735_ (
    .A(\rf[29] [11]),
    .B(_06414_),
    .S(_06375_),
    .Z(_01227_)
  );
  MUX2_X1 _27736_ (
    .A(\rf[29] [12]),
    .B(_06415_),
    .S(_06375_),
    .Z(_01228_)
  );
  MUX2_X1 _27737_ (
    .A(\rf[29] [13]),
    .B(_06416_),
    .S(_06375_),
    .Z(_01229_)
  );
  MUX2_X1 _27738_ (
    .A(\rf[29] [14]),
    .B(_06417_),
    .S(_06375_),
    .Z(_01230_)
  );
  MUX2_X1 _27739_ (
    .A(\rf[29] [15]),
    .B(_06418_),
    .S(_06375_),
    .Z(_01231_)
  );
  MUX2_X1 _27740_ (
    .A(\rf[29] [16]),
    .B(_06419_),
    .S(_06375_),
    .Z(_01232_)
  );
  MUX2_X1 _27741_ (
    .A(\rf[29] [17]),
    .B(_06420_),
    .S(_06375_),
    .Z(_01233_)
  );
  MUX2_X1 _27742_ (
    .A(\rf[29] [18]),
    .B(_06421_),
    .S(_06375_),
    .Z(_01234_)
  );
  MUX2_X1 _27743_ (
    .A(\rf[29] [19]),
    .B(_06422_),
    .S(_06375_),
    .Z(_01235_)
  );
  MUX2_X1 _27744_ (
    .A(\rf[29] [20]),
    .B(_06423_),
    .S(_06375_),
    .Z(_01236_)
  );
  MUX2_X1 _27745_ (
    .A(\rf[29] [21]),
    .B(_06424_),
    .S(_06375_),
    .Z(_01237_)
  );
  MUX2_X1 _27746_ (
    .A(\rf[29] [22]),
    .B(_06425_),
    .S(_06375_),
    .Z(_01238_)
  );
  MUX2_X1 _27747_ (
    .A(\rf[29] [23]),
    .B(_06426_),
    .S(_06375_),
    .Z(_01239_)
  );
  MUX2_X1 _27748_ (
    .A(\rf[29] [24]),
    .B(_06427_),
    .S(_06375_),
    .Z(_01240_)
  );
  MUX2_X1 _27749_ (
    .A(\rf[29] [25]),
    .B(_06428_),
    .S(_06375_),
    .Z(_01241_)
  );
  MUX2_X1 _27750_ (
    .A(\rf[29] [26]),
    .B(_06429_),
    .S(_06375_),
    .Z(_01242_)
  );
  MUX2_X1 _27751_ (
    .A(\rf[29] [27]),
    .B(_06430_),
    .S(_06375_),
    .Z(_01243_)
  );
  MUX2_X1 _27752_ (
    .A(\rf[29] [28]),
    .B(_06431_),
    .S(_06375_),
    .Z(_01244_)
  );
  MUX2_X1 _27753_ (
    .A(\rf[29] [29]),
    .B(_06432_),
    .S(_06375_),
    .Z(_01245_)
  );
  MUX2_X1 _27754_ (
    .A(\rf[29] [30]),
    .B(_06433_),
    .S(_06375_),
    .Z(_01246_)
  );
  MUX2_X1 _27755_ (
    .A(\rf[30] [0]),
    .B(_06403_),
    .S(_06373_),
    .Z(_01247_)
  );
  MUX2_X1 _27756_ (
    .A(\rf[30] [1]),
    .B(_06404_),
    .S(_06373_),
    .Z(_01248_)
  );
  MUX2_X1 _27757_ (
    .A(\rf[30] [2]),
    .B(_06405_),
    .S(_06373_),
    .Z(_01249_)
  );
  MUX2_X1 _27758_ (
    .A(\rf[30] [3]),
    .B(_06406_),
    .S(_06373_),
    .Z(_01250_)
  );
  MUX2_X1 _27759_ (
    .A(\rf[30] [4]),
    .B(_06407_),
    .S(_06373_),
    .Z(_01251_)
  );
  MUX2_X1 _27760_ (
    .A(\rf[30] [5]),
    .B(_06408_),
    .S(_06373_),
    .Z(_01252_)
  );
  MUX2_X1 _27761_ (
    .A(\rf[30] [6]),
    .B(_06409_),
    .S(_06373_),
    .Z(_01253_)
  );
  MUX2_X1 _27762_ (
    .A(\rf[30] [7]),
    .B(_06410_),
    .S(_06373_),
    .Z(_01254_)
  );
  MUX2_X1 _27763_ (
    .A(\rf[30] [8]),
    .B(_06411_),
    .S(_06373_),
    .Z(_01255_)
  );
  MUX2_X1 _27764_ (
    .A(\rf[30] [9]),
    .B(_06412_),
    .S(_06373_),
    .Z(_01256_)
  );
  MUX2_X1 _27765_ (
    .A(\rf[30] [10]),
    .B(_06413_),
    .S(_06373_),
    .Z(_01257_)
  );
  MUX2_X1 _27766_ (
    .A(\rf[30] [11]),
    .B(_06414_),
    .S(_06373_),
    .Z(_01258_)
  );
  MUX2_X1 _27767_ (
    .A(\rf[30] [12]),
    .B(_06415_),
    .S(_06373_),
    .Z(_01259_)
  );
  MUX2_X1 _27768_ (
    .A(\rf[30] [13]),
    .B(_06416_),
    .S(_06373_),
    .Z(_01260_)
  );
  MUX2_X1 _27769_ (
    .A(\rf[30] [14]),
    .B(_06417_),
    .S(_06373_),
    .Z(_01261_)
  );
  MUX2_X1 _27770_ (
    .A(\rf[30] [15]),
    .B(_06418_),
    .S(_06373_),
    .Z(_01262_)
  );
  MUX2_X1 _27771_ (
    .A(\rf[30] [16]),
    .B(_06419_),
    .S(_06373_),
    .Z(_01263_)
  );
  MUX2_X1 _27772_ (
    .A(\rf[30] [17]),
    .B(_06420_),
    .S(_06373_),
    .Z(_01264_)
  );
  MUX2_X1 _27773_ (
    .A(\rf[30] [18]),
    .B(_06421_),
    .S(_06373_),
    .Z(_01265_)
  );
  MUX2_X1 _27774_ (
    .A(\rf[30] [19]),
    .B(_06422_),
    .S(_06373_),
    .Z(_01266_)
  );
  MUX2_X1 _27775_ (
    .A(\rf[30] [20]),
    .B(_06423_),
    .S(_06373_),
    .Z(_01267_)
  );
  MUX2_X1 _27776_ (
    .A(\rf[30] [21]),
    .B(_06424_),
    .S(_06373_),
    .Z(_01268_)
  );
  MUX2_X1 _27777_ (
    .A(\rf[30] [22]),
    .B(_06425_),
    .S(_06373_),
    .Z(_01269_)
  );
  MUX2_X1 _27778_ (
    .A(\rf[30] [23]),
    .B(_06426_),
    .S(_06373_),
    .Z(_01270_)
  );
  MUX2_X1 _27779_ (
    .A(\rf[30] [24]),
    .B(_06427_),
    .S(_06373_),
    .Z(_01271_)
  );
  MUX2_X1 _27780_ (
    .A(\rf[30] [25]),
    .B(_06428_),
    .S(_06373_),
    .Z(_01272_)
  );
  MUX2_X1 _27781_ (
    .A(\rf[30] [26]),
    .B(_06429_),
    .S(_06373_),
    .Z(_01273_)
  );
  MUX2_X1 _27782_ (
    .A(\rf[30] [27]),
    .B(_06430_),
    .S(_06373_),
    .Z(_01274_)
  );
  MUX2_X1 _27783_ (
    .A(\rf[30] [28]),
    .B(_06431_),
    .S(_06373_),
    .Z(_01275_)
  );
  MUX2_X1 _27784_ (
    .A(\rf[30] [29]),
    .B(_06432_),
    .S(_06373_),
    .Z(_01276_)
  );
  MUX2_X1 _27785_ (
    .A(\rf[30] [30]),
    .B(_06433_),
    .S(_06373_),
    .Z(_01277_)
  );
  MUX2_X1 _27786_ (
    .A(\rf[14] [0]),
    .B(_06403_),
    .S(_06397_),
    .Z(_01278_)
  );
  MUX2_X1 _27787_ (
    .A(\rf[14] [1]),
    .B(_06404_),
    .S(_06397_),
    .Z(_01279_)
  );
  MUX2_X1 _27788_ (
    .A(\rf[14] [2]),
    .B(_06405_),
    .S(_06397_),
    .Z(_01280_)
  );
  MUX2_X1 _27789_ (
    .A(\rf[14] [3]),
    .B(_06406_),
    .S(_06397_),
    .Z(_01281_)
  );
  MUX2_X1 _27790_ (
    .A(\rf[14] [4]),
    .B(_06407_),
    .S(_06397_),
    .Z(_01282_)
  );
  MUX2_X1 _27791_ (
    .A(\rf[14] [5]),
    .B(_06408_),
    .S(_06397_),
    .Z(_01283_)
  );
  MUX2_X1 _27792_ (
    .A(\rf[14] [6]),
    .B(_06409_),
    .S(_06397_),
    .Z(_01284_)
  );
  MUX2_X1 _27793_ (
    .A(\rf[14] [7]),
    .B(_06410_),
    .S(_06397_),
    .Z(_01285_)
  );
  MUX2_X1 _27794_ (
    .A(\rf[14] [8]),
    .B(_06411_),
    .S(_06397_),
    .Z(_01286_)
  );
  MUX2_X1 _27795_ (
    .A(\rf[14] [9]),
    .B(_06412_),
    .S(_06397_),
    .Z(_01287_)
  );
  MUX2_X1 _27796_ (
    .A(\rf[14] [10]),
    .B(_06413_),
    .S(_06397_),
    .Z(_01288_)
  );
  MUX2_X1 _27797_ (
    .A(\rf[14] [11]),
    .B(_06414_),
    .S(_06397_),
    .Z(_01289_)
  );
  MUX2_X1 _27798_ (
    .A(\rf[14] [12]),
    .B(_06415_),
    .S(_06397_),
    .Z(_01290_)
  );
  MUX2_X1 _27799_ (
    .A(\rf[14] [13]),
    .B(_06416_),
    .S(_06397_),
    .Z(_01291_)
  );
  MUX2_X1 _27800_ (
    .A(\rf[14] [14]),
    .B(_06417_),
    .S(_06397_),
    .Z(_01292_)
  );
  MUX2_X1 _27801_ (
    .A(\rf[14] [15]),
    .B(_06418_),
    .S(_06397_),
    .Z(_01293_)
  );
  MUX2_X1 _27802_ (
    .A(\rf[14] [16]),
    .B(_06419_),
    .S(_06397_),
    .Z(_01294_)
  );
  MUX2_X1 _27803_ (
    .A(\rf[14] [17]),
    .B(_06420_),
    .S(_06397_),
    .Z(_01295_)
  );
  MUX2_X1 _27804_ (
    .A(\rf[14] [18]),
    .B(_06421_),
    .S(_06397_),
    .Z(_01296_)
  );
  MUX2_X1 _27805_ (
    .A(\rf[14] [19]),
    .B(_06422_),
    .S(_06397_),
    .Z(_01297_)
  );
  MUX2_X1 _27806_ (
    .A(\rf[14] [20]),
    .B(_06423_),
    .S(_06397_),
    .Z(_01298_)
  );
  MUX2_X1 _27807_ (
    .A(\rf[14] [21]),
    .B(_06424_),
    .S(_06397_),
    .Z(_01299_)
  );
  MUX2_X1 _27808_ (
    .A(\rf[14] [22]),
    .B(_06425_),
    .S(_06397_),
    .Z(_01300_)
  );
  MUX2_X1 _27809_ (
    .A(\rf[14] [23]),
    .B(_06426_),
    .S(_06397_),
    .Z(_01301_)
  );
  MUX2_X1 _27810_ (
    .A(\rf[14] [24]),
    .B(_06427_),
    .S(_06397_),
    .Z(_01302_)
  );
  MUX2_X1 _27811_ (
    .A(\rf[14] [25]),
    .B(_06428_),
    .S(_06397_),
    .Z(_01303_)
  );
  MUX2_X1 _27812_ (
    .A(\rf[14] [26]),
    .B(_06429_),
    .S(_06397_),
    .Z(_01304_)
  );
  MUX2_X1 _27813_ (
    .A(\rf[14] [27]),
    .B(_06430_),
    .S(_06397_),
    .Z(_01305_)
  );
  MUX2_X1 _27814_ (
    .A(\rf[14] [28]),
    .B(_06431_),
    .S(_06397_),
    .Z(_01306_)
  );
  MUX2_X1 _27815_ (
    .A(\rf[14] [29]),
    .B(_06432_),
    .S(_06397_),
    .Z(_01307_)
  );
  MUX2_X1 _27816_ (
    .A(\rf[14] [30]),
    .B(_06433_),
    .S(_06397_),
    .Z(_01308_)
  );
  MUX2_X1 _27817_ (
    .A(\rf[22] [0]),
    .B(_06403_),
    .S(_06386_),
    .Z(_01309_)
  );
  MUX2_X1 _27818_ (
    .A(\rf[22] [1]),
    .B(_06404_),
    .S(_06386_),
    .Z(_01310_)
  );
  MUX2_X1 _27819_ (
    .A(\rf[22] [2]),
    .B(_06405_),
    .S(_06386_),
    .Z(_01311_)
  );
  MUX2_X1 _27820_ (
    .A(\rf[22] [3]),
    .B(_06406_),
    .S(_06386_),
    .Z(_01312_)
  );
  MUX2_X1 _27821_ (
    .A(\rf[22] [4]),
    .B(_06407_),
    .S(_06386_),
    .Z(_01313_)
  );
  MUX2_X1 _27822_ (
    .A(\rf[22] [5]),
    .B(_06408_),
    .S(_06386_),
    .Z(_01314_)
  );
  MUX2_X1 _27823_ (
    .A(\rf[22] [6]),
    .B(_06409_),
    .S(_06386_),
    .Z(_01315_)
  );
  MUX2_X1 _27824_ (
    .A(\rf[22] [7]),
    .B(_06410_),
    .S(_06386_),
    .Z(_01316_)
  );
  MUX2_X1 _27825_ (
    .A(\rf[22] [8]),
    .B(_06411_),
    .S(_06386_),
    .Z(_01317_)
  );
  MUX2_X1 _27826_ (
    .A(\rf[22] [9]),
    .B(_06412_),
    .S(_06386_),
    .Z(_01318_)
  );
  MUX2_X1 _27827_ (
    .A(\rf[22] [10]),
    .B(_06413_),
    .S(_06386_),
    .Z(_01319_)
  );
  MUX2_X1 _27828_ (
    .A(\rf[22] [11]),
    .B(_06414_),
    .S(_06386_),
    .Z(_01320_)
  );
  MUX2_X1 _27829_ (
    .A(\rf[22] [12]),
    .B(_06415_),
    .S(_06386_),
    .Z(_01321_)
  );
  MUX2_X1 _27830_ (
    .A(\rf[22] [13]),
    .B(_06416_),
    .S(_06386_),
    .Z(_01322_)
  );
  MUX2_X1 _27831_ (
    .A(\rf[22] [14]),
    .B(_06417_),
    .S(_06386_),
    .Z(_01323_)
  );
  MUX2_X1 _27832_ (
    .A(\rf[22] [15]),
    .B(_06418_),
    .S(_06386_),
    .Z(_01324_)
  );
  MUX2_X1 _27833_ (
    .A(\rf[22] [16]),
    .B(_06419_),
    .S(_06386_),
    .Z(_01325_)
  );
  MUX2_X1 _27834_ (
    .A(\rf[22] [17]),
    .B(_06420_),
    .S(_06386_),
    .Z(_01326_)
  );
  MUX2_X1 _27835_ (
    .A(\rf[22] [18]),
    .B(_06421_),
    .S(_06386_),
    .Z(_01327_)
  );
  MUX2_X1 _27836_ (
    .A(\rf[22] [19]),
    .B(_06422_),
    .S(_06386_),
    .Z(_01328_)
  );
  MUX2_X1 _27837_ (
    .A(\rf[22] [20]),
    .B(_06423_),
    .S(_06386_),
    .Z(_01329_)
  );
  MUX2_X1 _27838_ (
    .A(\rf[22] [21]),
    .B(_06424_),
    .S(_06386_),
    .Z(_01330_)
  );
  MUX2_X1 _27839_ (
    .A(\rf[22] [22]),
    .B(_06425_),
    .S(_06386_),
    .Z(_01331_)
  );
  MUX2_X1 _27840_ (
    .A(\rf[22] [23]),
    .B(_06426_),
    .S(_06386_),
    .Z(_01332_)
  );
  MUX2_X1 _27841_ (
    .A(\rf[22] [24]),
    .B(_06427_),
    .S(_06386_),
    .Z(_01333_)
  );
  MUX2_X1 _27842_ (
    .A(\rf[22] [25]),
    .B(_06428_),
    .S(_06386_),
    .Z(_01334_)
  );
  MUX2_X1 _27843_ (
    .A(\rf[22] [26]),
    .B(_06429_),
    .S(_06386_),
    .Z(_01335_)
  );
  MUX2_X1 _27844_ (
    .A(\rf[22] [27]),
    .B(_06430_),
    .S(_06386_),
    .Z(_01336_)
  );
  MUX2_X1 _27845_ (
    .A(\rf[22] [28]),
    .B(_06431_),
    .S(_06386_),
    .Z(_01337_)
  );
  MUX2_X1 _27846_ (
    .A(\rf[22] [29]),
    .B(_06432_),
    .S(_06386_),
    .Z(_01338_)
  );
  MUX2_X1 _27847_ (
    .A(\rf[22] [30]),
    .B(_06433_),
    .S(_06386_),
    .Z(_01339_)
  );
  MUX2_X1 _27848_ (
    .A(\rf[26] [0]),
    .B(_06403_),
    .S(_06380_),
    .Z(_01340_)
  );
  MUX2_X1 _27849_ (
    .A(\rf[26] [1]),
    .B(_06404_),
    .S(_06380_),
    .Z(_01341_)
  );
  MUX2_X1 _27850_ (
    .A(\rf[26] [2]),
    .B(_06405_),
    .S(_06380_),
    .Z(_01342_)
  );
  MUX2_X1 _27851_ (
    .A(\rf[26] [3]),
    .B(_06406_),
    .S(_06380_),
    .Z(_01343_)
  );
  MUX2_X1 _27852_ (
    .A(\rf[26] [4]),
    .B(_06407_),
    .S(_06380_),
    .Z(_01344_)
  );
  MUX2_X1 _27853_ (
    .A(\rf[26] [5]),
    .B(_06408_),
    .S(_06380_),
    .Z(_01345_)
  );
  MUX2_X1 _27854_ (
    .A(\rf[26] [6]),
    .B(_06409_),
    .S(_06380_),
    .Z(_01346_)
  );
  MUX2_X1 _27855_ (
    .A(\rf[26] [7]),
    .B(_06410_),
    .S(_06380_),
    .Z(_01347_)
  );
  MUX2_X1 _27856_ (
    .A(\rf[26] [8]),
    .B(_06411_),
    .S(_06380_),
    .Z(_01348_)
  );
  MUX2_X1 _27857_ (
    .A(\rf[26] [9]),
    .B(_06412_),
    .S(_06380_),
    .Z(_01349_)
  );
  MUX2_X1 _27858_ (
    .A(\rf[26] [10]),
    .B(_06413_),
    .S(_06380_),
    .Z(_01350_)
  );
  MUX2_X1 _27859_ (
    .A(\rf[26] [11]),
    .B(_06414_),
    .S(_06380_),
    .Z(_01351_)
  );
  MUX2_X1 _27860_ (
    .A(\rf[26] [12]),
    .B(_06415_),
    .S(_06380_),
    .Z(_01352_)
  );
  MUX2_X1 _27861_ (
    .A(\rf[26] [13]),
    .B(_06416_),
    .S(_06380_),
    .Z(_01353_)
  );
  MUX2_X1 _27862_ (
    .A(\rf[26] [14]),
    .B(_06417_),
    .S(_06380_),
    .Z(_01354_)
  );
  MUX2_X1 _27863_ (
    .A(\rf[26] [15]),
    .B(_06418_),
    .S(_06380_),
    .Z(_01355_)
  );
  MUX2_X1 _27864_ (
    .A(\rf[26] [16]),
    .B(_06419_),
    .S(_06380_),
    .Z(_01356_)
  );
  MUX2_X1 _27865_ (
    .A(\rf[26] [17]),
    .B(_06420_),
    .S(_06380_),
    .Z(_01357_)
  );
  MUX2_X1 _27866_ (
    .A(\rf[26] [18]),
    .B(_06421_),
    .S(_06380_),
    .Z(_01358_)
  );
  MUX2_X1 _27867_ (
    .A(\rf[26] [19]),
    .B(_06422_),
    .S(_06380_),
    .Z(_01359_)
  );
  MUX2_X1 _27868_ (
    .A(\rf[26] [20]),
    .B(_06423_),
    .S(_06380_),
    .Z(_01360_)
  );
  MUX2_X1 _27869_ (
    .A(\rf[26] [21]),
    .B(_06424_),
    .S(_06380_),
    .Z(_01361_)
  );
  MUX2_X1 _27870_ (
    .A(\rf[26] [22]),
    .B(_06425_),
    .S(_06380_),
    .Z(_01362_)
  );
  MUX2_X1 _27871_ (
    .A(\rf[26] [23]),
    .B(_06426_),
    .S(_06380_),
    .Z(_01363_)
  );
  MUX2_X1 _27872_ (
    .A(\rf[26] [24]),
    .B(_06427_),
    .S(_06380_),
    .Z(_01364_)
  );
  MUX2_X1 _27873_ (
    .A(\rf[26] [25]),
    .B(_06428_),
    .S(_06380_),
    .Z(_01365_)
  );
  MUX2_X1 _27874_ (
    .A(\rf[26] [26]),
    .B(_06429_),
    .S(_06380_),
    .Z(_01366_)
  );
  MUX2_X1 _27875_ (
    .A(\rf[26] [27]),
    .B(_06430_),
    .S(_06380_),
    .Z(_01367_)
  );
  MUX2_X1 _27876_ (
    .A(\rf[26] [28]),
    .B(_06431_),
    .S(_06380_),
    .Z(_01368_)
  );
  MUX2_X1 _27877_ (
    .A(\rf[26] [29]),
    .B(_06432_),
    .S(_06380_),
    .Z(_01369_)
  );
  MUX2_X1 _27878_ (
    .A(\rf[26] [30]),
    .B(_06433_),
    .S(_06380_),
    .Z(_01370_)
  );
  MUX2_X1 _27879_ (
    .A(\rf[2] [0]),
    .B(_06403_),
    .S(_06374_),
    .Z(_01371_)
  );
  MUX2_X1 _27880_ (
    .A(\rf[2] [1]),
    .B(_06404_),
    .S(_06374_),
    .Z(_01372_)
  );
  MUX2_X1 _27881_ (
    .A(\rf[2] [2]),
    .B(_06405_),
    .S(_06374_),
    .Z(_01373_)
  );
  MUX2_X1 _27882_ (
    .A(\rf[2] [3]),
    .B(_06406_),
    .S(_06374_),
    .Z(_01374_)
  );
  MUX2_X1 _27883_ (
    .A(\rf[2] [4]),
    .B(_06407_),
    .S(_06374_),
    .Z(_01375_)
  );
  MUX2_X1 _27884_ (
    .A(\rf[2] [5]),
    .B(_06408_),
    .S(_06374_),
    .Z(_01376_)
  );
  MUX2_X1 _27885_ (
    .A(\rf[2] [6]),
    .B(_06409_),
    .S(_06374_),
    .Z(_01377_)
  );
  MUX2_X1 _27886_ (
    .A(\rf[2] [7]),
    .B(_06410_),
    .S(_06374_),
    .Z(_01378_)
  );
  MUX2_X1 _27887_ (
    .A(\rf[2] [8]),
    .B(_06411_),
    .S(_06374_),
    .Z(_01379_)
  );
  MUX2_X1 _27888_ (
    .A(\rf[2] [9]),
    .B(_06412_),
    .S(_06374_),
    .Z(_01380_)
  );
  MUX2_X1 _27889_ (
    .A(\rf[2] [10]),
    .B(_06413_),
    .S(_06374_),
    .Z(_01381_)
  );
  MUX2_X1 _27890_ (
    .A(\rf[2] [11]),
    .B(_06414_),
    .S(_06374_),
    .Z(_01382_)
  );
  MUX2_X1 _27891_ (
    .A(\rf[2] [12]),
    .B(_06415_),
    .S(_06374_),
    .Z(_01383_)
  );
  MUX2_X1 _27892_ (
    .A(\rf[2] [13]),
    .B(_06416_),
    .S(_06374_),
    .Z(_01384_)
  );
  MUX2_X1 _27893_ (
    .A(\rf[2] [14]),
    .B(_06417_),
    .S(_06374_),
    .Z(_01385_)
  );
  MUX2_X1 _27894_ (
    .A(\rf[2] [15]),
    .B(_06418_),
    .S(_06374_),
    .Z(_01386_)
  );
  MUX2_X1 _27895_ (
    .A(\rf[2] [16]),
    .B(_06419_),
    .S(_06374_),
    .Z(_01387_)
  );
  MUX2_X1 _27896_ (
    .A(\rf[2] [17]),
    .B(_06420_),
    .S(_06374_),
    .Z(_01388_)
  );
  MUX2_X1 _27897_ (
    .A(\rf[2] [18]),
    .B(_06421_),
    .S(_06374_),
    .Z(_01389_)
  );
  MUX2_X1 _27898_ (
    .A(\rf[2] [19]),
    .B(_06422_),
    .S(_06374_),
    .Z(_01390_)
  );
  MUX2_X1 _27899_ (
    .A(\rf[2] [20]),
    .B(_06423_),
    .S(_06374_),
    .Z(_01391_)
  );
  MUX2_X1 _27900_ (
    .A(\rf[2] [21]),
    .B(_06424_),
    .S(_06374_),
    .Z(_01392_)
  );
  MUX2_X1 _27901_ (
    .A(\rf[2] [22]),
    .B(_06425_),
    .S(_06374_),
    .Z(_01393_)
  );
  MUX2_X1 _27902_ (
    .A(\rf[2] [23]),
    .B(_06426_),
    .S(_06374_),
    .Z(_01394_)
  );
  MUX2_X1 _27903_ (
    .A(\rf[2] [24]),
    .B(_06427_),
    .S(_06374_),
    .Z(_01395_)
  );
  MUX2_X1 _27904_ (
    .A(\rf[2] [25]),
    .B(_06428_),
    .S(_06374_),
    .Z(_01396_)
  );
  MUX2_X1 _27905_ (
    .A(\rf[2] [26]),
    .B(_06429_),
    .S(_06374_),
    .Z(_01397_)
  );
  MUX2_X1 _27906_ (
    .A(\rf[2] [27]),
    .B(_06430_),
    .S(_06374_),
    .Z(_01398_)
  );
  MUX2_X1 _27907_ (
    .A(\rf[2] [28]),
    .B(_06431_),
    .S(_06374_),
    .Z(_01399_)
  );
  MUX2_X1 _27908_ (
    .A(\rf[2] [29]),
    .B(_06432_),
    .S(_06374_),
    .Z(_01400_)
  );
  MUX2_X1 _27909_ (
    .A(\rf[2] [30]),
    .B(_06433_),
    .S(_06374_),
    .Z(_01401_)
  );
  MUX2_X1 _27910_ (
    .A(\rf[27] [0]),
    .B(_06403_),
    .S(_06379_),
    .Z(_01402_)
  );
  MUX2_X1 _27911_ (
    .A(\rf[27] [1]),
    .B(_06404_),
    .S(_06379_),
    .Z(_01403_)
  );
  MUX2_X1 _27912_ (
    .A(\rf[27] [2]),
    .B(_06405_),
    .S(_06379_),
    .Z(_01404_)
  );
  MUX2_X1 _27913_ (
    .A(\rf[27] [3]),
    .B(_06406_),
    .S(_06379_),
    .Z(_01405_)
  );
  MUX2_X1 _27914_ (
    .A(\rf[27] [4]),
    .B(_06407_),
    .S(_06379_),
    .Z(_01406_)
  );
  MUX2_X1 _27915_ (
    .A(\rf[27] [5]),
    .B(_06408_),
    .S(_06379_),
    .Z(_01407_)
  );
  MUX2_X1 _27916_ (
    .A(\rf[27] [6]),
    .B(_06409_),
    .S(_06379_),
    .Z(_01408_)
  );
  MUX2_X1 _27917_ (
    .A(\rf[27] [7]),
    .B(_06410_),
    .S(_06379_),
    .Z(_01409_)
  );
  MUX2_X1 _27918_ (
    .A(\rf[27] [8]),
    .B(_06411_),
    .S(_06379_),
    .Z(_01410_)
  );
  MUX2_X1 _27919_ (
    .A(\rf[27] [9]),
    .B(_06412_),
    .S(_06379_),
    .Z(_01411_)
  );
  MUX2_X1 _27920_ (
    .A(\rf[27] [10]),
    .B(_06413_),
    .S(_06379_),
    .Z(_01412_)
  );
  MUX2_X1 _27921_ (
    .A(\rf[27] [11]),
    .B(_06414_),
    .S(_06379_),
    .Z(_01413_)
  );
  MUX2_X1 _27922_ (
    .A(\rf[27] [12]),
    .B(_06415_),
    .S(_06379_),
    .Z(_01414_)
  );
  MUX2_X1 _27923_ (
    .A(\rf[27] [13]),
    .B(_06416_),
    .S(_06379_),
    .Z(_01415_)
  );
  MUX2_X1 _27924_ (
    .A(\rf[27] [14]),
    .B(_06417_),
    .S(_06379_),
    .Z(_01416_)
  );
  MUX2_X1 _27925_ (
    .A(\rf[27] [15]),
    .B(_06418_),
    .S(_06379_),
    .Z(_01417_)
  );
  MUX2_X1 _27926_ (
    .A(\rf[27] [16]),
    .B(_06419_),
    .S(_06379_),
    .Z(_01418_)
  );
  MUX2_X1 _27927_ (
    .A(\rf[27] [17]),
    .B(_06420_),
    .S(_06379_),
    .Z(_01419_)
  );
  MUX2_X1 _27928_ (
    .A(\rf[27] [18]),
    .B(_06421_),
    .S(_06379_),
    .Z(_01420_)
  );
  MUX2_X1 _27929_ (
    .A(\rf[27] [19]),
    .B(_06422_),
    .S(_06379_),
    .Z(_01421_)
  );
  MUX2_X1 _27930_ (
    .A(\rf[27] [20]),
    .B(_06423_),
    .S(_06379_),
    .Z(_01422_)
  );
  MUX2_X1 _27931_ (
    .A(\rf[27] [21]),
    .B(_06424_),
    .S(_06379_),
    .Z(_01423_)
  );
  MUX2_X1 _27932_ (
    .A(\rf[27] [22]),
    .B(_06425_),
    .S(_06379_),
    .Z(_01424_)
  );
  MUX2_X1 _27933_ (
    .A(\rf[27] [23]),
    .B(_06426_),
    .S(_06379_),
    .Z(_01425_)
  );
  MUX2_X1 _27934_ (
    .A(\rf[27] [24]),
    .B(_06427_),
    .S(_06379_),
    .Z(_01426_)
  );
  MUX2_X1 _27935_ (
    .A(\rf[27] [25]),
    .B(_06428_),
    .S(_06379_),
    .Z(_01427_)
  );
  MUX2_X1 _27936_ (
    .A(\rf[27] [26]),
    .B(_06429_),
    .S(_06379_),
    .Z(_01428_)
  );
  MUX2_X1 _27937_ (
    .A(\rf[27] [27]),
    .B(_06430_),
    .S(_06379_),
    .Z(_01429_)
  );
  MUX2_X1 _27938_ (
    .A(\rf[27] [28]),
    .B(_06431_),
    .S(_06379_),
    .Z(_01430_)
  );
  MUX2_X1 _27939_ (
    .A(\rf[27] [29]),
    .B(_06432_),
    .S(_06379_),
    .Z(_01431_)
  );
  MUX2_X1 _27940_ (
    .A(\rf[27] [30]),
    .B(_06433_),
    .S(_06379_),
    .Z(_01432_)
  );
  MUX2_X1 _27941_ (
    .A(\rf[24] [0]),
    .B(_13580_),
    .S(_06382_),
    .Z(_01433_)
  );
  MUX2_X1 _27942_ (
    .A(\rf[24] [1]),
    .B(_13820_),
    .S(_06382_),
    .Z(_01434_)
  );
  MUX2_X1 _27943_ (
    .A(\rf[24] [2]),
    .B(_10137_),
    .S(_06382_),
    .Z(_01435_)
  );
  MUX2_X1 _27944_ (
    .A(\rf[24] [3]),
    .B(_10250_),
    .S(_06382_),
    .Z(_01436_)
  );
  MUX2_X1 _27945_ (
    .A(\rf[24] [4]),
    .B(_10389_),
    .S(_06382_),
    .Z(_01437_)
  );
  MUX2_X1 _27946_ (
    .A(\rf[24] [5]),
    .B(_10505_),
    .S(_06382_),
    .Z(_01438_)
  );
  MUX2_X1 _27947_ (
    .A(\rf[24] [6]),
    .B(_10620_),
    .S(_06382_),
    .Z(_01439_)
  );
  MUX2_X1 _27948_ (
    .A(\rf[24] [7]),
    .B(_10733_),
    .S(_06382_),
    .Z(_01440_)
  );
  MUX2_X1 _27949_ (
    .A(\rf[24] [8]),
    .B(_10846_),
    .S(_06382_),
    .Z(_01441_)
  );
  MUX2_X1 _27950_ (
    .A(\rf[24] [9]),
    .B(_10956_),
    .S(_06382_),
    .Z(_01442_)
  );
  MUX2_X1 _27951_ (
    .A(\rf[24] [10]),
    .B(_11066_),
    .S(_06382_),
    .Z(_01443_)
  );
  MUX2_X1 _27952_ (
    .A(\rf[24] [11]),
    .B(_11205_),
    .S(_06382_),
    .Z(_01444_)
  );
  MUX2_X1 _27953_ (
    .A(\rf[24] [12]),
    .B(_11315_),
    .S(_06382_),
    .Z(_01445_)
  );
  MUX2_X1 _27954_ (
    .A(\rf[24] [13]),
    .B(_11428_),
    .S(_06382_),
    .Z(_01446_)
  );
  MUX2_X1 _27955_ (
    .A(\rf[24] [14]),
    .B(_11541_),
    .S(_06382_),
    .Z(_01447_)
  );
  MUX2_X1 _27956_ (
    .A(\rf[24] [15]),
    .B(_11656_),
    .S(_06382_),
    .Z(_01448_)
  );
  MUX2_X1 _27957_ (
    .A(\rf[24] [16]),
    .B(_11766_),
    .S(_06382_),
    .Z(_01449_)
  );
  MUX2_X1 _27958_ (
    .A(\rf[24] [17]),
    .B(_11882_),
    .S(_06382_),
    .Z(_01450_)
  );
  MUX2_X1 _27959_ (
    .A(\rf[24] [18]),
    .B(_12088_),
    .S(_06382_),
    .Z(_01451_)
  );
  MUX2_X1 _27960_ (
    .A(\rf[24] [19]),
    .B(_12099_),
    .S(_06382_),
    .Z(_01452_)
  );
  MUX2_X1 _27961_ (
    .A(\rf[24] [20]),
    .B(_12305_),
    .S(_06382_),
    .Z(_01453_)
  );
  MUX2_X1 _27962_ (
    .A(\rf[24] [21]),
    .B(_12316_),
    .S(_06382_),
    .Z(_01454_)
  );
  MUX2_X1 _27963_ (
    .A(\rf[24] [22]),
    .B(_12537_),
    .S(_06382_),
    .Z(_01455_)
  );
  MUX2_X1 _27964_ (
    .A(\rf[24] [23]),
    .B(_12638_),
    .S(_06382_),
    .Z(_01456_)
  );
  MUX2_X1 _27965_ (
    .A(\rf[24] [24]),
    .B(_12649_),
    .S(_06382_),
    .Z(_01457_)
  );
  MUX2_X1 _27966_ (
    .A(\rf[24] [25]),
    .B(_12765_),
    .S(_06382_),
    .Z(_01458_)
  );
  MUX2_X1 _27967_ (
    .A(\rf[24] [26]),
    .B(_12986_),
    .S(_06382_),
    .Z(_01459_)
  );
  MUX2_X1 _27968_ (
    .A(\rf[24] [27]),
    .B(_13102_),
    .S(_06382_),
    .Z(_01460_)
  );
  MUX2_X1 _27969_ (
    .A(\rf[24] [28]),
    .B(_13218_),
    .S(_06382_),
    .Z(_01461_)
  );
  MUX2_X1 _27970_ (
    .A(\rf[24] [29]),
    .B(_13338_),
    .S(_06382_),
    .Z(_01462_)
  );
  MUX2_X1 _27971_ (
    .A(\rf[24] [30]),
    .B(_13349_),
    .S(_06382_),
    .Z(_01463_)
  );
  MUX2_X1 _27972_ (
    .A(\rf[5] [0]),
    .B(_06403_),
    .S(_06369_),
    .Z(_01464_)
  );
  MUX2_X1 _27973_ (
    .A(\rf[5] [1]),
    .B(_06404_),
    .S(_06369_),
    .Z(_01465_)
  );
  MUX2_X1 _27974_ (
    .A(\rf[5] [2]),
    .B(_06405_),
    .S(_06369_),
    .Z(_01466_)
  );
  MUX2_X1 _27975_ (
    .A(\rf[5] [3]),
    .B(_06406_),
    .S(_06369_),
    .Z(_01467_)
  );
  MUX2_X1 _27976_ (
    .A(\rf[5] [4]),
    .B(_06407_),
    .S(_06369_),
    .Z(_01468_)
  );
  MUX2_X1 _27977_ (
    .A(\rf[5] [5]),
    .B(_06408_),
    .S(_06369_),
    .Z(_01469_)
  );
  MUX2_X1 _27978_ (
    .A(\rf[5] [6]),
    .B(_06409_),
    .S(_06369_),
    .Z(_01470_)
  );
  MUX2_X1 _27979_ (
    .A(\rf[5] [7]),
    .B(_06410_),
    .S(_06369_),
    .Z(_01471_)
  );
  MUX2_X1 _27980_ (
    .A(\rf[5] [8]),
    .B(_06411_),
    .S(_06369_),
    .Z(_01472_)
  );
  MUX2_X1 _27981_ (
    .A(\rf[5] [9]),
    .B(_06412_),
    .S(_06369_),
    .Z(_01473_)
  );
  MUX2_X1 _27982_ (
    .A(\rf[5] [10]),
    .B(_06413_),
    .S(_06369_),
    .Z(_01474_)
  );
  MUX2_X1 _27983_ (
    .A(\rf[5] [11]),
    .B(_06414_),
    .S(_06369_),
    .Z(_01475_)
  );
  MUX2_X1 _27984_ (
    .A(\rf[5] [12]),
    .B(_06415_),
    .S(_06369_),
    .Z(_01476_)
  );
  MUX2_X1 _27985_ (
    .A(\rf[5] [13]),
    .B(_06416_),
    .S(_06369_),
    .Z(_01477_)
  );
  MUX2_X1 _27986_ (
    .A(\rf[5] [14]),
    .B(_06417_),
    .S(_06369_),
    .Z(_01478_)
  );
  MUX2_X1 _27987_ (
    .A(\rf[5] [15]),
    .B(_06418_),
    .S(_06369_),
    .Z(_01479_)
  );
  MUX2_X1 _27988_ (
    .A(\rf[5] [16]),
    .B(_06419_),
    .S(_06369_),
    .Z(_01480_)
  );
  MUX2_X1 _27989_ (
    .A(\rf[5] [17]),
    .B(_06420_),
    .S(_06369_),
    .Z(_01481_)
  );
  MUX2_X1 _27990_ (
    .A(\rf[5] [18]),
    .B(_06421_),
    .S(_06369_),
    .Z(_01482_)
  );
  MUX2_X1 _27991_ (
    .A(\rf[5] [19]),
    .B(_06422_),
    .S(_06369_),
    .Z(_01483_)
  );
  MUX2_X1 _27992_ (
    .A(\rf[5] [20]),
    .B(_06423_),
    .S(_06369_),
    .Z(_01484_)
  );
  MUX2_X1 _27993_ (
    .A(\rf[5] [21]),
    .B(_06424_),
    .S(_06369_),
    .Z(_01485_)
  );
  MUX2_X1 _27994_ (
    .A(\rf[5] [22]),
    .B(_06425_),
    .S(_06369_),
    .Z(_01486_)
  );
  MUX2_X1 _27995_ (
    .A(\rf[5] [23]),
    .B(_06426_),
    .S(_06369_),
    .Z(_01487_)
  );
  MUX2_X1 _27996_ (
    .A(\rf[5] [24]),
    .B(_06427_),
    .S(_06369_),
    .Z(_01488_)
  );
  MUX2_X1 _27997_ (
    .A(\rf[5] [25]),
    .B(_06428_),
    .S(_06369_),
    .Z(_01489_)
  );
  MUX2_X1 _27998_ (
    .A(\rf[5] [26]),
    .B(_06429_),
    .S(_06369_),
    .Z(_01490_)
  );
  MUX2_X1 _27999_ (
    .A(\rf[5] [27]),
    .B(_06430_),
    .S(_06369_),
    .Z(_01491_)
  );
  MUX2_X1 _28000_ (
    .A(\rf[5] [28]),
    .B(_06431_),
    .S(_06369_),
    .Z(_01492_)
  );
  MUX2_X1 _28001_ (
    .A(\rf[5] [29]),
    .B(_06432_),
    .S(_06369_),
    .Z(_01493_)
  );
  MUX2_X1 _28002_ (
    .A(\rf[5] [30]),
    .B(_06433_),
    .S(_06369_),
    .Z(_01494_)
  );
  MUX2_X1 _28003_ (
    .A(\rf[7] [0]),
    .B(_13580_),
    .S(_06366_),
    .Z(_01495_)
  );
  MUX2_X1 _28004_ (
    .A(\rf[7] [1]),
    .B(_06404_),
    .S(_06366_),
    .Z(_01496_)
  );
  MUX2_X1 _28005_ (
    .A(\rf[7] [2]),
    .B(_10137_),
    .S(_06366_),
    .Z(_01497_)
  );
  MUX2_X1 _28006_ (
    .A(\rf[7] [3]),
    .B(_10250_),
    .S(_06366_),
    .Z(_01498_)
  );
  MUX2_X1 _28007_ (
    .A(\rf[7] [4]),
    .B(_10389_),
    .S(_06366_),
    .Z(_01499_)
  );
  MUX2_X1 _28008_ (
    .A(\rf[7] [5]),
    .B(_10505_),
    .S(_06366_),
    .Z(_01500_)
  );
  MUX2_X1 _28009_ (
    .A(\rf[7] [6]),
    .B(_10620_),
    .S(_06366_),
    .Z(_01501_)
  );
  MUX2_X1 _28010_ (
    .A(\rf[7] [7]),
    .B(_06410_),
    .S(_06366_),
    .Z(_01502_)
  );
  MUX2_X1 _28011_ (
    .A(\rf[7] [8]),
    .B(_10846_),
    .S(_06366_),
    .Z(_01503_)
  );
  MUX2_X1 _28012_ (
    .A(\rf[7] [9]),
    .B(_10956_),
    .S(_06366_),
    .Z(_01504_)
  );
  MUX2_X1 _28013_ (
    .A(\rf[7] [10]),
    .B(_11066_),
    .S(_06366_),
    .Z(_01505_)
  );
  MUX2_X1 _28014_ (
    .A(\rf[7] [11]),
    .B(_11205_),
    .S(_06366_),
    .Z(_01506_)
  );
  MUX2_X1 _28015_ (
    .A(\rf[7] [12]),
    .B(_11315_),
    .S(_06366_),
    .Z(_01507_)
  );
  MUX2_X1 _28016_ (
    .A(\rf[7] [13]),
    .B(_11428_),
    .S(_06366_),
    .Z(_01508_)
  );
  MUX2_X1 _28017_ (
    .A(\rf[7] [14]),
    .B(_06417_),
    .S(_06366_),
    .Z(_01509_)
  );
  MUX2_X1 _28018_ (
    .A(\rf[7] [15]),
    .B(_11656_),
    .S(_06366_),
    .Z(_01510_)
  );
  MUX2_X1 _28019_ (
    .A(\rf[7] [16]),
    .B(_06419_),
    .S(_06366_),
    .Z(_01511_)
  );
  MUX2_X1 _28020_ (
    .A(\rf[7] [17]),
    .B(_11882_),
    .S(_06366_),
    .Z(_01512_)
  );
  MUX2_X1 _28021_ (
    .A(\rf[7] [18]),
    .B(_06421_),
    .S(_06366_),
    .Z(_01513_)
  );
  MUX2_X1 _28022_ (
    .A(\rf[7] [19]),
    .B(_06422_),
    .S(_06366_),
    .Z(_01514_)
  );
  MUX2_X1 _28023_ (
    .A(\rf[7] [20]),
    .B(_12305_),
    .S(_06366_),
    .Z(_01515_)
  );
  MUX2_X1 _28024_ (
    .A(\rf[7] [21]),
    .B(_12316_),
    .S(_06366_),
    .Z(_01516_)
  );
  MUX2_X1 _28025_ (
    .A(\rf[7] [22]),
    .B(_12537_),
    .S(_06366_),
    .Z(_01517_)
  );
  MUX2_X1 _28026_ (
    .A(\rf[7] [23]),
    .B(_12638_),
    .S(_06366_),
    .Z(_01518_)
  );
  MUX2_X1 _28027_ (
    .A(\rf[7] [24]),
    .B(_12649_),
    .S(_06366_),
    .Z(_01519_)
  );
  MUX2_X1 _28028_ (
    .A(\rf[7] [25]),
    .B(_12765_),
    .S(_06366_),
    .Z(_01520_)
  );
  MUX2_X1 _28029_ (
    .A(\rf[7] [26]),
    .B(_12986_),
    .S(_06366_),
    .Z(_01521_)
  );
  MUX2_X1 _28030_ (
    .A(\rf[7] [27]),
    .B(_06430_),
    .S(_06366_),
    .Z(_01522_)
  );
  MUX2_X1 _28031_ (
    .A(\rf[7] [28]),
    .B(_06431_),
    .S(_06366_),
    .Z(_01523_)
  );
  MUX2_X1 _28032_ (
    .A(\rf[7] [29]),
    .B(_06432_),
    .S(_06366_),
    .Z(_01524_)
  );
  MUX2_X1 _28033_ (
    .A(\rf[7] [30]),
    .B(_13349_),
    .S(_06366_),
    .Z(_01525_)
  );
  MUX2_X1 _28034_ (
    .A(\rf[3] [0]),
    .B(_13580_),
    .S(_06372_),
    .Z(_01526_)
  );
  MUX2_X1 _28035_ (
    .A(\rf[3] [1]),
    .B(_13820_),
    .S(_06372_),
    .Z(_01527_)
  );
  MUX2_X1 _28036_ (
    .A(\rf[3] [2]),
    .B(_10137_),
    .S(_06372_),
    .Z(_01528_)
  );
  MUX2_X1 _28037_ (
    .A(\rf[3] [3]),
    .B(_10250_),
    .S(_06372_),
    .Z(_01529_)
  );
  MUX2_X1 _28038_ (
    .A(\rf[3] [4]),
    .B(_10389_),
    .S(_06372_),
    .Z(_01530_)
  );
  MUX2_X1 _28039_ (
    .A(\rf[3] [5]),
    .B(_10505_),
    .S(_06372_),
    .Z(_01531_)
  );
  MUX2_X1 _28040_ (
    .A(\rf[3] [6]),
    .B(_10620_),
    .S(_06372_),
    .Z(_01532_)
  );
  MUX2_X1 _28041_ (
    .A(\rf[3] [7]),
    .B(_06410_),
    .S(_06372_),
    .Z(_01533_)
  );
  MUX2_X1 _28042_ (
    .A(\rf[3] [8]),
    .B(_10846_),
    .S(_06372_),
    .Z(_01534_)
  );
  MUX2_X1 _28043_ (
    .A(\rf[3] [9]),
    .B(_10956_),
    .S(_06372_),
    .Z(_01535_)
  );
  MUX2_X1 _28044_ (
    .A(\rf[3] [10]),
    .B(_11066_),
    .S(_06372_),
    .Z(_01536_)
  );
  MUX2_X1 _28045_ (
    .A(\rf[3] [11]),
    .B(_11205_),
    .S(_06372_),
    .Z(_01537_)
  );
  MUX2_X1 _28046_ (
    .A(\rf[3] [12]),
    .B(_11315_),
    .S(_06372_),
    .Z(_01538_)
  );
  MUX2_X1 _28047_ (
    .A(\rf[3] [13]),
    .B(_11428_),
    .S(_06372_),
    .Z(_01539_)
  );
  MUX2_X1 _28048_ (
    .A(\rf[3] [14]),
    .B(_11541_),
    .S(_06372_),
    .Z(_01540_)
  );
  MUX2_X1 _28049_ (
    .A(\rf[3] [15]),
    .B(_11656_),
    .S(_06372_),
    .Z(_01541_)
  );
  MUX2_X1 _28050_ (
    .A(\rf[3] [16]),
    .B(_06419_),
    .S(_06372_),
    .Z(_01542_)
  );
  MUX2_X1 _28051_ (
    .A(\rf[3] [17]),
    .B(_11882_),
    .S(_06372_),
    .Z(_01543_)
  );
  MUX2_X1 _28052_ (
    .A(\rf[3] [18]),
    .B(_06421_),
    .S(_06372_),
    .Z(_01544_)
  );
  MUX2_X1 _28053_ (
    .A(\rf[3] [19]),
    .B(_06422_),
    .S(_06372_),
    .Z(_01545_)
  );
  MUX2_X1 _28054_ (
    .A(\rf[3] [20]),
    .B(_12305_),
    .S(_06372_),
    .Z(_01546_)
  );
  MUX2_X1 _28055_ (
    .A(\rf[3] [21]),
    .B(_12316_),
    .S(_06372_),
    .Z(_01547_)
  );
  MUX2_X1 _28056_ (
    .A(\rf[3] [22]),
    .B(_12537_),
    .S(_06372_),
    .Z(_01548_)
  );
  MUX2_X1 _28057_ (
    .A(\rf[3] [23]),
    .B(_12638_),
    .S(_06372_),
    .Z(_01549_)
  );
  MUX2_X1 _28058_ (
    .A(\rf[3] [24]),
    .B(_12649_),
    .S(_06372_),
    .Z(_01550_)
  );
  MUX2_X1 _28059_ (
    .A(\rf[3] [25]),
    .B(_12765_),
    .S(_06372_),
    .Z(_01551_)
  );
  MUX2_X1 _28060_ (
    .A(\rf[3] [26]),
    .B(_12986_),
    .S(_06372_),
    .Z(_01552_)
  );
  MUX2_X1 _28061_ (
    .A(\rf[3] [27]),
    .B(_13102_),
    .S(_06372_),
    .Z(_01553_)
  );
  MUX2_X1 _28062_ (
    .A(\rf[3] [28]),
    .B(_06431_),
    .S(_06372_),
    .Z(_01554_)
  );
  MUX2_X1 _28063_ (
    .A(\rf[3] [29]),
    .B(_06432_),
    .S(_06372_),
    .Z(_01555_)
  );
  MUX2_X1 _28064_ (
    .A(\rf[3] [30]),
    .B(_13349_),
    .S(_06372_),
    .Z(_01556_)
  );
  MUX2_X1 _28065_ (
    .A(\rf[1] [0]),
    .B(_06403_),
    .S(_06389_),
    .Z(_01557_)
  );
  MUX2_X1 _28066_ (
    .A(\rf[1] [1]),
    .B(_06404_),
    .S(_06389_),
    .Z(_01558_)
  );
  MUX2_X1 _28067_ (
    .A(\rf[1] [2]),
    .B(_06405_),
    .S(_06389_),
    .Z(_01559_)
  );
  MUX2_X1 _28068_ (
    .A(\rf[1] [3]),
    .B(_06406_),
    .S(_06389_),
    .Z(_01560_)
  );
  MUX2_X1 _28069_ (
    .A(\rf[1] [4]),
    .B(_06407_),
    .S(_06389_),
    .Z(_01561_)
  );
  MUX2_X1 _28070_ (
    .A(\rf[1] [5]),
    .B(_06408_),
    .S(_06389_),
    .Z(_01562_)
  );
  MUX2_X1 _28071_ (
    .A(\rf[1] [6]),
    .B(_06409_),
    .S(_06389_),
    .Z(_01563_)
  );
  MUX2_X1 _28072_ (
    .A(\rf[1] [7]),
    .B(_06410_),
    .S(_06389_),
    .Z(_01564_)
  );
  MUX2_X1 _28073_ (
    .A(\rf[1] [8]),
    .B(_06411_),
    .S(_06389_),
    .Z(_01565_)
  );
  MUX2_X1 _28074_ (
    .A(\rf[1] [9]),
    .B(_06412_),
    .S(_06389_),
    .Z(_01566_)
  );
  MUX2_X1 _28075_ (
    .A(\rf[1] [10]),
    .B(_06413_),
    .S(_06389_),
    .Z(_01567_)
  );
  MUX2_X1 _28076_ (
    .A(\rf[1] [11]),
    .B(_06414_),
    .S(_06389_),
    .Z(_01568_)
  );
  MUX2_X1 _28077_ (
    .A(\rf[1] [12]),
    .B(_06415_),
    .S(_06389_),
    .Z(_01569_)
  );
  MUX2_X1 _28078_ (
    .A(\rf[1] [13]),
    .B(_06416_),
    .S(_06389_),
    .Z(_01570_)
  );
  MUX2_X1 _28079_ (
    .A(\rf[1] [14]),
    .B(_06417_),
    .S(_06389_),
    .Z(_01571_)
  );
  MUX2_X1 _28080_ (
    .A(\rf[1] [15]),
    .B(_06418_),
    .S(_06389_),
    .Z(_01572_)
  );
  MUX2_X1 _28081_ (
    .A(\rf[1] [16]),
    .B(_06419_),
    .S(_06389_),
    .Z(_01573_)
  );
  MUX2_X1 _28082_ (
    .A(\rf[1] [17]),
    .B(_06420_),
    .S(_06389_),
    .Z(_01574_)
  );
  MUX2_X1 _28083_ (
    .A(\rf[1] [18]),
    .B(_06421_),
    .S(_06389_),
    .Z(_01575_)
  );
  MUX2_X1 _28084_ (
    .A(\rf[1] [19]),
    .B(_06422_),
    .S(_06389_),
    .Z(_01576_)
  );
  MUX2_X1 _28085_ (
    .A(\rf[1] [20]),
    .B(_06423_),
    .S(_06389_),
    .Z(_01577_)
  );
  MUX2_X1 _28086_ (
    .A(\rf[1] [21]),
    .B(_06424_),
    .S(_06389_),
    .Z(_01578_)
  );
  MUX2_X1 _28087_ (
    .A(\rf[1] [22]),
    .B(_06425_),
    .S(_06389_),
    .Z(_01579_)
  );
  MUX2_X1 _28088_ (
    .A(\rf[1] [23]),
    .B(_06426_),
    .S(_06389_),
    .Z(_01580_)
  );
  MUX2_X1 _28089_ (
    .A(\rf[1] [24]),
    .B(_06427_),
    .S(_06389_),
    .Z(_01581_)
  );
  MUX2_X1 _28090_ (
    .A(\rf[1] [25]),
    .B(_06428_),
    .S(_06389_),
    .Z(_01582_)
  );
  MUX2_X1 _28091_ (
    .A(\rf[1] [26]),
    .B(_06429_),
    .S(_06389_),
    .Z(_01583_)
  );
  MUX2_X1 _28092_ (
    .A(\rf[1] [27]),
    .B(_06430_),
    .S(_06389_),
    .Z(_01584_)
  );
  MUX2_X1 _28093_ (
    .A(\rf[1] [28]),
    .B(_06431_),
    .S(_06389_),
    .Z(_01585_)
  );
  MUX2_X1 _28094_ (
    .A(\rf[1] [29]),
    .B(_06432_),
    .S(_06389_),
    .Z(_01586_)
  );
  MUX2_X1 _28095_ (
    .A(\rf[1] [30]),
    .B(_06433_),
    .S(_06389_),
    .Z(_01587_)
  );
  AND2_X1 _28096_ (
    .A1(_08567_),
    .A2(_08568_),
    .ZN(_06440_)
  );
  AND2_X1 _28097_ (
    .A1(_07955_),
    .A2(_08568_),
    .ZN(_06441_)
  );
  INV_X1 _28098_ (
    .A(_06441_),
    .ZN(_06442_)
  );
  AND2_X1 _28099_ (
    .A1(_07956_),
    .A2(_08567_),
    .ZN(_06443_)
  );
  AND2_X1 _28100_ (
    .A1(_06442_),
    .A2(_06443_),
    .ZN(_06444_)
  );
  AND2_X1 _28101_ (
    .A1(mem_reg_wdata[0]),
    .A2(_06444_),
    .ZN(_06445_)
  );
  INV_X1 _28102_ (
    .A(_06445_),
    .ZN(_06446_)
  );
  AND2_X1 _28103_ (
    .A1(wb_reg_wdata[0]),
    .A2(_06441_),
    .ZN(_06447_)
  );
  INV_X1 _28104_ (
    .A(_06447_),
    .ZN(_06448_)
  );
  AND2_X1 _28105_ (
    .A1(_06446_),
    .A2(_06448_),
    .ZN(_06449_)
  );
  INV_X1 _28106_ (
    .A(_06449_),
    .ZN(_06450_)
  );
  MUX2_X1 _28107_ (
    .A(_06450_),
    .B(io_dmem_resp_bits_data_word_bypass[0]),
    .S(_06440_),
    .Z(_06451_)
  );
  MUX2_X1 _28108_ (
    .A(ex_reg_rs_lsb_0[0]),
    .B(_06451_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[0])
  );
  AND2_X1 _28109_ (
    .A1(mem_reg_wdata[1]),
    .A2(_06444_),
    .ZN(_06452_)
  );
  INV_X1 _28110_ (
    .A(_06452_),
    .ZN(_06453_)
  );
  AND2_X1 _28111_ (
    .A1(wb_reg_wdata[1]),
    .A2(_06441_),
    .ZN(_06454_)
  );
  INV_X1 _28112_ (
    .A(_06454_),
    .ZN(_06455_)
  );
  AND2_X1 _28113_ (
    .A1(_06453_),
    .A2(_06455_),
    .ZN(_06456_)
  );
  INV_X1 _28114_ (
    .A(_06456_),
    .ZN(_06457_)
  );
  MUX2_X1 _28115_ (
    .A(_06457_),
    .B(io_dmem_resp_bits_data_word_bypass[1]),
    .S(_06440_),
    .Z(_06458_)
  );
  MUX2_X1 _28116_ (
    .A(ex_reg_rs_lsb_0[1]),
    .B(_06458_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[1])
  );
  AND2_X1 _28117_ (
    .A1(mem_reg_wdata[2]),
    .A2(_06444_),
    .ZN(_06459_)
  );
  INV_X1 _28118_ (
    .A(_06459_),
    .ZN(_06460_)
  );
  AND2_X1 _28119_ (
    .A1(wb_reg_wdata[2]),
    .A2(_06441_),
    .ZN(_06461_)
  );
  INV_X1 _28120_ (
    .A(_06461_),
    .ZN(_06462_)
  );
  AND2_X1 _28121_ (
    .A1(_06460_),
    .A2(_06462_),
    .ZN(_06463_)
  );
  INV_X1 _28122_ (
    .A(_06463_),
    .ZN(_06464_)
  );
  MUX2_X1 _28123_ (
    .A(_06464_),
    .B(io_dmem_resp_bits_data_word_bypass[2]),
    .S(_06440_),
    .Z(_06465_)
  );
  MUX2_X1 _28124_ (
    .A(ex_reg_rs_msb_0[0]),
    .B(_06465_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[2])
  );
  AND2_X1 _28125_ (
    .A1(mem_reg_wdata[3]),
    .A2(_06444_),
    .ZN(_06466_)
  );
  INV_X1 _28126_ (
    .A(_06466_),
    .ZN(_06467_)
  );
  AND2_X1 _28127_ (
    .A1(wb_reg_wdata[3]),
    .A2(_06441_),
    .ZN(_06468_)
  );
  INV_X1 _28128_ (
    .A(_06468_),
    .ZN(_06469_)
  );
  AND2_X1 _28129_ (
    .A1(_06467_),
    .A2(_06469_),
    .ZN(_06470_)
  );
  INV_X1 _28130_ (
    .A(_06470_),
    .ZN(_06471_)
  );
  MUX2_X1 _28131_ (
    .A(_06471_),
    .B(io_dmem_resp_bits_data_word_bypass[3]),
    .S(_06440_),
    .Z(_06472_)
  );
  MUX2_X1 _28132_ (
    .A(ex_reg_rs_msb_0[1]),
    .B(_06472_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[3])
  );
  AND2_X1 _28133_ (
    .A1(mem_reg_wdata[4]),
    .A2(_06444_),
    .ZN(_06473_)
  );
  INV_X1 _28134_ (
    .A(_06473_),
    .ZN(_06474_)
  );
  AND2_X1 _28135_ (
    .A1(wb_reg_wdata[4]),
    .A2(_06441_),
    .ZN(_06475_)
  );
  INV_X1 _28136_ (
    .A(_06475_),
    .ZN(_06476_)
  );
  AND2_X1 _28137_ (
    .A1(_06474_),
    .A2(_06476_),
    .ZN(_06477_)
  );
  INV_X1 _28138_ (
    .A(_06477_),
    .ZN(_06478_)
  );
  MUX2_X1 _28139_ (
    .A(_06478_),
    .B(io_dmem_resp_bits_data_word_bypass[4]),
    .S(_06440_),
    .Z(_06479_)
  );
  MUX2_X1 _28140_ (
    .A(ex_reg_rs_msb_0[2]),
    .B(_06479_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[4])
  );
  AND2_X1 _28141_ (
    .A1(mem_reg_wdata[5]),
    .A2(_06444_),
    .ZN(_06480_)
  );
  INV_X1 _28142_ (
    .A(_06480_),
    .ZN(_06481_)
  );
  AND2_X1 _28143_ (
    .A1(wb_reg_wdata[5]),
    .A2(_06441_),
    .ZN(_06482_)
  );
  INV_X1 _28144_ (
    .A(_06482_),
    .ZN(_06483_)
  );
  AND2_X1 _28145_ (
    .A1(_06481_),
    .A2(_06483_),
    .ZN(_06484_)
  );
  INV_X1 _28146_ (
    .A(_06484_),
    .ZN(_06485_)
  );
  MUX2_X1 _28147_ (
    .A(_06485_),
    .B(io_dmem_resp_bits_data_word_bypass[5]),
    .S(_06440_),
    .Z(_06486_)
  );
  MUX2_X1 _28148_ (
    .A(ex_reg_rs_msb_0[3]),
    .B(_06486_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[5])
  );
  AND2_X1 _28149_ (
    .A1(mem_reg_wdata[6]),
    .A2(_06444_),
    .ZN(_06487_)
  );
  INV_X1 _28150_ (
    .A(_06487_),
    .ZN(_06488_)
  );
  AND2_X1 _28151_ (
    .A1(wb_reg_wdata[6]),
    .A2(_06441_),
    .ZN(_06489_)
  );
  INV_X1 _28152_ (
    .A(_06489_),
    .ZN(_06490_)
  );
  AND2_X1 _28153_ (
    .A1(_06488_),
    .A2(_06490_),
    .ZN(_06491_)
  );
  INV_X1 _28154_ (
    .A(_06491_),
    .ZN(_06492_)
  );
  MUX2_X1 _28155_ (
    .A(_06492_),
    .B(io_dmem_resp_bits_data_word_bypass[6]),
    .S(_06440_),
    .Z(_06493_)
  );
  MUX2_X1 _28156_ (
    .A(ex_reg_rs_msb_0[4]),
    .B(_06493_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[6])
  );
  AND2_X1 _28157_ (
    .A1(mem_reg_wdata[7]),
    .A2(_06444_),
    .ZN(_06494_)
  );
  INV_X1 _28158_ (
    .A(_06494_),
    .ZN(_06495_)
  );
  AND2_X1 _28159_ (
    .A1(wb_reg_wdata[7]),
    .A2(_06441_),
    .ZN(_06496_)
  );
  INV_X1 _28160_ (
    .A(_06496_),
    .ZN(_06497_)
  );
  AND2_X1 _28161_ (
    .A1(_06495_),
    .A2(_06497_),
    .ZN(_06498_)
  );
  INV_X1 _28162_ (
    .A(_06498_),
    .ZN(_06499_)
  );
  MUX2_X1 _28163_ (
    .A(_06499_),
    .B(io_dmem_resp_bits_data_word_bypass[7]),
    .S(_06440_),
    .Z(_06500_)
  );
  MUX2_X1 _28164_ (
    .A(ex_reg_rs_msb_0[5]),
    .B(_06500_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[7])
  );
  AND2_X1 _28165_ (
    .A1(mem_reg_wdata[8]),
    .A2(_06444_),
    .ZN(_06501_)
  );
  INV_X1 _28166_ (
    .A(_06501_),
    .ZN(_06502_)
  );
  AND2_X1 _28167_ (
    .A1(wb_reg_wdata[8]),
    .A2(_06441_),
    .ZN(_06503_)
  );
  INV_X1 _28168_ (
    .A(_06503_),
    .ZN(_06504_)
  );
  AND2_X1 _28169_ (
    .A1(_06502_),
    .A2(_06504_),
    .ZN(_06505_)
  );
  INV_X1 _28170_ (
    .A(_06505_),
    .ZN(_06506_)
  );
  MUX2_X1 _28171_ (
    .A(_06506_),
    .B(io_dmem_resp_bits_data_word_bypass[8]),
    .S(_06440_),
    .Z(_06507_)
  );
  MUX2_X1 _28172_ (
    .A(ex_reg_rs_msb_0[6]),
    .B(_06507_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[8])
  );
  AND2_X1 _28173_ (
    .A1(mem_reg_wdata[9]),
    .A2(_06444_),
    .ZN(_06508_)
  );
  INV_X1 _28174_ (
    .A(_06508_),
    .ZN(_06509_)
  );
  AND2_X1 _28175_ (
    .A1(wb_reg_wdata[9]),
    .A2(_06441_),
    .ZN(_06510_)
  );
  INV_X1 _28176_ (
    .A(_06510_),
    .ZN(_06511_)
  );
  AND2_X1 _28177_ (
    .A1(_06509_),
    .A2(_06511_),
    .ZN(_06512_)
  );
  INV_X1 _28178_ (
    .A(_06512_),
    .ZN(_06513_)
  );
  MUX2_X1 _28179_ (
    .A(_06513_),
    .B(io_dmem_resp_bits_data_word_bypass[9]),
    .S(_06440_),
    .Z(_06514_)
  );
  MUX2_X1 _28180_ (
    .A(ex_reg_rs_msb_0[7]),
    .B(_06514_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[9])
  );
  AND2_X1 _28181_ (
    .A1(mem_reg_wdata[10]),
    .A2(_06444_),
    .ZN(_06515_)
  );
  INV_X1 _28182_ (
    .A(_06515_),
    .ZN(_06516_)
  );
  AND2_X1 _28183_ (
    .A1(wb_reg_wdata[10]),
    .A2(_06441_),
    .ZN(_06517_)
  );
  INV_X1 _28184_ (
    .A(_06517_),
    .ZN(_06518_)
  );
  AND2_X1 _28185_ (
    .A1(_06516_),
    .A2(_06518_),
    .ZN(_06519_)
  );
  INV_X1 _28186_ (
    .A(_06519_),
    .ZN(_06520_)
  );
  MUX2_X1 _28187_ (
    .A(_06520_),
    .B(io_dmem_resp_bits_data_word_bypass[10]),
    .S(_06440_),
    .Z(_06521_)
  );
  MUX2_X1 _28188_ (
    .A(ex_reg_rs_msb_0[8]),
    .B(_06521_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[10])
  );
  AND2_X1 _28189_ (
    .A1(mem_reg_wdata[11]),
    .A2(_06444_),
    .ZN(_06522_)
  );
  INV_X1 _28190_ (
    .A(_06522_),
    .ZN(_06523_)
  );
  AND2_X1 _28191_ (
    .A1(wb_reg_wdata[11]),
    .A2(_06441_),
    .ZN(_06524_)
  );
  INV_X1 _28192_ (
    .A(_06524_),
    .ZN(_06525_)
  );
  AND2_X1 _28193_ (
    .A1(_06523_),
    .A2(_06525_),
    .ZN(_06526_)
  );
  INV_X1 _28194_ (
    .A(_06526_),
    .ZN(_06527_)
  );
  MUX2_X1 _28195_ (
    .A(_06527_),
    .B(io_dmem_resp_bits_data_word_bypass[11]),
    .S(_06440_),
    .Z(_06528_)
  );
  MUX2_X1 _28196_ (
    .A(ex_reg_rs_msb_0[9]),
    .B(_06528_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[11])
  );
  AND2_X1 _28197_ (
    .A1(mem_reg_wdata[12]),
    .A2(_06444_),
    .ZN(_06529_)
  );
  INV_X1 _28198_ (
    .A(_06529_),
    .ZN(_06530_)
  );
  AND2_X1 _28199_ (
    .A1(wb_reg_wdata[12]),
    .A2(_06441_),
    .ZN(_06531_)
  );
  INV_X1 _28200_ (
    .A(_06531_),
    .ZN(_06532_)
  );
  AND2_X1 _28201_ (
    .A1(_06530_),
    .A2(_06532_),
    .ZN(_06533_)
  );
  INV_X1 _28202_ (
    .A(_06533_),
    .ZN(_06534_)
  );
  MUX2_X1 _28203_ (
    .A(_06534_),
    .B(io_dmem_resp_bits_data_word_bypass[12]),
    .S(_06440_),
    .Z(_06535_)
  );
  MUX2_X1 _28204_ (
    .A(ex_reg_rs_msb_0[10]),
    .B(_06535_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[12])
  );
  AND2_X1 _28205_ (
    .A1(mem_reg_wdata[13]),
    .A2(_06444_),
    .ZN(_06536_)
  );
  INV_X1 _28206_ (
    .A(_06536_),
    .ZN(_06537_)
  );
  AND2_X1 _28207_ (
    .A1(wb_reg_wdata[13]),
    .A2(_06441_),
    .ZN(_06538_)
  );
  INV_X1 _28208_ (
    .A(_06538_),
    .ZN(_06539_)
  );
  AND2_X1 _28209_ (
    .A1(_06537_),
    .A2(_06539_),
    .ZN(_06540_)
  );
  INV_X1 _28210_ (
    .A(_06540_),
    .ZN(_06541_)
  );
  MUX2_X1 _28211_ (
    .A(_06541_),
    .B(io_dmem_resp_bits_data_word_bypass[13]),
    .S(_06440_),
    .Z(_06542_)
  );
  MUX2_X1 _28212_ (
    .A(ex_reg_rs_msb_0[11]),
    .B(_06542_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[13])
  );
  AND2_X1 _28213_ (
    .A1(mem_reg_wdata[14]),
    .A2(_06444_),
    .ZN(_06543_)
  );
  INV_X1 _28214_ (
    .A(_06543_),
    .ZN(_06544_)
  );
  AND2_X1 _28215_ (
    .A1(wb_reg_wdata[14]),
    .A2(_06441_),
    .ZN(_06545_)
  );
  INV_X1 _28216_ (
    .A(_06545_),
    .ZN(_06546_)
  );
  AND2_X1 _28217_ (
    .A1(_06544_),
    .A2(_06546_),
    .ZN(_06547_)
  );
  INV_X1 _28218_ (
    .A(_06547_),
    .ZN(_06548_)
  );
  MUX2_X1 _28219_ (
    .A(_06548_),
    .B(io_dmem_resp_bits_data_word_bypass[14]),
    .S(_06440_),
    .Z(_06549_)
  );
  MUX2_X1 _28220_ (
    .A(ex_reg_rs_msb_0[12]),
    .B(_06549_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[14])
  );
  AND2_X1 _28221_ (
    .A1(mem_reg_wdata[15]),
    .A2(_06444_),
    .ZN(_06550_)
  );
  INV_X1 _28222_ (
    .A(_06550_),
    .ZN(_06551_)
  );
  AND2_X1 _28223_ (
    .A1(wb_reg_wdata[15]),
    .A2(_06441_),
    .ZN(_06552_)
  );
  INV_X1 _28224_ (
    .A(_06552_),
    .ZN(_06553_)
  );
  AND2_X1 _28225_ (
    .A1(_06551_),
    .A2(_06553_),
    .ZN(_06554_)
  );
  INV_X1 _28226_ (
    .A(_06554_),
    .ZN(_06555_)
  );
  MUX2_X1 _28227_ (
    .A(_06555_),
    .B(io_dmem_resp_bits_data_word_bypass[15]),
    .S(_06440_),
    .Z(_06556_)
  );
  MUX2_X1 _28228_ (
    .A(ex_reg_rs_msb_0[13]),
    .B(_06556_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[15])
  );
  AND2_X1 _28229_ (
    .A1(mem_reg_wdata[16]),
    .A2(_06444_),
    .ZN(_06557_)
  );
  INV_X1 _28230_ (
    .A(_06557_),
    .ZN(_06558_)
  );
  AND2_X1 _28231_ (
    .A1(wb_reg_wdata[16]),
    .A2(_06441_),
    .ZN(_06559_)
  );
  INV_X1 _28232_ (
    .A(_06559_),
    .ZN(_06560_)
  );
  AND2_X1 _28233_ (
    .A1(_06558_),
    .A2(_06560_),
    .ZN(_06561_)
  );
  INV_X1 _28234_ (
    .A(_06561_),
    .ZN(_06562_)
  );
  MUX2_X1 _28235_ (
    .A(_06562_),
    .B(io_dmem_resp_bits_data_word_bypass[16]),
    .S(_06440_),
    .Z(_06563_)
  );
  MUX2_X1 _28236_ (
    .A(ex_reg_rs_msb_0[14]),
    .B(_06563_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[16])
  );
  AND2_X1 _28237_ (
    .A1(mem_reg_wdata[17]),
    .A2(_06444_),
    .ZN(_06564_)
  );
  INV_X1 _28238_ (
    .A(_06564_),
    .ZN(_06565_)
  );
  AND2_X1 _28239_ (
    .A1(wb_reg_wdata[17]),
    .A2(_06441_),
    .ZN(_06566_)
  );
  INV_X1 _28240_ (
    .A(_06566_),
    .ZN(_06567_)
  );
  AND2_X1 _28241_ (
    .A1(_06565_),
    .A2(_06567_),
    .ZN(_06568_)
  );
  INV_X1 _28242_ (
    .A(_06568_),
    .ZN(_06569_)
  );
  MUX2_X1 _28243_ (
    .A(_06569_),
    .B(io_dmem_resp_bits_data_word_bypass[17]),
    .S(_06440_),
    .Z(_06570_)
  );
  MUX2_X1 _28244_ (
    .A(ex_reg_rs_msb_0[15]),
    .B(_06570_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[17])
  );
  AND2_X1 _28245_ (
    .A1(mem_reg_wdata[18]),
    .A2(_06444_),
    .ZN(_06571_)
  );
  INV_X1 _28246_ (
    .A(_06571_),
    .ZN(_06572_)
  );
  AND2_X1 _28247_ (
    .A1(wb_reg_wdata[18]),
    .A2(_06441_),
    .ZN(_06573_)
  );
  INV_X1 _28248_ (
    .A(_06573_),
    .ZN(_06574_)
  );
  AND2_X1 _28249_ (
    .A1(_06572_),
    .A2(_06574_),
    .ZN(_06575_)
  );
  INV_X1 _28250_ (
    .A(_06575_),
    .ZN(_06576_)
  );
  MUX2_X1 _28251_ (
    .A(_06576_),
    .B(io_dmem_resp_bits_data_word_bypass[18]),
    .S(_06440_),
    .Z(_06577_)
  );
  MUX2_X1 _28252_ (
    .A(ex_reg_rs_msb_0[16]),
    .B(_06577_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[18])
  );
  AND2_X1 _28253_ (
    .A1(mem_reg_wdata[19]),
    .A2(_06444_),
    .ZN(_06578_)
  );
  INV_X1 _28254_ (
    .A(_06578_),
    .ZN(_06579_)
  );
  AND2_X1 _28255_ (
    .A1(wb_reg_wdata[19]),
    .A2(_06441_),
    .ZN(_06580_)
  );
  INV_X1 _28256_ (
    .A(_06580_),
    .ZN(_06581_)
  );
  AND2_X1 _28257_ (
    .A1(_06579_),
    .A2(_06581_),
    .ZN(_06582_)
  );
  INV_X1 _28258_ (
    .A(_06582_),
    .ZN(_06583_)
  );
  MUX2_X1 _28259_ (
    .A(_06583_),
    .B(io_dmem_resp_bits_data_word_bypass[19]),
    .S(_06440_),
    .Z(_06584_)
  );
  MUX2_X1 _28260_ (
    .A(ex_reg_rs_msb_0[17]),
    .B(_06584_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[19])
  );
  AND2_X1 _28261_ (
    .A1(mem_reg_wdata[20]),
    .A2(_06444_),
    .ZN(_06585_)
  );
  INV_X1 _28262_ (
    .A(_06585_),
    .ZN(_06586_)
  );
  AND2_X1 _28263_ (
    .A1(wb_reg_wdata[20]),
    .A2(_06441_),
    .ZN(_06587_)
  );
  INV_X1 _28264_ (
    .A(_06587_),
    .ZN(_06588_)
  );
  AND2_X1 _28265_ (
    .A1(_06586_),
    .A2(_06588_),
    .ZN(_06589_)
  );
  INV_X1 _28266_ (
    .A(_06589_),
    .ZN(_06590_)
  );
  MUX2_X1 _28267_ (
    .A(_06590_),
    .B(io_dmem_resp_bits_data_word_bypass[20]),
    .S(_06440_),
    .Z(_06591_)
  );
  MUX2_X1 _28268_ (
    .A(ex_reg_rs_msb_0[18]),
    .B(_06591_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[20])
  );
  AND2_X1 _28269_ (
    .A1(mem_reg_wdata[21]),
    .A2(_06444_),
    .ZN(_06592_)
  );
  INV_X1 _28270_ (
    .A(_06592_),
    .ZN(_06593_)
  );
  AND2_X1 _28271_ (
    .A1(wb_reg_wdata[21]),
    .A2(_06441_),
    .ZN(_06594_)
  );
  INV_X1 _28272_ (
    .A(_06594_),
    .ZN(_06595_)
  );
  AND2_X1 _28273_ (
    .A1(_06593_),
    .A2(_06595_),
    .ZN(_06596_)
  );
  INV_X1 _28274_ (
    .A(_06596_),
    .ZN(_06597_)
  );
  MUX2_X1 _28275_ (
    .A(_06597_),
    .B(io_dmem_resp_bits_data_word_bypass[21]),
    .S(_06440_),
    .Z(_06598_)
  );
  MUX2_X1 _28276_ (
    .A(ex_reg_rs_msb_0[19]),
    .B(_06598_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[21])
  );
  AND2_X1 _28277_ (
    .A1(mem_reg_wdata[22]),
    .A2(_06444_),
    .ZN(_06599_)
  );
  INV_X1 _28278_ (
    .A(_06599_),
    .ZN(_06600_)
  );
  AND2_X1 _28279_ (
    .A1(wb_reg_wdata[22]),
    .A2(_06441_),
    .ZN(_06601_)
  );
  INV_X1 _28280_ (
    .A(_06601_),
    .ZN(_06602_)
  );
  AND2_X1 _28281_ (
    .A1(_06600_),
    .A2(_06602_),
    .ZN(_06603_)
  );
  INV_X1 _28282_ (
    .A(_06603_),
    .ZN(_06604_)
  );
  MUX2_X1 _28283_ (
    .A(_06604_),
    .B(io_dmem_resp_bits_data_word_bypass[22]),
    .S(_06440_),
    .Z(_06605_)
  );
  MUX2_X1 _28284_ (
    .A(ex_reg_rs_msb_0[20]),
    .B(_06605_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[22])
  );
  AND2_X1 _28285_ (
    .A1(mem_reg_wdata[23]),
    .A2(_06444_),
    .ZN(_06606_)
  );
  INV_X1 _28286_ (
    .A(_06606_),
    .ZN(_06607_)
  );
  AND2_X1 _28287_ (
    .A1(wb_reg_wdata[23]),
    .A2(_06441_),
    .ZN(_06608_)
  );
  INV_X1 _28288_ (
    .A(_06608_),
    .ZN(_06609_)
  );
  AND2_X1 _28289_ (
    .A1(_06607_),
    .A2(_06609_),
    .ZN(_06610_)
  );
  INV_X1 _28290_ (
    .A(_06610_),
    .ZN(_06611_)
  );
  MUX2_X1 _28291_ (
    .A(_06611_),
    .B(io_dmem_resp_bits_data_word_bypass[23]),
    .S(_06440_),
    .Z(_06612_)
  );
  MUX2_X1 _28292_ (
    .A(ex_reg_rs_msb_0[21]),
    .B(_06612_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[23])
  );
  AND2_X1 _28293_ (
    .A1(mem_reg_wdata[24]),
    .A2(_06444_),
    .ZN(_06613_)
  );
  INV_X1 _28294_ (
    .A(_06613_),
    .ZN(_06614_)
  );
  AND2_X1 _28295_ (
    .A1(wb_reg_wdata[24]),
    .A2(_06441_),
    .ZN(_06615_)
  );
  INV_X1 _28296_ (
    .A(_06615_),
    .ZN(_06616_)
  );
  AND2_X1 _28297_ (
    .A1(_06614_),
    .A2(_06616_),
    .ZN(_06617_)
  );
  INV_X1 _28298_ (
    .A(_06617_),
    .ZN(_06618_)
  );
  MUX2_X1 _28299_ (
    .A(_06618_),
    .B(io_dmem_resp_bits_data_word_bypass[24]),
    .S(_06440_),
    .Z(_06619_)
  );
  MUX2_X1 _28300_ (
    .A(ex_reg_rs_msb_0[22]),
    .B(_06619_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[24])
  );
  AND2_X1 _28301_ (
    .A1(mem_reg_wdata[25]),
    .A2(_06444_),
    .ZN(_06620_)
  );
  INV_X1 _28302_ (
    .A(_06620_),
    .ZN(_06621_)
  );
  AND2_X1 _28303_ (
    .A1(wb_reg_wdata[25]),
    .A2(_06441_),
    .ZN(_06622_)
  );
  INV_X1 _28304_ (
    .A(_06622_),
    .ZN(_06623_)
  );
  AND2_X1 _28305_ (
    .A1(_06621_),
    .A2(_06623_),
    .ZN(_06624_)
  );
  INV_X1 _28306_ (
    .A(_06624_),
    .ZN(_06625_)
  );
  MUX2_X1 _28307_ (
    .A(_06625_),
    .B(io_dmem_resp_bits_data_word_bypass[25]),
    .S(_06440_),
    .Z(_06626_)
  );
  MUX2_X1 _28308_ (
    .A(ex_reg_rs_msb_0[23]),
    .B(_06626_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[25])
  );
  AND2_X1 _28309_ (
    .A1(mem_reg_wdata[26]),
    .A2(_06444_),
    .ZN(_06627_)
  );
  INV_X1 _28310_ (
    .A(_06627_),
    .ZN(_06628_)
  );
  AND2_X1 _28311_ (
    .A1(wb_reg_wdata[26]),
    .A2(_06441_),
    .ZN(_06629_)
  );
  INV_X1 _28312_ (
    .A(_06629_),
    .ZN(_06630_)
  );
  AND2_X1 _28313_ (
    .A1(_06628_),
    .A2(_06630_),
    .ZN(_06631_)
  );
  INV_X1 _28314_ (
    .A(_06631_),
    .ZN(_06632_)
  );
  MUX2_X1 _28315_ (
    .A(_06632_),
    .B(io_dmem_resp_bits_data_word_bypass[26]),
    .S(_06440_),
    .Z(_06633_)
  );
  MUX2_X1 _28316_ (
    .A(ex_reg_rs_msb_0[24]),
    .B(_06633_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[26])
  );
  AND2_X1 _28317_ (
    .A1(mem_reg_wdata[27]),
    .A2(_06444_),
    .ZN(_06634_)
  );
  INV_X1 _28318_ (
    .A(_06634_),
    .ZN(_06635_)
  );
  AND2_X1 _28319_ (
    .A1(wb_reg_wdata[27]),
    .A2(_06441_),
    .ZN(_06636_)
  );
  INV_X1 _28320_ (
    .A(_06636_),
    .ZN(_06637_)
  );
  AND2_X1 _28321_ (
    .A1(_06635_),
    .A2(_06637_),
    .ZN(_06638_)
  );
  INV_X1 _28322_ (
    .A(_06638_),
    .ZN(_06639_)
  );
  MUX2_X1 _28323_ (
    .A(_06639_),
    .B(io_dmem_resp_bits_data_word_bypass[27]),
    .S(_06440_),
    .Z(_06640_)
  );
  MUX2_X1 _28324_ (
    .A(ex_reg_rs_msb_0[25]),
    .B(_06640_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[27])
  );
  AND2_X1 _28325_ (
    .A1(mem_reg_wdata[28]),
    .A2(_06444_),
    .ZN(_06641_)
  );
  INV_X1 _28326_ (
    .A(_06641_),
    .ZN(_06642_)
  );
  AND2_X1 _28327_ (
    .A1(wb_reg_wdata[28]),
    .A2(_06441_),
    .ZN(_06643_)
  );
  INV_X1 _28328_ (
    .A(_06643_),
    .ZN(_06644_)
  );
  AND2_X1 _28329_ (
    .A1(_06642_),
    .A2(_06644_),
    .ZN(_06645_)
  );
  INV_X1 _28330_ (
    .A(_06645_),
    .ZN(_06646_)
  );
  MUX2_X1 _28331_ (
    .A(_06646_),
    .B(io_dmem_resp_bits_data_word_bypass[28]),
    .S(_06440_),
    .Z(_06647_)
  );
  MUX2_X1 _28332_ (
    .A(ex_reg_rs_msb_0[26]),
    .B(_06647_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[28])
  );
  AND2_X1 _28333_ (
    .A1(mem_reg_wdata[29]),
    .A2(_06444_),
    .ZN(_06648_)
  );
  INV_X1 _28334_ (
    .A(_06648_),
    .ZN(_06649_)
  );
  AND2_X1 _28335_ (
    .A1(wb_reg_wdata[29]),
    .A2(_06441_),
    .ZN(_06650_)
  );
  INV_X1 _28336_ (
    .A(_06650_),
    .ZN(_06651_)
  );
  AND2_X1 _28337_ (
    .A1(_06649_),
    .A2(_06651_),
    .ZN(_06652_)
  );
  INV_X1 _28338_ (
    .A(_06652_),
    .ZN(_06653_)
  );
  MUX2_X1 _28339_ (
    .A(_06653_),
    .B(io_dmem_resp_bits_data_word_bypass[29]),
    .S(_06440_),
    .Z(_06654_)
  );
  MUX2_X1 _28340_ (
    .A(ex_reg_rs_msb_0[27]),
    .B(_06654_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[29])
  );
  AND2_X1 _28341_ (
    .A1(mem_reg_wdata[30]),
    .A2(_06444_),
    .ZN(_06655_)
  );
  INV_X1 _28342_ (
    .A(_06655_),
    .ZN(_06656_)
  );
  AND2_X1 _28343_ (
    .A1(wb_reg_wdata[30]),
    .A2(_06441_),
    .ZN(_06657_)
  );
  INV_X1 _28344_ (
    .A(_06657_),
    .ZN(_06658_)
  );
  AND2_X1 _28345_ (
    .A1(_06656_),
    .A2(_06658_),
    .ZN(_06659_)
  );
  INV_X1 _28346_ (
    .A(_06659_),
    .ZN(_06660_)
  );
  MUX2_X1 _28347_ (
    .A(_06660_),
    .B(io_dmem_resp_bits_data_word_bypass[30]),
    .S(_06440_),
    .Z(_06661_)
  );
  MUX2_X1 _28348_ (
    .A(ex_reg_rs_msb_0[28]),
    .B(_06661_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[30])
  );
  AND2_X1 _28349_ (
    .A1(mem_reg_wdata[31]),
    .A2(_06444_),
    .ZN(_06662_)
  );
  INV_X1 _28350_ (
    .A(_06662_),
    .ZN(_06663_)
  );
  AND2_X1 _28351_ (
    .A1(wb_reg_wdata[31]),
    .A2(_06441_),
    .ZN(_06664_)
  );
  INV_X1 _28352_ (
    .A(_06664_),
    .ZN(_06665_)
  );
  AND2_X1 _28353_ (
    .A1(_06663_),
    .A2(_06665_),
    .ZN(_06666_)
  );
  INV_X1 _28354_ (
    .A(_06666_),
    .ZN(_06667_)
  );
  MUX2_X1 _28355_ (
    .A(_06667_),
    .B(io_dmem_resp_bits_data_word_bypass[31]),
    .S(_06440_),
    .Z(_06668_)
  );
  MUX2_X1 _28356_ (
    .A(ex_reg_rs_msb_0[29]),
    .B(_06668_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[31])
  );
  AND2_X1 _28357_ (
    .A1(wb_reg_raw_inst[0]),
    .A2(wb_reg_raw_inst[1]),
    .ZN(_06669_)
  );
  AND2_X1 _28358_ (
    .A1(wb_reg_inst[16]),
    .A2(_06669_),
    .ZN(_csr_io_inst_0_T_3[0])
  );
  AND2_X1 _28359_ (
    .A1(wb_reg_inst[17]),
    .A2(_06669_),
    .ZN(_csr_io_inst_0_T_3[1])
  );
  AND2_X1 _28360_ (
    .A1(wb_reg_inst[18]),
    .A2(_06669_),
    .ZN(_csr_io_inst_0_T_3[2])
  );
  AND2_X1 _28361_ (
    .A1(wb_reg_inst[19]),
    .A2(_06669_),
    .ZN(_csr_io_inst_0_T_3[3])
  );
  AND2_X1 _28362_ (
    .A1(wb_reg_inst[20]),
    .A2(_06669_),
    .ZN(_csr_io_inst_0_T_3[4])
  );
  AND2_X1 _28363_ (
    .A1(wb_reg_inst[21]),
    .A2(_06669_),
    .ZN(_csr_io_inst_0_T_3[5])
  );
  AND2_X1 _28364_ (
    .A1(wb_reg_inst[22]),
    .A2(_06669_),
    .ZN(_csr_io_inst_0_T_3[6])
  );
  AND2_X1 _28365_ (
    .A1(wb_reg_inst[23]),
    .A2(_06669_),
    .ZN(_csr_io_inst_0_T_3[7])
  );
  AND2_X1 _28366_ (
    .A1(wb_reg_inst[24]),
    .A2(_06669_),
    .ZN(_csr_io_inst_0_T_3[8])
  );
  AND2_X1 _28367_ (
    .A1(wb_reg_inst[25]),
    .A2(_06669_),
    .ZN(_csr_io_inst_0_T_3[9])
  );
  AND2_X1 _28368_ (
    .A1(wb_reg_inst[26]),
    .A2(_06669_),
    .ZN(_csr_io_inst_0_T_3[10])
  );
  AND2_X1 _28369_ (
    .A1(wb_reg_inst[27]),
    .A2(_06669_),
    .ZN(_csr_io_inst_0_T_3[11])
  );
  AND2_X1 _28370_ (
    .A1(wb_reg_inst[28]),
    .A2(_06669_),
    .ZN(_csr_io_inst_0_T_3[12])
  );
  AND2_X1 _28371_ (
    .A1(wb_reg_inst[29]),
    .A2(_06669_),
    .ZN(_csr_io_inst_0_T_3[13])
  );
  AND2_X1 _28372_ (
    .A1(wb_reg_inst[30]),
    .A2(_06669_),
    .ZN(_csr_io_inst_0_T_3[14])
  );
  AND2_X1 _28373_ (
    .A1(wb_reg_inst[31]),
    .A2(_06669_),
    .ZN(_csr_io_inst_0_T_3[15])
  );
  AND2_X1 _28374_ (
    .A1(wb_reg_pc[0]),
    .A2(_08687_),
    .ZN(_06670_)
  );
  MUX2_X1 _28375_ (
    .A(csr_io_evec[0]),
    .B(_06670_),
    .S(_10063_),
    .Z(io_imem_req_bits_pc[0])
  );
  AND2_X1 _28376_ (
    .A1(_08686_),
    .A2(_13843_),
    .ZN(_06671_)
  );
  INV_X1 _28377_ (
    .A(_06671_),
    .ZN(_06672_)
  );
  AND2_X1 _28378_ (
    .A1(wb_reg_pc[1]),
    .A2(_08687_),
    .ZN(_06673_)
  );
  INV_X1 _28379_ (
    .A(_06673_),
    .ZN(_06674_)
  );
  AND2_X1 _28380_ (
    .A1(_10063_),
    .A2(_06674_),
    .ZN(_06675_)
  );
  AND2_X1 _28381_ (
    .A1(_06672_),
    .A2(_06675_),
    .ZN(_06676_)
  );
  INV_X1 _28382_ (
    .A(_06676_),
    .ZN(_06677_)
  );
  AND2_X1 _28383_ (
    .A1(_08594_),
    .A2(_10064_),
    .ZN(_06678_)
  );
  INV_X1 _28384_ (
    .A(_06678_),
    .ZN(_06679_)
  );
  AND2_X1 _28385_ (
    .A1(_06677_),
    .A2(_06679_),
    .ZN(io_imem_req_bits_pc[1])
  );
  MUX2_X1 _28386_ (
    .A(mem_reg_wdata[2]),
    .B(_13869_),
    .S(_08206_),
    .Z(_06680_)
  );
  INV_X1 _28387_ (
    .A(_06680_),
    .ZN(_06681_)
  );
  MUX2_X1 _28388_ (
    .A(wb_reg_pc[2]),
    .B(_06680_),
    .S(_08686_),
    .Z(_06682_)
  );
  MUX2_X1 _28389_ (
    .A(csr_io_evec[2]),
    .B(_06682_),
    .S(_10063_),
    .Z(io_imem_req_bits_pc[2])
  );
  MUX2_X1 _28390_ (
    .A(mem_reg_wdata[3]),
    .B(_13886_),
    .S(_08206_),
    .Z(_06683_)
  );
  INV_X1 _28391_ (
    .A(_06683_),
    .ZN(_06684_)
  );
  MUX2_X1 _28392_ (
    .A(wb_reg_pc[3]),
    .B(_06683_),
    .S(_08686_),
    .Z(_06685_)
  );
  MUX2_X1 _28393_ (
    .A(csr_io_evec[3]),
    .B(_06685_),
    .S(_10063_),
    .Z(io_imem_req_bits_pc[3])
  );
  MUX2_X1 _28394_ (
    .A(mem_reg_wdata[4]),
    .B(_13907_),
    .S(_08206_),
    .Z(_06686_)
  );
  INV_X1 _28395_ (
    .A(_06686_),
    .ZN(_06687_)
  );
  MUX2_X1 _28396_ (
    .A(wb_reg_pc[4]),
    .B(_06686_),
    .S(_08686_),
    .Z(_06688_)
  );
  MUX2_X1 _28397_ (
    .A(csr_io_evec[4]),
    .B(_06688_),
    .S(_10063_),
    .Z(io_imem_req_bits_pc[4])
  );
  AND2_X1 _28398_ (
    .A1(csr_io_evec[5]),
    .A2(_10064_),
    .ZN(_06689_)
  );
  INV_X1 _28399_ (
    .A(_06689_),
    .ZN(_06690_)
  );
  MUX2_X1 _28400_ (
    .A(_08057_),
    .B(_13926_),
    .S(_08206_),
    .Z(_06691_)
  );
  INV_X1 _28401_ (
    .A(_06691_),
    .ZN(_06692_)
  );
  AND2_X1 _28402_ (
    .A1(_08686_),
    .A2(_06691_),
    .ZN(_06693_)
  );
  INV_X1 _28403_ (
    .A(_06693_),
    .ZN(_06694_)
  );
  AND2_X1 _28404_ (
    .A1(_07989_),
    .A2(_08687_),
    .ZN(_06695_)
  );
  INV_X1 _28405_ (
    .A(_06695_),
    .ZN(_06696_)
  );
  AND2_X1 _28406_ (
    .A1(_10063_),
    .A2(_06696_),
    .ZN(_06697_)
  );
  AND2_X1 _28407_ (
    .A1(_06694_),
    .A2(_06697_),
    .ZN(_06698_)
  );
  INV_X1 _28408_ (
    .A(_06698_),
    .ZN(_06699_)
  );
  AND2_X1 _28409_ (
    .A1(_06690_),
    .A2(_06699_),
    .ZN(_06700_)
  );
  INV_X1 _28410_ (
    .A(_06700_),
    .ZN(io_imem_req_bits_pc[5])
  );
  AND2_X1 _28411_ (
    .A1(csr_io_evec[6]),
    .A2(_10064_),
    .ZN(_06701_)
  );
  INV_X1 _28412_ (
    .A(_06701_),
    .ZN(_06702_)
  );
  MUX2_X1 _28413_ (
    .A(_08058_),
    .B(_13952_),
    .S(_08206_),
    .Z(_06703_)
  );
  INV_X1 _28414_ (
    .A(_06703_),
    .ZN(_06704_)
  );
  AND2_X1 _28415_ (
    .A1(_08686_),
    .A2(_06703_),
    .ZN(_06705_)
  );
  INV_X1 _28416_ (
    .A(_06705_),
    .ZN(_06706_)
  );
  AND2_X1 _28417_ (
    .A1(_07991_),
    .A2(_08687_),
    .ZN(_06707_)
  );
  INV_X1 _28418_ (
    .A(_06707_),
    .ZN(_06708_)
  );
  AND2_X1 _28419_ (
    .A1(_10063_),
    .A2(_06708_),
    .ZN(_06709_)
  );
  AND2_X1 _28420_ (
    .A1(_06706_),
    .A2(_06709_),
    .ZN(_06710_)
  );
  INV_X1 _28421_ (
    .A(_06710_),
    .ZN(_06711_)
  );
  AND2_X1 _28422_ (
    .A1(_06702_),
    .A2(_06711_),
    .ZN(_06712_)
  );
  INV_X1 _28423_ (
    .A(_06712_),
    .ZN(io_imem_req_bits_pc[6])
  );
  AND2_X1 _28424_ (
    .A1(csr_io_evec[7]),
    .A2(_10064_),
    .ZN(_06713_)
  );
  INV_X1 _28425_ (
    .A(_06713_),
    .ZN(_06714_)
  );
  MUX2_X1 _28426_ (
    .A(_08059_),
    .B(_13977_),
    .S(_08206_),
    .Z(_06715_)
  );
  INV_X1 _28427_ (
    .A(_06715_),
    .ZN(_06716_)
  );
  AND2_X1 _28428_ (
    .A1(_08686_),
    .A2(_06715_),
    .ZN(_06717_)
  );
  INV_X1 _28429_ (
    .A(_06717_),
    .ZN(_06718_)
  );
  AND2_X1 _28430_ (
    .A1(_07993_),
    .A2(_08687_),
    .ZN(_06719_)
  );
  INV_X1 _28431_ (
    .A(_06719_),
    .ZN(_06720_)
  );
  AND2_X1 _28432_ (
    .A1(_10063_),
    .A2(_06720_),
    .ZN(_06721_)
  );
  AND2_X1 _28433_ (
    .A1(_06718_),
    .A2(_06721_),
    .ZN(_06722_)
  );
  INV_X1 _28434_ (
    .A(_06722_),
    .ZN(_06723_)
  );
  AND2_X1 _28435_ (
    .A1(_06714_),
    .A2(_06723_),
    .ZN(_06724_)
  );
  INV_X1 _28436_ (
    .A(_06724_),
    .ZN(io_imem_req_bits_pc[7])
  );
  AND2_X1 _28437_ (
    .A1(csr_io_evec[8]),
    .A2(_10064_),
    .ZN(_06725_)
  );
  INV_X1 _28438_ (
    .A(_06725_),
    .ZN(_06726_)
  );
  MUX2_X1 _28439_ (
    .A(_08060_),
    .B(_14005_),
    .S(_08206_),
    .Z(_06727_)
  );
  INV_X1 _28440_ (
    .A(_06727_),
    .ZN(_06728_)
  );
  AND2_X1 _28441_ (
    .A1(_08686_),
    .A2(_06727_),
    .ZN(_06729_)
  );
  INV_X1 _28442_ (
    .A(_06729_),
    .ZN(_06730_)
  );
  AND2_X1 _28443_ (
    .A1(_07995_),
    .A2(_08687_),
    .ZN(_06731_)
  );
  INV_X1 _28444_ (
    .A(_06731_),
    .ZN(_06732_)
  );
  AND2_X1 _28445_ (
    .A1(_10063_),
    .A2(_06732_),
    .ZN(_06733_)
  );
  AND2_X1 _28446_ (
    .A1(_06730_),
    .A2(_06733_),
    .ZN(_06734_)
  );
  INV_X1 _28447_ (
    .A(_06734_),
    .ZN(_06735_)
  );
  AND2_X1 _28448_ (
    .A1(_06726_),
    .A2(_06735_),
    .ZN(_06736_)
  );
  INV_X1 _28449_ (
    .A(_06736_),
    .ZN(io_imem_req_bits_pc[8])
  );
  AND2_X1 _28450_ (
    .A1(csr_io_evec[9]),
    .A2(_10064_),
    .ZN(_06737_)
  );
  INV_X1 _28451_ (
    .A(_06737_),
    .ZN(_06738_)
  );
  MUX2_X1 _28452_ (
    .A(_08061_),
    .B(_14023_),
    .S(_08206_),
    .Z(_06739_)
  );
  INV_X1 _28453_ (
    .A(_06739_),
    .ZN(_06740_)
  );
  AND2_X1 _28454_ (
    .A1(_08686_),
    .A2(_06739_),
    .ZN(_06741_)
  );
  INV_X1 _28455_ (
    .A(_06741_),
    .ZN(_06742_)
  );
  AND2_X1 _28456_ (
    .A1(_07997_),
    .A2(_08687_),
    .ZN(_06743_)
  );
  INV_X1 _28457_ (
    .A(_06743_),
    .ZN(_06744_)
  );
  AND2_X1 _28458_ (
    .A1(_10063_),
    .A2(_06744_),
    .ZN(_06745_)
  );
  AND2_X1 _28459_ (
    .A1(_06742_),
    .A2(_06745_),
    .ZN(_06746_)
  );
  INV_X1 _28460_ (
    .A(_06746_),
    .ZN(_06747_)
  );
  AND2_X1 _28461_ (
    .A1(_06738_),
    .A2(_06747_),
    .ZN(_06748_)
  );
  INV_X1 _28462_ (
    .A(_06748_),
    .ZN(io_imem_req_bits_pc[9])
  );
  AND2_X1 _28463_ (
    .A1(csr_io_evec[10]),
    .A2(_10064_),
    .ZN(_06749_)
  );
  INV_X1 _28464_ (
    .A(_06749_),
    .ZN(_06750_)
  );
  MUX2_X1 _28465_ (
    .A(_08062_),
    .B(_01614_),
    .S(_08206_),
    .Z(_06751_)
  );
  INV_X1 _28466_ (
    .A(_06751_),
    .ZN(_06752_)
  );
  AND2_X1 _28467_ (
    .A1(_08686_),
    .A2(_06751_),
    .ZN(_06753_)
  );
  INV_X1 _28468_ (
    .A(_06753_),
    .ZN(_06754_)
  );
  AND2_X1 _28469_ (
    .A1(_07999_),
    .A2(_08687_),
    .ZN(_06755_)
  );
  INV_X1 _28470_ (
    .A(_06755_),
    .ZN(_06756_)
  );
  AND2_X1 _28471_ (
    .A1(_10063_),
    .A2(_06756_),
    .ZN(_06757_)
  );
  AND2_X1 _28472_ (
    .A1(_06754_),
    .A2(_06757_),
    .ZN(_06758_)
  );
  INV_X1 _28473_ (
    .A(_06758_),
    .ZN(_06759_)
  );
  AND2_X1 _28474_ (
    .A1(_06750_),
    .A2(_06759_),
    .ZN(_06760_)
  );
  INV_X1 _28475_ (
    .A(_06760_),
    .ZN(io_imem_req_bits_pc[10])
  );
  AND2_X1 _28476_ (
    .A1(csr_io_evec[11]),
    .A2(_10064_),
    .ZN(_06761_)
  );
  INV_X1 _28477_ (
    .A(_06761_),
    .ZN(_06762_)
  );
  MUX2_X1 _28478_ (
    .A(_08063_),
    .B(_01640_),
    .S(_08206_),
    .Z(_06763_)
  );
  INV_X1 _28479_ (
    .A(_06763_),
    .ZN(_06764_)
  );
  AND2_X1 _28480_ (
    .A1(_08686_),
    .A2(_06763_),
    .ZN(_06765_)
  );
  INV_X1 _28481_ (
    .A(_06765_),
    .ZN(_06766_)
  );
  AND2_X1 _28482_ (
    .A1(_08001_),
    .A2(_08687_),
    .ZN(_06767_)
  );
  INV_X1 _28483_ (
    .A(_06767_),
    .ZN(_06768_)
  );
  AND2_X1 _28484_ (
    .A1(_10063_),
    .A2(_06768_),
    .ZN(_06769_)
  );
  AND2_X1 _28485_ (
    .A1(_06766_),
    .A2(_06769_),
    .ZN(_06770_)
  );
  INV_X1 _28486_ (
    .A(_06770_),
    .ZN(_06771_)
  );
  AND2_X1 _28487_ (
    .A1(_06762_),
    .A2(_06771_),
    .ZN(_06772_)
  );
  INV_X1 _28488_ (
    .A(_06772_),
    .ZN(io_imem_req_bits_pc[11])
  );
  AND2_X1 _28489_ (
    .A1(csr_io_evec[12]),
    .A2(_10064_),
    .ZN(_06773_)
  );
  INV_X1 _28490_ (
    .A(_06773_),
    .ZN(_06774_)
  );
  MUX2_X1 _28491_ (
    .A(_08064_),
    .B(_01671_),
    .S(_08206_),
    .Z(_06775_)
  );
  INV_X1 _28492_ (
    .A(_06775_),
    .ZN(_06776_)
  );
  AND2_X1 _28493_ (
    .A1(_08686_),
    .A2(_06775_),
    .ZN(_06777_)
  );
  INV_X1 _28494_ (
    .A(_06777_),
    .ZN(_06778_)
  );
  AND2_X1 _28495_ (
    .A1(_08003_),
    .A2(_08687_),
    .ZN(_06779_)
  );
  INV_X1 _28496_ (
    .A(_06779_),
    .ZN(_06780_)
  );
  AND2_X1 _28497_ (
    .A1(_10063_),
    .A2(_06780_),
    .ZN(_06781_)
  );
  AND2_X1 _28498_ (
    .A1(_06778_),
    .A2(_06781_),
    .ZN(_06782_)
  );
  INV_X1 _28499_ (
    .A(_06782_),
    .ZN(_06783_)
  );
  AND2_X1 _28500_ (
    .A1(_06774_),
    .A2(_06783_),
    .ZN(_06784_)
  );
  INV_X1 _28501_ (
    .A(_06784_),
    .ZN(io_imem_req_bits_pc[12])
  );
  AND2_X1 _28502_ (
    .A1(csr_io_evec[13]),
    .A2(_10064_),
    .ZN(_06785_)
  );
  INV_X1 _28503_ (
    .A(_06785_),
    .ZN(_06786_)
  );
  MUX2_X1 _28504_ (
    .A(_08065_),
    .B(_01697_),
    .S(_08206_),
    .Z(_06787_)
  );
  INV_X1 _28505_ (
    .A(_06787_),
    .ZN(_06788_)
  );
  AND2_X1 _28506_ (
    .A1(_08686_),
    .A2(_06787_),
    .ZN(_06789_)
  );
  INV_X1 _28507_ (
    .A(_06789_),
    .ZN(_06790_)
  );
  AND2_X1 _28508_ (
    .A1(_08005_),
    .A2(_08687_),
    .ZN(_06791_)
  );
  INV_X1 _28509_ (
    .A(_06791_),
    .ZN(_06792_)
  );
  AND2_X1 _28510_ (
    .A1(_10063_),
    .A2(_06792_),
    .ZN(_06793_)
  );
  AND2_X1 _28511_ (
    .A1(_06790_),
    .A2(_06793_),
    .ZN(_06794_)
  );
  INV_X1 _28512_ (
    .A(_06794_),
    .ZN(_06795_)
  );
  AND2_X1 _28513_ (
    .A1(_06786_),
    .A2(_06795_),
    .ZN(_06796_)
  );
  INV_X1 _28514_ (
    .A(_06796_),
    .ZN(io_imem_req_bits_pc[13])
  );
  AND2_X1 _28515_ (
    .A1(csr_io_evec[14]),
    .A2(_10064_),
    .ZN(_06797_)
  );
  INV_X1 _28516_ (
    .A(_06797_),
    .ZN(_06798_)
  );
  MUX2_X1 _28517_ (
    .A(_08066_),
    .B(_01728_),
    .S(_08206_),
    .Z(_06799_)
  );
  INV_X1 _28518_ (
    .A(_06799_),
    .ZN(_06800_)
  );
  AND2_X1 _28519_ (
    .A1(_08686_),
    .A2(_06799_),
    .ZN(_06801_)
  );
  INV_X1 _28520_ (
    .A(_06801_),
    .ZN(_06802_)
  );
  AND2_X1 _28521_ (
    .A1(_08007_),
    .A2(_08687_),
    .ZN(_06803_)
  );
  INV_X1 _28522_ (
    .A(_06803_),
    .ZN(_06804_)
  );
  AND2_X1 _28523_ (
    .A1(_10063_),
    .A2(_06804_),
    .ZN(_06805_)
  );
  AND2_X1 _28524_ (
    .A1(_06802_),
    .A2(_06805_),
    .ZN(_06806_)
  );
  INV_X1 _28525_ (
    .A(_06806_),
    .ZN(_06807_)
  );
  AND2_X1 _28526_ (
    .A1(_06798_),
    .A2(_06807_),
    .ZN(_06808_)
  );
  INV_X1 _28527_ (
    .A(_06808_),
    .ZN(io_imem_req_bits_pc[14])
  );
  AND2_X1 _28528_ (
    .A1(csr_io_evec[15]),
    .A2(_10064_),
    .ZN(_06809_)
  );
  INV_X1 _28529_ (
    .A(_06809_),
    .ZN(_06810_)
  );
  MUX2_X1 _28530_ (
    .A(_08067_),
    .B(_01754_),
    .S(_08206_),
    .Z(_06811_)
  );
  INV_X1 _28531_ (
    .A(_06811_),
    .ZN(_06812_)
  );
  AND2_X1 _28532_ (
    .A1(_08686_),
    .A2(_06811_),
    .ZN(_06813_)
  );
  INV_X1 _28533_ (
    .A(_06813_),
    .ZN(_06814_)
  );
  AND2_X1 _28534_ (
    .A1(_08009_),
    .A2(_08687_),
    .ZN(_06815_)
  );
  INV_X1 _28535_ (
    .A(_06815_),
    .ZN(_06816_)
  );
  AND2_X1 _28536_ (
    .A1(_10063_),
    .A2(_06816_),
    .ZN(_06817_)
  );
  AND2_X1 _28537_ (
    .A1(_06814_),
    .A2(_06817_),
    .ZN(_06818_)
  );
  INV_X1 _28538_ (
    .A(_06818_),
    .ZN(_06819_)
  );
  AND2_X1 _28539_ (
    .A1(_06810_),
    .A2(_06819_),
    .ZN(_06820_)
  );
  INV_X1 _28540_ (
    .A(_06820_),
    .ZN(io_imem_req_bits_pc[15])
  );
  AND2_X1 _28541_ (
    .A1(csr_io_evec[16]),
    .A2(_10064_),
    .ZN(_06821_)
  );
  INV_X1 _28542_ (
    .A(_06821_),
    .ZN(_06822_)
  );
  MUX2_X1 _28543_ (
    .A(_08068_),
    .B(_01785_),
    .S(_08206_),
    .Z(_06823_)
  );
  INV_X1 _28544_ (
    .A(_06823_),
    .ZN(_06824_)
  );
  AND2_X1 _28545_ (
    .A1(_08686_),
    .A2(_06823_),
    .ZN(_06825_)
  );
  INV_X1 _28546_ (
    .A(_06825_),
    .ZN(_06826_)
  );
  AND2_X1 _28547_ (
    .A1(_08011_),
    .A2(_08687_),
    .ZN(_06827_)
  );
  INV_X1 _28548_ (
    .A(_06827_),
    .ZN(_06828_)
  );
  AND2_X1 _28549_ (
    .A1(_10063_),
    .A2(_06828_),
    .ZN(_06829_)
  );
  AND2_X1 _28550_ (
    .A1(_06826_),
    .A2(_06829_),
    .ZN(_06830_)
  );
  INV_X1 _28551_ (
    .A(_06830_),
    .ZN(_06831_)
  );
  AND2_X1 _28552_ (
    .A1(_06822_),
    .A2(_06831_),
    .ZN(_06832_)
  );
  INV_X1 _28553_ (
    .A(_06832_),
    .ZN(io_imem_req_bits_pc[16])
  );
  AND2_X1 _28554_ (
    .A1(csr_io_evec[17]),
    .A2(_10064_),
    .ZN(_06833_)
  );
  INV_X1 _28555_ (
    .A(_06833_),
    .ZN(_06834_)
  );
  MUX2_X1 _28556_ (
    .A(_08069_),
    .B(_01811_),
    .S(_08206_),
    .Z(_06835_)
  );
  INV_X1 _28557_ (
    .A(_06835_),
    .ZN(_06836_)
  );
  AND2_X1 _28558_ (
    .A1(_08686_),
    .A2(_06835_),
    .ZN(_06837_)
  );
  INV_X1 _28559_ (
    .A(_06837_),
    .ZN(_06838_)
  );
  AND2_X1 _28560_ (
    .A1(_08013_),
    .A2(_08687_),
    .ZN(_06839_)
  );
  INV_X1 _28561_ (
    .A(_06839_),
    .ZN(_06840_)
  );
  AND2_X1 _28562_ (
    .A1(_10063_),
    .A2(_06840_),
    .ZN(_06841_)
  );
  AND2_X1 _28563_ (
    .A1(_06838_),
    .A2(_06841_),
    .ZN(_06842_)
  );
  INV_X1 _28564_ (
    .A(_06842_),
    .ZN(_06843_)
  );
  AND2_X1 _28565_ (
    .A1(_06834_),
    .A2(_06843_),
    .ZN(_06844_)
  );
  INV_X1 _28566_ (
    .A(_06844_),
    .ZN(io_imem_req_bits_pc[17])
  );
  AND2_X1 _28567_ (
    .A1(csr_io_evec[18]),
    .A2(_10064_),
    .ZN(_06845_)
  );
  INV_X1 _28568_ (
    .A(_06845_),
    .ZN(_06846_)
  );
  MUX2_X1 _28569_ (
    .A(_08070_),
    .B(_01842_),
    .S(_08206_),
    .Z(_06847_)
  );
  INV_X1 _28570_ (
    .A(_06847_),
    .ZN(_06848_)
  );
  AND2_X1 _28571_ (
    .A1(_08686_),
    .A2(_06847_),
    .ZN(_06849_)
  );
  INV_X1 _28572_ (
    .A(_06849_),
    .ZN(_06850_)
  );
  AND2_X1 _28573_ (
    .A1(_08015_),
    .A2(_08687_),
    .ZN(_06851_)
  );
  INV_X1 _28574_ (
    .A(_06851_),
    .ZN(_06852_)
  );
  AND2_X1 _28575_ (
    .A1(_10063_),
    .A2(_06852_),
    .ZN(_06853_)
  );
  AND2_X1 _28576_ (
    .A1(_06850_),
    .A2(_06853_),
    .ZN(_06854_)
  );
  INV_X1 _28577_ (
    .A(_06854_),
    .ZN(_06855_)
  );
  AND2_X1 _28578_ (
    .A1(_06846_),
    .A2(_06855_),
    .ZN(_06856_)
  );
  INV_X1 _28579_ (
    .A(_06856_),
    .ZN(io_imem_req_bits_pc[18])
  );
  AND2_X1 _28580_ (
    .A1(csr_io_evec[19]),
    .A2(_10064_),
    .ZN(_06857_)
  );
  INV_X1 _28581_ (
    .A(_06857_),
    .ZN(_06858_)
  );
  MUX2_X1 _28582_ (
    .A(_08071_),
    .B(_01868_),
    .S(_08206_),
    .Z(_06859_)
  );
  INV_X1 _28583_ (
    .A(_06859_),
    .ZN(_06860_)
  );
  AND2_X1 _28584_ (
    .A1(_08686_),
    .A2(_06859_),
    .ZN(_06861_)
  );
  INV_X1 _28585_ (
    .A(_06861_),
    .ZN(_06862_)
  );
  AND2_X1 _28586_ (
    .A1(_08017_),
    .A2(_08687_),
    .ZN(_06863_)
  );
  INV_X1 _28587_ (
    .A(_06863_),
    .ZN(_06864_)
  );
  AND2_X1 _28588_ (
    .A1(_10063_),
    .A2(_06864_),
    .ZN(_06865_)
  );
  AND2_X1 _28589_ (
    .A1(_06862_),
    .A2(_06865_),
    .ZN(_06866_)
  );
  INV_X1 _28590_ (
    .A(_06866_),
    .ZN(_06867_)
  );
  AND2_X1 _28591_ (
    .A1(_06858_),
    .A2(_06867_),
    .ZN(_06868_)
  );
  INV_X1 _28592_ (
    .A(_06868_),
    .ZN(io_imem_req_bits_pc[19])
  );
  AND2_X1 _28593_ (
    .A1(csr_io_evec[20]),
    .A2(_10064_),
    .ZN(_06869_)
  );
  INV_X1 _28594_ (
    .A(_06869_),
    .ZN(_06870_)
  );
  MUX2_X1 _28595_ (
    .A(_08072_),
    .B(_01898_),
    .S(_08206_),
    .Z(_06871_)
  );
  INV_X1 _28596_ (
    .A(_06871_),
    .ZN(_06872_)
  );
  AND2_X1 _28597_ (
    .A1(_08686_),
    .A2(_06871_),
    .ZN(_06873_)
  );
  INV_X1 _28598_ (
    .A(_06873_),
    .ZN(_06874_)
  );
  AND2_X1 _28599_ (
    .A1(_08019_),
    .A2(_08687_),
    .ZN(_06875_)
  );
  INV_X1 _28600_ (
    .A(_06875_),
    .ZN(_06876_)
  );
  AND2_X1 _28601_ (
    .A1(_10063_),
    .A2(_06876_),
    .ZN(_06877_)
  );
  AND2_X1 _28602_ (
    .A1(_06874_),
    .A2(_06877_),
    .ZN(_06878_)
  );
  INV_X1 _28603_ (
    .A(_06878_),
    .ZN(_06879_)
  );
  AND2_X1 _28604_ (
    .A1(_06870_),
    .A2(_06879_),
    .ZN(_06880_)
  );
  INV_X1 _28605_ (
    .A(_06880_),
    .ZN(io_imem_req_bits_pc[20])
  );
  AND2_X1 _28606_ (
    .A1(csr_io_evec[21]),
    .A2(_10064_),
    .ZN(_06881_)
  );
  INV_X1 _28607_ (
    .A(_06881_),
    .ZN(_06882_)
  );
  MUX2_X1 _28608_ (
    .A(_08073_),
    .B(_01921_),
    .S(_08206_),
    .Z(_06883_)
  );
  INV_X1 _28609_ (
    .A(_06883_),
    .ZN(_06884_)
  );
  AND2_X1 _28610_ (
    .A1(_08686_),
    .A2(_06883_),
    .ZN(_06885_)
  );
  INV_X1 _28611_ (
    .A(_06885_),
    .ZN(_06886_)
  );
  AND2_X1 _28612_ (
    .A1(_08021_),
    .A2(_08687_),
    .ZN(_06887_)
  );
  INV_X1 _28613_ (
    .A(_06887_),
    .ZN(_06888_)
  );
  AND2_X1 _28614_ (
    .A1(_10063_),
    .A2(_06888_),
    .ZN(_06889_)
  );
  AND2_X1 _28615_ (
    .A1(_06886_),
    .A2(_06889_),
    .ZN(_06890_)
  );
  INV_X1 _28616_ (
    .A(_06890_),
    .ZN(_06891_)
  );
  AND2_X1 _28617_ (
    .A1(_06882_),
    .A2(_06891_),
    .ZN(_06892_)
  );
  INV_X1 _28618_ (
    .A(_06892_),
    .ZN(io_imem_req_bits_pc[21])
  );
  AND2_X1 _28619_ (
    .A1(csr_io_evec[22]),
    .A2(_10064_),
    .ZN(_06893_)
  );
  INV_X1 _28620_ (
    .A(_06893_),
    .ZN(_06894_)
  );
  MUX2_X1 _28621_ (
    .A(_08074_),
    .B(_01949_),
    .S(_08206_),
    .Z(_06895_)
  );
  INV_X1 _28622_ (
    .A(_06895_),
    .ZN(_06896_)
  );
  AND2_X1 _28623_ (
    .A1(_08686_),
    .A2(_06895_),
    .ZN(_06897_)
  );
  INV_X1 _28624_ (
    .A(_06897_),
    .ZN(_06898_)
  );
  AND2_X1 _28625_ (
    .A1(_08023_),
    .A2(_08687_),
    .ZN(_06899_)
  );
  INV_X1 _28626_ (
    .A(_06899_),
    .ZN(_06900_)
  );
  AND2_X1 _28627_ (
    .A1(_10063_),
    .A2(_06900_),
    .ZN(_06901_)
  );
  AND2_X1 _28628_ (
    .A1(_06898_),
    .A2(_06901_),
    .ZN(_06902_)
  );
  INV_X1 _28629_ (
    .A(_06902_),
    .ZN(_06903_)
  );
  AND2_X1 _28630_ (
    .A1(_06894_),
    .A2(_06903_),
    .ZN(_06904_)
  );
  INV_X1 _28631_ (
    .A(_06904_),
    .ZN(io_imem_req_bits_pc[22])
  );
  AND2_X1 _28632_ (
    .A1(csr_io_evec[23]),
    .A2(_10064_),
    .ZN(_06905_)
  );
  INV_X1 _28633_ (
    .A(_06905_),
    .ZN(_06906_)
  );
  MUX2_X1 _28634_ (
    .A(_08075_),
    .B(_01972_),
    .S(_08206_),
    .Z(_06907_)
  );
  INV_X1 _28635_ (
    .A(_06907_),
    .ZN(_06908_)
  );
  AND2_X1 _28636_ (
    .A1(_08686_),
    .A2(_06907_),
    .ZN(_06909_)
  );
  INV_X1 _28637_ (
    .A(_06909_),
    .ZN(_06910_)
  );
  AND2_X1 _28638_ (
    .A1(_08025_),
    .A2(_08687_),
    .ZN(_06911_)
  );
  INV_X1 _28639_ (
    .A(_06911_),
    .ZN(_06912_)
  );
  AND2_X1 _28640_ (
    .A1(_10063_),
    .A2(_06912_),
    .ZN(_06913_)
  );
  AND2_X1 _28641_ (
    .A1(_06910_),
    .A2(_06913_),
    .ZN(_06914_)
  );
  INV_X1 _28642_ (
    .A(_06914_),
    .ZN(_06915_)
  );
  AND2_X1 _28643_ (
    .A1(_06906_),
    .A2(_06915_),
    .ZN(_06916_)
  );
  INV_X1 _28644_ (
    .A(_06916_),
    .ZN(io_imem_req_bits_pc[23])
  );
  AND2_X1 _28645_ (
    .A1(csr_io_evec[24]),
    .A2(_10064_),
    .ZN(_06917_)
  );
  INV_X1 _28646_ (
    .A(_06917_),
    .ZN(_06918_)
  );
  MUX2_X1 _28647_ (
    .A(_08076_),
    .B(_02003_),
    .S(_08206_),
    .Z(_06919_)
  );
  INV_X1 _28648_ (
    .A(_06919_),
    .ZN(_06920_)
  );
  AND2_X1 _28649_ (
    .A1(_08686_),
    .A2(_06919_),
    .ZN(_06921_)
  );
  INV_X1 _28650_ (
    .A(_06921_),
    .ZN(_06922_)
  );
  AND2_X1 _28651_ (
    .A1(_08027_),
    .A2(_08687_),
    .ZN(_06923_)
  );
  INV_X1 _28652_ (
    .A(_06923_),
    .ZN(_06924_)
  );
  AND2_X1 _28653_ (
    .A1(_10063_),
    .A2(_06924_),
    .ZN(_06925_)
  );
  AND2_X1 _28654_ (
    .A1(_06922_),
    .A2(_06925_),
    .ZN(_06926_)
  );
  INV_X1 _28655_ (
    .A(_06926_),
    .ZN(_06927_)
  );
  AND2_X1 _28656_ (
    .A1(_06918_),
    .A2(_06927_),
    .ZN(_06928_)
  );
  INV_X1 _28657_ (
    .A(_06928_),
    .ZN(io_imem_req_bits_pc[24])
  );
  AND2_X1 _28658_ (
    .A1(csr_io_evec[25]),
    .A2(_10064_),
    .ZN(_06929_)
  );
  INV_X1 _28659_ (
    .A(_06929_),
    .ZN(_06930_)
  );
  MUX2_X1 _28660_ (
    .A(_08077_),
    .B(_02026_),
    .S(_08206_),
    .Z(_06931_)
  );
  INV_X1 _28661_ (
    .A(_06931_),
    .ZN(_06932_)
  );
  AND2_X1 _28662_ (
    .A1(_08686_),
    .A2(_06931_),
    .ZN(_06933_)
  );
  INV_X1 _28663_ (
    .A(_06933_),
    .ZN(_06934_)
  );
  AND2_X1 _28664_ (
    .A1(_08029_),
    .A2(_08687_),
    .ZN(_06935_)
  );
  INV_X1 _28665_ (
    .A(_06935_),
    .ZN(_06936_)
  );
  AND2_X1 _28666_ (
    .A1(_10063_),
    .A2(_06936_),
    .ZN(_06937_)
  );
  AND2_X1 _28667_ (
    .A1(_06934_),
    .A2(_06937_),
    .ZN(_06938_)
  );
  INV_X1 _28668_ (
    .A(_06938_),
    .ZN(_06939_)
  );
  AND2_X1 _28669_ (
    .A1(_06930_),
    .A2(_06939_),
    .ZN(_06940_)
  );
  INV_X1 _28670_ (
    .A(_06940_),
    .ZN(io_imem_req_bits_pc[25])
  );
  AND2_X1 _28671_ (
    .A1(csr_io_evec[26]),
    .A2(_10064_),
    .ZN(_06941_)
  );
  INV_X1 _28672_ (
    .A(_06941_),
    .ZN(_06942_)
  );
  MUX2_X1 _28673_ (
    .A(_08078_),
    .B(_02054_),
    .S(_08206_),
    .Z(_06943_)
  );
  INV_X1 _28674_ (
    .A(_06943_),
    .ZN(_06944_)
  );
  AND2_X1 _28675_ (
    .A1(_08686_),
    .A2(_06943_),
    .ZN(_06945_)
  );
  INV_X1 _28676_ (
    .A(_06945_),
    .ZN(_06946_)
  );
  AND2_X1 _28677_ (
    .A1(_08031_),
    .A2(_08687_),
    .ZN(_06947_)
  );
  INV_X1 _28678_ (
    .A(_06947_),
    .ZN(_06948_)
  );
  AND2_X1 _28679_ (
    .A1(_10063_),
    .A2(_06948_),
    .ZN(_06949_)
  );
  AND2_X1 _28680_ (
    .A1(_06946_),
    .A2(_06949_),
    .ZN(_06950_)
  );
  INV_X1 _28681_ (
    .A(_06950_),
    .ZN(_06951_)
  );
  AND2_X1 _28682_ (
    .A1(_06942_),
    .A2(_06951_),
    .ZN(_06952_)
  );
  INV_X1 _28683_ (
    .A(_06952_),
    .ZN(io_imem_req_bits_pc[26])
  );
  AND2_X1 _28684_ (
    .A1(csr_io_evec[27]),
    .A2(_10064_),
    .ZN(_06953_)
  );
  INV_X1 _28685_ (
    .A(_06953_),
    .ZN(_06954_)
  );
  MUX2_X1 _28686_ (
    .A(_08079_),
    .B(_02077_),
    .S(_08206_),
    .Z(_06955_)
  );
  INV_X1 _28687_ (
    .A(_06955_),
    .ZN(_06956_)
  );
  AND2_X1 _28688_ (
    .A1(_08686_),
    .A2(_06955_),
    .ZN(_06957_)
  );
  INV_X1 _28689_ (
    .A(_06957_),
    .ZN(_06958_)
  );
  AND2_X1 _28690_ (
    .A1(_08033_),
    .A2(_08687_),
    .ZN(_06959_)
  );
  INV_X1 _28691_ (
    .A(_06959_),
    .ZN(_06960_)
  );
  AND2_X1 _28692_ (
    .A1(_10063_),
    .A2(_06960_),
    .ZN(_06961_)
  );
  AND2_X1 _28693_ (
    .A1(_06958_),
    .A2(_06961_),
    .ZN(_06962_)
  );
  INV_X1 _28694_ (
    .A(_06962_),
    .ZN(_06963_)
  );
  AND2_X1 _28695_ (
    .A1(_06954_),
    .A2(_06963_),
    .ZN(_06964_)
  );
  INV_X1 _28696_ (
    .A(_06964_),
    .ZN(io_imem_req_bits_pc[27])
  );
  AND2_X1 _28697_ (
    .A1(csr_io_evec[28]),
    .A2(_10064_),
    .ZN(_06965_)
  );
  INV_X1 _28698_ (
    .A(_06965_),
    .ZN(_06966_)
  );
  MUX2_X1 _28699_ (
    .A(_08080_),
    .B(_02108_),
    .S(_08206_),
    .Z(_06967_)
  );
  INV_X1 _28700_ (
    .A(_06967_),
    .ZN(_06968_)
  );
  AND2_X1 _28701_ (
    .A1(_08686_),
    .A2(_06967_),
    .ZN(_06969_)
  );
  INV_X1 _28702_ (
    .A(_06969_),
    .ZN(_06970_)
  );
  AND2_X1 _28703_ (
    .A1(_08035_),
    .A2(_08687_),
    .ZN(_06971_)
  );
  INV_X1 _28704_ (
    .A(_06971_),
    .ZN(_06972_)
  );
  AND2_X1 _28705_ (
    .A1(_10063_),
    .A2(_06972_),
    .ZN(_06973_)
  );
  AND2_X1 _28706_ (
    .A1(_06970_),
    .A2(_06973_),
    .ZN(_06974_)
  );
  INV_X1 _28707_ (
    .A(_06974_),
    .ZN(_06975_)
  );
  AND2_X1 _28708_ (
    .A1(_06966_),
    .A2(_06975_),
    .ZN(_06976_)
  );
  INV_X1 _28709_ (
    .A(_06976_),
    .ZN(io_imem_req_bits_pc[28])
  );
  AND2_X1 _28710_ (
    .A1(csr_io_evec[29]),
    .A2(_10064_),
    .ZN(_06977_)
  );
  INV_X1 _28711_ (
    .A(_06977_),
    .ZN(_06978_)
  );
  MUX2_X1 _28712_ (
    .A(_08081_),
    .B(_02132_),
    .S(_08206_),
    .Z(_06979_)
  );
  INV_X1 _28713_ (
    .A(_06979_),
    .ZN(_06980_)
  );
  AND2_X1 _28714_ (
    .A1(_08686_),
    .A2(_06979_),
    .ZN(_06981_)
  );
  INV_X1 _28715_ (
    .A(_06981_),
    .ZN(_06982_)
  );
  AND2_X1 _28716_ (
    .A1(_08037_),
    .A2(_08687_),
    .ZN(_06983_)
  );
  INV_X1 _28717_ (
    .A(_06983_),
    .ZN(_06984_)
  );
  AND2_X1 _28718_ (
    .A1(_10063_),
    .A2(_06984_),
    .ZN(_06985_)
  );
  AND2_X1 _28719_ (
    .A1(_06982_),
    .A2(_06985_),
    .ZN(_06986_)
  );
  INV_X1 _28720_ (
    .A(_06986_),
    .ZN(_06987_)
  );
  AND2_X1 _28721_ (
    .A1(_06978_),
    .A2(_06987_),
    .ZN(_06988_)
  );
  INV_X1 _28722_ (
    .A(_06988_),
    .ZN(io_imem_req_bits_pc[29])
  );
  AND2_X1 _28723_ (
    .A1(csr_io_evec[30]),
    .A2(_10064_),
    .ZN(_06989_)
  );
  INV_X1 _28724_ (
    .A(_06989_),
    .ZN(_06990_)
  );
  MUX2_X1 _28725_ (
    .A(_08082_),
    .B(_02160_),
    .S(_08206_),
    .Z(_06991_)
  );
  INV_X1 _28726_ (
    .A(_06991_),
    .ZN(_06992_)
  );
  AND2_X1 _28727_ (
    .A1(_08686_),
    .A2(_06991_),
    .ZN(_06993_)
  );
  INV_X1 _28728_ (
    .A(_06993_),
    .ZN(_06994_)
  );
  AND2_X1 _28729_ (
    .A1(_08039_),
    .A2(_08687_),
    .ZN(_06995_)
  );
  INV_X1 _28730_ (
    .A(_06995_),
    .ZN(_06996_)
  );
  AND2_X1 _28731_ (
    .A1(_10063_),
    .A2(_06996_),
    .ZN(_06997_)
  );
  AND2_X1 _28732_ (
    .A1(_06994_),
    .A2(_06997_),
    .ZN(_06998_)
  );
  INV_X1 _28733_ (
    .A(_06998_),
    .ZN(_06999_)
  );
  AND2_X1 _28734_ (
    .A1(_06990_),
    .A2(_06999_),
    .ZN(_07000_)
  );
  INV_X1 _28735_ (
    .A(_07000_),
    .ZN(io_imem_req_bits_pc[30])
  );
  AND2_X1 _28736_ (
    .A1(csr_io_evec[31]),
    .A2(_10064_),
    .ZN(_07001_)
  );
  INV_X1 _28737_ (
    .A(_07001_),
    .ZN(_07002_)
  );
  MUX2_X1 _28738_ (
    .A(_08083_),
    .B(_02191_),
    .S(_08206_),
    .Z(_07003_)
  );
  MUX2_X1 _28739_ (
    .A(mem_reg_wdata[31]),
    .B(_02192_),
    .S(_08206_),
    .Z(_07004_)
  );
  AND2_X1 _28740_ (
    .A1(_08686_),
    .A2(_07003_),
    .ZN(_07005_)
  );
  INV_X1 _28741_ (
    .A(_07005_),
    .ZN(_07006_)
  );
  AND2_X1 _28742_ (
    .A1(_08041_),
    .A2(_08687_),
    .ZN(_07007_)
  );
  INV_X1 _28743_ (
    .A(_07007_),
    .ZN(_07008_)
  );
  AND2_X1 _28744_ (
    .A1(_10063_),
    .A2(_07008_),
    .ZN(_07009_)
  );
  AND2_X1 _28745_ (
    .A1(_07006_),
    .A2(_07009_),
    .ZN(_07010_)
  );
  INV_X1 _28746_ (
    .A(_07010_),
    .ZN(_07011_)
  );
  AND2_X1 _28747_ (
    .A1(_07002_),
    .A2(_07011_),
    .ZN(_07012_)
  );
  INV_X1 _28748_ (
    .A(_07012_),
    .ZN(io_imem_req_bits_pc[31])
  );
  AND2_X1 _28749_ (
    .A1(_08222_),
    .A2(wb_reg_xcpt),
    .ZN(_07013_)
  );
  INV_X1 _28750_ (
    .A(_07013_),
    .ZN(_07014_)
  );
  AND2_X1 _28751_ (
    .A1(_08679_),
    .A2(_07014_),
    .ZN(csr_io_cause[0])
  );
  AND2_X1 _28752_ (
    .A1(_08611_),
    .A2(_08682_),
    .ZN(_07015_)
  );
  INV_X1 _28753_ (
    .A(_07015_),
    .ZN(_07016_)
  );
  AND2_X1 _28754_ (
    .A1(_08676_),
    .A2(_07016_),
    .ZN(_07017_)
  );
  INV_X1 _28755_ (
    .A(_07017_),
    .ZN(_07018_)
  );
  AND2_X1 _28756_ (
    .A1(_08670_),
    .A2(_07018_),
    .ZN(_07019_)
  );
  INV_X1 _28757_ (
    .A(_07019_),
    .ZN(_07020_)
  );
  MUX2_X1 _28758_ (
    .A(wb_reg_cause[1]),
    .B(_08666_),
    .S(_08595_),
    .Z(_07021_)
  );
  INV_X1 _28759_ (
    .A(_07021_),
    .ZN(_07022_)
  );
  AND2_X1 _28760_ (
    .A1(_07020_),
    .A2(_07022_),
    .ZN(_07023_)
  );
  INV_X1 _28761_ (
    .A(_07023_),
    .ZN(csr_io_cause[1])
  );
  AND2_X1 _28762_ (
    .A1(_08224_),
    .A2(wb_reg_xcpt),
    .ZN(_07024_)
  );
  INV_X1 _28763_ (
    .A(_07024_),
    .ZN(csr_io_cause[2])
  );
  AND2_X1 _28764_ (
    .A1(_08225_),
    .A2(wb_reg_xcpt),
    .ZN(_07025_)
  );
  INV_X1 _28765_ (
    .A(_07025_),
    .ZN(_07026_)
  );
  AND2_X1 _28766_ (
    .A1(_08672_),
    .A2(_07026_),
    .ZN(csr_io_cause[3])
  );
  AND2_X1 _28767_ (
    .A1(wb_reg_cause[4]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[4])
  );
  AND2_X1 _28768_ (
    .A1(wb_reg_cause[5]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[5])
  );
  AND2_X1 _28769_ (
    .A1(wb_reg_cause[6]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[6])
  );
  AND2_X1 _28770_ (
    .A1(wb_reg_cause[7]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[7])
  );
  AND2_X1 _28771_ (
    .A1(wb_reg_cause[8]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[8])
  );
  AND2_X1 _28772_ (
    .A1(wb_reg_cause[9]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[9])
  );
  AND2_X1 _28773_ (
    .A1(wb_reg_cause[10]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[10])
  );
  AND2_X1 _28774_ (
    .A1(wb_reg_cause[11]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[11])
  );
  AND2_X1 _28775_ (
    .A1(wb_reg_cause[12]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[12])
  );
  AND2_X1 _28776_ (
    .A1(wb_reg_cause[13]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[13])
  );
  AND2_X1 _28777_ (
    .A1(wb_reg_cause[14]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[14])
  );
  AND2_X1 _28778_ (
    .A1(wb_reg_cause[15]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[15])
  );
  AND2_X1 _28779_ (
    .A1(wb_reg_cause[16]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[16])
  );
  AND2_X1 _28780_ (
    .A1(wb_reg_cause[17]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[17])
  );
  AND2_X1 _28781_ (
    .A1(wb_reg_cause[18]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[18])
  );
  AND2_X1 _28782_ (
    .A1(wb_reg_cause[19]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[19])
  );
  AND2_X1 _28783_ (
    .A1(wb_reg_cause[20]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[20])
  );
  AND2_X1 _28784_ (
    .A1(wb_reg_cause[21]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[21])
  );
  AND2_X1 _28785_ (
    .A1(wb_reg_cause[22]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[22])
  );
  AND2_X1 _28786_ (
    .A1(wb_reg_cause[23]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[23])
  );
  AND2_X1 _28787_ (
    .A1(wb_reg_cause[24]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[24])
  );
  AND2_X1 _28788_ (
    .A1(wb_reg_cause[25]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[25])
  );
  AND2_X1 _28789_ (
    .A1(wb_reg_cause[26]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[26])
  );
  AND2_X1 _28790_ (
    .A1(wb_reg_cause[27]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[27])
  );
  AND2_X1 _28791_ (
    .A1(wb_reg_cause[28]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[28])
  );
  AND2_X1 _28792_ (
    .A1(wb_reg_cause[29]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[29])
  );
  AND2_X1 _28793_ (
    .A1(wb_reg_cause[30]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[30])
  );
  AND2_X1 _28794_ (
    .A1(wb_reg_cause[31]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[31])
  );
  AND2_X1 _28795_ (
    .A1(_07957_),
    .A2(_08224_),
    .ZN(_07027_)
  );
  AND2_X1 _28796_ (
    .A1(_08225_),
    .A2(_07027_),
    .ZN(_07028_)
  );
  AND2_X1 _28797_ (
    .A1(_08559_),
    .A2(_07028_),
    .ZN(_07029_)
  );
  INV_X1 _28798_ (
    .A(_07029_),
    .ZN(_07030_)
  );
  AND2_X1 _28799_ (
    .A1(_08225_),
    .A2(_08562_),
    .ZN(_07031_)
  );
  INV_X1 _28800_ (
    .A(_07031_),
    .ZN(_07032_)
  );
  AND2_X1 _28801_ (
    .A1(_07957_),
    .A2(_08561_),
    .ZN(_07033_)
  );
  INV_X1 _28802_ (
    .A(_07033_),
    .ZN(_07034_)
  );
  AND2_X1 _28803_ (
    .A1(_07032_),
    .A2(_07034_),
    .ZN(_07035_)
  );
  INV_X1 _28804_ (
    .A(_07035_),
    .ZN(_07036_)
  );
  AND2_X1 _28805_ (
    .A1(_08223_),
    .A2(_08560_),
    .ZN(_07037_)
  );
  AND2_X1 _28806_ (
    .A1(_07036_),
    .A2(_07037_),
    .ZN(_07038_)
  );
  INV_X1 _28807_ (
    .A(_07038_),
    .ZN(_07039_)
  );
  AND2_X1 _28808_ (
    .A1(_07030_),
    .A2(_07039_),
    .ZN(_07040_)
  );
  INV_X1 _28809_ (
    .A(_07040_),
    .ZN(_07041_)
  );
  AND2_X1 _28810_ (
    .A1(_08222_),
    .A2(_07041_),
    .ZN(_07042_)
  );
  INV_X1 _28811_ (
    .A(_07042_),
    .ZN(_07043_)
  );
  AND2_X1 _28812_ (
    .A1(wb_reg_cause[1]),
    .A2(_00015_),
    .ZN(_07044_)
  );
  INV_X1 _28813_ (
    .A(_07044_),
    .ZN(_07045_)
  );
  AND2_X1 _28814_ (
    .A1(_08558_),
    .A2(_07045_),
    .ZN(_07046_)
  );
  AND2_X1 _28815_ (
    .A1(_07028_),
    .A2(_07046_),
    .ZN(_07047_)
  );
  INV_X1 _28816_ (
    .A(_07047_),
    .ZN(_07048_)
  );
  AND2_X1 _28817_ (
    .A1(_07043_),
    .A2(_07048_),
    .ZN(_07049_)
  );
  INV_X1 _28818_ (
    .A(_07049_),
    .ZN(_07050_)
  );
  AND2_X1 _28819_ (
    .A1(_07982_),
    .A2(_07983_),
    .ZN(_07051_)
  );
  AND2_X1 _28820_ (
    .A1(_07984_),
    .A2(_07051_),
    .ZN(_07052_)
  );
  AND2_X1 _28821_ (
    .A1(_07978_),
    .A2(_07979_),
    .ZN(_07053_)
  );
  AND2_X1 _28822_ (
    .A1(_07980_),
    .A2(_07981_),
    .ZN(_07054_)
  );
  AND2_X1 _28823_ (
    .A1(_07053_),
    .A2(_07054_),
    .ZN(_07055_)
  );
  AND2_X1 _28824_ (
    .A1(_07974_),
    .A2(_07975_),
    .ZN(_07056_)
  );
  AND2_X1 _28825_ (
    .A1(_07976_),
    .A2(_07977_),
    .ZN(_07057_)
  );
  AND2_X1 _28826_ (
    .A1(_07056_),
    .A2(_07057_),
    .ZN(_07058_)
  );
  AND2_X1 _28827_ (
    .A1(_07055_),
    .A2(_07058_),
    .ZN(_07059_)
  );
  AND2_X1 _28828_ (
    .A1(_07052_),
    .A2(_07059_),
    .ZN(_07060_)
  );
  AND2_X1 _28829_ (
    .A1(_07972_),
    .A2(_07973_),
    .ZN(_07061_)
  );
  AND2_X1 _28830_ (
    .A1(_07970_),
    .A2(_07971_),
    .ZN(_07062_)
  );
  AND2_X1 _28831_ (
    .A1(_07061_),
    .A2(_07062_),
    .ZN(_07063_)
  );
  AND2_X1 _28832_ (
    .A1(_07966_),
    .A2(_07967_),
    .ZN(_07064_)
  );
  AND2_X1 _28833_ (
    .A1(_07968_),
    .A2(_07969_),
    .ZN(_07065_)
  );
  AND2_X1 _28834_ (
    .A1(_07064_),
    .A2(_07065_),
    .ZN(_07066_)
  );
  AND2_X1 _28835_ (
    .A1(_07063_),
    .A2(_07066_),
    .ZN(_07067_)
  );
  AND2_X1 _28836_ (
    .A1(_07964_),
    .A2(_07965_),
    .ZN(_07068_)
  );
  AND2_X1 _28837_ (
    .A1(_07962_),
    .A2(_07963_),
    .ZN(_07069_)
  );
  AND2_X1 _28838_ (
    .A1(_07068_),
    .A2(_07069_),
    .ZN(_07070_)
  );
  AND2_X1 _28839_ (
    .A1(_07958_),
    .A2(_07959_),
    .ZN(_07071_)
  );
  AND2_X1 _28840_ (
    .A1(_07960_),
    .A2(_07961_),
    .ZN(_07072_)
  );
  AND2_X1 _28841_ (
    .A1(_07071_),
    .A2(_07072_),
    .ZN(_07073_)
  );
  AND2_X1 _28842_ (
    .A1(_07070_),
    .A2(_07073_),
    .ZN(_07074_)
  );
  AND2_X1 _28843_ (
    .A1(_07067_),
    .A2(_07074_),
    .ZN(_07075_)
  );
  AND2_X1 _28844_ (
    .A1(_07060_),
    .A2(_07075_),
    .ZN(_07076_)
  );
  AND2_X1 _28845_ (
    .A1(_07050_),
    .A2(_07076_),
    .ZN(_07077_)
  );
  INV_X1 _28846_ (
    .A(_07077_),
    .ZN(_07078_)
  );
  AND2_X1 _28847_ (
    .A1(_08627_),
    .A2(_07078_),
    .ZN(_07079_)
  );
  INV_X1 _28848_ (
    .A(_07079_),
    .ZN(_07080_)
  );
  AND2_X1 _28849_ (
    .A1(csr_io_exception),
    .A2(_07080_),
    .ZN(_07081_)
  );
  AND2_X1 _28850_ (
    .A1(wb_reg_wdata[0]),
    .A2(_07081_),
    .ZN(csr_io_tval[0])
  );
  AND2_X1 _28851_ (
    .A1(wb_reg_wdata[1]),
    .A2(_07081_),
    .ZN(csr_io_tval[1])
  );
  AND2_X1 _28852_ (
    .A1(wb_reg_wdata[2]),
    .A2(_07081_),
    .ZN(csr_io_tval[2])
  );
  AND2_X1 _28853_ (
    .A1(wb_reg_wdata[3]),
    .A2(_07081_),
    .ZN(csr_io_tval[3])
  );
  AND2_X1 _28854_ (
    .A1(wb_reg_wdata[4]),
    .A2(_07081_),
    .ZN(csr_io_tval[4])
  );
  AND2_X1 _28855_ (
    .A1(wb_reg_wdata[5]),
    .A2(_07081_),
    .ZN(csr_io_tval[5])
  );
  AND2_X1 _28856_ (
    .A1(wb_reg_wdata[6]),
    .A2(_07081_),
    .ZN(csr_io_tval[6])
  );
  AND2_X1 _28857_ (
    .A1(wb_reg_wdata[7]),
    .A2(_07081_),
    .ZN(csr_io_tval[7])
  );
  AND2_X1 _28858_ (
    .A1(wb_reg_wdata[8]),
    .A2(_07081_),
    .ZN(csr_io_tval[8])
  );
  AND2_X1 _28859_ (
    .A1(wb_reg_wdata[9]),
    .A2(_07081_),
    .ZN(csr_io_tval[9])
  );
  AND2_X1 _28860_ (
    .A1(wb_reg_wdata[10]),
    .A2(_07081_),
    .ZN(csr_io_tval[10])
  );
  AND2_X1 _28861_ (
    .A1(wb_reg_wdata[11]),
    .A2(_07081_),
    .ZN(csr_io_tval[11])
  );
  AND2_X1 _28862_ (
    .A1(wb_reg_wdata[12]),
    .A2(_07081_),
    .ZN(csr_io_tval[12])
  );
  AND2_X1 _28863_ (
    .A1(wb_reg_wdata[13]),
    .A2(_07081_),
    .ZN(csr_io_tval[13])
  );
  AND2_X1 _28864_ (
    .A1(wb_reg_wdata[14]),
    .A2(_07081_),
    .ZN(csr_io_tval[14])
  );
  AND2_X1 _28865_ (
    .A1(wb_reg_wdata[15]),
    .A2(_07081_),
    .ZN(csr_io_tval[15])
  );
  AND2_X1 _28866_ (
    .A1(wb_reg_wdata[16]),
    .A2(_07081_),
    .ZN(csr_io_tval[16])
  );
  AND2_X1 _28867_ (
    .A1(wb_reg_wdata[17]),
    .A2(_07081_),
    .ZN(csr_io_tval[17])
  );
  AND2_X1 _28868_ (
    .A1(wb_reg_wdata[18]),
    .A2(_07081_),
    .ZN(csr_io_tval[18])
  );
  AND2_X1 _28869_ (
    .A1(wb_reg_wdata[19]),
    .A2(_07081_),
    .ZN(csr_io_tval[19])
  );
  AND2_X1 _28870_ (
    .A1(wb_reg_wdata[20]),
    .A2(_07081_),
    .ZN(csr_io_tval[20])
  );
  AND2_X1 _28871_ (
    .A1(wb_reg_wdata[21]),
    .A2(_07081_),
    .ZN(csr_io_tval[21])
  );
  AND2_X1 _28872_ (
    .A1(wb_reg_wdata[22]),
    .A2(_07081_),
    .ZN(csr_io_tval[22])
  );
  AND2_X1 _28873_ (
    .A1(wb_reg_wdata[23]),
    .A2(_07081_),
    .ZN(csr_io_tval[23])
  );
  AND2_X1 _28874_ (
    .A1(wb_reg_wdata[24]),
    .A2(_07081_),
    .ZN(csr_io_tval[24])
  );
  AND2_X1 _28875_ (
    .A1(wb_reg_wdata[25]),
    .A2(_07081_),
    .ZN(csr_io_tval[25])
  );
  AND2_X1 _28876_ (
    .A1(wb_reg_wdata[26]),
    .A2(_07081_),
    .ZN(csr_io_tval[26])
  );
  AND2_X1 _28877_ (
    .A1(wb_reg_wdata[27]),
    .A2(_07081_),
    .ZN(csr_io_tval[27])
  );
  AND2_X1 _28878_ (
    .A1(wb_reg_wdata[28]),
    .A2(_07081_),
    .ZN(csr_io_tval[28])
  );
  AND2_X1 _28879_ (
    .A1(wb_reg_wdata[29]),
    .A2(_07081_),
    .ZN(csr_io_tval[29])
  );
  AND2_X1 _28880_ (
    .A1(wb_reg_wdata[30]),
    .A2(_07081_),
    .ZN(csr_io_tval[30])
  );
  AND2_X1 _28881_ (
    .A1(wb_reg_wdata[31]),
    .A2(_07081_),
    .ZN(csr_io_tval[31])
  );
  AND2_X1 _28882_ (
    .A1(_08251_),
    .A2(_08539_),
    .ZN(_07082_)
  );
  INV_X1 _28883_ (
    .A(_07082_),
    .ZN(_07083_)
  );
  AND2_X1 _28884_ (
    .A1(_08219_),
    .A2(_08538_),
    .ZN(_07084_)
  );
  AND2_X1 _28885_ (
    .A1(_00018_),
    .A2(_07084_),
    .ZN(_07085_)
  );
  AND2_X1 _28886_ (
    .A1(_ex_op2_T[0]),
    .A2(_07085_),
    .ZN(_07086_)
  );
  INV_X1 _28887_ (
    .A(_07086_),
    .ZN(_07087_)
  );
  AND2_X1 _28888_ (
    .A1(_08538_),
    .A2(_08539_),
    .ZN(_07088_)
  );
  AND2_X1 _28889_ (
    .A1(_08214_),
    .A2(_08215_),
    .ZN(_07089_)
  );
  INV_X1 _28890_ (
    .A(_07089_),
    .ZN(_07090_)
  );
  AND2_X1 _28891_ (
    .A1(_08216_),
    .A2(_07089_),
    .ZN(_07091_)
  );
  INV_X1 _28892_ (
    .A(_07091_),
    .ZN(_07092_)
  );
  AND2_X1 _28893_ (
    .A1(_08215_),
    .A2(_08534_),
    .ZN(_07093_)
  );
  AND2_X1 _28894_ (
    .A1(_08536_),
    .A2(_07093_),
    .ZN(_07094_)
  );
  INV_X1 _28895_ (
    .A(_07094_),
    .ZN(_07095_)
  );
  AND2_X1 _28896_ (
    .A1(ex_reg_inst[15]),
    .A2(_07090_),
    .ZN(_07096_)
  );
  AND2_X1 _28897_ (
    .A1(_07094_),
    .A2(_07096_),
    .ZN(_07097_)
  );
  INV_X1 _28898_ (
    .A(_07097_),
    .ZN(_07098_)
  );
  AND2_X1 _28899_ (
    .A1(ex_reg_inst[20]),
    .A2(_08536_),
    .ZN(_07099_)
  );
  AND2_X1 _28900_ (
    .A1(_07089_),
    .A2(_07099_),
    .ZN(_07100_)
  );
  INV_X1 _28901_ (
    .A(_07100_),
    .ZN(_07101_)
  );
  AND2_X1 _28902_ (
    .A1(_07098_),
    .A2(_07101_),
    .ZN(_07102_)
  );
  INV_X1 _28903_ (
    .A(_07102_),
    .ZN(_07103_)
  );
  MUX2_X1 _28904_ (
    .A(ex_reg_inst[7]),
    .B(_07103_),
    .S(_07092_),
    .Z(_07104_)
  );
  AND2_X1 _28905_ (
    .A1(_07088_),
    .A2(_07104_),
    .ZN(_07105_)
  );
  INV_X1 _28906_ (
    .A(_07105_),
    .ZN(_07106_)
  );
  AND2_X1 _28907_ (
    .A1(_07087_),
    .A2(_07106_),
    .ZN(_07107_)
  );
  INV_X1 _28908_ (
    .A(_07107_),
    .ZN(_07108_)
  );
  AND2_X1 _28909_ (
    .A1(_07083_),
    .A2(_07108_),
    .ZN(alu_io_in2[0])
  );
  AND2_X1 _28910_ (
    .A1(_ex_op2_T[1]),
    .A2(_07085_),
    .ZN(_07109_)
  );
  INV_X1 _28911_ (
    .A(_07109_),
    .ZN(_07110_)
  );
  AND2_X1 _28912_ (
    .A1(_08216_),
    .A2(_08535_),
    .ZN(_07111_)
  );
  AND2_X1 _28913_ (
    .A1(_08214_),
    .A2(_07111_),
    .ZN(_07112_)
  );
  INV_X1 _28914_ (
    .A(_07112_),
    .ZN(_07113_)
  );
  AND2_X1 _28915_ (
    .A1(_07088_),
    .A2(_07113_),
    .ZN(_07114_)
  );
  AND2_X1 _28916_ (
    .A1(_08216_),
    .A2(_07093_),
    .ZN(_07115_)
  );
  INV_X1 _28917_ (
    .A(_07115_),
    .ZN(_07116_)
  );
  AND2_X1 _28918_ (
    .A1(_07092_),
    .A2(_07116_),
    .ZN(_07117_)
  );
  INV_X1 _28919_ (
    .A(_07117_),
    .ZN(_07118_)
  );
  MUX2_X1 _28920_ (
    .A(ex_reg_inst[21]),
    .B(ex_reg_inst[16]),
    .S(_07094_),
    .Z(_07119_)
  );
  MUX2_X1 _28921_ (
    .A(ex_reg_inst[8]),
    .B(_07119_),
    .S(_07117_),
    .Z(_07120_)
  );
  AND2_X1 _28922_ (
    .A1(_07114_),
    .A2(_07120_),
    .ZN(_07121_)
  );
  INV_X1 _28923_ (
    .A(_07121_),
    .ZN(_07122_)
  );
  AND2_X1 _28924_ (
    .A1(_07110_),
    .A2(_07122_),
    .ZN(_07123_)
  );
  INV_X1 _28925_ (
    .A(_07123_),
    .ZN(_07124_)
  );
  MUX2_X1 _28926_ (
    .A(ex_reg_rvc),
    .B(_07124_),
    .S(_07083_),
    .Z(alu_io_in2[1])
  );
  AND2_X1 _28927_ (
    .A1(_ex_op2_T[2]),
    .A2(_07085_),
    .ZN(_07125_)
  );
  INV_X1 _28928_ (
    .A(_07125_),
    .ZN(_07126_)
  );
  MUX2_X1 _28929_ (
    .A(ex_reg_inst[22]),
    .B(ex_reg_inst[17]),
    .S(_07094_),
    .Z(_07127_)
  );
  MUX2_X1 _28930_ (
    .A(ex_reg_inst[9]),
    .B(_07127_),
    .S(_07117_),
    .Z(_07128_)
  );
  AND2_X1 _28931_ (
    .A1(_07114_),
    .A2(_07128_),
    .ZN(_07129_)
  );
  INV_X1 _28932_ (
    .A(_07129_),
    .ZN(_07130_)
  );
  AND2_X1 _28933_ (
    .A1(_07126_),
    .A2(_07130_),
    .ZN(_07131_)
  );
  INV_X1 _28934_ (
    .A(_07131_),
    .ZN(_07132_)
  );
  MUX2_X1 _28935_ (
    .A(_ex_op2_T_1[2]),
    .B(_07132_),
    .S(_07083_),
    .Z(alu_io_in2[2])
  );
  AND2_X1 _28936_ (
    .A1(_ex_op2_T[3]),
    .A2(_07085_),
    .ZN(_07133_)
  );
  INV_X1 _28937_ (
    .A(_07133_),
    .ZN(_07134_)
  );
  MUX2_X1 _28938_ (
    .A(ex_reg_inst[23]),
    .B(ex_reg_inst[18]),
    .S(_07094_),
    .Z(_07135_)
  );
  MUX2_X1 _28939_ (
    .A(ex_reg_inst[10]),
    .B(_07135_),
    .S(_07117_),
    .Z(_07136_)
  );
  AND2_X1 _28940_ (
    .A1(_07114_),
    .A2(_07136_),
    .ZN(_07137_)
  );
  INV_X1 _28941_ (
    .A(_07137_),
    .ZN(_07138_)
  );
  AND2_X1 _28942_ (
    .A1(_07134_),
    .A2(_07138_),
    .ZN(_07139_)
  );
  INV_X1 _28943_ (
    .A(_07139_),
    .ZN(_07140_)
  );
  AND2_X1 _28944_ (
    .A1(_07083_),
    .A2(_07140_),
    .ZN(alu_io_in2[3])
  );
  AND2_X1 _28945_ (
    .A1(_ex_op2_T[4]),
    .A2(_07085_),
    .ZN(_07141_)
  );
  INV_X1 _28946_ (
    .A(_07141_),
    .ZN(_07142_)
  );
  MUX2_X1 _28947_ (
    .A(ex_reg_inst[24]),
    .B(ex_reg_inst[19]),
    .S(_07094_),
    .Z(_07143_)
  );
  INV_X1 _28948_ (
    .A(_07143_),
    .ZN(_07144_)
  );
  AND2_X1 _28949_ (
    .A1(_07117_),
    .A2(_07144_),
    .ZN(_07145_)
  );
  INV_X1 _28950_ (
    .A(_07145_),
    .ZN(_07146_)
  );
  AND2_X1 _28951_ (
    .A1(_08093_),
    .A2(_07118_),
    .ZN(_07147_)
  );
  INV_X1 _28952_ (
    .A(_07147_),
    .ZN(_07148_)
  );
  AND2_X1 _28953_ (
    .A1(_07114_),
    .A2(_07148_),
    .ZN(_07149_)
  );
  AND2_X1 _28954_ (
    .A1(_07146_),
    .A2(_07149_),
    .ZN(_07150_)
  );
  INV_X1 _28955_ (
    .A(_07150_),
    .ZN(_07151_)
  );
  AND2_X1 _28956_ (
    .A1(_07142_),
    .A2(_07151_),
    .ZN(_07152_)
  );
  INV_X1 _28957_ (
    .A(_07152_),
    .ZN(_07153_)
  );
  AND2_X1 _28958_ (
    .A1(_07083_),
    .A2(_07153_),
    .ZN(alu_io_in2[4])
  );
  AND2_X1 _28959_ (
    .A1(_07095_),
    .A2(_07114_),
    .ZN(_07154_)
  );
  AND2_X1 _28960_ (
    .A1(ex_reg_inst[25]),
    .A2(_07154_),
    .ZN(_07155_)
  );
  INV_X1 _28961_ (
    .A(_07155_),
    .ZN(_07156_)
  );
  AND2_X1 _28962_ (
    .A1(_ex_op2_T[5]),
    .A2(_07085_),
    .ZN(_07157_)
  );
  INV_X1 _28963_ (
    .A(_07157_),
    .ZN(_07158_)
  );
  AND2_X1 _28964_ (
    .A1(_07156_),
    .A2(_07158_),
    .ZN(_07159_)
  );
  INV_X1 _28965_ (
    .A(_07159_),
    .ZN(_07160_)
  );
  AND2_X1 _28966_ (
    .A1(_07083_),
    .A2(_07160_),
    .ZN(alu_io_in2[5])
  );
  AND2_X1 _28967_ (
    .A1(ex_reg_inst[26]),
    .A2(_07154_),
    .ZN(_07161_)
  );
  INV_X1 _28968_ (
    .A(_07161_),
    .ZN(_07162_)
  );
  AND2_X1 _28969_ (
    .A1(_ex_op2_T[6]),
    .A2(_07085_),
    .ZN(_07163_)
  );
  INV_X1 _28970_ (
    .A(_07163_),
    .ZN(_07164_)
  );
  AND2_X1 _28971_ (
    .A1(_07162_),
    .A2(_07164_),
    .ZN(_07165_)
  );
  INV_X1 _28972_ (
    .A(_07165_),
    .ZN(_07166_)
  );
  AND2_X1 _28973_ (
    .A1(_07083_),
    .A2(_07166_),
    .ZN(alu_io_in2[6])
  );
  AND2_X1 _28974_ (
    .A1(ex_reg_inst[27]),
    .A2(_07154_),
    .ZN(_07167_)
  );
  INV_X1 _28975_ (
    .A(_07167_),
    .ZN(_07168_)
  );
  AND2_X1 _28976_ (
    .A1(_ex_op2_T[7]),
    .A2(_07085_),
    .ZN(_07169_)
  );
  INV_X1 _28977_ (
    .A(_07169_),
    .ZN(_07170_)
  );
  AND2_X1 _28978_ (
    .A1(_07168_),
    .A2(_07170_),
    .ZN(_07171_)
  );
  INV_X1 _28979_ (
    .A(_07171_),
    .ZN(_07172_)
  );
  AND2_X1 _28980_ (
    .A1(_07083_),
    .A2(_07172_),
    .ZN(alu_io_in2[7])
  );
  AND2_X1 _28981_ (
    .A1(ex_reg_inst[28]),
    .A2(_07154_),
    .ZN(_07173_)
  );
  INV_X1 _28982_ (
    .A(_07173_),
    .ZN(_07174_)
  );
  AND2_X1 _28983_ (
    .A1(_ex_op2_T[8]),
    .A2(_07085_),
    .ZN(_07175_)
  );
  INV_X1 _28984_ (
    .A(_07175_),
    .ZN(_07176_)
  );
  AND2_X1 _28985_ (
    .A1(_07174_),
    .A2(_07176_),
    .ZN(_07177_)
  );
  INV_X1 _28986_ (
    .A(_07177_),
    .ZN(_07178_)
  );
  AND2_X1 _28987_ (
    .A1(_07083_),
    .A2(_07178_),
    .ZN(alu_io_in2[8])
  );
  AND2_X1 _28988_ (
    .A1(ex_reg_inst[29]),
    .A2(_07154_),
    .ZN(_07179_)
  );
  INV_X1 _28989_ (
    .A(_07179_),
    .ZN(_07180_)
  );
  AND2_X1 _28990_ (
    .A1(_ex_op2_T[9]),
    .A2(_07085_),
    .ZN(_07181_)
  );
  INV_X1 _28991_ (
    .A(_07181_),
    .ZN(_07182_)
  );
  AND2_X1 _28992_ (
    .A1(_07180_),
    .A2(_07182_),
    .ZN(_07183_)
  );
  INV_X1 _28993_ (
    .A(_07183_),
    .ZN(_07184_)
  );
  AND2_X1 _28994_ (
    .A1(_07083_),
    .A2(_07184_),
    .ZN(alu_io_in2[9])
  );
  AND2_X1 _28995_ (
    .A1(ex_reg_inst[30]),
    .A2(_07154_),
    .ZN(_07185_)
  );
  INV_X1 _28996_ (
    .A(_07185_),
    .ZN(_07186_)
  );
  AND2_X1 _28997_ (
    .A1(_ex_op2_T[10]),
    .A2(_07085_),
    .ZN(_07187_)
  );
  INV_X1 _28998_ (
    .A(_07187_),
    .ZN(_07188_)
  );
  AND2_X1 _28999_ (
    .A1(_07186_),
    .A2(_07188_),
    .ZN(_07189_)
  );
  INV_X1 _29000_ (
    .A(_07189_),
    .ZN(_07190_)
  );
  AND2_X1 _29001_ (
    .A1(_07083_),
    .A2(_07190_),
    .ZN(alu_io_in2[10])
  );
  AND2_X1 _29002_ (
    .A1(_ex_op2_T[11]),
    .A2(_07085_),
    .ZN(_07191_)
  );
  INV_X1 _29003_ (
    .A(_07191_),
    .ZN(_07192_)
  );
  AND2_X1 _29004_ (
    .A1(_08534_),
    .A2(_07111_),
    .ZN(_07193_)
  );
  INV_X1 _29005_ (
    .A(_07193_),
    .ZN(_07194_)
  );
  AND2_X1 _29006_ (
    .A1(ex_reg_inst[31]),
    .A2(_07095_),
    .ZN(_07195_)
  );
  MUX2_X1 _29007_ (
    .A(ex_reg_inst[7]),
    .B(_07195_),
    .S(_07116_),
    .Z(_07196_)
  );
  INV_X1 _29008_ (
    .A(_07196_),
    .ZN(_07197_)
  );
  AND2_X1 _29009_ (
    .A1(_07194_),
    .A2(_07197_),
    .ZN(_07198_)
  );
  INV_X1 _29010_ (
    .A(_07198_),
    .ZN(_07199_)
  );
  AND2_X1 _29011_ (
    .A1(_08094_),
    .A2(_07193_),
    .ZN(_07200_)
  );
  INV_X1 _29012_ (
    .A(_07200_),
    .ZN(_07201_)
  );
  AND2_X1 _29013_ (
    .A1(_07154_),
    .A2(_07201_),
    .ZN(_07202_)
  );
  AND2_X1 _29014_ (
    .A1(_07199_),
    .A2(_07202_),
    .ZN(_07203_)
  );
  INV_X1 _29015_ (
    .A(_07203_),
    .ZN(_07204_)
  );
  AND2_X1 _29016_ (
    .A1(_07192_),
    .A2(_07204_),
    .ZN(_07205_)
  );
  INV_X1 _29017_ (
    .A(_07205_),
    .ZN(_07206_)
  );
  AND2_X1 _29018_ (
    .A1(_07083_),
    .A2(_07206_),
    .ZN(alu_io_in2[11])
  );
  AND2_X1 _29019_ (
    .A1(_07113_),
    .A2(_07194_),
    .ZN(_07207_)
  );
  MUX2_X1 _29020_ (
    .A(ex_reg_inst[12]),
    .B(_07195_),
    .S(_07207_),
    .Z(_07208_)
  );
  AND2_X1 _29021_ (
    .A1(_07088_),
    .A2(_07208_),
    .ZN(_07209_)
  );
  INV_X1 _29022_ (
    .A(_07209_),
    .ZN(_07210_)
  );
  AND2_X1 _29023_ (
    .A1(_ex_op2_T[12]),
    .A2(_07085_),
    .ZN(_07211_)
  );
  INV_X1 _29024_ (
    .A(_07211_),
    .ZN(_07212_)
  );
  AND2_X1 _29025_ (
    .A1(_07210_),
    .A2(_07212_),
    .ZN(_07213_)
  );
  INV_X1 _29026_ (
    .A(_07213_),
    .ZN(_07214_)
  );
  AND2_X1 _29027_ (
    .A1(_07083_),
    .A2(_07214_),
    .ZN(alu_io_in2[12])
  );
  MUX2_X1 _29028_ (
    .A(ex_reg_inst[13]),
    .B(_07195_),
    .S(_07207_),
    .Z(_07215_)
  );
  AND2_X1 _29029_ (
    .A1(_07088_),
    .A2(_07215_),
    .ZN(_07216_)
  );
  INV_X1 _29030_ (
    .A(_07216_),
    .ZN(_07217_)
  );
  AND2_X1 _29031_ (
    .A1(_ex_op2_T[13]),
    .A2(_07085_),
    .ZN(_07218_)
  );
  INV_X1 _29032_ (
    .A(_07218_),
    .ZN(_07219_)
  );
  AND2_X1 _29033_ (
    .A1(_07217_),
    .A2(_07219_),
    .ZN(_07220_)
  );
  INV_X1 _29034_ (
    .A(_07220_),
    .ZN(_07221_)
  );
  AND2_X1 _29035_ (
    .A1(_07083_),
    .A2(_07221_),
    .ZN(alu_io_in2[13])
  );
  MUX2_X1 _29036_ (
    .A(ex_reg_inst[14]),
    .B(_07195_),
    .S(_07207_),
    .Z(_07222_)
  );
  AND2_X1 _29037_ (
    .A1(_07088_),
    .A2(_07222_),
    .ZN(_07223_)
  );
  INV_X1 _29038_ (
    .A(_07223_),
    .ZN(_07224_)
  );
  AND2_X1 _29039_ (
    .A1(_ex_op2_T[14]),
    .A2(_07085_),
    .ZN(_07225_)
  );
  INV_X1 _29040_ (
    .A(_07225_),
    .ZN(_07226_)
  );
  AND2_X1 _29041_ (
    .A1(_07224_),
    .A2(_07226_),
    .ZN(_07227_)
  );
  INV_X1 _29042_ (
    .A(_07227_),
    .ZN(_07228_)
  );
  AND2_X1 _29043_ (
    .A1(_07083_),
    .A2(_07228_),
    .ZN(alu_io_in2[14])
  );
  MUX2_X1 _29044_ (
    .A(ex_reg_inst[15]),
    .B(_07195_),
    .S(_07207_),
    .Z(_07229_)
  );
  AND2_X1 _29045_ (
    .A1(_07088_),
    .A2(_07229_),
    .ZN(_07230_)
  );
  INV_X1 _29046_ (
    .A(_07230_),
    .ZN(_07231_)
  );
  AND2_X1 _29047_ (
    .A1(_ex_op2_T[15]),
    .A2(_07085_),
    .ZN(_07232_)
  );
  INV_X1 _29048_ (
    .A(_07232_),
    .ZN(_07233_)
  );
  AND2_X1 _29049_ (
    .A1(_07231_),
    .A2(_07233_),
    .ZN(_07234_)
  );
  INV_X1 _29050_ (
    .A(_07234_),
    .ZN(_07235_)
  );
  AND2_X1 _29051_ (
    .A1(_07083_),
    .A2(_07235_),
    .ZN(alu_io_in2[15])
  );
  MUX2_X1 _29052_ (
    .A(ex_reg_inst[16]),
    .B(_07195_),
    .S(_07207_),
    .Z(_07236_)
  );
  AND2_X1 _29053_ (
    .A1(_07088_),
    .A2(_07236_),
    .ZN(_07237_)
  );
  INV_X1 _29054_ (
    .A(_07237_),
    .ZN(_07238_)
  );
  AND2_X1 _29055_ (
    .A1(_ex_op2_T[16]),
    .A2(_07085_),
    .ZN(_07239_)
  );
  INV_X1 _29056_ (
    .A(_07239_),
    .ZN(_07240_)
  );
  AND2_X1 _29057_ (
    .A1(_07238_),
    .A2(_07240_),
    .ZN(_07241_)
  );
  INV_X1 _29058_ (
    .A(_07241_),
    .ZN(_07242_)
  );
  AND2_X1 _29059_ (
    .A1(_07083_),
    .A2(_07242_),
    .ZN(alu_io_in2[16])
  );
  MUX2_X1 _29060_ (
    .A(ex_reg_inst[17]),
    .B(_07195_),
    .S(_07207_),
    .Z(_07243_)
  );
  AND2_X1 _29061_ (
    .A1(_07088_),
    .A2(_07243_),
    .ZN(_07244_)
  );
  INV_X1 _29062_ (
    .A(_07244_),
    .ZN(_07245_)
  );
  AND2_X1 _29063_ (
    .A1(_ex_op2_T[17]),
    .A2(_07085_),
    .ZN(_07246_)
  );
  INV_X1 _29064_ (
    .A(_07246_),
    .ZN(_07247_)
  );
  AND2_X1 _29065_ (
    .A1(_07245_),
    .A2(_07247_),
    .ZN(_07248_)
  );
  INV_X1 _29066_ (
    .A(_07248_),
    .ZN(_07249_)
  );
  AND2_X1 _29067_ (
    .A1(_07083_),
    .A2(_07249_),
    .ZN(alu_io_in2[17])
  );
  MUX2_X1 _29068_ (
    .A(ex_reg_inst[18]),
    .B(_07195_),
    .S(_07207_),
    .Z(_07250_)
  );
  AND2_X1 _29069_ (
    .A1(_07088_),
    .A2(_07250_),
    .ZN(_07251_)
  );
  INV_X1 _29070_ (
    .A(_07251_),
    .ZN(_07252_)
  );
  AND2_X1 _29071_ (
    .A1(_ex_op2_T[18]),
    .A2(_07085_),
    .ZN(_07253_)
  );
  INV_X1 _29072_ (
    .A(_07253_),
    .ZN(_07254_)
  );
  AND2_X1 _29073_ (
    .A1(_07252_),
    .A2(_07254_),
    .ZN(_07255_)
  );
  INV_X1 _29074_ (
    .A(_07255_),
    .ZN(_07256_)
  );
  AND2_X1 _29075_ (
    .A1(_07083_),
    .A2(_07256_),
    .ZN(alu_io_in2[18])
  );
  MUX2_X1 _29076_ (
    .A(ex_reg_inst[19]),
    .B(_07195_),
    .S(_07207_),
    .Z(_07257_)
  );
  AND2_X1 _29077_ (
    .A1(_07088_),
    .A2(_07257_),
    .ZN(_07258_)
  );
  INV_X1 _29078_ (
    .A(_07258_),
    .ZN(_07259_)
  );
  AND2_X1 _29079_ (
    .A1(_ex_op2_T[19]),
    .A2(_07085_),
    .ZN(_07260_)
  );
  INV_X1 _29080_ (
    .A(_07260_),
    .ZN(_07261_)
  );
  AND2_X1 _29081_ (
    .A1(_07259_),
    .A2(_07261_),
    .ZN(_07262_)
  );
  INV_X1 _29082_ (
    .A(_07262_),
    .ZN(_07263_)
  );
  AND2_X1 _29083_ (
    .A1(_07083_),
    .A2(_07263_),
    .ZN(alu_io_in2[19])
  );
  MUX2_X1 _29084_ (
    .A(ex_reg_inst[20]),
    .B(_07195_),
    .S(_07113_),
    .Z(_07264_)
  );
  AND2_X1 _29085_ (
    .A1(_07088_),
    .A2(_07264_),
    .ZN(_07265_)
  );
  INV_X1 _29086_ (
    .A(_07265_),
    .ZN(_07266_)
  );
  AND2_X1 _29087_ (
    .A1(_ex_op2_T[20]),
    .A2(_07085_),
    .ZN(_07267_)
  );
  INV_X1 _29088_ (
    .A(_07267_),
    .ZN(_07268_)
  );
  AND2_X1 _29089_ (
    .A1(_07266_),
    .A2(_07268_),
    .ZN(_07269_)
  );
  INV_X1 _29090_ (
    .A(_07269_),
    .ZN(_07270_)
  );
  AND2_X1 _29091_ (
    .A1(_07083_),
    .A2(_07270_),
    .ZN(alu_io_in2[20])
  );
  MUX2_X1 _29092_ (
    .A(ex_reg_inst[21]),
    .B(_07195_),
    .S(_07113_),
    .Z(_07271_)
  );
  AND2_X1 _29093_ (
    .A1(_07088_),
    .A2(_07271_),
    .ZN(_07272_)
  );
  INV_X1 _29094_ (
    .A(_07272_),
    .ZN(_07273_)
  );
  AND2_X1 _29095_ (
    .A1(_ex_op2_T[21]),
    .A2(_07085_),
    .ZN(_07274_)
  );
  INV_X1 _29096_ (
    .A(_07274_),
    .ZN(_07275_)
  );
  AND2_X1 _29097_ (
    .A1(_07273_),
    .A2(_07275_),
    .ZN(_07276_)
  );
  INV_X1 _29098_ (
    .A(_07276_),
    .ZN(_07277_)
  );
  AND2_X1 _29099_ (
    .A1(_07083_),
    .A2(_07277_),
    .ZN(alu_io_in2[21])
  );
  MUX2_X1 _29100_ (
    .A(ex_reg_inst[22]),
    .B(_07195_),
    .S(_07113_),
    .Z(_07278_)
  );
  AND2_X1 _29101_ (
    .A1(_07088_),
    .A2(_07278_),
    .ZN(_07279_)
  );
  INV_X1 _29102_ (
    .A(_07279_),
    .ZN(_07280_)
  );
  AND2_X1 _29103_ (
    .A1(_ex_op2_T[22]),
    .A2(_07085_),
    .ZN(_07281_)
  );
  INV_X1 _29104_ (
    .A(_07281_),
    .ZN(_07282_)
  );
  AND2_X1 _29105_ (
    .A1(_07280_),
    .A2(_07282_),
    .ZN(_07283_)
  );
  INV_X1 _29106_ (
    .A(_07283_),
    .ZN(_07284_)
  );
  AND2_X1 _29107_ (
    .A1(_07083_),
    .A2(_07284_),
    .ZN(alu_io_in2[22])
  );
  MUX2_X1 _29108_ (
    .A(ex_reg_inst[23]),
    .B(_07195_),
    .S(_07113_),
    .Z(_07285_)
  );
  AND2_X1 _29109_ (
    .A1(_07088_),
    .A2(_07285_),
    .ZN(_07286_)
  );
  INV_X1 _29110_ (
    .A(_07286_),
    .ZN(_07287_)
  );
  AND2_X1 _29111_ (
    .A1(_ex_op2_T[23]),
    .A2(_07085_),
    .ZN(_07288_)
  );
  INV_X1 _29112_ (
    .A(_07288_),
    .ZN(_07289_)
  );
  AND2_X1 _29113_ (
    .A1(_07287_),
    .A2(_07289_),
    .ZN(_07290_)
  );
  INV_X1 _29114_ (
    .A(_07290_),
    .ZN(_07291_)
  );
  AND2_X1 _29115_ (
    .A1(_07083_),
    .A2(_07291_),
    .ZN(alu_io_in2[23])
  );
  MUX2_X1 _29116_ (
    .A(ex_reg_inst[24]),
    .B(_07195_),
    .S(_07113_),
    .Z(_07292_)
  );
  AND2_X1 _29117_ (
    .A1(_07088_),
    .A2(_07292_),
    .ZN(_07293_)
  );
  INV_X1 _29118_ (
    .A(_07293_),
    .ZN(_07294_)
  );
  AND2_X1 _29119_ (
    .A1(_ex_op2_T[24]),
    .A2(_07085_),
    .ZN(_07295_)
  );
  INV_X1 _29120_ (
    .A(_07295_),
    .ZN(_07296_)
  );
  AND2_X1 _29121_ (
    .A1(_07294_),
    .A2(_07296_),
    .ZN(_07297_)
  );
  INV_X1 _29122_ (
    .A(_07297_),
    .ZN(_07298_)
  );
  AND2_X1 _29123_ (
    .A1(_07083_),
    .A2(_07298_),
    .ZN(alu_io_in2[24])
  );
  MUX2_X1 _29124_ (
    .A(ex_reg_inst[25]),
    .B(_07195_),
    .S(_07113_),
    .Z(_07299_)
  );
  AND2_X1 _29125_ (
    .A1(_07088_),
    .A2(_07299_),
    .ZN(_07300_)
  );
  INV_X1 _29126_ (
    .A(_07300_),
    .ZN(_07301_)
  );
  AND2_X1 _29127_ (
    .A1(_ex_op2_T[25]),
    .A2(_07085_),
    .ZN(_07302_)
  );
  INV_X1 _29128_ (
    .A(_07302_),
    .ZN(_07303_)
  );
  AND2_X1 _29129_ (
    .A1(_07301_),
    .A2(_07303_),
    .ZN(_07304_)
  );
  INV_X1 _29130_ (
    .A(_07304_),
    .ZN(_07305_)
  );
  AND2_X1 _29131_ (
    .A1(_07083_),
    .A2(_07305_),
    .ZN(alu_io_in2[25])
  );
  MUX2_X1 _29132_ (
    .A(ex_reg_inst[26]),
    .B(_07195_),
    .S(_07113_),
    .Z(_07306_)
  );
  AND2_X1 _29133_ (
    .A1(_07088_),
    .A2(_07306_),
    .ZN(_07307_)
  );
  INV_X1 _29134_ (
    .A(_07307_),
    .ZN(_07308_)
  );
  AND2_X1 _29135_ (
    .A1(_ex_op2_T[26]),
    .A2(_07085_),
    .ZN(_07309_)
  );
  INV_X1 _29136_ (
    .A(_07309_),
    .ZN(_07310_)
  );
  AND2_X1 _29137_ (
    .A1(_07308_),
    .A2(_07310_),
    .ZN(_07311_)
  );
  INV_X1 _29138_ (
    .A(_07311_),
    .ZN(_07312_)
  );
  AND2_X1 _29139_ (
    .A1(_07083_),
    .A2(_07312_),
    .ZN(alu_io_in2[26])
  );
  MUX2_X1 _29140_ (
    .A(ex_reg_inst[27]),
    .B(_07195_),
    .S(_07113_),
    .Z(_07313_)
  );
  AND2_X1 _29141_ (
    .A1(_07088_),
    .A2(_07313_),
    .ZN(_07314_)
  );
  INV_X1 _29142_ (
    .A(_07314_),
    .ZN(_07315_)
  );
  AND2_X1 _29143_ (
    .A1(_ex_op2_T[27]),
    .A2(_07085_),
    .ZN(_07316_)
  );
  INV_X1 _29144_ (
    .A(_07316_),
    .ZN(_07317_)
  );
  AND2_X1 _29145_ (
    .A1(_07315_),
    .A2(_07317_),
    .ZN(_07318_)
  );
  INV_X1 _29146_ (
    .A(_07318_),
    .ZN(_07319_)
  );
  AND2_X1 _29147_ (
    .A1(_07083_),
    .A2(_07319_),
    .ZN(alu_io_in2[27])
  );
  MUX2_X1 _29148_ (
    .A(ex_reg_inst[28]),
    .B(_07195_),
    .S(_07113_),
    .Z(_07320_)
  );
  AND2_X1 _29149_ (
    .A1(_07088_),
    .A2(_07320_),
    .ZN(_07321_)
  );
  INV_X1 _29150_ (
    .A(_07321_),
    .ZN(_07322_)
  );
  AND2_X1 _29151_ (
    .A1(_ex_op2_T[28]),
    .A2(_07085_),
    .ZN(_07323_)
  );
  INV_X1 _29152_ (
    .A(_07323_),
    .ZN(_07324_)
  );
  AND2_X1 _29153_ (
    .A1(_07322_),
    .A2(_07324_),
    .ZN(_07325_)
  );
  INV_X1 _29154_ (
    .A(_07325_),
    .ZN(_07326_)
  );
  AND2_X1 _29155_ (
    .A1(_07083_),
    .A2(_07326_),
    .ZN(alu_io_in2[28])
  );
  MUX2_X1 _29156_ (
    .A(ex_reg_inst[29]),
    .B(_07195_),
    .S(_07113_),
    .Z(_07327_)
  );
  AND2_X1 _29157_ (
    .A1(_07088_),
    .A2(_07327_),
    .ZN(_07328_)
  );
  INV_X1 _29158_ (
    .A(_07328_),
    .ZN(_07329_)
  );
  AND2_X1 _29159_ (
    .A1(_ex_op2_T[29]),
    .A2(_07085_),
    .ZN(_07330_)
  );
  INV_X1 _29160_ (
    .A(_07330_),
    .ZN(_07331_)
  );
  AND2_X1 _29161_ (
    .A1(_07329_),
    .A2(_07331_),
    .ZN(_07332_)
  );
  INV_X1 _29162_ (
    .A(_07332_),
    .ZN(_07333_)
  );
  AND2_X1 _29163_ (
    .A1(_07083_),
    .A2(_07333_),
    .ZN(alu_io_in2[29])
  );
  MUX2_X1 _29164_ (
    .A(ex_reg_inst[30]),
    .B(_07195_),
    .S(_07113_),
    .Z(_07334_)
  );
  AND2_X1 _29165_ (
    .A1(_07088_),
    .A2(_07334_),
    .ZN(_07335_)
  );
  INV_X1 _29166_ (
    .A(_07335_),
    .ZN(_07336_)
  );
  AND2_X1 _29167_ (
    .A1(_ex_op2_T[30]),
    .A2(_07085_),
    .ZN(_07337_)
  );
  INV_X1 _29168_ (
    .A(_07337_),
    .ZN(_07338_)
  );
  AND2_X1 _29169_ (
    .A1(_07336_),
    .A2(_07338_),
    .ZN(_07339_)
  );
  INV_X1 _29170_ (
    .A(_07339_),
    .ZN(_07340_)
  );
  AND2_X1 _29171_ (
    .A1(_07083_),
    .A2(_07340_),
    .ZN(alu_io_in2[30])
  );
  AND2_X1 _29172_ (
    .A1(_07088_),
    .A2(_07195_),
    .ZN(_07341_)
  );
  INV_X1 _29173_ (
    .A(_07341_),
    .ZN(_07342_)
  );
  AND2_X1 _29174_ (
    .A1(_ex_op2_T[31]),
    .A2(_07085_),
    .ZN(_07343_)
  );
  INV_X1 _29175_ (
    .A(_07343_),
    .ZN(_07344_)
  );
  AND2_X1 _29176_ (
    .A1(_07342_),
    .A2(_07344_),
    .ZN(_07345_)
  );
  INV_X1 _29177_ (
    .A(_07345_),
    .ZN(_07346_)
  );
  AND2_X1 _29178_ (
    .A1(_07083_),
    .A2(_07346_),
    .ZN(alu_io_in2[31])
  );
  AND2_X1 _29179_ (
    .A1(_08217_),
    .A2(_08563_),
    .ZN(_07347_)
  );
  INV_X1 _29180_ (
    .A(_07347_),
    .ZN(_07348_)
  );
  AND2_X1 _29181_ (
    .A1(ex_reg_pc[0]),
    .A2(_07347_),
    .ZN(_07349_)
  );
  INV_X1 _29182_ (
    .A(_07349_),
    .ZN(_07350_)
  );
  AND2_X1 _29183_ (
    .A1(_08218_),
    .A2(_08537_),
    .ZN(_07351_)
  );
  AND2_X1 _29184_ (
    .A1(_07348_),
    .A2(_07351_),
    .ZN(_07352_)
  );
  AND2_X1 _29185_ (
    .A1(_ex_op1_T[0]),
    .A2(_07352_),
    .ZN(_07353_)
  );
  INV_X1 _29186_ (
    .A(_07353_),
    .ZN(_07354_)
  );
  AND2_X1 _29187_ (
    .A1(_07350_),
    .A2(_07354_),
    .ZN(_07355_)
  );
  INV_X1 _29188_ (
    .A(_07355_),
    .ZN(alu_io_in1[0])
  );
  AND2_X1 _29189_ (
    .A1(ex_reg_pc[1]),
    .A2(_07347_),
    .ZN(_07356_)
  );
  INV_X1 _29190_ (
    .A(_07356_),
    .ZN(_07357_)
  );
  AND2_X1 _29191_ (
    .A1(_ex_op1_T[1]),
    .A2(_07352_),
    .ZN(_07358_)
  );
  INV_X1 _29192_ (
    .A(_07358_),
    .ZN(_07359_)
  );
  AND2_X1 _29193_ (
    .A1(_07357_),
    .A2(_07359_),
    .ZN(_07360_)
  );
  INV_X1 _29194_ (
    .A(_07360_),
    .ZN(alu_io_in1[1])
  );
  AND2_X1 _29195_ (
    .A1(ex_reg_pc[2]),
    .A2(_07347_),
    .ZN(_07361_)
  );
  INV_X1 _29196_ (
    .A(_07361_),
    .ZN(_07362_)
  );
  AND2_X1 _29197_ (
    .A1(_ex_op1_T[2]),
    .A2(_07352_),
    .ZN(_07363_)
  );
  INV_X1 _29198_ (
    .A(_07363_),
    .ZN(_07364_)
  );
  AND2_X1 _29199_ (
    .A1(_07362_),
    .A2(_07364_),
    .ZN(_07365_)
  );
  INV_X1 _29200_ (
    .A(_07365_),
    .ZN(alu_io_in1[2])
  );
  AND2_X1 _29201_ (
    .A1(ex_reg_pc[3]),
    .A2(_07347_),
    .ZN(_07366_)
  );
  INV_X1 _29202_ (
    .A(_07366_),
    .ZN(_07367_)
  );
  AND2_X1 _29203_ (
    .A1(_ex_op1_T[3]),
    .A2(_07352_),
    .ZN(_07368_)
  );
  INV_X1 _29204_ (
    .A(_07368_),
    .ZN(_07369_)
  );
  AND2_X1 _29205_ (
    .A1(_07367_),
    .A2(_07369_),
    .ZN(_07370_)
  );
  INV_X1 _29206_ (
    .A(_07370_),
    .ZN(alu_io_in1[3])
  );
  AND2_X1 _29207_ (
    .A1(ex_reg_pc[4]),
    .A2(_07347_),
    .ZN(_07371_)
  );
  INV_X1 _29208_ (
    .A(_07371_),
    .ZN(_07372_)
  );
  AND2_X1 _29209_ (
    .A1(_ex_op1_T[4]),
    .A2(_07352_),
    .ZN(_07373_)
  );
  INV_X1 _29210_ (
    .A(_07373_),
    .ZN(_07374_)
  );
  AND2_X1 _29211_ (
    .A1(_07372_),
    .A2(_07374_),
    .ZN(_07375_)
  );
  INV_X1 _29212_ (
    .A(_07375_),
    .ZN(alu_io_in1[4])
  );
  AND2_X1 _29213_ (
    .A1(ex_reg_pc[5]),
    .A2(_07347_),
    .ZN(_07376_)
  );
  INV_X1 _29214_ (
    .A(_07376_),
    .ZN(_07377_)
  );
  AND2_X1 _29215_ (
    .A1(_ex_op1_T[5]),
    .A2(_07352_),
    .ZN(_07378_)
  );
  INV_X1 _29216_ (
    .A(_07378_),
    .ZN(_07379_)
  );
  AND2_X1 _29217_ (
    .A1(_07377_),
    .A2(_07379_),
    .ZN(_07380_)
  );
  INV_X1 _29218_ (
    .A(_07380_),
    .ZN(alu_io_in1[5])
  );
  AND2_X1 _29219_ (
    .A1(ex_reg_pc[6]),
    .A2(_07347_),
    .ZN(_07381_)
  );
  INV_X1 _29220_ (
    .A(_07381_),
    .ZN(_07382_)
  );
  AND2_X1 _29221_ (
    .A1(_ex_op1_T[6]),
    .A2(_07352_),
    .ZN(_07383_)
  );
  INV_X1 _29222_ (
    .A(_07383_),
    .ZN(_07384_)
  );
  AND2_X1 _29223_ (
    .A1(_07382_),
    .A2(_07384_),
    .ZN(_07385_)
  );
  INV_X1 _29224_ (
    .A(_07385_),
    .ZN(alu_io_in1[6])
  );
  AND2_X1 _29225_ (
    .A1(ex_reg_pc[7]),
    .A2(_07347_),
    .ZN(_07386_)
  );
  INV_X1 _29226_ (
    .A(_07386_),
    .ZN(_07387_)
  );
  AND2_X1 _29227_ (
    .A1(_ex_op1_T[7]),
    .A2(_07352_),
    .ZN(_07388_)
  );
  INV_X1 _29228_ (
    .A(_07388_),
    .ZN(_07389_)
  );
  AND2_X1 _29229_ (
    .A1(_07387_),
    .A2(_07389_),
    .ZN(_07390_)
  );
  INV_X1 _29230_ (
    .A(_07390_),
    .ZN(alu_io_in1[7])
  );
  AND2_X1 _29231_ (
    .A1(ex_reg_pc[8]),
    .A2(_07347_),
    .ZN(_07391_)
  );
  INV_X1 _29232_ (
    .A(_07391_),
    .ZN(_07392_)
  );
  AND2_X1 _29233_ (
    .A1(_ex_op1_T[8]),
    .A2(_07352_),
    .ZN(_07393_)
  );
  INV_X1 _29234_ (
    .A(_07393_),
    .ZN(_07394_)
  );
  AND2_X1 _29235_ (
    .A1(_07392_),
    .A2(_07394_),
    .ZN(_07395_)
  );
  INV_X1 _29236_ (
    .A(_07395_),
    .ZN(alu_io_in1[8])
  );
  AND2_X1 _29237_ (
    .A1(ex_reg_pc[9]),
    .A2(_07347_),
    .ZN(_07396_)
  );
  INV_X1 _29238_ (
    .A(_07396_),
    .ZN(_07397_)
  );
  AND2_X1 _29239_ (
    .A1(_ex_op1_T[9]),
    .A2(_07352_),
    .ZN(_07398_)
  );
  INV_X1 _29240_ (
    .A(_07398_),
    .ZN(_07399_)
  );
  AND2_X1 _29241_ (
    .A1(_07397_),
    .A2(_07399_),
    .ZN(_07400_)
  );
  INV_X1 _29242_ (
    .A(_07400_),
    .ZN(alu_io_in1[9])
  );
  AND2_X1 _29243_ (
    .A1(ex_reg_pc[10]),
    .A2(_07347_),
    .ZN(_07401_)
  );
  INV_X1 _29244_ (
    .A(_07401_),
    .ZN(_07402_)
  );
  AND2_X1 _29245_ (
    .A1(_ex_op1_T[10]),
    .A2(_07352_),
    .ZN(_07403_)
  );
  INV_X1 _29246_ (
    .A(_07403_),
    .ZN(_07404_)
  );
  AND2_X1 _29247_ (
    .A1(_07402_),
    .A2(_07404_),
    .ZN(_07405_)
  );
  INV_X1 _29248_ (
    .A(_07405_),
    .ZN(alu_io_in1[10])
  );
  AND2_X1 _29249_ (
    .A1(ex_reg_pc[11]),
    .A2(_07347_),
    .ZN(_07406_)
  );
  INV_X1 _29250_ (
    .A(_07406_),
    .ZN(_07407_)
  );
  AND2_X1 _29251_ (
    .A1(_ex_op1_T[11]),
    .A2(_07352_),
    .ZN(_07408_)
  );
  INV_X1 _29252_ (
    .A(_07408_),
    .ZN(_07409_)
  );
  AND2_X1 _29253_ (
    .A1(_07407_),
    .A2(_07409_),
    .ZN(_07410_)
  );
  INV_X1 _29254_ (
    .A(_07410_),
    .ZN(alu_io_in1[11])
  );
  AND2_X1 _29255_ (
    .A1(ex_reg_pc[12]),
    .A2(_07347_),
    .ZN(_07411_)
  );
  INV_X1 _29256_ (
    .A(_07411_),
    .ZN(_07412_)
  );
  AND2_X1 _29257_ (
    .A1(_ex_op1_T[12]),
    .A2(_07352_),
    .ZN(_07413_)
  );
  INV_X1 _29258_ (
    .A(_07413_),
    .ZN(_07414_)
  );
  AND2_X1 _29259_ (
    .A1(_07412_),
    .A2(_07414_),
    .ZN(_07415_)
  );
  INV_X1 _29260_ (
    .A(_07415_),
    .ZN(alu_io_in1[12])
  );
  AND2_X1 _29261_ (
    .A1(ex_reg_pc[13]),
    .A2(_07347_),
    .ZN(_07416_)
  );
  INV_X1 _29262_ (
    .A(_07416_),
    .ZN(_07417_)
  );
  AND2_X1 _29263_ (
    .A1(_ex_op1_T[13]),
    .A2(_07352_),
    .ZN(_07418_)
  );
  INV_X1 _29264_ (
    .A(_07418_),
    .ZN(_07419_)
  );
  AND2_X1 _29265_ (
    .A1(_07417_),
    .A2(_07419_),
    .ZN(_07420_)
  );
  INV_X1 _29266_ (
    .A(_07420_),
    .ZN(alu_io_in1[13])
  );
  AND2_X1 _29267_ (
    .A1(ex_reg_pc[14]),
    .A2(_07347_),
    .ZN(_07421_)
  );
  INV_X1 _29268_ (
    .A(_07421_),
    .ZN(_07422_)
  );
  AND2_X1 _29269_ (
    .A1(_ex_op1_T[14]),
    .A2(_07352_),
    .ZN(_07423_)
  );
  INV_X1 _29270_ (
    .A(_07423_),
    .ZN(_07424_)
  );
  AND2_X1 _29271_ (
    .A1(_07422_),
    .A2(_07424_),
    .ZN(_07425_)
  );
  INV_X1 _29272_ (
    .A(_07425_),
    .ZN(alu_io_in1[14])
  );
  AND2_X1 _29273_ (
    .A1(ex_reg_pc[15]),
    .A2(_07347_),
    .ZN(_07426_)
  );
  INV_X1 _29274_ (
    .A(_07426_),
    .ZN(_07427_)
  );
  AND2_X1 _29275_ (
    .A1(_ex_op1_T[15]),
    .A2(_07352_),
    .ZN(_07428_)
  );
  INV_X1 _29276_ (
    .A(_07428_),
    .ZN(_07429_)
  );
  AND2_X1 _29277_ (
    .A1(_07427_),
    .A2(_07429_),
    .ZN(_07430_)
  );
  INV_X1 _29278_ (
    .A(_07430_),
    .ZN(alu_io_in1[15])
  );
  AND2_X1 _29279_ (
    .A1(ex_reg_pc[16]),
    .A2(_07347_),
    .ZN(_07431_)
  );
  INV_X1 _29280_ (
    .A(_07431_),
    .ZN(_07432_)
  );
  AND2_X1 _29281_ (
    .A1(_ex_op1_T[16]),
    .A2(_07352_),
    .ZN(_07433_)
  );
  INV_X1 _29282_ (
    .A(_07433_),
    .ZN(_07434_)
  );
  AND2_X1 _29283_ (
    .A1(_07432_),
    .A2(_07434_),
    .ZN(_07435_)
  );
  INV_X1 _29284_ (
    .A(_07435_),
    .ZN(alu_io_in1[16])
  );
  AND2_X1 _29285_ (
    .A1(ex_reg_pc[17]),
    .A2(_07347_),
    .ZN(_07436_)
  );
  INV_X1 _29286_ (
    .A(_07436_),
    .ZN(_07437_)
  );
  AND2_X1 _29287_ (
    .A1(_ex_op1_T[17]),
    .A2(_07352_),
    .ZN(_07438_)
  );
  INV_X1 _29288_ (
    .A(_07438_),
    .ZN(_07439_)
  );
  AND2_X1 _29289_ (
    .A1(_07437_),
    .A2(_07439_),
    .ZN(_07440_)
  );
  INV_X1 _29290_ (
    .A(_07440_),
    .ZN(alu_io_in1[17])
  );
  AND2_X1 _29291_ (
    .A1(ex_reg_pc[18]),
    .A2(_07347_),
    .ZN(_07441_)
  );
  INV_X1 _29292_ (
    .A(_07441_),
    .ZN(_07442_)
  );
  AND2_X1 _29293_ (
    .A1(_ex_op1_T[18]),
    .A2(_07352_),
    .ZN(_07443_)
  );
  INV_X1 _29294_ (
    .A(_07443_),
    .ZN(_07444_)
  );
  AND2_X1 _29295_ (
    .A1(_07442_),
    .A2(_07444_),
    .ZN(_07445_)
  );
  INV_X1 _29296_ (
    .A(_07445_),
    .ZN(alu_io_in1[18])
  );
  AND2_X1 _29297_ (
    .A1(ex_reg_pc[19]),
    .A2(_07347_),
    .ZN(_07446_)
  );
  INV_X1 _29298_ (
    .A(_07446_),
    .ZN(_07447_)
  );
  AND2_X1 _29299_ (
    .A1(_ex_op1_T[19]),
    .A2(_07352_),
    .ZN(_07448_)
  );
  INV_X1 _29300_ (
    .A(_07448_),
    .ZN(_07449_)
  );
  AND2_X1 _29301_ (
    .A1(_07447_),
    .A2(_07449_),
    .ZN(_07450_)
  );
  INV_X1 _29302_ (
    .A(_07450_),
    .ZN(alu_io_in1[19])
  );
  AND2_X1 _29303_ (
    .A1(ex_reg_pc[20]),
    .A2(_07347_),
    .ZN(_07451_)
  );
  INV_X1 _29304_ (
    .A(_07451_),
    .ZN(_07452_)
  );
  AND2_X1 _29305_ (
    .A1(_ex_op1_T[20]),
    .A2(_07352_),
    .ZN(_07453_)
  );
  INV_X1 _29306_ (
    .A(_07453_),
    .ZN(_07454_)
  );
  AND2_X1 _29307_ (
    .A1(_07452_),
    .A2(_07454_),
    .ZN(_07455_)
  );
  INV_X1 _29308_ (
    .A(_07455_),
    .ZN(alu_io_in1[20])
  );
  AND2_X1 _29309_ (
    .A1(ex_reg_pc[21]),
    .A2(_07347_),
    .ZN(_07456_)
  );
  INV_X1 _29310_ (
    .A(_07456_),
    .ZN(_07457_)
  );
  AND2_X1 _29311_ (
    .A1(_ex_op1_T[21]),
    .A2(_07352_),
    .ZN(_07458_)
  );
  INV_X1 _29312_ (
    .A(_07458_),
    .ZN(_07459_)
  );
  AND2_X1 _29313_ (
    .A1(_07457_),
    .A2(_07459_),
    .ZN(_07460_)
  );
  INV_X1 _29314_ (
    .A(_07460_),
    .ZN(alu_io_in1[21])
  );
  AND2_X1 _29315_ (
    .A1(ex_reg_pc[22]),
    .A2(_07347_),
    .ZN(_07461_)
  );
  INV_X1 _29316_ (
    .A(_07461_),
    .ZN(_07462_)
  );
  AND2_X1 _29317_ (
    .A1(_ex_op1_T[22]),
    .A2(_07352_),
    .ZN(_07463_)
  );
  INV_X1 _29318_ (
    .A(_07463_),
    .ZN(_07464_)
  );
  AND2_X1 _29319_ (
    .A1(_07462_),
    .A2(_07464_),
    .ZN(_07465_)
  );
  INV_X1 _29320_ (
    .A(_07465_),
    .ZN(alu_io_in1[22])
  );
  AND2_X1 _29321_ (
    .A1(ex_reg_pc[23]),
    .A2(_07347_),
    .ZN(_07466_)
  );
  INV_X1 _29322_ (
    .A(_07466_),
    .ZN(_07467_)
  );
  AND2_X1 _29323_ (
    .A1(_ex_op1_T[23]),
    .A2(_07352_),
    .ZN(_07468_)
  );
  INV_X1 _29324_ (
    .A(_07468_),
    .ZN(_07469_)
  );
  AND2_X1 _29325_ (
    .A1(_07467_),
    .A2(_07469_),
    .ZN(_07470_)
  );
  INV_X1 _29326_ (
    .A(_07470_),
    .ZN(alu_io_in1[23])
  );
  AND2_X1 _29327_ (
    .A1(ex_reg_pc[24]),
    .A2(_07347_),
    .ZN(_07471_)
  );
  INV_X1 _29328_ (
    .A(_07471_),
    .ZN(_07472_)
  );
  AND2_X1 _29329_ (
    .A1(_ex_op1_T[24]),
    .A2(_07352_),
    .ZN(_07473_)
  );
  INV_X1 _29330_ (
    .A(_07473_),
    .ZN(_07474_)
  );
  AND2_X1 _29331_ (
    .A1(_07472_),
    .A2(_07474_),
    .ZN(_07475_)
  );
  INV_X1 _29332_ (
    .A(_07475_),
    .ZN(alu_io_in1[24])
  );
  AND2_X1 _29333_ (
    .A1(ex_reg_pc[25]),
    .A2(_07347_),
    .ZN(_07476_)
  );
  INV_X1 _29334_ (
    .A(_07476_),
    .ZN(_07477_)
  );
  AND2_X1 _29335_ (
    .A1(_ex_op1_T[25]),
    .A2(_07352_),
    .ZN(_07478_)
  );
  INV_X1 _29336_ (
    .A(_07478_),
    .ZN(_07479_)
  );
  AND2_X1 _29337_ (
    .A1(_07477_),
    .A2(_07479_),
    .ZN(_07480_)
  );
  INV_X1 _29338_ (
    .A(_07480_),
    .ZN(alu_io_in1[25])
  );
  AND2_X1 _29339_ (
    .A1(ex_reg_pc[26]),
    .A2(_07347_),
    .ZN(_07481_)
  );
  INV_X1 _29340_ (
    .A(_07481_),
    .ZN(_07482_)
  );
  AND2_X1 _29341_ (
    .A1(_ex_op1_T[26]),
    .A2(_07352_),
    .ZN(_07483_)
  );
  INV_X1 _29342_ (
    .A(_07483_),
    .ZN(_07484_)
  );
  AND2_X1 _29343_ (
    .A1(_07482_),
    .A2(_07484_),
    .ZN(_07485_)
  );
  INV_X1 _29344_ (
    .A(_07485_),
    .ZN(alu_io_in1[26])
  );
  AND2_X1 _29345_ (
    .A1(ex_reg_pc[27]),
    .A2(_07347_),
    .ZN(_07486_)
  );
  INV_X1 _29346_ (
    .A(_07486_),
    .ZN(_07487_)
  );
  AND2_X1 _29347_ (
    .A1(_ex_op1_T[27]),
    .A2(_07352_),
    .ZN(_07488_)
  );
  INV_X1 _29348_ (
    .A(_07488_),
    .ZN(_07489_)
  );
  AND2_X1 _29349_ (
    .A1(_07487_),
    .A2(_07489_),
    .ZN(_07490_)
  );
  INV_X1 _29350_ (
    .A(_07490_),
    .ZN(alu_io_in1[27])
  );
  AND2_X1 _29351_ (
    .A1(ex_reg_pc[28]),
    .A2(_07347_),
    .ZN(_07491_)
  );
  INV_X1 _29352_ (
    .A(_07491_),
    .ZN(_07492_)
  );
  AND2_X1 _29353_ (
    .A1(_ex_op1_T[28]),
    .A2(_07352_),
    .ZN(_07493_)
  );
  INV_X1 _29354_ (
    .A(_07493_),
    .ZN(_07494_)
  );
  AND2_X1 _29355_ (
    .A1(_07492_),
    .A2(_07494_),
    .ZN(_07495_)
  );
  INV_X1 _29356_ (
    .A(_07495_),
    .ZN(alu_io_in1[28])
  );
  AND2_X1 _29357_ (
    .A1(ex_reg_pc[29]),
    .A2(_07347_),
    .ZN(_07496_)
  );
  INV_X1 _29358_ (
    .A(_07496_),
    .ZN(_07497_)
  );
  AND2_X1 _29359_ (
    .A1(_ex_op1_T[29]),
    .A2(_07352_),
    .ZN(_07498_)
  );
  INV_X1 _29360_ (
    .A(_07498_),
    .ZN(_07499_)
  );
  AND2_X1 _29361_ (
    .A1(_07497_),
    .A2(_07499_),
    .ZN(_07500_)
  );
  INV_X1 _29362_ (
    .A(_07500_),
    .ZN(alu_io_in1[29])
  );
  AND2_X1 _29363_ (
    .A1(ex_reg_pc[30]),
    .A2(_07347_),
    .ZN(_07501_)
  );
  INV_X1 _29364_ (
    .A(_07501_),
    .ZN(_07502_)
  );
  AND2_X1 _29365_ (
    .A1(_ex_op1_T[30]),
    .A2(_07352_),
    .ZN(_07503_)
  );
  INV_X1 _29366_ (
    .A(_07503_),
    .ZN(_07504_)
  );
  AND2_X1 _29367_ (
    .A1(_07502_),
    .A2(_07504_),
    .ZN(_07505_)
  );
  INV_X1 _29368_ (
    .A(_07505_),
    .ZN(alu_io_in1[30])
  );
  AND2_X1 _29369_ (
    .A1(ex_reg_pc[31]),
    .A2(_07347_),
    .ZN(_07506_)
  );
  INV_X1 _29370_ (
    .A(_07506_),
    .ZN(_07507_)
  );
  AND2_X1 _29371_ (
    .A1(_ex_op1_T[31]),
    .A2(_07352_),
    .ZN(_07508_)
  );
  INV_X1 _29372_ (
    .A(_07508_),
    .ZN(_07509_)
  );
  AND2_X1 _29373_ (
    .A1(_07507_),
    .A2(_07509_),
    .ZN(_07510_)
  );
  INV_X1 _29374_ (
    .A(_07510_),
    .ZN(alu_io_in1[31])
  );
  AND2_X1 _29375_ (
    .A1(_08633_),
    .A2(_08647_),
    .ZN(div_io_resp_ready)
  );
  AND2_X1 _29376_ (
    .A1(ex_reg_load_use),
    .A2(_08661_),
    .ZN(_07511_)
  );
  INV_X1 _29377_ (
    .A(_07511_),
    .ZN(_07512_)
  );
  AND2_X1 _29378_ (
    .A1(ex_ctrl_mem),
    .A2(_08605_),
    .ZN(_07513_)
  );
  INV_X1 _29379_ (
    .A(_07513_),
    .ZN(_07514_)
  );
  AND2_X1 _29380_ (
    .A1(ex_ctrl_div),
    .A2(_08604_),
    .ZN(_07515_)
  );
  INV_X1 _29381_ (
    .A(_07515_),
    .ZN(_07516_)
  );
  AND2_X1 _29382_ (
    .A1(_07514_),
    .A2(_07516_),
    .ZN(_07517_)
  );
  AND2_X1 _29383_ (
    .A1(_07512_),
    .A2(_07517_),
    .ZN(_07518_)
  );
  INV_X1 _29384_ (
    .A(_07518_),
    .ZN(_07519_)
  );
  AND2_X1 _29385_ (
    .A1(ex_reg_valid),
    .A2(_07519_),
    .ZN(_07520_)
  );
  INV_X1 _29386_ (
    .A(_07520_),
    .ZN(_07521_)
  );
  AND2_X1 _29387_ (
    .A1(_08618_),
    .A2(_07521_),
    .ZN(_07522_)
  );
  INV_X1 _29388_ (
    .A(_07522_),
    .ZN(_07523_)
  );
  AND2_X1 _29389_ (
    .A1(_08620_),
    .A2(_07522_),
    .ZN(_07524_)
  );
  AND2_X1 _29390_ (
    .A1(_10075_),
    .A2(_07524_),
    .ZN(_mem_reg_valid_T)
  );
  AND2_X1 _29391_ (
    .A1(io_dmem_replay_next),
    .A2(_09148_),
    .ZN(_07525_)
  );
  INV_X1 _29392_ (
    .A(_07525_),
    .ZN(_07526_)
  );
  AND2_X1 _29393_ (
    .A1(_08596_),
    .A2(_08626_),
    .ZN(_07527_)
  );
  AND2_X1 _29394_ (
    .A1(_07526_),
    .A2(_07527_),
    .ZN(_07528_)
  );
  AND2_X1 _29395_ (
    .A1(io_imem_req_bits_speculative),
    .A2(_07528_),
    .ZN(_07529_)
  );
  INV_X1 _29396_ (
    .A(_07529_),
    .ZN(_07530_)
  );
  AND2_X1 _29397_ (
    .A1(mem_reg_load),
    .A2(bpu_io_xcpt_ld),
    .ZN(_07531_)
  );
  INV_X1 _29398_ (
    .A(_07531_),
    .ZN(_07532_)
  );
  AND2_X1 _29399_ (
    .A1(mem_reg_store),
    .A2(bpu_io_xcpt_st),
    .ZN(_07533_)
  );
  INV_X1 _29400_ (
    .A(_07533_),
    .ZN(_07534_)
  );
  AND2_X1 _29401_ (
    .A1(_07532_),
    .A2(_07534_),
    .ZN(_07535_)
  );
  AND2_X1 _29402_ (
    .A1(_06310_),
    .A2(_07535_),
    .ZN(_07536_)
  );
  INV_X1 _29403_ (
    .A(_07536_),
    .ZN(_07537_)
  );
  AND2_X1 _29404_ (
    .A1(mem_reg_valid),
    .A2(_07537_),
    .ZN(_07538_)
  );
  INV_X1 _29405_ (
    .A(_07538_),
    .ZN(_07539_)
  );
  AND2_X1 _29406_ (
    .A1(_06314_),
    .A2(_07539_),
    .ZN(_07540_)
  );
  INV_X1 _29407_ (
    .A(_07540_),
    .ZN(_07541_)
  );
  AND2_X1 _29408_ (
    .A1(_07529_),
    .A2(_07540_),
    .ZN(_wb_reg_valid_T)
  );
  AND2_X1 _29409_ (
    .A1(mem_reg_valid),
    .A2(io_imem_req_bits_speculative),
    .ZN(io_imem_bht_update_valid)
  );
  AND2_X1 _29410_ (
    .A1(bpu_io_pc[31]),
    .A2(_07003_),
    .ZN(_07542_)
  );
  INV_X1 _29411_ (
    .A(_07542_),
    .ZN(_07543_)
  );
  AND2_X1 _29412_ (
    .A1(_08186_),
    .A2(_07004_),
    .ZN(_07544_)
  );
  INV_X1 _29413_ (
    .A(_07544_),
    .ZN(_07545_)
  );
  AND2_X1 _29414_ (
    .A1(bpu_io_pc[30]),
    .A2(_06991_),
    .ZN(_07546_)
  );
  INV_X1 _29415_ (
    .A(_07546_),
    .ZN(_07547_)
  );
  AND2_X1 _29416_ (
    .A1(_08185_),
    .A2(_06992_),
    .ZN(_07548_)
  );
  INV_X1 _29417_ (
    .A(_07548_),
    .ZN(_07549_)
  );
  AND2_X1 _29418_ (
    .A1(bpu_io_pc[29]),
    .A2(_06980_),
    .ZN(_07550_)
  );
  INV_X1 _29419_ (
    .A(_07550_),
    .ZN(_07551_)
  );
  AND2_X1 _29420_ (
    .A1(_08184_),
    .A2(_06979_),
    .ZN(_07552_)
  );
  INV_X1 _29421_ (
    .A(_07552_),
    .ZN(_07553_)
  );
  AND2_X1 _29422_ (
    .A1(_07551_),
    .A2(_07553_),
    .ZN(_07554_)
  );
  INV_X1 _29423_ (
    .A(_07554_),
    .ZN(_07555_)
  );
  AND2_X1 _29424_ (
    .A1(_08182_),
    .A2(_06956_),
    .ZN(_07556_)
  );
  INV_X1 _29425_ (
    .A(_07556_),
    .ZN(_07557_)
  );
  AND2_X1 _29426_ (
    .A1(bpu_io_pc[27]),
    .A2(_06955_),
    .ZN(_07558_)
  );
  INV_X1 _29427_ (
    .A(_07558_),
    .ZN(_07559_)
  );
  AND2_X1 _29428_ (
    .A1(_07557_),
    .A2(_07559_),
    .ZN(_07560_)
  );
  AND2_X1 _29429_ (
    .A1(_08181_),
    .A2(_06944_),
    .ZN(_07561_)
  );
  INV_X1 _29430_ (
    .A(_07561_),
    .ZN(_07562_)
  );
  AND2_X1 _29431_ (
    .A1(bpu_io_pc[26]),
    .A2(_06943_),
    .ZN(_07563_)
  );
  INV_X1 _29432_ (
    .A(_07563_),
    .ZN(_07564_)
  );
  AND2_X1 _29433_ (
    .A1(_07562_),
    .A2(_07564_),
    .ZN(_07565_)
  );
  AND2_X1 _29434_ (
    .A1(bpu_io_pc[25]),
    .A2(_06931_),
    .ZN(_07566_)
  );
  INV_X1 _29435_ (
    .A(_07566_),
    .ZN(_07567_)
  );
  AND2_X1 _29436_ (
    .A1(_08179_),
    .A2(_06920_),
    .ZN(_07568_)
  );
  INV_X1 _29437_ (
    .A(_07568_),
    .ZN(_07569_)
  );
  AND2_X1 _29438_ (
    .A1(bpu_io_pc[24]),
    .A2(_06919_),
    .ZN(_07570_)
  );
  INV_X1 _29439_ (
    .A(_07570_),
    .ZN(_07571_)
  );
  AND2_X1 _29440_ (
    .A1(_07569_),
    .A2(_07571_),
    .ZN(_07572_)
  );
  AND2_X1 _29441_ (
    .A1(_08177_),
    .A2(_06896_),
    .ZN(_07573_)
  );
  INV_X1 _29442_ (
    .A(_07573_),
    .ZN(_07574_)
  );
  AND2_X1 _29443_ (
    .A1(bpu_io_pc[22]),
    .A2(_06895_),
    .ZN(_07575_)
  );
  INV_X1 _29444_ (
    .A(_07575_),
    .ZN(_07576_)
  );
  AND2_X1 _29445_ (
    .A1(_07574_),
    .A2(_07576_),
    .ZN(_07577_)
  );
  AND2_X1 _29446_ (
    .A1(_08176_),
    .A2(_06884_),
    .ZN(_07578_)
  );
  INV_X1 _29447_ (
    .A(_07578_),
    .ZN(_07579_)
  );
  AND2_X1 _29448_ (
    .A1(bpu_io_pc[21]),
    .A2(_06883_),
    .ZN(_07580_)
  );
  INV_X1 _29449_ (
    .A(_07580_),
    .ZN(_07581_)
  );
  AND2_X1 _29450_ (
    .A1(bpu_io_pc[20]),
    .A2(_06871_),
    .ZN(_07582_)
  );
  INV_X1 _29451_ (
    .A(_07582_),
    .ZN(_07583_)
  );
  AND2_X1 _29452_ (
    .A1(_08175_),
    .A2(_06872_),
    .ZN(_07584_)
  );
  INV_X1 _29453_ (
    .A(_07584_),
    .ZN(_07585_)
  );
  AND2_X1 _29454_ (
    .A1(bpu_io_pc[19]),
    .A2(_06859_),
    .ZN(_07586_)
  );
  INV_X1 _29455_ (
    .A(_07586_),
    .ZN(_07587_)
  );
  AND2_X1 _29456_ (
    .A1(_08174_),
    .A2(_06860_),
    .ZN(_07588_)
  );
  INV_X1 _29457_ (
    .A(_07588_),
    .ZN(_07589_)
  );
  AND2_X1 _29458_ (
    .A1(bpu_io_pc[18]),
    .A2(_06847_),
    .ZN(_07590_)
  );
  INV_X1 _29459_ (
    .A(_07590_),
    .ZN(_07591_)
  );
  AND2_X1 _29460_ (
    .A1(_08173_),
    .A2(_06848_),
    .ZN(_07592_)
  );
  INV_X1 _29461_ (
    .A(_07592_),
    .ZN(_07593_)
  );
  AND2_X1 _29462_ (
    .A1(bpu_io_pc[17]),
    .A2(_06835_),
    .ZN(_07594_)
  );
  INV_X1 _29463_ (
    .A(_07594_),
    .ZN(_07595_)
  );
  AND2_X1 _29464_ (
    .A1(_08172_),
    .A2(_06836_),
    .ZN(_07596_)
  );
  INV_X1 _29465_ (
    .A(_07596_),
    .ZN(_07597_)
  );
  AND2_X1 _29466_ (
    .A1(bpu_io_pc[16]),
    .A2(_06823_),
    .ZN(_07598_)
  );
  INV_X1 _29467_ (
    .A(_07598_),
    .ZN(_07599_)
  );
  AND2_X1 _29468_ (
    .A1(_08171_),
    .A2(_06824_),
    .ZN(_07600_)
  );
  INV_X1 _29469_ (
    .A(_07600_),
    .ZN(_07601_)
  );
  AND2_X1 _29470_ (
    .A1(bpu_io_pc[15]),
    .A2(_06811_),
    .ZN(_07602_)
  );
  INV_X1 _29471_ (
    .A(_07602_),
    .ZN(_07603_)
  );
  AND2_X1 _29472_ (
    .A1(_08170_),
    .A2(_06812_),
    .ZN(_07604_)
  );
  INV_X1 _29473_ (
    .A(_07604_),
    .ZN(_07605_)
  );
  AND2_X1 _29474_ (
    .A1(_08169_),
    .A2(_06800_),
    .ZN(_07606_)
  );
  INV_X1 _29475_ (
    .A(_07606_),
    .ZN(_07607_)
  );
  AND2_X1 _29476_ (
    .A1(bpu_io_pc[14]),
    .A2(_06799_),
    .ZN(_07608_)
  );
  INV_X1 _29477_ (
    .A(_07608_),
    .ZN(_07609_)
  );
  AND2_X1 _29478_ (
    .A1(_08168_),
    .A2(_06788_),
    .ZN(_07610_)
  );
  INV_X1 _29479_ (
    .A(_07610_),
    .ZN(_07611_)
  );
  AND2_X1 _29480_ (
    .A1(bpu_io_pc[13]),
    .A2(_06787_),
    .ZN(_07612_)
  );
  INV_X1 _29481_ (
    .A(_07612_),
    .ZN(_07613_)
  );
  AND2_X1 _29482_ (
    .A1(bpu_io_pc[12]),
    .A2(_06775_),
    .ZN(_07614_)
  );
  INV_X1 _29483_ (
    .A(_07614_),
    .ZN(_07615_)
  );
  AND2_X1 _29484_ (
    .A1(_08167_),
    .A2(_06776_),
    .ZN(_07616_)
  );
  INV_X1 _29485_ (
    .A(_07616_),
    .ZN(_07617_)
  );
  AND2_X1 _29486_ (
    .A1(_08166_),
    .A2(_06764_),
    .ZN(_07618_)
  );
  INV_X1 _29487_ (
    .A(_07618_),
    .ZN(_07619_)
  );
  AND2_X1 _29488_ (
    .A1(bpu_io_pc[11]),
    .A2(_06763_),
    .ZN(_07620_)
  );
  INV_X1 _29489_ (
    .A(_07620_),
    .ZN(_07621_)
  );
  AND2_X1 _29490_ (
    .A1(_08165_),
    .A2(_06752_),
    .ZN(_07622_)
  );
  INV_X1 _29491_ (
    .A(_07622_),
    .ZN(_07623_)
  );
  AND2_X1 _29492_ (
    .A1(bpu_io_pc[10]),
    .A2(_06751_),
    .ZN(_07624_)
  );
  INV_X1 _29493_ (
    .A(_07624_),
    .ZN(_07625_)
  );
  AND2_X1 _29494_ (
    .A1(_08164_),
    .A2(_06740_),
    .ZN(_07626_)
  );
  INV_X1 _29495_ (
    .A(_07626_),
    .ZN(_07627_)
  );
  AND2_X1 _29496_ (
    .A1(bpu_io_pc[9]),
    .A2(_06739_),
    .ZN(_07628_)
  );
  INV_X1 _29497_ (
    .A(_07628_),
    .ZN(_07629_)
  );
  AND2_X1 _29498_ (
    .A1(_08163_),
    .A2(_06728_),
    .ZN(_07630_)
  );
  INV_X1 _29499_ (
    .A(_07630_),
    .ZN(_07631_)
  );
  AND2_X1 _29500_ (
    .A1(bpu_io_pc[8]),
    .A2(_06727_),
    .ZN(_07632_)
  );
  INV_X1 _29501_ (
    .A(_07632_),
    .ZN(_07633_)
  );
  AND2_X1 _29502_ (
    .A1(bpu_io_pc[7]),
    .A2(_06715_),
    .ZN(_07634_)
  );
  INV_X1 _29503_ (
    .A(_07634_),
    .ZN(_07635_)
  );
  AND2_X1 _29504_ (
    .A1(_08162_),
    .A2(_06716_),
    .ZN(_07636_)
  );
  INV_X1 _29505_ (
    .A(_07636_),
    .ZN(_07637_)
  );
  AND2_X1 _29506_ (
    .A1(bpu_io_pc[6]),
    .A2(_06703_),
    .ZN(_07638_)
  );
  INV_X1 _29507_ (
    .A(_07638_),
    .ZN(_07639_)
  );
  AND2_X1 _29508_ (
    .A1(_08161_),
    .A2(_06704_),
    .ZN(_07640_)
  );
  INV_X1 _29509_ (
    .A(_07640_),
    .ZN(_07641_)
  );
  AND2_X1 _29510_ (
    .A1(_08160_),
    .A2(_06692_),
    .ZN(_07642_)
  );
  INV_X1 _29511_ (
    .A(_07642_),
    .ZN(_07643_)
  );
  AND2_X1 _29512_ (
    .A1(bpu_io_pc[5]),
    .A2(_06691_),
    .ZN(_07644_)
  );
  INV_X1 _29513_ (
    .A(_07644_),
    .ZN(_07645_)
  );
  AND2_X1 _29514_ (
    .A1(_08159_),
    .A2(_06686_),
    .ZN(_07646_)
  );
  INV_X1 _29515_ (
    .A(_07646_),
    .ZN(_07647_)
  );
  AND2_X1 _29516_ (
    .A1(bpu_io_pc[4]),
    .A2(_06687_),
    .ZN(_07648_)
  );
  INV_X1 _29517_ (
    .A(_07648_),
    .ZN(_07649_)
  );
  AND2_X1 _29518_ (
    .A1(bpu_io_pc[3]),
    .A2(_06684_),
    .ZN(_07650_)
  );
  INV_X1 _29519_ (
    .A(_07650_),
    .ZN(_07651_)
  );
  AND2_X1 _29520_ (
    .A1(_08158_),
    .A2(_06683_),
    .ZN(_07652_)
  );
  INV_X1 _29521_ (
    .A(_07652_),
    .ZN(_07653_)
  );
  AND2_X1 _29522_ (
    .A1(_08157_),
    .A2(_06680_),
    .ZN(_07654_)
  );
  INV_X1 _29523_ (
    .A(_07654_),
    .ZN(_07655_)
  );
  AND2_X1 _29524_ (
    .A1(bpu_io_pc[2]),
    .A2(_06681_),
    .ZN(_07656_)
  );
  INV_X1 _29525_ (
    .A(_07656_),
    .ZN(_07657_)
  );
  AND2_X1 _29526_ (
    .A1(_08156_),
    .A2(_13843_),
    .ZN(_07658_)
  );
  INV_X1 _29527_ (
    .A(_07658_),
    .ZN(_07659_)
  );
  AND2_X1 _29528_ (
    .A1(bpu_io_pc[1]),
    .A2(_13844_),
    .ZN(_07660_)
  );
  INV_X1 _29529_ (
    .A(_07660_),
    .ZN(_07661_)
  );
  AND2_X1 _29530_ (
    .A1(_07659_),
    .A2(_07661_),
    .ZN(_07662_)
  );
  AND2_X1 _29531_ (
    .A1(_08603_),
    .A2(_08625_),
    .ZN(_07663_)
  );
  INV_X1 _29532_ (
    .A(_07663_),
    .ZN(_07664_)
  );
  AND2_X1 _29533_ (
    .A1(_08155_),
    .A2(_07664_),
    .ZN(_07665_)
  );
  AND2_X1 _29534_ (
    .A1(_05249_),
    .A2(_07665_),
    .ZN(_07666_)
  );
  AND2_X1 _29535_ (
    .A1(_07662_),
    .A2(_07666_),
    .ZN(_07667_)
  );
  AND2_X1 _29536_ (
    .A1(bpu_io_pc[23]),
    .A2(_06908_),
    .ZN(_07668_)
  );
  INV_X1 _29537_ (
    .A(_07668_),
    .ZN(_07669_)
  );
  AND2_X1 _29538_ (
    .A1(_08178_),
    .A2(_06907_),
    .ZN(_07670_)
  );
  INV_X1 _29539_ (
    .A(_07670_),
    .ZN(_07671_)
  );
  AND2_X1 _29540_ (
    .A1(_07669_),
    .A2(_07671_),
    .ZN(_07672_)
  );
  INV_X1 _29541_ (
    .A(_07672_),
    .ZN(_07673_)
  );
  AND2_X1 _29542_ (
    .A1(_08180_),
    .A2(_06932_),
    .ZN(_07674_)
  );
  INV_X1 _29543_ (
    .A(_07674_),
    .ZN(_07675_)
  );
  AND2_X1 _29544_ (
    .A1(_08183_),
    .A2(_06968_),
    .ZN(_07676_)
  );
  INV_X1 _29545_ (
    .A(_07676_),
    .ZN(_07677_)
  );
  AND2_X1 _29546_ (
    .A1(bpu_io_pc[28]),
    .A2(_06967_),
    .ZN(_07678_)
  );
  INV_X1 _29547_ (
    .A(_07678_),
    .ZN(_07679_)
  );
  AND2_X1 _29548_ (
    .A1(mem_ctrl_branch),
    .A2(_10070_),
    .ZN(_07680_)
  );
  INV_X1 _29549_ (
    .A(_07680_),
    .ZN(_07681_)
  );
  AND2_X1 _29550_ (
    .A1(io_imem_bht_update_valid),
    .A2(_07681_),
    .ZN(_07682_)
  );
  AND2_X1 _29551_ (
    .A1(ex_reg_pc[31]),
    .A2(_07004_),
    .ZN(_07683_)
  );
  INV_X1 _29552_ (
    .A(_07683_),
    .ZN(_07684_)
  );
  AND2_X1 _29553_ (
    .A1(_08126_),
    .A2(_07003_),
    .ZN(_07685_)
  );
  INV_X1 _29554_ (
    .A(_07685_),
    .ZN(_07686_)
  );
  AND2_X1 _29555_ (
    .A1(_07684_),
    .A2(_07686_),
    .ZN(_07687_)
  );
  INV_X1 _29556_ (
    .A(_07687_),
    .ZN(_07688_)
  );
  AND2_X1 _29557_ (
    .A1(ex_reg_pc[30]),
    .A2(_06991_),
    .ZN(_07689_)
  );
  INV_X1 _29558_ (
    .A(_07689_),
    .ZN(_07690_)
  );
  AND2_X1 _29559_ (
    .A1(_08125_),
    .A2(_06992_),
    .ZN(_07691_)
  );
  INV_X1 _29560_ (
    .A(_07691_),
    .ZN(_07692_)
  );
  AND2_X1 _29561_ (
    .A1(ex_reg_pc[29]),
    .A2(_06979_),
    .ZN(_07693_)
  );
  INV_X1 _29562_ (
    .A(_07693_),
    .ZN(_07694_)
  );
  AND2_X1 _29563_ (
    .A1(_08124_),
    .A2(_06980_),
    .ZN(_07695_)
  );
  INV_X1 _29564_ (
    .A(_07695_),
    .ZN(_07696_)
  );
  AND2_X1 _29565_ (
    .A1(_07694_),
    .A2(_07696_),
    .ZN(_07697_)
  );
  AND2_X1 _29566_ (
    .A1(ex_reg_pc[27]),
    .A2(_06955_),
    .ZN(_07698_)
  );
  INV_X1 _29567_ (
    .A(_07698_),
    .ZN(_07699_)
  );
  AND2_X1 _29568_ (
    .A1(_08122_),
    .A2(_06956_),
    .ZN(_07700_)
  );
  INV_X1 _29569_ (
    .A(_07700_),
    .ZN(_07701_)
  );
  AND2_X1 _29570_ (
    .A1(_07699_),
    .A2(_07701_),
    .ZN(_07702_)
  );
  AND2_X1 _29571_ (
    .A1(ex_reg_pc[28]),
    .A2(_06967_),
    .ZN(_07703_)
  );
  INV_X1 _29572_ (
    .A(_07703_),
    .ZN(_07704_)
  );
  AND2_X1 _29573_ (
    .A1(_08123_),
    .A2(_06968_),
    .ZN(_07705_)
  );
  INV_X1 _29574_ (
    .A(_07705_),
    .ZN(_07706_)
  );
  AND2_X1 _29575_ (
    .A1(_07704_),
    .A2(_07706_),
    .ZN(_07707_)
  );
  AND2_X1 _29576_ (
    .A1(ex_reg_pc[26]),
    .A2(_06943_),
    .ZN(_07708_)
  );
  INV_X1 _29577_ (
    .A(_07708_),
    .ZN(_07709_)
  );
  AND2_X1 _29578_ (
    .A1(_08121_),
    .A2(_06944_),
    .ZN(_07710_)
  );
  INV_X1 _29579_ (
    .A(_07710_),
    .ZN(_07711_)
  );
  AND2_X1 _29580_ (
    .A1(_07709_),
    .A2(_07711_),
    .ZN(_07712_)
  );
  AND2_X1 _29581_ (
    .A1(_08120_),
    .A2(_06932_),
    .ZN(_07713_)
  );
  INV_X1 _29582_ (
    .A(_07713_),
    .ZN(_07714_)
  );
  AND2_X1 _29583_ (
    .A1(ex_reg_pc[25]),
    .A2(_06931_),
    .ZN(_07715_)
  );
  INV_X1 _29584_ (
    .A(_07715_),
    .ZN(_07716_)
  );
  AND2_X1 _29585_ (
    .A1(_07714_),
    .A2(_07716_),
    .ZN(_07717_)
  );
  AND2_X1 _29586_ (
    .A1(ex_reg_pc[23]),
    .A2(_06907_),
    .ZN(_07718_)
  );
  INV_X1 _29587_ (
    .A(_07718_),
    .ZN(_07719_)
  );
  AND2_X1 _29588_ (
    .A1(_08118_),
    .A2(_06908_),
    .ZN(_07720_)
  );
  INV_X1 _29589_ (
    .A(_07720_),
    .ZN(_07721_)
  );
  AND2_X1 _29590_ (
    .A1(_07719_),
    .A2(_07721_),
    .ZN(_07722_)
  );
  AND2_X1 _29591_ (
    .A1(_08119_),
    .A2(_06920_),
    .ZN(_07723_)
  );
  INV_X1 _29592_ (
    .A(_07723_),
    .ZN(_07724_)
  );
  AND2_X1 _29593_ (
    .A1(ex_reg_pc[24]),
    .A2(_06919_),
    .ZN(_07725_)
  );
  INV_X1 _29594_ (
    .A(_07725_),
    .ZN(_07726_)
  );
  AND2_X1 _29595_ (
    .A1(_07724_),
    .A2(_07726_),
    .ZN(_07727_)
  );
  AND2_X1 _29596_ (
    .A1(_08117_),
    .A2(_06896_),
    .ZN(_07728_)
  );
  INV_X1 _29597_ (
    .A(_07728_),
    .ZN(_07729_)
  );
  AND2_X1 _29598_ (
    .A1(ex_reg_pc[22]),
    .A2(_06895_),
    .ZN(_07730_)
  );
  INV_X1 _29599_ (
    .A(_07730_),
    .ZN(_07731_)
  );
  AND2_X1 _29600_ (
    .A1(_07729_),
    .A2(_07731_),
    .ZN(_07732_)
  );
  AND2_X1 _29601_ (
    .A1(_08116_),
    .A2(_06884_),
    .ZN(_07733_)
  );
  INV_X1 _29602_ (
    .A(_07733_),
    .ZN(_07734_)
  );
  AND2_X1 _29603_ (
    .A1(ex_reg_pc[21]),
    .A2(_06883_),
    .ZN(_07735_)
  );
  INV_X1 _29604_ (
    .A(_07735_),
    .ZN(_07736_)
  );
  AND2_X1 _29605_ (
    .A1(_08115_),
    .A2(_06872_),
    .ZN(_07737_)
  );
  INV_X1 _29606_ (
    .A(_07737_),
    .ZN(_07738_)
  );
  AND2_X1 _29607_ (
    .A1(ex_reg_pc[20]),
    .A2(_06871_),
    .ZN(_07739_)
  );
  INV_X1 _29608_ (
    .A(_07739_),
    .ZN(_07740_)
  );
  AND2_X1 _29609_ (
    .A1(_08114_),
    .A2(_06860_),
    .ZN(_07741_)
  );
  INV_X1 _29610_ (
    .A(_07741_),
    .ZN(_07742_)
  );
  AND2_X1 _29611_ (
    .A1(ex_reg_pc[19]),
    .A2(_06859_),
    .ZN(_07743_)
  );
  INV_X1 _29612_ (
    .A(_07743_),
    .ZN(_07744_)
  );
  AND2_X1 _29613_ (
    .A1(_08113_),
    .A2(_06848_),
    .ZN(_07745_)
  );
  INV_X1 _29614_ (
    .A(_07745_),
    .ZN(_07746_)
  );
  AND2_X1 _29615_ (
    .A1(ex_reg_pc[18]),
    .A2(_06847_),
    .ZN(_07747_)
  );
  INV_X1 _29616_ (
    .A(_07747_),
    .ZN(_07748_)
  );
  AND2_X1 _29617_ (
    .A1(ex_reg_pc[17]),
    .A2(_06835_),
    .ZN(_07749_)
  );
  INV_X1 _29618_ (
    .A(_07749_),
    .ZN(_07750_)
  );
  AND2_X1 _29619_ (
    .A1(_08112_),
    .A2(_06836_),
    .ZN(_07751_)
  );
  INV_X1 _29620_ (
    .A(_07751_),
    .ZN(_07752_)
  );
  AND2_X1 _29621_ (
    .A1(_08111_),
    .A2(_06824_),
    .ZN(_07753_)
  );
  INV_X1 _29622_ (
    .A(_07753_),
    .ZN(_07754_)
  );
  AND2_X1 _29623_ (
    .A1(ex_reg_pc[16]),
    .A2(_06823_),
    .ZN(_07755_)
  );
  INV_X1 _29624_ (
    .A(_07755_),
    .ZN(_07756_)
  );
  AND2_X1 _29625_ (
    .A1(ex_reg_pc[15]),
    .A2(_06811_),
    .ZN(_07757_)
  );
  INV_X1 _29626_ (
    .A(_07757_),
    .ZN(_07758_)
  );
  AND2_X1 _29627_ (
    .A1(_08110_),
    .A2(_06812_),
    .ZN(_07759_)
  );
  INV_X1 _29628_ (
    .A(_07759_),
    .ZN(_07760_)
  );
  AND2_X1 _29629_ (
    .A1(_08109_),
    .A2(_06800_),
    .ZN(_07761_)
  );
  INV_X1 _29630_ (
    .A(_07761_),
    .ZN(_07762_)
  );
  AND2_X1 _29631_ (
    .A1(ex_reg_pc[14]),
    .A2(_06799_),
    .ZN(_07763_)
  );
  INV_X1 _29632_ (
    .A(_07763_),
    .ZN(_07764_)
  );
  AND2_X1 _29633_ (
    .A1(ex_reg_pc[13]),
    .A2(_06787_),
    .ZN(_07765_)
  );
  INV_X1 _29634_ (
    .A(_07765_),
    .ZN(_07766_)
  );
  AND2_X1 _29635_ (
    .A1(_08108_),
    .A2(_06788_),
    .ZN(_07767_)
  );
  INV_X1 _29636_ (
    .A(_07767_),
    .ZN(_07768_)
  );
  AND2_X1 _29637_ (
    .A1(_08107_),
    .A2(_06776_),
    .ZN(_07769_)
  );
  INV_X1 _29638_ (
    .A(_07769_),
    .ZN(_07770_)
  );
  AND2_X1 _29639_ (
    .A1(ex_reg_pc[12]),
    .A2(_06775_),
    .ZN(_07771_)
  );
  INV_X1 _29640_ (
    .A(_07771_),
    .ZN(_07772_)
  );
  AND2_X1 _29641_ (
    .A1(_08106_),
    .A2(_06764_),
    .ZN(_07773_)
  );
  INV_X1 _29642_ (
    .A(_07773_),
    .ZN(_07774_)
  );
  AND2_X1 _29643_ (
    .A1(ex_reg_pc[11]),
    .A2(_06763_),
    .ZN(_07775_)
  );
  INV_X1 _29644_ (
    .A(_07775_),
    .ZN(_07776_)
  );
  AND2_X1 _29645_ (
    .A1(_08105_),
    .A2(_06752_),
    .ZN(_07777_)
  );
  INV_X1 _29646_ (
    .A(_07777_),
    .ZN(_07778_)
  );
  AND2_X1 _29647_ (
    .A1(ex_reg_pc[10]),
    .A2(_06751_),
    .ZN(_07779_)
  );
  INV_X1 _29648_ (
    .A(_07779_),
    .ZN(_07780_)
  );
  AND2_X1 _29649_ (
    .A1(ex_reg_pc[9]),
    .A2(_06739_),
    .ZN(_07781_)
  );
  INV_X1 _29650_ (
    .A(_07781_),
    .ZN(_07782_)
  );
  AND2_X1 _29651_ (
    .A1(_08104_),
    .A2(_06740_),
    .ZN(_07783_)
  );
  INV_X1 _29652_ (
    .A(_07783_),
    .ZN(_07784_)
  );
  AND2_X1 _29653_ (
    .A1(_08103_),
    .A2(_06728_),
    .ZN(_07785_)
  );
  INV_X1 _29654_ (
    .A(_07785_),
    .ZN(_07786_)
  );
  AND2_X1 _29655_ (
    .A1(ex_reg_pc[8]),
    .A2(_06727_),
    .ZN(_07787_)
  );
  INV_X1 _29656_ (
    .A(_07787_),
    .ZN(_07788_)
  );
  AND2_X1 _29657_ (
    .A1(ex_reg_pc[7]),
    .A2(_06715_),
    .ZN(_07789_)
  );
  INV_X1 _29658_ (
    .A(_07789_),
    .ZN(_07790_)
  );
  AND2_X1 _29659_ (
    .A1(_08102_),
    .A2(_06716_),
    .ZN(_07791_)
  );
  INV_X1 _29660_ (
    .A(_07791_),
    .ZN(_07792_)
  );
  AND2_X1 _29661_ (
    .A1(_08101_),
    .A2(_06704_),
    .ZN(_07793_)
  );
  INV_X1 _29662_ (
    .A(_07793_),
    .ZN(_07794_)
  );
  AND2_X1 _29663_ (
    .A1(ex_reg_pc[6]),
    .A2(_06703_),
    .ZN(_07795_)
  );
  INV_X1 _29664_ (
    .A(_07795_),
    .ZN(_07796_)
  );
  AND2_X1 _29665_ (
    .A1(_07794_),
    .A2(_07796_),
    .ZN(_07797_)
  );
  AND2_X1 _29666_ (
    .A1(ex_reg_pc[5]),
    .A2(_06691_),
    .ZN(_07798_)
  );
  INV_X1 _29667_ (
    .A(_07798_),
    .ZN(_07799_)
  );
  AND2_X1 _29668_ (
    .A1(ex_reg_pc[4]),
    .A2(_06687_),
    .ZN(_07800_)
  );
  INV_X1 _29669_ (
    .A(_07800_),
    .ZN(_07801_)
  );
  AND2_X1 _29670_ (
    .A1(_08099_),
    .A2(_06686_),
    .ZN(_07802_)
  );
  INV_X1 _29671_ (
    .A(_07802_),
    .ZN(_07803_)
  );
  AND2_X1 _29672_ (
    .A1(_08098_),
    .A2(_06683_),
    .ZN(_07804_)
  );
  INV_X1 _29673_ (
    .A(_07804_),
    .ZN(_07805_)
  );
  AND2_X1 _29674_ (
    .A1(ex_reg_pc[3]),
    .A2(_06684_),
    .ZN(_07806_)
  );
  INV_X1 _29675_ (
    .A(_07806_),
    .ZN(_07807_)
  );
  AND2_X1 _29676_ (
    .A1(ex_reg_pc[2]),
    .A2(_06681_),
    .ZN(_07808_)
  );
  INV_X1 _29677_ (
    .A(_07808_),
    .ZN(_07809_)
  );
  AND2_X1 _29678_ (
    .A1(_08097_),
    .A2(_06680_),
    .ZN(_07810_)
  );
  INV_X1 _29679_ (
    .A(_07810_),
    .ZN(_07811_)
  );
  AND2_X1 _29680_ (
    .A1(_08096_),
    .A2(_13843_),
    .ZN(_07812_)
  );
  INV_X1 _29681_ (
    .A(_07812_),
    .ZN(_07813_)
  );
  AND2_X1 _29682_ (
    .A1(ex_reg_pc[1]),
    .A2(_13844_),
    .ZN(_07814_)
  );
  INV_X1 _29683_ (
    .A(_07814_),
    .ZN(_07815_)
  );
  AND2_X1 _29684_ (
    .A1(_08095_),
    .A2(_05250_),
    .ZN(_07816_)
  );
  AND2_X1 _29685_ (
    .A1(_07813_),
    .A2(_07815_),
    .ZN(_07817_)
  );
  AND2_X1 _29686_ (
    .A1(_07816_),
    .A2(_07817_),
    .ZN(_07818_)
  );
  AND2_X1 _29687_ (
    .A1(_07811_),
    .A2(_07818_),
    .ZN(_07819_)
  );
  AND2_X1 _29688_ (
    .A1(_07809_),
    .A2(_07819_),
    .ZN(_07820_)
  );
  AND2_X1 _29689_ (
    .A1(_07805_),
    .A2(_07807_),
    .ZN(_07821_)
  );
  AND2_X1 _29690_ (
    .A1(_07820_),
    .A2(_07821_),
    .ZN(_07822_)
  );
  AND2_X1 _29691_ (
    .A1(_07803_),
    .A2(_07822_),
    .ZN(_07823_)
  );
  AND2_X1 _29692_ (
    .A1(_07801_),
    .A2(_07823_),
    .ZN(_07824_)
  );
  AND2_X1 _29693_ (
    .A1(_08100_),
    .A2(_06692_),
    .ZN(_07825_)
  );
  INV_X1 _29694_ (
    .A(_07825_),
    .ZN(_07826_)
  );
  AND2_X1 _29695_ (
    .A1(_07824_),
    .A2(_07826_),
    .ZN(_07827_)
  );
  AND2_X1 _29696_ (
    .A1(_07799_),
    .A2(_07827_),
    .ZN(_07828_)
  );
  AND2_X1 _29697_ (
    .A1(_07797_),
    .A2(_07828_),
    .ZN(_07829_)
  );
  AND2_X1 _29698_ (
    .A1(_07547_),
    .A2(_07549_),
    .ZN(_07830_)
  );
  AND2_X1 _29699_ (
    .A1(_07567_),
    .A2(_07675_),
    .ZN(_07831_)
  );
  AND2_X1 _29700_ (
    .A1(_07565_),
    .A2(_07679_),
    .ZN(_07832_)
  );
  AND2_X1 _29701_ (
    .A1(_07587_),
    .A2(_07589_),
    .ZN(_07833_)
  );
  AND2_X1 _29702_ (
    .A1(_07591_),
    .A2(_07593_),
    .ZN(_07834_)
  );
  AND2_X1 _29703_ (
    .A1(_07603_),
    .A2(_07605_),
    .ZN(_07835_)
  );
  AND2_X1 _29704_ (
    .A1(_07653_),
    .A2(_07667_),
    .ZN(_07836_)
  );
  AND2_X1 _29705_ (
    .A1(_07649_),
    .A2(_07836_),
    .ZN(_07837_)
  );
  AND2_X1 _29706_ (
    .A1(_07645_),
    .A2(_07837_),
    .ZN(_07838_)
  );
  AND2_X1 _29707_ (
    .A1(_07641_),
    .A2(_07838_),
    .ZN(_07839_)
  );
  AND2_X1 _29708_ (
    .A1(_07637_),
    .A2(_07839_),
    .ZN(_07840_)
  );
  AND2_X1 _29709_ (
    .A1(_07633_),
    .A2(_07840_),
    .ZN(_07841_)
  );
  AND2_X1 _29710_ (
    .A1(_07629_),
    .A2(_07841_),
    .ZN(_07842_)
  );
  AND2_X1 _29711_ (
    .A1(_07625_),
    .A2(_07842_),
    .ZN(_07843_)
  );
  AND2_X1 _29712_ (
    .A1(_07621_),
    .A2(_07843_),
    .ZN(_07844_)
  );
  AND2_X1 _29713_ (
    .A1(_07617_),
    .A2(_07844_),
    .ZN(_07845_)
  );
  AND2_X1 _29714_ (
    .A1(_07613_),
    .A2(_07845_),
    .ZN(_07846_)
  );
  AND2_X1 _29715_ (
    .A1(_07609_),
    .A2(_07846_),
    .ZN(_07847_)
  );
  AND2_X1 _29716_ (
    .A1(_07655_),
    .A2(_07657_),
    .ZN(_07848_)
  );
  AND2_X1 _29717_ (
    .A1(_07651_),
    .A2(_07848_),
    .ZN(_07849_)
  );
  AND2_X1 _29718_ (
    .A1(_07647_),
    .A2(_07849_),
    .ZN(_07850_)
  );
  AND2_X1 _29719_ (
    .A1(_07643_),
    .A2(_07850_),
    .ZN(_07851_)
  );
  AND2_X1 _29720_ (
    .A1(_07639_),
    .A2(_07851_),
    .ZN(_07852_)
  );
  AND2_X1 _29721_ (
    .A1(_07635_),
    .A2(_07852_),
    .ZN(_07853_)
  );
  AND2_X1 _29722_ (
    .A1(_07631_),
    .A2(_07853_),
    .ZN(_07854_)
  );
  AND2_X1 _29723_ (
    .A1(_07627_),
    .A2(_07854_),
    .ZN(_07855_)
  );
  AND2_X1 _29724_ (
    .A1(_07623_),
    .A2(_07855_),
    .ZN(_07856_)
  );
  AND2_X1 _29725_ (
    .A1(_07619_),
    .A2(_07856_),
    .ZN(_07857_)
  );
  AND2_X1 _29726_ (
    .A1(_07615_),
    .A2(_07857_),
    .ZN(_07858_)
  );
  AND2_X1 _29727_ (
    .A1(_07611_),
    .A2(_07858_),
    .ZN(_07859_)
  );
  AND2_X1 _29728_ (
    .A1(_07607_),
    .A2(_07859_),
    .ZN(_07860_)
  );
  AND2_X1 _29729_ (
    .A1(_07847_),
    .A2(_07860_),
    .ZN(_07861_)
  );
  AND2_X1 _29730_ (
    .A1(_07835_),
    .A2(_07861_),
    .ZN(_07862_)
  );
  AND2_X1 _29731_ (
    .A1(_07599_),
    .A2(_07601_),
    .ZN(_07863_)
  );
  AND2_X1 _29732_ (
    .A1(_07862_),
    .A2(_07863_),
    .ZN(_07864_)
  );
  AND2_X1 _29733_ (
    .A1(_07595_),
    .A2(_07864_),
    .ZN(_07865_)
  );
  AND2_X1 _29734_ (
    .A1(_07597_),
    .A2(_07865_),
    .ZN(_07866_)
  );
  AND2_X1 _29735_ (
    .A1(_07834_),
    .A2(_07866_),
    .ZN(_07867_)
  );
  AND2_X1 _29736_ (
    .A1(_07833_),
    .A2(_07867_),
    .ZN(_07868_)
  );
  AND2_X1 _29737_ (
    .A1(_07583_),
    .A2(_07585_),
    .ZN(_07869_)
  );
  AND2_X1 _29738_ (
    .A1(_07868_),
    .A2(_07869_),
    .ZN(_07870_)
  );
  AND2_X1 _29739_ (
    .A1(_07579_),
    .A2(_07581_),
    .ZN(_07871_)
  );
  AND2_X1 _29740_ (
    .A1(_07870_),
    .A2(_07871_),
    .ZN(_07872_)
  );
  AND2_X1 _29741_ (
    .A1(_07577_),
    .A2(_07872_),
    .ZN(_07873_)
  );
  AND2_X1 _29742_ (
    .A1(_07572_),
    .A2(_07873_),
    .ZN(_07874_)
  );
  AND2_X1 _29743_ (
    .A1(_07673_),
    .A2(_07874_),
    .ZN(_07875_)
  );
  AND2_X1 _29744_ (
    .A1(_07677_),
    .A2(_07875_),
    .ZN(_07876_)
  );
  AND2_X1 _29745_ (
    .A1(_07832_),
    .A2(_07876_),
    .ZN(_07877_)
  );
  AND2_X1 _29746_ (
    .A1(_07560_),
    .A2(_07877_),
    .ZN(_07878_)
  );
  AND2_X1 _29747_ (
    .A1(_07831_),
    .A2(_07878_),
    .ZN(_07879_)
  );
  AND2_X1 _29748_ (
    .A1(_07555_),
    .A2(_07879_),
    .ZN(_07880_)
  );
  AND2_X1 _29749_ (
    .A1(_07830_),
    .A2(_07880_),
    .ZN(_07881_)
  );
  AND2_X1 _29750_ (
    .A1(_07543_),
    .A2(_07545_),
    .ZN(_07882_)
  );
  AND2_X1 _29751_ (
    .A1(_07881_),
    .A2(_07882_),
    .ZN(_07883_)
  );
  INV_X1 _29752_ (
    .A(_07883_),
    .ZN(_07884_)
  );
  AND2_X1 _29753_ (
    .A1(_07682_),
    .A2(_07884_),
    .ZN(_07885_)
  );
  AND2_X1 _29754_ (
    .A1(_07690_),
    .A2(_07692_),
    .ZN(_07886_)
  );
  AND2_X1 _29755_ (
    .A1(_07742_),
    .A2(_07744_),
    .ZN(_07887_)
  );
  AND2_X1 _29756_ (
    .A1(_07746_),
    .A2(_07748_),
    .ZN(_07888_)
  );
  AND2_X1 _29757_ (
    .A1(_07790_),
    .A2(_07792_),
    .ZN(_07889_)
  );
  AND2_X1 _29758_ (
    .A1(_07829_),
    .A2(_07889_),
    .ZN(_07890_)
  );
  AND2_X1 _29759_ (
    .A1(_07786_),
    .A2(_07788_),
    .ZN(_07891_)
  );
  AND2_X1 _29760_ (
    .A1(_07890_),
    .A2(_07891_),
    .ZN(_07892_)
  );
  AND2_X1 _29761_ (
    .A1(_07780_),
    .A2(_07892_),
    .ZN(_07893_)
  );
  AND2_X1 _29762_ (
    .A1(_07776_),
    .A2(_07893_),
    .ZN(_07894_)
  );
  AND2_X1 _29763_ (
    .A1(_07772_),
    .A2(_07894_),
    .ZN(_07895_)
  );
  AND2_X1 _29764_ (
    .A1(_07768_),
    .A2(_07895_),
    .ZN(_07896_)
  );
  AND2_X1 _29765_ (
    .A1(_07764_),
    .A2(_07896_),
    .ZN(_07897_)
  );
  AND2_X1 _29766_ (
    .A1(_07758_),
    .A2(_07897_),
    .ZN(_07898_)
  );
  AND2_X1 _29767_ (
    .A1(_07756_),
    .A2(_07898_),
    .ZN(_07899_)
  );
  AND2_X1 _29768_ (
    .A1(_07752_),
    .A2(_07899_),
    .ZN(_07900_)
  );
  AND2_X1 _29769_ (
    .A1(_07782_),
    .A2(_07784_),
    .ZN(_07901_)
  );
  AND2_X1 _29770_ (
    .A1(_07778_),
    .A2(_07901_),
    .ZN(_07902_)
  );
  AND2_X1 _29771_ (
    .A1(_07774_),
    .A2(_07902_),
    .ZN(_07903_)
  );
  AND2_X1 _29772_ (
    .A1(_07770_),
    .A2(_07903_),
    .ZN(_07904_)
  );
  AND2_X1 _29773_ (
    .A1(_07766_),
    .A2(_07904_),
    .ZN(_07905_)
  );
  AND2_X1 _29774_ (
    .A1(_07762_),
    .A2(_07905_),
    .ZN(_07906_)
  );
  AND2_X1 _29775_ (
    .A1(_07760_),
    .A2(_07906_),
    .ZN(_07907_)
  );
  AND2_X1 _29776_ (
    .A1(_07754_),
    .A2(_07907_),
    .ZN(_07908_)
  );
  AND2_X1 _29777_ (
    .A1(_07750_),
    .A2(_07908_),
    .ZN(_07909_)
  );
  AND2_X1 _29778_ (
    .A1(_07900_),
    .A2(_07909_),
    .ZN(_07910_)
  );
  AND2_X1 _29779_ (
    .A1(_07888_),
    .A2(_07910_),
    .ZN(_07911_)
  );
  AND2_X1 _29780_ (
    .A1(_07887_),
    .A2(_07911_),
    .ZN(_07912_)
  );
  AND2_X1 _29781_ (
    .A1(_07738_),
    .A2(_07740_),
    .ZN(_07913_)
  );
  AND2_X1 _29782_ (
    .A1(_07912_),
    .A2(_07913_),
    .ZN(_07914_)
  );
  AND2_X1 _29783_ (
    .A1(_07734_),
    .A2(_07736_),
    .ZN(_07915_)
  );
  AND2_X1 _29784_ (
    .A1(_07914_),
    .A2(_07915_),
    .ZN(_07916_)
  );
  AND2_X1 _29785_ (
    .A1(_07732_),
    .A2(_07916_),
    .ZN(_07917_)
  );
  AND2_X1 _29786_ (
    .A1(_07727_),
    .A2(_07917_),
    .ZN(_07918_)
  );
  AND2_X1 _29787_ (
    .A1(_07722_),
    .A2(_07918_),
    .ZN(_07919_)
  );
  AND2_X1 _29788_ (
    .A1(_07717_),
    .A2(_07919_),
    .ZN(_07920_)
  );
  AND2_X1 _29789_ (
    .A1(_07712_),
    .A2(_07920_),
    .ZN(_07921_)
  );
  AND2_X1 _29790_ (
    .A1(_07707_),
    .A2(_07921_),
    .ZN(_07922_)
  );
  AND2_X1 _29791_ (
    .A1(_07702_),
    .A2(_07922_),
    .ZN(_07923_)
  );
  AND2_X1 _29792_ (
    .A1(_07697_),
    .A2(_07923_),
    .ZN(_07924_)
  );
  AND2_X1 _29793_ (
    .A1(_07886_),
    .A2(_07924_),
    .ZN(_07925_)
  );
  AND2_X1 _29794_ (
    .A1(_07688_),
    .A2(_07925_),
    .ZN(_07926_)
  );
  INV_X1 _29795_ (
    .A(_07926_),
    .ZN(_07927_)
  );
  AND2_X1 _29796_ (
    .A1(_07885_),
    .A2(_07927_),
    .ZN(io_imem_btb_update_valid)
  );
  AND2_X1 _29797_ (
    .A1(wb_ctrl_fence_i),
    .A2(wb_reg_valid),
    .ZN(_07928_)
  );
  AND2_X1 _29798_ (
    .A1(_08608_),
    .A2(_07928_),
    .ZN(io_imem_flush_icache)
  );
  AND2_X1 _29799_ (
    .A1(_07529_),
    .A2(_07536_),
    .ZN(_07929_)
  );
  INV_X1 _29800_ (
    .A(_07929_),
    .ZN(io_dmem_s1_kill)
  );
  AND2_X1 _29801_ (
    .A1(wb_ctrl_csr[2]),
    .A2(wb_reg_valid),
    .ZN(csr_io_rw_cmd[2])
  );
  AND2_X1 _29802_ (
    .A1(div_io_kill_REG),
    .A2(_07530_),
    .ZN(div_io_kill)
  );
  AND2_X1 _29803_ (
    .A1(_13833_),
    .A2(_05249_),
    .ZN(_07930_)
  );
  AND2_X1 _29804_ (
    .A1(_08629_),
    .A2(_07930_),
    .ZN(_07931_)
  );
  INV_X1 _29805_ (
    .A(_07931_),
    .ZN(_00005_)
  );
  AND2_X1 _29806_ (
    .A1(csr_io_interrupt),
    .A2(_10076_),
    .ZN(_00004_)
  );
  AND2_X1 _29807_ (
    .A1(_ex_reg_valid_T),
    .A2(_05897_),
    .ZN(_00003_)
  );
  AND2_X1 _29808_ (
    .A1(ibuf_io_inst_0_bits_replay),
    .A2(_10076_),
    .ZN(_00002_)
  );
  AND2_X1 _29809_ (
    .A1(ex_reg_xcpt_interrupt),
    .A2(_10075_),
    .ZN(_00008_)
  );
  AND2_X1 _29810_ (
    .A1(_08619_),
    .A2(_08622_),
    .ZN(_07932_)
  );
  INV_X1 _29811_ (
    .A(_07932_),
    .ZN(_07933_)
  );
  AND2_X1 _29812_ (
    .A1(_mem_reg_valid_T),
    .A2(_07933_),
    .ZN(_00007_)
  );
  AND2_X1 _29813_ (
    .A1(_10075_),
    .A2(_07523_),
    .ZN(_00006_)
  );
  AND2_X1 _29814_ (
    .A1(io_imem_req_bits_speculative),
    .A2(_07541_),
    .ZN(_00011_)
  );
  AND2_X1 _29815_ (
    .A1(_08623_),
    .A2(_07526_),
    .ZN(_07934_)
  );
  INV_X1 _29816_ (
    .A(_07934_),
    .ZN(_07935_)
  );
  AND2_X1 _29817_ (
    .A1(io_imem_req_bits_speculative),
    .A2(_07935_),
    .ZN(_00010_)
  );
  AND2_X1 _29818_ (
    .A1(mem_reg_flush_pipe),
    .A2(_wb_reg_valid_T),
    .ZN(_00009_)
  );
  AND2_X1 _29819_ (
    .A1(_08608_),
    .A2(_08615_),
    .ZN(_07936_)
  );
  AND2_X1 _29820_ (
    .A1(_09466_),
    .A2(_07936_),
    .ZN(_07937_)
  );
  INV_X1 _29821_ (
    .A(_07937_),
    .ZN(_07938_)
  );
  AND2_X1 _29822_ (
    .A1(_08602_),
    .A2(_08605_),
    .ZN(_07939_)
  );
  AND2_X1 _29823_ (
    .A1(_07938_),
    .A2(_07939_),
    .ZN(_00000_)
  );
  AND2_X1 _29824_ (
    .A1(div_io_req_ready),
    .A2(div_io_req_valid),
    .ZN(_00001_)
  );
  DFF_X1 \_r[10]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00045_),
    .Q(_r[10]),
    .QN(_15543_)
  );
  DFF_X1 \_r[11]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00046_),
    .Q(_r[11]),
    .QN(_15542_)
  );
  DFF_X1 \_r[12]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00047_),
    .Q(_r[12]),
    .QN(_15541_)
  );
  DFF_X1 \_r[13]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00048_),
    .Q(_r[13]),
    .QN(_15540_)
  );
  DFF_X1 \_r[14]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00049_),
    .Q(_r[14]),
    .QN(_15539_)
  );
  DFF_X1 \_r[15]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00050_),
    .Q(_r[15]),
    .QN(_15538_)
  );
  DFF_X1 \_r[16]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00051_),
    .Q(_r[16]),
    .QN(_15537_)
  );
  DFF_X1 \_r[17]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00052_),
    .Q(_r[17]),
    .QN(_15536_)
  );
  DFF_X1 \_r[18]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00053_),
    .Q(_r[18]),
    .QN(_15535_)
  );
  DFF_X1 \_r[19]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00054_),
    .Q(_r[19]),
    .QN(_15534_)
  );
  DFF_X1 \_r[1]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00036_),
    .Q(_r[1]),
    .QN(_15552_)
  );
  DFF_X1 \_r[20]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00055_),
    .Q(_r[20]),
    .QN(_15533_)
  );
  DFF_X1 \_r[21]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00056_),
    .Q(_r[21]),
    .QN(_15532_)
  );
  DFF_X1 \_r[22]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00057_),
    .Q(_r[22]),
    .QN(_15531_)
  );
  DFF_X1 \_r[23]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00058_),
    .Q(_r[23]),
    .QN(_15530_)
  );
  DFF_X1 \_r[24]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00059_),
    .Q(_r[24]),
    .QN(_15529_)
  );
  DFF_X1 \_r[25]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00060_),
    .Q(_r[25]),
    .QN(_15528_)
  );
  DFF_X1 \_r[26]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00061_),
    .Q(_r[26]),
    .QN(_15527_)
  );
  DFF_X1 \_r[27]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00062_),
    .Q(_r[27]),
    .QN(_15526_)
  );
  DFF_X1 \_r[28]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00063_),
    .Q(_r[28]),
    .QN(_15525_)
  );
  DFF_X1 \_r[29]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00064_),
    .Q(_r[29]),
    .QN(_15524_)
  );
  DFF_X1 \_r[2]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00037_),
    .Q(_r[2]),
    .QN(_15551_)
  );
  DFF_X1 \_r[30]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00065_),
    .Q(_r[30]),
    .QN(_15523_)
  );
  DFF_X1 \_r[31]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00066_),
    .Q(_r[31]),
    .QN(_15522_)
  );
  DFF_X1 \_r[3]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00038_),
    .Q(_r[3]),
    .QN(_15550_)
  );
  DFF_X1 \_r[4]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00039_),
    .Q(_r[4]),
    .QN(_15549_)
  );
  DFF_X1 \_r[5]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00040_),
    .Q(_r[5]),
    .QN(_15548_)
  );
  DFF_X1 \_r[6]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00041_),
    .Q(_r[6]),
    .QN(_15547_)
  );
  DFF_X1 \_r[7]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00042_),
    .Q(_r[7]),
    .QN(_15546_)
  );
  DFF_X1 \_r[8]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00043_),
    .Q(_r[8]),
    .QN(_15545_)
  );
  DFF_X1 \_r[9]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00044_),
    .Q(_r[9]),
    .QN(_15544_)
  );
  ALU alu (
    .io_adder_out(alu_io_adder_out),
    .io_cmp_out(alu_io_cmp_out),
    .io_fn(ex_ctrl_alu_fn),
    .io_in1(alu_io_in1),
    .io_in2(alu_io_in2),
    .io_out(alu_io_out)
  );
  DFF_X1 \blocked$_DFF_P_  (
    .CK(clock),
    .D(_00000_),
    .Q(blocked),
    .QN(_14027_)
  );
  BreakpointUnit bpu (
    .io_bp_0_address(bpu_io_bp_0_address),
    .io_bp_0_control_action(bpu_io_bp_0_control_action),
    .io_bp_0_control_r(bpu_io_bp_0_control_r),
    .io_bp_0_control_tmatch(bpu_io_bp_0_control_tmatch),
    .io_bp_0_control_w(bpu_io_bp_0_control_w),
    .io_bp_0_control_x(bpu_io_bp_0_control_x),
    .io_debug_if(bpu_io_debug_if),
    .io_debug_ld(bpu_io_debug_ld),
    .io_debug_st(bpu_io_debug_st),
    .io_ea(mem_reg_wdata),
    .io_pc(bpu_io_pc),
    .io_status_debug(bpu_io_status_debug),
    .io_xcpt_if(bpu_io_xcpt_if),
    .io_xcpt_ld(bpu_io_xcpt_ld),
    .io_xcpt_st(bpu_io_xcpt_st)
  );
  CSRFile csr (
    .clock(clock),
    .io_bp_0_address(bpu_io_bp_0_address),
    .io_bp_0_control_action(bpu_io_bp_0_control_action),
    .io_bp_0_control_r(bpu_io_bp_0_control_r),
    .io_bp_0_control_tmatch(bpu_io_bp_0_control_tmatch),
    .io_bp_0_control_w(bpu_io_bp_0_control_w),
    .io_bp_0_control_x(bpu_io_bp_0_control_x),
    .io_cause(csr_io_cause),
    .io_csr_stall(csr_io_csr_stall),
    .io_customCSRs_0_value({ csr_io_customCSRs_0_value[31:2], io_ptw_customCSRs_csrs_0_value[1], csr_io_customCSRs_0_value[0] }),
    .io_decode_0_fp_csr(csr_io_decode_0_fp_csr),
    .io_decode_0_fp_illegal(csr_io_decode_0_fp_illegal),
    .io_decode_0_inst(csr_io_decode_0_inst),
    .io_decode_0_read_illegal(csr_io_decode_0_read_illegal),
    .io_decode_0_rocc_illegal(csr_io_decode_0_rocc_illegal),
    .io_decode_0_system_illegal(csr_io_decode_0_system_illegal),
    .io_decode_0_write_flush(csr_io_decode_0_write_flush),
    .io_decode_0_write_illegal(csr_io_decode_0_write_illegal),
    .io_eret(csr_io_eret),
    .io_evec(csr_io_evec),
    .io_exception(csr_io_exception),
    .io_gva(1'h0),
    .io_hartid(io_hartid),
    .io_inhibit_cycle(csr_io_inhibit_cycle),
    .io_inst_0({ _csr_io_inst_0_T_3, wb_reg_raw_inst[15:0] }),
    .io_interrupt(csr_io_interrupt),
    .io_interrupt_cause(csr_io_interrupt_cause),
    .io_interrupts_debug(io_interrupts_debug),
    .io_interrupts_meip(io_interrupts_meip),
    .io_interrupts_msip(io_interrupts_msip),
    .io_interrupts_mtip(io_interrupts_mtip),
    .io_pc(wb_reg_pc),
    .io_pmp_0_addr(csr_io_pmp_0_addr),
    .io_pmp_0_cfg_a(csr_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_l(csr_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_r(csr_io_pmp_0_cfg_r),
    .io_pmp_0_cfg_w(csr_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_x(csr_io_pmp_0_cfg_x),
    .io_pmp_0_mask(csr_io_pmp_0_mask),
    .io_pmp_1_addr(csr_io_pmp_1_addr),
    .io_pmp_1_cfg_a(csr_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_l(csr_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_r(csr_io_pmp_1_cfg_r),
    .io_pmp_1_cfg_w(csr_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_x(csr_io_pmp_1_cfg_x),
    .io_pmp_1_mask(csr_io_pmp_1_mask),
    .io_pmp_2_addr(csr_io_pmp_2_addr),
    .io_pmp_2_cfg_a(csr_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_l(csr_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_r(csr_io_pmp_2_cfg_r),
    .io_pmp_2_cfg_w(csr_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_x(csr_io_pmp_2_cfg_x),
    .io_pmp_2_mask(csr_io_pmp_2_mask),
    .io_pmp_3_addr(csr_io_pmp_3_addr),
    .io_pmp_3_cfg_a(csr_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_l(csr_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_r(csr_io_pmp_3_cfg_r),
    .io_pmp_3_cfg_w(csr_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_x(csr_io_pmp_3_cfg_x),
    .io_pmp_3_mask(csr_io_pmp_3_mask),
    .io_pmp_4_addr(csr_io_pmp_4_addr),
    .io_pmp_4_cfg_a(csr_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_l(csr_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_r(csr_io_pmp_4_cfg_r),
    .io_pmp_4_cfg_w(csr_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_x(csr_io_pmp_4_cfg_x),
    .io_pmp_4_mask(csr_io_pmp_4_mask),
    .io_pmp_5_addr(csr_io_pmp_5_addr),
    .io_pmp_5_cfg_a(csr_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_l(csr_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_r(csr_io_pmp_5_cfg_r),
    .io_pmp_5_cfg_w(csr_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_x(csr_io_pmp_5_cfg_x),
    .io_pmp_5_mask(csr_io_pmp_5_mask),
    .io_pmp_6_addr(csr_io_pmp_6_addr),
    .io_pmp_6_cfg_a(csr_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_l(csr_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_r(csr_io_pmp_6_cfg_r),
    .io_pmp_6_cfg_w(csr_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_x(csr_io_pmp_6_cfg_x),
    .io_pmp_6_mask(csr_io_pmp_6_mask),
    .io_pmp_7_addr(csr_io_pmp_7_addr),
    .io_pmp_7_cfg_a(csr_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_l(csr_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_r(csr_io_pmp_7_cfg_r),
    .io_pmp_7_cfg_w(csr_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_x(csr_io_pmp_7_cfg_x),
    .io_pmp_7_mask(csr_io_pmp_7_mask),
    .io_retire(csr_io_retire),
    .io_rw_addr(wb_reg_inst[31:20]),
    .io_rw_cmd({ csr_io_rw_cmd[2], wb_ctrl_csr[1:0] }),
    .io_rw_rdata(csr_io_rw_rdata),
    .io_rw_wdata(wb_reg_wdata),
    .io_singleStep(csr_io_singleStep),
    .io_status_cease(csr_io_status_cease),
    .io_status_debug(bpu_io_status_debug),
    .io_status_dprv(csr_io_status_dprv),
    .io_status_dv(csr_io_status_dv),
    .io_status_fs(csr_io_status_fs),
    .io_status_gva(csr_io_status_gva),
    .io_status_hie(csr_io_status_hie),
    .io_status_isa(csr_io_status_isa),
    .io_status_mbe(csr_io_status_mbe),
    .io_status_mie(csr_io_status_mie),
    .io_status_mpie(csr_io_status_mpie),
    .io_status_mpp(csr_io_status_mpp),
    .io_status_mprv(csr_io_status_mprv),
    .io_status_mpv(csr_io_status_mpv),
    .io_status_mxr(csr_io_status_mxr),
    .io_status_prv(csr_io_status_prv),
    .io_status_sbe(csr_io_status_sbe),
    .io_status_sd(csr_io_status_sd),
    .io_status_sd_rv32(csr_io_status_sd_rv32),
    .io_status_sie(csr_io_status_sie),
    .io_status_spie(csr_io_status_spie),
    .io_status_spp(csr_io_status_spp),
    .io_status_sum(csr_io_status_sum),
    .io_status_sxl(csr_io_status_sxl),
    .io_status_tsr(csr_io_status_tsr),
    .io_status_tvm(csr_io_status_tvm),
    .io_status_tw(csr_io_status_tw),
    .io_status_ube(csr_io_status_ube),
    .io_status_uie(csr_io_status_uie),
    .io_status_upie(csr_io_status_upie),
    .io_status_uxl(csr_io_status_uxl),
    .io_status_v(csr_io_status_v),
    .io_status_vs(csr_io_status_vs),
    .io_status_wfi(csr_io_status_wfi),
    .io_status_xs(csr_io_status_xs),
    .io_status_zero1(csr_io_status_zero1),
    .io_status_zero2(csr_io_status_zero2),
    .io_time(csr_io_time),
    .io_trace_0_exception(csr_io_trace_0_exception),
    .io_trace_0_iaddr(csr_io_trace_0_iaddr),
    .io_trace_0_insn(csr_io_trace_0_insn),
    .io_trace_0_valid(csr_io_trace_0_valid),
    .io_tval(csr_io_tval),
    .io_ungated_clock(clock),
    .reset(reset)
  );
  MulDiv div (
    .clock(clock),
    .io_kill(div_io_kill),
    .io_req_bits_fn(ex_ctrl_alu_fn),
    .io_req_bits_in1(_ex_op1_T),
    .io_req_bits_in2(_ex_op2_T),
    .io_req_bits_tag(ex_reg_inst[11:7]),
    .io_req_ready(div_io_req_ready),
    .io_req_valid(div_io_req_valid),
    .io_resp_bits_data(div_io_resp_bits_data),
    .io_resp_bits_tag(div_io_resp_bits_tag),
    .io_resp_ready(div_io_resp_ready),
    .io_resp_valid(div_io_resp_valid),
    .reset(reset)
  );
  DFF_X1 \div_io_kill_REG$_DFF_P_  (
    .CK(clock),
    .D(_00001_),
    .Q(div_io_kill_REG),
    .QN(_15553_)
  );
  DFF_X1 \ex_ctrl_alu_fn[0]$_SDFFCE_PP0N_  (
    .CK(clock),
    .D(_00565_),
    .Q(ex_ctrl_alu_fn[0]),
    .QN(_15037_)
  );
  DFF_X1 \ex_ctrl_alu_fn[1]$_SDFFCE_PP0N_  (
    .CK(clock),
    .D(_00566_),
    .Q(ex_ctrl_alu_fn[1]),
    .QN(_15036_)
  );
  DFF_X1 \ex_ctrl_alu_fn[2]$_SDFFCE_PP0N_  (
    .CK(clock),
    .D(_00567_),
    .Q(ex_ctrl_alu_fn[2]),
    .QN(_15035_)
  );
  DFF_X1 \ex_ctrl_alu_fn[3]$_SDFFCE_PP0N_  (
    .CK(clock),
    .D(_00568_),
    .Q(ex_ctrl_alu_fn[3]),
    .QN(_15034_)
  );
  DFF_X1 \ex_ctrl_branch$_DFFE_PN_  (
    .CK(clock),
    .D(_00579_),
    .Q(ex_ctrl_branch),
    .QN(_15029_)
  );
  DFF_X1 \ex_ctrl_csr[0]$_SDFFCE_PP0N_  (
    .CK(clock),
    .D(_00589_),
    .Q(ex_ctrl_csr[0]),
    .QN(_15020_)
  );
  DFF_X1 \ex_ctrl_csr[1]$_SDFFCE_PP0N_  (
    .CK(clock),
    .D(_00557_),
    .Q(ex_ctrl_csr[1]),
    .QN(_15041_)
  );
  DFF_X1 \ex_ctrl_csr[2]$_SDFFCE_PP0N_  (
    .CK(clock),
    .D(_00590_),
    .Q(ex_ctrl_csr[2]),
    .QN(_15019_)
  );
  DFF_X1 \ex_ctrl_div$_DFFE_PN_  (
    .CK(clock),
    .D(_00560_),
    .Q(ex_ctrl_div),
    .QN(_15038_)
  );
  DFF_X1 \ex_ctrl_fence_i$_DFFE_PN_  (
    .CK(clock),
    .D(_00558_),
    .Q(ex_ctrl_fence_i),
    .QN(_15040_)
  );
  DFF_X1 \ex_ctrl_jal$_DFFE_PN_  (
    .CK(clock),
    .D(_00578_),
    .Q(ex_ctrl_jal),
    .QN(_15030_)
  );
  DFF_X1 \ex_ctrl_jalr$_DFFE_PN_  (
    .CK(clock),
    .D(_00577_),
    .Q(ex_ctrl_jalr),
    .QN(_15031_)
  );
  DFF_X1 \ex_ctrl_mem$_DFFE_PN_  (
    .CK(clock),
    .D(_00569_),
    .Q(ex_ctrl_mem),
    .QN(_15033_)
  );
  DFF_X1 \ex_ctrl_mem_cmd[0]$_DFFE_PN_  (
    .CK(clock),
    .D(_00561_),
    .Q(ex_ctrl_mem_cmd[0]),
    .QN(_00027_)
  );
  DFF_X1 \ex_ctrl_mem_cmd[1]$_DFFE_PN_  (
    .CK(clock),
    .D(_00562_),
    .Q(ex_ctrl_mem_cmd[1]),
    .QN(_00026_)
  );
  DFF_X1 \ex_ctrl_mem_cmd[2]$_DFFE_PN_  (
    .CK(clock),
    .D(_00563_),
    .Q(ex_ctrl_mem_cmd[2]),
    .QN(_00025_)
  );
  DFF_X1 \ex_ctrl_mem_cmd[3]$_DFFE_PN_  (
    .CK(clock),
    .D(_00564_),
    .Q(ex_ctrl_mem_cmd[3]),
    .QN(_00024_)
  );
  DFF_X1 \ex_ctrl_rxs2$_DFFE_PN_  (
    .CK(clock),
    .D(_00576_),
    .Q(ex_ctrl_rxs2),
    .QN(_15032_)
  );
  DFF_X1 \ex_ctrl_sel_alu1[0]$_DFFE_PN_  (
    .CK(clock),
    .D(_00573_),
    .Q(ex_ctrl_sel_alu1[0]),
    .QN(_00020_)
  );
  DFF_X1 \ex_ctrl_sel_alu1[1]$_DFFE_PN_  (
    .CK(clock),
    .D(_00574_),
    .Q(ex_ctrl_sel_alu1[1]),
    .QN(_00019_)
  );
  DFF_X1 \ex_ctrl_sel_alu2[0]$_DFFE_PN_  (
    .CK(clock),
    .D(_00575_),
    .Q(ex_ctrl_sel_alu2[0]),
    .QN(_00018_)
  );
  DFF_X1 \ex_ctrl_sel_alu2[1]$_SDFFCE_PP0N_  (
    .CK(clock),
    .D(_00747_),
    .Q(ex_ctrl_sel_alu2[1]),
    .QN(_00012_)
  );
  DFF_X1 \ex_ctrl_sel_imm[0]$_DFFE_PN_  (
    .CK(clock),
    .D(_00570_),
    .Q(ex_ctrl_sel_imm[0]),
    .QN(_00023_)
  );
  DFF_X1 \ex_ctrl_sel_imm[1]$_DFFE_PN_  (
    .CK(clock),
    .D(_00571_),
    .Q(ex_ctrl_sel_imm[1]),
    .QN(_00022_)
  );
  DFF_X1 \ex_ctrl_sel_imm[2]$_DFFE_PN_  (
    .CK(clock),
    .D(_00572_),
    .Q(ex_ctrl_sel_imm[2]),
    .QN(_00021_)
  );
  DFF_X1 \ex_ctrl_wxd$_DFFE_PN_  (
    .CK(clock),
    .D(_00559_),
    .Q(ex_ctrl_wxd),
    .QN(_15039_)
  );
  DFF_X1 \ex_reg_cause[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00584_),
    .Q(ex_reg_cause[0]),
    .QN(_15025_)
  );
  DFF_X1 \ex_reg_cause[10]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00463_),
    .Q(ex_reg_cause[10]),
    .QN(_15133_)
  );
  DFF_X1 \ex_reg_cause[11]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00464_),
    .Q(ex_reg_cause[11]),
    .QN(_15132_)
  );
  DFF_X1 \ex_reg_cause[12]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00465_),
    .Q(ex_reg_cause[12]),
    .QN(_15131_)
  );
  DFF_X1 \ex_reg_cause[13]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00466_),
    .Q(ex_reg_cause[13]),
    .QN(_15130_)
  );
  DFF_X1 \ex_reg_cause[14]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00467_),
    .Q(ex_reg_cause[14]),
    .QN(_15129_)
  );
  DFF_X1 \ex_reg_cause[15]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00468_),
    .Q(ex_reg_cause[15]),
    .QN(_15128_)
  );
  DFF_X1 \ex_reg_cause[16]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00469_),
    .Q(ex_reg_cause[16]),
    .QN(_15127_)
  );
  DFF_X1 \ex_reg_cause[17]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00470_),
    .Q(ex_reg_cause[17]),
    .QN(_15126_)
  );
  DFF_X1 \ex_reg_cause[18]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00471_),
    .Q(ex_reg_cause[18]),
    .QN(_15125_)
  );
  DFF_X1 \ex_reg_cause[19]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00472_),
    .Q(ex_reg_cause[19]),
    .QN(_15124_)
  );
  DFF_X1 \ex_reg_cause[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00585_),
    .Q(ex_reg_cause[1]),
    .QN(_15024_)
  );
  DFF_X1 \ex_reg_cause[20]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00473_),
    .Q(ex_reg_cause[20]),
    .QN(_15123_)
  );
  DFF_X1 \ex_reg_cause[21]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00474_),
    .Q(ex_reg_cause[21]),
    .QN(_15122_)
  );
  DFF_X1 \ex_reg_cause[22]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00475_),
    .Q(ex_reg_cause[22]),
    .QN(_15121_)
  );
  DFF_X1 \ex_reg_cause[23]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00476_),
    .Q(ex_reg_cause[23]),
    .QN(_15120_)
  );
  DFF_X1 \ex_reg_cause[24]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00477_),
    .Q(ex_reg_cause[24]),
    .QN(_15119_)
  );
  DFF_X1 \ex_reg_cause[25]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00478_),
    .Q(ex_reg_cause[25]),
    .QN(_15118_)
  );
  DFF_X1 \ex_reg_cause[26]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00479_),
    .Q(ex_reg_cause[26]),
    .QN(_15117_)
  );
  DFF_X1 \ex_reg_cause[27]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00480_),
    .Q(ex_reg_cause[27]),
    .QN(_15116_)
  );
  DFF_X1 \ex_reg_cause[28]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00481_),
    .Q(ex_reg_cause[28]),
    .QN(_15115_)
  );
  DFF_X1 \ex_reg_cause[29]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00482_),
    .Q(ex_reg_cause[29]),
    .QN(_15114_)
  );
  DFF_X1 \ex_reg_cause[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00586_),
    .Q(ex_reg_cause[2]),
    .QN(_15023_)
  );
  DFF_X1 \ex_reg_cause[30]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00483_),
    .Q(ex_reg_cause[30]),
    .QN(_15113_)
  );
  DFF_X1 \ex_reg_cause[31]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00484_),
    .Q(ex_reg_cause[31]),
    .QN(_15112_)
  );
  DFF_X1 \ex_reg_cause[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00587_),
    .Q(ex_reg_cause[3]),
    .QN(_15022_)
  );
  DFF_X1 \ex_reg_cause[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00588_),
    .Q(ex_reg_cause[4]),
    .QN(_15021_)
  );
  DFF_X1 \ex_reg_cause[5]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00458_),
    .Q(ex_reg_cause[5]),
    .QN(_15138_)
  );
  DFF_X1 \ex_reg_cause[6]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00459_),
    .Q(ex_reg_cause[6]),
    .QN(_15137_)
  );
  DFF_X1 \ex_reg_cause[7]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00460_),
    .Q(ex_reg_cause[7]),
    .QN(_15136_)
  );
  DFF_X1 \ex_reg_cause[8]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00461_),
    .Q(ex_reg_cause[8]),
    .QN(_15135_)
  );
  DFF_X1 \ex_reg_cause[9]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00462_),
    .Q(ex_reg_cause[9]),
    .QN(_15134_)
  );
  DFF_X1 \ex_reg_flush_pipe$_DFFE_PN_  (
    .CK(clock),
    .D(_00518_),
    .Q(ex_reg_flush_pipe),
    .QN(_15561_)
  );
  DFF_X1 \ex_reg_inst[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00434_),
    .Q(ex_reg_inst[10]),
    .QN(_15160_)
  );
  DFF_X1 \ex_reg_inst[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00435_),
    .Q(ex_reg_inst[11]),
    .QN(_15159_)
  );
  DFF_X1 \ex_reg_inst[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00436_),
    .Q(ex_reg_inst[12]),
    .QN(_15158_)
  );
  DFF_X1 \ex_reg_inst[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00437_),
    .Q(ex_reg_inst[13]),
    .QN(_15157_)
  );
  DFF_X1 \ex_reg_inst[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00438_),
    .Q(ex_reg_inst[14]),
    .QN(io_dmem_req_bits_signed)
  );
  DFF_X1 \ex_reg_inst[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00439_),
    .Q(ex_reg_inst[15]),
    .QN(_15156_)
  );
  DFF_X1 \ex_reg_inst[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00440_),
    .Q(ex_reg_inst[16]),
    .QN(_15155_)
  );
  DFF_X1 \ex_reg_inst[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00441_),
    .Q(ex_reg_inst[17]),
    .QN(_15154_)
  );
  DFF_X1 \ex_reg_inst[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00442_),
    .Q(ex_reg_inst[18]),
    .QN(_15153_)
  );
  DFF_X1 \ex_reg_inst[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00443_),
    .Q(ex_reg_inst[19]),
    .QN(_15152_)
  );
  DFF_X1 \ex_reg_inst[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00444_),
    .Q(ex_reg_inst[20]),
    .QN(_15151_)
  );
  DFF_X1 \ex_reg_inst[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00445_),
    .Q(ex_reg_inst[21]),
    .QN(_15150_)
  );
  DFF_X1 \ex_reg_inst[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00446_),
    .Q(ex_reg_inst[22]),
    .QN(_15149_)
  );
  DFF_X1 \ex_reg_inst[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00447_),
    .Q(ex_reg_inst[23]),
    .QN(_15148_)
  );
  DFF_X1 \ex_reg_inst[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00448_),
    .Q(ex_reg_inst[24]),
    .QN(_15147_)
  );
  DFF_X1 \ex_reg_inst[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00449_),
    .Q(ex_reg_inst[25]),
    .QN(_15146_)
  );
  DFF_X1 \ex_reg_inst[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00450_),
    .Q(ex_reg_inst[26]),
    .QN(_15145_)
  );
  DFF_X1 \ex_reg_inst[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00451_),
    .Q(ex_reg_inst[27]),
    .QN(_15144_)
  );
  DFF_X1 \ex_reg_inst[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00452_),
    .Q(ex_reg_inst[28]),
    .QN(_15143_)
  );
  DFF_X1 \ex_reg_inst[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00453_),
    .Q(ex_reg_inst[29]),
    .QN(_15142_)
  );
  DFF_X1 \ex_reg_inst[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00454_),
    .Q(ex_reg_inst[30]),
    .QN(_15141_)
  );
  DFF_X1 \ex_reg_inst[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00455_),
    .Q(ex_reg_inst[31]),
    .QN(_15140_)
  );
  DFF_X1 \ex_reg_inst[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00431_),
    .Q(ex_reg_inst[7]),
    .QN(_15163_)
  );
  DFF_X1 \ex_reg_inst[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00432_),
    .Q(ex_reg_inst[8]),
    .QN(_15162_)
  );
  DFF_X1 \ex_reg_inst[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00433_),
    .Q(ex_reg_inst[9]),
    .QN(_15161_)
  );
  DFF_X1 \ex_reg_load_use$_DFFE_PN_  (
    .CK(clock),
    .D(_00517_),
    .Q(ex_reg_load_use),
    .QN(_15560_)
  );
  DFF_X1 \ex_reg_mem_size[0]$_DFFE_PN_  (
    .CK(clock),
    .D(_00456_),
    .Q(ex_reg_mem_size[0]),
    .QN(_15563_[0])
  );
  DFF_X1 \ex_reg_mem_size[1]$_DFFE_PN_  (
    .CK(clock),
    .D(_00457_),
    .Q(ex_reg_mem_size[1]),
    .QN(_15564_[1])
  );
  DFF_X1 \ex_reg_pc[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00485_),
    .Q(ex_reg_pc[0]),
    .QN(_15111_)
  );
  DFF_X1 \ex_reg_pc[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00495_),
    .Q(ex_reg_pc[10]),
    .QN(_15101_)
  );
  DFF_X1 \ex_reg_pc[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00496_),
    .Q(ex_reg_pc[11]),
    .QN(_15100_)
  );
  DFF_X1 \ex_reg_pc[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00497_),
    .Q(ex_reg_pc[12]),
    .QN(_15099_)
  );
  DFF_X1 \ex_reg_pc[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00498_),
    .Q(ex_reg_pc[13]),
    .QN(_15098_)
  );
  DFF_X1 \ex_reg_pc[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00499_),
    .Q(ex_reg_pc[14]),
    .QN(_15097_)
  );
  DFF_X1 \ex_reg_pc[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00500_),
    .Q(ex_reg_pc[15]),
    .QN(_15096_)
  );
  DFF_X1 \ex_reg_pc[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00501_),
    .Q(ex_reg_pc[16]),
    .QN(_15095_)
  );
  DFF_X1 \ex_reg_pc[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00502_),
    .Q(ex_reg_pc[17]),
    .QN(_15094_)
  );
  DFF_X1 \ex_reg_pc[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00503_),
    .Q(ex_reg_pc[18]),
    .QN(_15093_)
  );
  DFF_X1 \ex_reg_pc[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00504_),
    .Q(ex_reg_pc[19]),
    .QN(_15092_)
  );
  DFF_X1 \ex_reg_pc[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00486_),
    .Q(ex_reg_pc[1]),
    .QN(_15110_)
  );
  DFF_X1 \ex_reg_pc[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00505_),
    .Q(ex_reg_pc[20]),
    .QN(_15091_)
  );
  DFF_X1 \ex_reg_pc[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00506_),
    .Q(ex_reg_pc[21]),
    .QN(_15090_)
  );
  DFF_X1 \ex_reg_pc[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00507_),
    .Q(ex_reg_pc[22]),
    .QN(_15089_)
  );
  DFF_X1 \ex_reg_pc[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00508_),
    .Q(ex_reg_pc[23]),
    .QN(_15088_)
  );
  DFF_X1 \ex_reg_pc[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00509_),
    .Q(ex_reg_pc[24]),
    .QN(_15087_)
  );
  DFF_X1 \ex_reg_pc[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00510_),
    .Q(ex_reg_pc[25]),
    .QN(_15086_)
  );
  DFF_X1 \ex_reg_pc[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00511_),
    .Q(ex_reg_pc[26]),
    .QN(_15085_)
  );
  DFF_X1 \ex_reg_pc[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00512_),
    .Q(ex_reg_pc[27]),
    .QN(_15084_)
  );
  DFF_X1 \ex_reg_pc[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00513_),
    .Q(ex_reg_pc[28]),
    .QN(_15083_)
  );
  DFF_X1 \ex_reg_pc[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00514_),
    .Q(ex_reg_pc[29]),
    .QN(_15082_)
  );
  DFF_X1 \ex_reg_pc[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00487_),
    .Q(ex_reg_pc[2]),
    .QN(_15109_)
  );
  DFF_X1 \ex_reg_pc[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00515_),
    .Q(ex_reg_pc[30]),
    .QN(_15081_)
  );
  DFF_X1 \ex_reg_pc[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00516_),
    .Q(ex_reg_pc[31]),
    .QN(_15080_)
  );
  DFF_X1 \ex_reg_pc[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00488_),
    .Q(ex_reg_pc[3]),
    .QN(_15108_)
  );
  DFF_X1 \ex_reg_pc[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00489_),
    .Q(ex_reg_pc[4]),
    .QN(_15107_)
  );
  DFF_X1 \ex_reg_pc[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00490_),
    .Q(ex_reg_pc[5]),
    .QN(_15106_)
  );
  DFF_X1 \ex_reg_pc[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00491_),
    .Q(ex_reg_pc[6]),
    .QN(_15105_)
  );
  DFF_X1 \ex_reg_pc[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00492_),
    .Q(ex_reg_pc[7]),
    .QN(_15104_)
  );
  DFF_X1 \ex_reg_pc[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00493_),
    .Q(ex_reg_pc[8]),
    .QN(_15103_)
  );
  DFF_X1 \ex_reg_pc[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00494_),
    .Q(ex_reg_pc[9]),
    .QN(_15102_)
  );
  DFF_X1 \ex_reg_raw_inst[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00415_),
    .Q(ex_reg_raw_inst[0]),
    .QN(_15179_)
  );
  DFF_X1 \ex_reg_raw_inst[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00425_),
    .Q(ex_reg_raw_inst[10]),
    .QN(_15169_)
  );
  DFF_X1 \ex_reg_raw_inst[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00426_),
    .Q(ex_reg_raw_inst[11]),
    .QN(_15168_)
  );
  DFF_X1 \ex_reg_raw_inst[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00427_),
    .Q(ex_reg_raw_inst[12]),
    .QN(_15167_)
  );
  DFF_X1 \ex_reg_raw_inst[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00428_),
    .Q(ex_reg_raw_inst[13]),
    .QN(_15166_)
  );
  DFF_X1 \ex_reg_raw_inst[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00429_),
    .Q(ex_reg_raw_inst[14]),
    .QN(_15165_)
  );
  DFF_X1 \ex_reg_raw_inst[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00430_),
    .Q(ex_reg_raw_inst[15]),
    .QN(_15164_)
  );
  DFF_X1 \ex_reg_raw_inst[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00416_),
    .Q(ex_reg_raw_inst[1]),
    .QN(_15178_)
  );
  DFF_X1 \ex_reg_raw_inst[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00417_),
    .Q(ex_reg_raw_inst[2]),
    .QN(_15177_)
  );
  DFF_X1 \ex_reg_raw_inst[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00418_),
    .Q(ex_reg_raw_inst[3]),
    .QN(_15176_)
  );
  DFF_X1 \ex_reg_raw_inst[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00419_),
    .Q(ex_reg_raw_inst[4]),
    .QN(_15175_)
  );
  DFF_X1 \ex_reg_raw_inst[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00420_),
    .Q(ex_reg_raw_inst[5]),
    .QN(_15174_)
  );
  DFF_X1 \ex_reg_raw_inst[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00421_),
    .Q(ex_reg_raw_inst[6]),
    .QN(_15173_)
  );
  DFF_X1 \ex_reg_raw_inst[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00422_),
    .Q(ex_reg_raw_inst[7]),
    .QN(_15172_)
  );
  DFF_X1 \ex_reg_raw_inst[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00423_),
    .Q(ex_reg_raw_inst[8]),
    .QN(_15171_)
  );
  DFF_X1 \ex_reg_raw_inst[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00424_),
    .Q(ex_reg_raw_inst[9]),
    .QN(_15170_)
  );
  DFF_X1 \ex_reg_replay$_DFF_P_  (
    .CK(clock),
    .D(_00002_),
    .Q(ex_reg_replay),
    .QN(_15139_)
  );
  DFF_X1 \ex_reg_rs_bypass_0$_SDFFCE_PP0N_  (
    .CK(clock),
    .D(_00100_),
    .Q(ex_reg_rs_bypass_0),
    .QN(_15490_)
  );
  DFF_X1 \ex_reg_rs_bypass_1$_DFFE_PN_  (
    .CK(clock),
    .D(_00099_),
    .Q(ex_reg_rs_bypass_1),
    .QN(_15491_)
  );
  DFF_X1 \ex_reg_rs_lsb_0[0]$_DFFE_PN_  (
    .CK(clock),
    .D(_00097_),
    .Q(ex_reg_rs_lsb_0[0]),
    .QN(_00032_)
  );
  DFF_X1 \ex_reg_rs_lsb_0[1]$_DFFE_PN_  (
    .CK(clock),
    .D(_00098_),
    .Q(ex_reg_rs_lsb_0[1]),
    .QN(_00031_)
  );
  DFF_X1 \ex_reg_rs_lsb_1[0]$_DFFE_PN_  (
    .CK(clock),
    .D(_00580_),
    .Q(ex_reg_rs_lsb_1[0]),
    .QN(_00017_)
  );
  DFF_X1 \ex_reg_rs_lsb_1[1]$_DFFE_PN_  (
    .CK(clock),
    .D(_00581_),
    .Q(ex_reg_rs_lsb_1[1]),
    .QN(_00035_)
  );
  DFF_X1 \ex_reg_rs_msb_0[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00067_),
    .Q(ex_reg_rs_msb_0[0]),
    .QN(_15521_)
  );
  DFF_X1 \ex_reg_rs_msb_0[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00077_),
    .Q(ex_reg_rs_msb_0[10]),
    .QN(_15511_)
  );
  DFF_X1 \ex_reg_rs_msb_0[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00078_),
    .Q(ex_reg_rs_msb_0[11]),
    .QN(_15510_)
  );
  DFF_X1 \ex_reg_rs_msb_0[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00079_),
    .Q(ex_reg_rs_msb_0[12]),
    .QN(_15509_)
  );
  DFF_X1 \ex_reg_rs_msb_0[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00080_),
    .Q(ex_reg_rs_msb_0[13]),
    .QN(_15508_)
  );
  DFF_X1 \ex_reg_rs_msb_0[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00081_),
    .Q(ex_reg_rs_msb_0[14]),
    .QN(_15507_)
  );
  DFF_X1 \ex_reg_rs_msb_0[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00082_),
    .Q(ex_reg_rs_msb_0[15]),
    .QN(_15506_)
  );
  DFF_X1 \ex_reg_rs_msb_0[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00083_),
    .Q(ex_reg_rs_msb_0[16]),
    .QN(_15505_)
  );
  DFF_X1 \ex_reg_rs_msb_0[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00084_),
    .Q(ex_reg_rs_msb_0[17]),
    .QN(_15504_)
  );
  DFF_X1 \ex_reg_rs_msb_0[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00085_),
    .Q(ex_reg_rs_msb_0[18]),
    .QN(_15503_)
  );
  DFF_X1 \ex_reg_rs_msb_0[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00086_),
    .Q(ex_reg_rs_msb_0[19]),
    .QN(_15502_)
  );
  DFF_X1 \ex_reg_rs_msb_0[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00068_),
    .Q(ex_reg_rs_msb_0[1]),
    .QN(_15520_)
  );
  DFF_X1 \ex_reg_rs_msb_0[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00087_),
    .Q(ex_reg_rs_msb_0[20]),
    .QN(_15501_)
  );
  DFF_X1 \ex_reg_rs_msb_0[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00088_),
    .Q(ex_reg_rs_msb_0[21]),
    .QN(_15500_)
  );
  DFF_X1 \ex_reg_rs_msb_0[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00089_),
    .Q(ex_reg_rs_msb_0[22]),
    .QN(_15499_)
  );
  DFF_X1 \ex_reg_rs_msb_0[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00090_),
    .Q(ex_reg_rs_msb_0[23]),
    .QN(_15498_)
  );
  DFF_X1 \ex_reg_rs_msb_0[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00091_),
    .Q(ex_reg_rs_msb_0[24]),
    .QN(_15497_)
  );
  DFF_X1 \ex_reg_rs_msb_0[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00092_),
    .Q(ex_reg_rs_msb_0[25]),
    .QN(_15496_)
  );
  DFF_X1 \ex_reg_rs_msb_0[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00093_),
    .Q(ex_reg_rs_msb_0[26]),
    .QN(_15495_)
  );
  DFF_X1 \ex_reg_rs_msb_0[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00094_),
    .Q(ex_reg_rs_msb_0[27]),
    .QN(_15494_)
  );
  DFF_X1 \ex_reg_rs_msb_0[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00095_),
    .Q(ex_reg_rs_msb_0[28]),
    .QN(_15493_)
  );
  DFF_X1 \ex_reg_rs_msb_0[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00096_),
    .Q(ex_reg_rs_msb_0[29]),
    .QN(_15492_)
  );
  DFF_X1 \ex_reg_rs_msb_0[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00069_),
    .Q(ex_reg_rs_msb_0[2]),
    .QN(_15519_)
  );
  DFF_X1 \ex_reg_rs_msb_0[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00070_),
    .Q(ex_reg_rs_msb_0[3]),
    .QN(_15518_)
  );
  DFF_X1 \ex_reg_rs_msb_0[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00071_),
    .Q(ex_reg_rs_msb_0[4]),
    .QN(_15517_)
  );
  DFF_X1 \ex_reg_rs_msb_0[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00072_),
    .Q(ex_reg_rs_msb_0[5]),
    .QN(_15516_)
  );
  DFF_X1 \ex_reg_rs_msb_0[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00073_),
    .Q(ex_reg_rs_msb_0[6]),
    .QN(_15515_)
  );
  DFF_X1 \ex_reg_rs_msb_0[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00074_),
    .Q(ex_reg_rs_msb_0[7]),
    .QN(_15514_)
  );
  DFF_X1 \ex_reg_rs_msb_0[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00075_),
    .Q(ex_reg_rs_msb_0[8]),
    .QN(_15513_)
  );
  DFF_X1 \ex_reg_rs_msb_0[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00076_),
    .Q(ex_reg_rs_msb_0[9]),
    .QN(_15512_)
  );
  DFF_X1 \ex_reg_rs_msb_1[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00149_),
    .Q(ex_reg_rs_msb_1[0]),
    .QN(_15441_)
  );
  DFF_X1 \ex_reg_rs_msb_1[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00159_),
    .Q(ex_reg_rs_msb_1[10]),
    .QN(_15431_)
  );
  DFF_X1 \ex_reg_rs_msb_1[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00160_),
    .Q(ex_reg_rs_msb_1[11]),
    .QN(_15430_)
  );
  DFF_X1 \ex_reg_rs_msb_1[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00161_),
    .Q(ex_reg_rs_msb_1[12]),
    .QN(_15429_)
  );
  DFF_X1 \ex_reg_rs_msb_1[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00162_),
    .Q(ex_reg_rs_msb_1[13]),
    .QN(_15428_)
  );
  DFF_X1 \ex_reg_rs_msb_1[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00163_),
    .Q(ex_reg_rs_msb_1[14]),
    .QN(_15427_)
  );
  DFF_X1 \ex_reg_rs_msb_1[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00164_),
    .Q(ex_reg_rs_msb_1[15]),
    .QN(_15426_)
  );
  DFF_X1 \ex_reg_rs_msb_1[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00165_),
    .Q(ex_reg_rs_msb_1[16]),
    .QN(_15425_)
  );
  DFF_X1 \ex_reg_rs_msb_1[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00166_),
    .Q(ex_reg_rs_msb_1[17]),
    .QN(_15424_)
  );
  DFF_X1 \ex_reg_rs_msb_1[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00167_),
    .Q(ex_reg_rs_msb_1[18]),
    .QN(_15423_)
  );
  DFF_X1 \ex_reg_rs_msb_1[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00168_),
    .Q(ex_reg_rs_msb_1[19]),
    .QN(_15422_)
  );
  DFF_X1 \ex_reg_rs_msb_1[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00150_),
    .Q(ex_reg_rs_msb_1[1]),
    .QN(_15440_)
  );
  DFF_X1 \ex_reg_rs_msb_1[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00169_),
    .Q(ex_reg_rs_msb_1[20]),
    .QN(_15421_)
  );
  DFF_X1 \ex_reg_rs_msb_1[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00170_),
    .Q(ex_reg_rs_msb_1[21]),
    .QN(_15420_)
  );
  DFF_X1 \ex_reg_rs_msb_1[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00171_),
    .Q(ex_reg_rs_msb_1[22]),
    .QN(_15419_)
  );
  DFF_X1 \ex_reg_rs_msb_1[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00172_),
    .Q(ex_reg_rs_msb_1[23]),
    .QN(_15418_)
  );
  DFF_X1 \ex_reg_rs_msb_1[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00173_),
    .Q(ex_reg_rs_msb_1[24]),
    .QN(_15417_)
  );
  DFF_X1 \ex_reg_rs_msb_1[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00174_),
    .Q(ex_reg_rs_msb_1[25]),
    .QN(_15416_)
  );
  DFF_X1 \ex_reg_rs_msb_1[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00175_),
    .Q(ex_reg_rs_msb_1[26]),
    .QN(_15415_)
  );
  DFF_X1 \ex_reg_rs_msb_1[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00176_),
    .Q(ex_reg_rs_msb_1[27]),
    .QN(_15414_)
  );
  DFF_X1 \ex_reg_rs_msb_1[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00177_),
    .Q(ex_reg_rs_msb_1[28]),
    .QN(_15413_)
  );
  DFF_X1 \ex_reg_rs_msb_1[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00178_),
    .Q(ex_reg_rs_msb_1[29]),
    .QN(_15412_)
  );
  DFF_X1 \ex_reg_rs_msb_1[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00151_),
    .Q(ex_reg_rs_msb_1[2]),
    .QN(_15439_)
  );
  DFF_X1 \ex_reg_rs_msb_1[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00152_),
    .Q(ex_reg_rs_msb_1[3]),
    .QN(_15438_)
  );
  DFF_X1 \ex_reg_rs_msb_1[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00153_),
    .Q(ex_reg_rs_msb_1[4]),
    .QN(_15437_)
  );
  DFF_X1 \ex_reg_rs_msb_1[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00154_),
    .Q(ex_reg_rs_msb_1[5]),
    .QN(_15436_)
  );
  DFF_X1 \ex_reg_rs_msb_1[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00155_),
    .Q(ex_reg_rs_msb_1[6]),
    .QN(_15435_)
  );
  DFF_X1 \ex_reg_rs_msb_1[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00156_),
    .Q(ex_reg_rs_msb_1[7]),
    .QN(_15434_)
  );
  DFF_X1 \ex_reg_rs_msb_1[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00157_),
    .Q(ex_reg_rs_msb_1[8]),
    .QN(_15433_)
  );
  DFF_X1 \ex_reg_rs_msb_1[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00158_),
    .Q(ex_reg_rs_msb_1[9]),
    .QN(_15432_)
  );
  DFF_X1 \ex_reg_rvc$_DFFE_PN_  (
    .CK(clock),
    .D(_00179_),
    .Q(ex_reg_rvc),
    .QN(_ex_op2_T_1[2])
  );
  DFF_X1 \ex_reg_valid$_DFF_P_  (
    .CK(clock),
    .D(_ex_reg_valid_T),
    .Q(ex_reg_valid),
    .QN(_00034_)
  );
  DFF_X1 \ex_reg_xcpt$_DFF_P_  (
    .CK(clock),
    .D(_00003_),
    .Q(ex_reg_xcpt),
    .QN(_15079_)
  );
  DFF_X1 \ex_reg_xcpt_interrupt$_DFF_P_  (
    .CK(clock),
    .D(_00004_),
    .Q(ex_reg_xcpt_interrupt),
    .QN(_15078_)
  );
  IBuf ibuf (
    .clock(clock),
    .io_imem_bits_data(io_imem_resp_bits_data),
    .io_imem_bits_pc(io_imem_resp_bits_pc),
    .io_imem_bits_replay(io_imem_resp_bits_replay),
    .io_imem_bits_xcpt_ae_inst(io_imem_resp_bits_xcpt_ae_inst),
    .io_imem_ready(ibuf_io_imem_ready),
    .io_imem_valid(io_imem_resp_valid),
    .io_inst_0_bits_inst_bits(csr_io_decode_0_inst),
    .io_inst_0_bits_inst_rd(ibuf_io_inst_0_bits_inst_rd),
    .io_inst_0_bits_inst_rs1(ibuf_io_inst_0_bits_inst_rs1),
    .io_inst_0_bits_inst_rs2(ibuf_io_inst_0_bits_inst_rs2),
    .io_inst_0_bits_raw(ibuf_io_inst_0_bits_raw),
    .io_inst_0_bits_replay(ibuf_io_inst_0_bits_replay),
    .io_inst_0_bits_rvc(ibuf_io_inst_0_bits_rvc),
    .io_inst_0_bits_xcpt0_ae_inst(ibuf_io_inst_0_bits_xcpt0_ae_inst),
    .io_inst_0_bits_xcpt1_ae_inst(ibuf_io_inst_0_bits_xcpt1_ae_inst),
    .io_inst_0_bits_xcpt1_gf_inst(ibuf_io_inst_0_bits_xcpt1_gf_inst),
    .io_inst_0_bits_xcpt1_pf_inst(ibuf_io_inst_0_bits_xcpt1_pf_inst),
    .io_inst_0_ready(ibuf_io_inst_0_ready),
    .io_inst_0_valid(ibuf_io_inst_0_valid),
    .io_kill(ibuf_io_kill),
    .io_pc(bpu_io_pc),
    .reset(reset)
  );
  DFF_X1 \id_reg_fence$_SDFF_PP0_  (
    .CK(clock),
    .D(_00583_),
    .Q(id_reg_fence),
    .QN(_15026_)
  );
  DFF_X1 \id_reg_pause$_SDFFE_PP0N_  (
    .CK(clock),
    .D(_00582_),
    .Q(id_reg_pause),
    .QN(_15027_)
  );
  DFF_X1 \imem_might_request_reg$_DFF_P_  (
    .CK(clock),
    .D(_00005_),
    .Q(imem_might_request_reg),
    .QN(_15028_)
  );
  DFF_X1 \mem_br_taken$_DFFE_PP_  (
    .CK(clock),
    .D(_00240_),
    .Q(mem_br_taken),
    .QN(_15352_)
  );
  DFF_X1 \mem_ctrl_branch$_DFFE_PP_  (
    .CK(clock),
    .D(_00556_),
    .Q(mem_ctrl_branch),
    .QN(_15042_)
  );
  DFF_X1 \mem_ctrl_csr[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00548_),
    .Q(mem_ctrl_csr[0]),
    .QN(_15049_)
  );
  DFF_X1 \mem_ctrl_csr[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00549_),
    .Q(mem_ctrl_csr[1]),
    .QN(_15048_)
  );
  DFF_X1 \mem_ctrl_csr[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00550_),
    .Q(mem_ctrl_csr[2]),
    .QN(_15047_)
  );
  DFF_X1 \mem_ctrl_div$_DFFE_PP_  (
    .CK(clock),
    .D(_00552_),
    .Q(mem_ctrl_div),
    .QN(_15045_)
  );
  DFF_X1 \mem_ctrl_fence_i$_DFFE_PP_  (
    .CK(clock),
    .D(_00547_),
    .Q(mem_ctrl_fence_i),
    .QN(_15050_)
  );
  DFF_X1 \mem_ctrl_jal$_DFFE_PP_  (
    .CK(clock),
    .D(_00555_),
    .Q(mem_ctrl_jal),
    .QN(_15043_)
  );
  DFF_X1 \mem_ctrl_jalr$_DFFE_PP_  (
    .CK(clock),
    .D(_00554_),
    .Q(mem_ctrl_jalr),
    .QN(_15044_)
  );
  DFF_X1 \mem_ctrl_mem$_DFFE_PP_  (
    .CK(clock),
    .D(_00553_),
    .Q(mem_ctrl_mem),
    .QN(_00028_)
  );
  DFF_X1 \mem_ctrl_wxd$_DFFE_PP_  (
    .CK(clock),
    .D(_00551_),
    .Q(mem_ctrl_wxd),
    .QN(_15046_)
  );
  DFF_X1 \mem_reg_cause[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00381_),
    .Q(mem_reg_cause[0]),
    .QN(_15211_)
  );
  DFF_X1 \mem_reg_cause[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00391_),
    .Q(mem_reg_cause[10]),
    .QN(_15201_)
  );
  DFF_X1 \mem_reg_cause[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00392_),
    .Q(mem_reg_cause[11]),
    .QN(_15200_)
  );
  DFF_X1 \mem_reg_cause[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00393_),
    .Q(mem_reg_cause[12]),
    .QN(_15199_)
  );
  DFF_X1 \mem_reg_cause[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00394_),
    .Q(mem_reg_cause[13]),
    .QN(_15198_)
  );
  DFF_X1 \mem_reg_cause[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00395_),
    .Q(mem_reg_cause[14]),
    .QN(_15197_)
  );
  DFF_X1 \mem_reg_cause[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00396_),
    .Q(mem_reg_cause[15]),
    .QN(_15196_)
  );
  DFF_X1 \mem_reg_cause[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00397_),
    .Q(mem_reg_cause[16]),
    .QN(_15195_)
  );
  DFF_X1 \mem_reg_cause[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00398_),
    .Q(mem_reg_cause[17]),
    .QN(_15194_)
  );
  DFF_X1 \mem_reg_cause[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00399_),
    .Q(mem_reg_cause[18]),
    .QN(_15193_)
  );
  DFF_X1 \mem_reg_cause[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00400_),
    .Q(mem_reg_cause[19]),
    .QN(_15192_)
  );
  DFF_X1 \mem_reg_cause[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00382_),
    .Q(mem_reg_cause[1]),
    .QN(_15210_)
  );
  DFF_X1 \mem_reg_cause[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00401_),
    .Q(mem_reg_cause[20]),
    .QN(_15191_)
  );
  DFF_X1 \mem_reg_cause[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00402_),
    .Q(mem_reg_cause[21]),
    .QN(_15190_)
  );
  DFF_X1 \mem_reg_cause[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00403_),
    .Q(mem_reg_cause[22]),
    .QN(_15189_)
  );
  DFF_X1 \mem_reg_cause[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00404_),
    .Q(mem_reg_cause[23]),
    .QN(_15188_)
  );
  DFF_X1 \mem_reg_cause[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00405_),
    .Q(mem_reg_cause[24]),
    .QN(_15187_)
  );
  DFF_X1 \mem_reg_cause[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00406_),
    .Q(mem_reg_cause[25]),
    .QN(_15186_)
  );
  DFF_X1 \mem_reg_cause[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00407_),
    .Q(mem_reg_cause[26]),
    .QN(_15185_)
  );
  DFF_X1 \mem_reg_cause[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00408_),
    .Q(mem_reg_cause[27]),
    .QN(_15184_)
  );
  DFF_X1 \mem_reg_cause[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00409_),
    .Q(mem_reg_cause[28]),
    .QN(_15183_)
  );
  DFF_X1 \mem_reg_cause[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00410_),
    .Q(mem_reg_cause[29]),
    .QN(_15182_)
  );
  DFF_X1 \mem_reg_cause[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00383_),
    .Q(mem_reg_cause[2]),
    .QN(_15209_)
  );
  DFF_X1 \mem_reg_cause[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00411_),
    .Q(mem_reg_cause[30]),
    .QN(_15181_)
  );
  DFF_X1 \mem_reg_cause[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00412_),
    .Q(mem_reg_cause[31]),
    .QN(_15557_)
  );
  DFF_X1 \mem_reg_cause[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00384_),
    .Q(mem_reg_cause[3]),
    .QN(_15208_)
  );
  DFF_X1 \mem_reg_cause[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00385_),
    .Q(mem_reg_cause[4]),
    .QN(_15207_)
  );
  DFF_X1 \mem_reg_cause[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00386_),
    .Q(mem_reg_cause[5]),
    .QN(_15206_)
  );
  DFF_X1 \mem_reg_cause[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00387_),
    .Q(mem_reg_cause[6]),
    .QN(_15205_)
  );
  DFF_X1 \mem_reg_cause[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00388_),
    .Q(mem_reg_cause[7]),
    .QN(_15204_)
  );
  DFF_X1 \mem_reg_cause[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00389_),
    .Q(mem_reg_cause[8]),
    .QN(_15203_)
  );
  DFF_X1 \mem_reg_cause[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00390_),
    .Q(mem_reg_cause[9]),
    .QN(_15202_)
  );
  DFF_X1 \mem_reg_flush_pipe$_DFFE_PP_  (
    .CK(clock),
    .D(_00413_),
    .Q(mem_reg_flush_pipe),
    .QN(_15559_)
  );
  DFF_X1 \mem_reg_inst[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00324_),
    .Q(mem_reg_inst[10]),
    .QN(_15268_)
  );
  DFF_X1 \mem_reg_inst[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00325_),
    .Q(mem_reg_inst[11]),
    .QN(_15267_)
  );
  DFF_X1 \mem_reg_inst[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00326_),
    .Q(mem_reg_inst[12]),
    .QN(_15266_)
  );
  DFF_X1 \mem_reg_inst[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00327_),
    .Q(mem_reg_inst[13]),
    .QN(_15265_)
  );
  DFF_X1 \mem_reg_inst[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00328_),
    .Q(mem_reg_inst[14]),
    .QN(_15264_)
  );
  DFF_X1 \mem_reg_inst[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00329_),
    .Q(mem_reg_inst[15]),
    .QN(_15263_)
  );
  DFF_X1 \mem_reg_inst[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00330_),
    .Q(mem_reg_inst[16]),
    .QN(_15262_)
  );
  DFF_X1 \mem_reg_inst[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00331_),
    .Q(mem_reg_inst[17]),
    .QN(_15261_)
  );
  DFF_X1 \mem_reg_inst[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00332_),
    .Q(mem_reg_inst[18]),
    .QN(_15260_)
  );
  DFF_X1 \mem_reg_inst[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00333_),
    .Q(mem_reg_inst[19]),
    .QN(_15259_)
  );
  DFF_X1 \mem_reg_inst[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00334_),
    .Q(mem_reg_inst[20]),
    .QN(_15258_)
  );
  DFF_X1 \mem_reg_inst[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00335_),
    .Q(mem_reg_inst[21]),
    .QN(_15257_)
  );
  DFF_X1 \mem_reg_inst[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00336_),
    .Q(mem_reg_inst[22]),
    .QN(_15256_)
  );
  DFF_X1 \mem_reg_inst[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00337_),
    .Q(mem_reg_inst[23]),
    .QN(_15255_)
  );
  DFF_X1 \mem_reg_inst[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00338_),
    .Q(mem_reg_inst[24]),
    .QN(_15254_)
  );
  DFF_X1 \mem_reg_inst[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00339_),
    .Q(mem_reg_inst[25]),
    .QN(_15253_)
  );
  DFF_X1 \mem_reg_inst[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00340_),
    .Q(mem_reg_inst[26]),
    .QN(_15252_)
  );
  DFF_X1 \mem_reg_inst[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00341_),
    .Q(mem_reg_inst[27]),
    .QN(_15251_)
  );
  DFF_X1 \mem_reg_inst[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00342_),
    .Q(mem_reg_inst[28]),
    .QN(_15250_)
  );
  DFF_X1 \mem_reg_inst[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00343_),
    .Q(mem_reg_inst[29]),
    .QN(_15249_)
  );
  DFF_X1 \mem_reg_inst[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00344_),
    .Q(mem_reg_inst[30]),
    .QN(_15248_)
  );
  DFF_X1 \mem_reg_inst[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00345_),
    .Q(mem_reg_inst[31]),
    .QN(_15247_)
  );
  DFF_X1 \mem_reg_inst[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00321_),
    .Q(mem_reg_inst[7]),
    .QN(_15271_)
  );
  DFF_X1 \mem_reg_inst[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00322_),
    .Q(mem_reg_inst[8]),
    .QN(_15270_)
  );
  DFF_X1 \mem_reg_inst[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00323_),
    .Q(mem_reg_inst[9]),
    .QN(_15269_)
  );
  DFF_X1 \mem_reg_load$_DFFE_PP_  (
    .CK(clock),
    .D(_00379_),
    .Q(mem_reg_load),
    .QN(_15213_)
  );
  DFF_X1 \mem_reg_pc[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00346_),
    .Q(mem_reg_pc[0]),
    .QN(_15246_)
  );
  DFF_X1 \mem_reg_pc[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00356_),
    .Q(mem_reg_pc[10]),
    .QN(_15236_)
  );
  DFF_X1 \mem_reg_pc[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00357_),
    .Q(mem_reg_pc[11]),
    .QN(_15235_)
  );
  DFF_X1 \mem_reg_pc[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00358_),
    .Q(mem_reg_pc[12]),
    .QN(_15234_)
  );
  DFF_X1 \mem_reg_pc[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00359_),
    .Q(mem_reg_pc[13]),
    .QN(_15233_)
  );
  DFF_X1 \mem_reg_pc[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00360_),
    .Q(mem_reg_pc[14]),
    .QN(_15232_)
  );
  DFF_X1 \mem_reg_pc[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00361_),
    .Q(mem_reg_pc[15]),
    .QN(_15231_)
  );
  DFF_X1 \mem_reg_pc[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00362_),
    .Q(mem_reg_pc[16]),
    .QN(_15230_)
  );
  DFF_X1 \mem_reg_pc[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00363_),
    .Q(mem_reg_pc[17]),
    .QN(_15229_)
  );
  DFF_X1 \mem_reg_pc[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00364_),
    .Q(mem_reg_pc[18]),
    .QN(_15228_)
  );
  DFF_X1 \mem_reg_pc[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00365_),
    .Q(mem_reg_pc[19]),
    .QN(_15227_)
  );
  DFF_X1 \mem_reg_pc[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00347_),
    .Q(mem_reg_pc[1]),
    .QN(_15245_)
  );
  DFF_X1 \mem_reg_pc[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00366_),
    .Q(mem_reg_pc[20]),
    .QN(_15226_)
  );
  DFF_X1 \mem_reg_pc[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00367_),
    .Q(mem_reg_pc[21]),
    .QN(_15225_)
  );
  DFF_X1 \mem_reg_pc[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00368_),
    .Q(mem_reg_pc[22]),
    .QN(_15224_)
  );
  DFF_X1 \mem_reg_pc[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00369_),
    .Q(mem_reg_pc[23]),
    .QN(_15223_)
  );
  DFF_X1 \mem_reg_pc[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00370_),
    .Q(mem_reg_pc[24]),
    .QN(_15222_)
  );
  DFF_X1 \mem_reg_pc[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00371_),
    .Q(mem_reg_pc[25]),
    .QN(_15221_)
  );
  DFF_X1 \mem_reg_pc[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00372_),
    .Q(mem_reg_pc[26]),
    .QN(_15220_)
  );
  DFF_X1 \mem_reg_pc[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00373_),
    .Q(mem_reg_pc[27]),
    .QN(_15219_)
  );
  DFF_X1 \mem_reg_pc[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00374_),
    .Q(mem_reg_pc[28]),
    .QN(_15218_)
  );
  DFF_X1 \mem_reg_pc[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00375_),
    .Q(mem_reg_pc[29]),
    .QN(_15217_)
  );
  DFF_X1 \mem_reg_pc[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00348_),
    .Q(mem_reg_pc[2]),
    .QN(_15244_)
  );
  DFF_X1 \mem_reg_pc[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00376_),
    .Q(mem_reg_pc[30]),
    .QN(_15216_)
  );
  DFF_X1 \mem_reg_pc[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00377_),
    .Q(mem_reg_pc[31]),
    .QN(_15215_)
  );
  DFF_X1 \mem_reg_pc[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00349_),
    .Q(mem_reg_pc[3]),
    .QN(_15243_)
  );
  DFF_X1 \mem_reg_pc[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00350_),
    .Q(mem_reg_pc[4]),
    .QN(_15242_)
  );
  DFF_X1 \mem_reg_pc[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00351_),
    .Q(mem_reg_pc[5]),
    .QN(_15241_)
  );
  DFF_X1 \mem_reg_pc[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00352_),
    .Q(mem_reg_pc[6]),
    .QN(_15240_)
  );
  DFF_X1 \mem_reg_pc[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00353_),
    .Q(mem_reg_pc[7]),
    .QN(_15239_)
  );
  DFF_X1 \mem_reg_pc[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00354_),
    .Q(mem_reg_pc[8]),
    .QN(_15238_)
  );
  DFF_X1 \mem_reg_pc[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00355_),
    .Q(mem_reg_pc[9]),
    .QN(_15237_)
  );
  DFF_X1 \mem_reg_raw_inst[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00305_),
    .Q(mem_reg_raw_inst[0]),
    .QN(_15287_)
  );
  DFF_X1 \mem_reg_raw_inst[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00315_),
    .Q(mem_reg_raw_inst[10]),
    .QN(_15277_)
  );
  DFF_X1 \mem_reg_raw_inst[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00316_),
    .Q(mem_reg_raw_inst[11]),
    .QN(_15276_)
  );
  DFF_X1 \mem_reg_raw_inst[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00317_),
    .Q(mem_reg_raw_inst[12]),
    .QN(_15275_)
  );
  DFF_X1 \mem_reg_raw_inst[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00318_),
    .Q(mem_reg_raw_inst[13]),
    .QN(_15274_)
  );
  DFF_X1 \mem_reg_raw_inst[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00319_),
    .Q(mem_reg_raw_inst[14]),
    .QN(_15273_)
  );
  DFF_X1 \mem_reg_raw_inst[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00320_),
    .Q(mem_reg_raw_inst[15]),
    .QN(_15272_)
  );
  DFF_X1 \mem_reg_raw_inst[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00306_),
    .Q(mem_reg_raw_inst[1]),
    .QN(_15286_)
  );
  DFF_X1 \mem_reg_raw_inst[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00307_),
    .Q(mem_reg_raw_inst[2]),
    .QN(_15285_)
  );
  DFF_X1 \mem_reg_raw_inst[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00308_),
    .Q(mem_reg_raw_inst[3]),
    .QN(_15284_)
  );
  DFF_X1 \mem_reg_raw_inst[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00309_),
    .Q(mem_reg_raw_inst[4]),
    .QN(_15283_)
  );
  DFF_X1 \mem_reg_raw_inst[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00310_),
    .Q(mem_reg_raw_inst[5]),
    .QN(_15282_)
  );
  DFF_X1 \mem_reg_raw_inst[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00311_),
    .Q(mem_reg_raw_inst[6]),
    .QN(_15281_)
  );
  DFF_X1 \mem_reg_raw_inst[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00312_),
    .Q(mem_reg_raw_inst[7]),
    .QN(_15280_)
  );
  DFF_X1 \mem_reg_raw_inst[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00313_),
    .Q(mem_reg_raw_inst[8]),
    .QN(_15279_)
  );
  DFF_X1 \mem_reg_raw_inst[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00314_),
    .Q(mem_reg_raw_inst[9]),
    .QN(_15278_)
  );
  DFF_X1 \mem_reg_replay$_DFF_P_  (
    .CK(clock),
    .D(_00006_),
    .Q(mem_reg_replay),
    .QN(_15558_)
  );
  DFF_X1 \mem_reg_rs2[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00241_),
    .Q(mem_reg_rs2[0]),
    .QN(_15351_)
  );
  DFF_X1 \mem_reg_rs2[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00251_),
    .Q(mem_reg_rs2[10]),
    .QN(_15341_)
  );
  DFF_X1 \mem_reg_rs2[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00252_),
    .Q(mem_reg_rs2[11]),
    .QN(_15340_)
  );
  DFF_X1 \mem_reg_rs2[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00253_),
    .Q(mem_reg_rs2[12]),
    .QN(_15339_)
  );
  DFF_X1 \mem_reg_rs2[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00254_),
    .Q(mem_reg_rs2[13]),
    .QN(_15338_)
  );
  DFF_X1 \mem_reg_rs2[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00255_),
    .Q(mem_reg_rs2[14]),
    .QN(_15337_)
  );
  DFF_X1 \mem_reg_rs2[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00256_),
    .Q(mem_reg_rs2[15]),
    .QN(_15336_)
  );
  DFF_X1 \mem_reg_rs2[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00257_),
    .Q(mem_reg_rs2[16]),
    .QN(_15335_)
  );
  DFF_X1 \mem_reg_rs2[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00258_),
    .Q(mem_reg_rs2[17]),
    .QN(_15334_)
  );
  DFF_X1 \mem_reg_rs2[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00259_),
    .Q(mem_reg_rs2[18]),
    .QN(_15333_)
  );
  DFF_X1 \mem_reg_rs2[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00260_),
    .Q(mem_reg_rs2[19]),
    .QN(_15332_)
  );
  DFF_X1 \mem_reg_rs2[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00242_),
    .Q(mem_reg_rs2[1]),
    .QN(_15350_)
  );
  DFF_X1 \mem_reg_rs2[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00261_),
    .Q(mem_reg_rs2[20]),
    .QN(_15331_)
  );
  DFF_X1 \mem_reg_rs2[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00262_),
    .Q(mem_reg_rs2[21]),
    .QN(_15330_)
  );
  DFF_X1 \mem_reg_rs2[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00263_),
    .Q(mem_reg_rs2[22]),
    .QN(_15329_)
  );
  DFF_X1 \mem_reg_rs2[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00264_),
    .Q(mem_reg_rs2[23]),
    .QN(_15328_)
  );
  DFF_X1 \mem_reg_rs2[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00265_),
    .Q(mem_reg_rs2[24]),
    .QN(_15327_)
  );
  DFF_X1 \mem_reg_rs2[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00266_),
    .Q(mem_reg_rs2[25]),
    .QN(_15326_)
  );
  DFF_X1 \mem_reg_rs2[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00267_),
    .Q(mem_reg_rs2[26]),
    .QN(_15325_)
  );
  DFF_X1 \mem_reg_rs2[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00268_),
    .Q(mem_reg_rs2[27]),
    .QN(_15324_)
  );
  DFF_X1 \mem_reg_rs2[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00269_),
    .Q(mem_reg_rs2[28]),
    .QN(_15323_)
  );
  DFF_X1 \mem_reg_rs2[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00270_),
    .Q(mem_reg_rs2[29]),
    .QN(_15322_)
  );
  DFF_X1 \mem_reg_rs2[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00243_),
    .Q(mem_reg_rs2[2]),
    .QN(_15349_)
  );
  DFF_X1 \mem_reg_rs2[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00271_),
    .Q(mem_reg_rs2[30]),
    .QN(_15321_)
  );
  DFF_X1 \mem_reg_rs2[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00272_),
    .Q(mem_reg_rs2[31]),
    .QN(_15320_)
  );
  DFF_X1 \mem_reg_rs2[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00244_),
    .Q(mem_reg_rs2[3]),
    .QN(_15348_)
  );
  DFF_X1 \mem_reg_rs2[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00245_),
    .Q(mem_reg_rs2[4]),
    .QN(_15347_)
  );
  DFF_X1 \mem_reg_rs2[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00246_),
    .Q(mem_reg_rs2[5]),
    .QN(_15346_)
  );
  DFF_X1 \mem_reg_rs2[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00247_),
    .Q(mem_reg_rs2[6]),
    .QN(_15345_)
  );
  DFF_X1 \mem_reg_rs2[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00248_),
    .Q(mem_reg_rs2[7]),
    .QN(_15344_)
  );
  DFF_X1 \mem_reg_rs2[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00249_),
    .Q(mem_reg_rs2[8]),
    .QN(_15343_)
  );
  DFF_X1 \mem_reg_rs2[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00250_),
    .Q(mem_reg_rs2[9]),
    .QN(_15342_)
  );
  DFF_X1 \mem_reg_rvc$_DFFE_PP_  (
    .CK(clock),
    .D(_00414_),
    .Q(mem_reg_rvc),
    .QN(_mem_br_target_T_6[2])
  );
  DFF_X1 \mem_reg_slow_bypass$_DFFE_PP_  (
    .CK(clock),
    .D(_00380_),
    .Q(mem_reg_slow_bypass),
    .QN(_15212_)
  );
  DFF_X1 \mem_reg_store$_DFFE_PP_  (
    .CK(clock),
    .D(_00378_),
    .Q(mem_reg_store),
    .QN(_15214_)
  );
  DFF_X1 \mem_reg_valid$_DFF_P_  (
    .CK(clock),
    .D(_mem_reg_valid_T),
    .Q(mem_reg_valid),
    .QN(_00033_)
  );
  DFF_X1 \mem_reg_wdata[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00273_),
    .Q(mem_reg_wdata[0]),
    .QN(_15319_)
  );
  DFF_X1 \mem_reg_wdata[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00283_),
    .Q(mem_reg_wdata[10]),
    .QN(_15309_)
  );
  DFF_X1 \mem_reg_wdata[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00284_),
    .Q(mem_reg_wdata[11]),
    .QN(_15308_)
  );
  DFF_X1 \mem_reg_wdata[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00285_),
    .Q(mem_reg_wdata[12]),
    .QN(_15307_)
  );
  DFF_X1 \mem_reg_wdata[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00286_),
    .Q(mem_reg_wdata[13]),
    .QN(_15306_)
  );
  DFF_X1 \mem_reg_wdata[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00287_),
    .Q(mem_reg_wdata[14]),
    .QN(_15305_)
  );
  DFF_X1 \mem_reg_wdata[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00288_),
    .Q(mem_reg_wdata[15]),
    .QN(_15304_)
  );
  DFF_X1 \mem_reg_wdata[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00289_),
    .Q(mem_reg_wdata[16]),
    .QN(_15303_)
  );
  DFF_X1 \mem_reg_wdata[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00290_),
    .Q(mem_reg_wdata[17]),
    .QN(_15302_)
  );
  DFF_X1 \mem_reg_wdata[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00291_),
    .Q(mem_reg_wdata[18]),
    .QN(_15301_)
  );
  DFF_X1 \mem_reg_wdata[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00292_),
    .Q(mem_reg_wdata[19]),
    .QN(_15300_)
  );
  DFF_X1 \mem_reg_wdata[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00274_),
    .Q(mem_reg_wdata[1]),
    .QN(_15318_)
  );
  DFF_X1 \mem_reg_wdata[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00293_),
    .Q(mem_reg_wdata[20]),
    .QN(_15299_)
  );
  DFF_X1 \mem_reg_wdata[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00294_),
    .Q(mem_reg_wdata[21]),
    .QN(_15298_)
  );
  DFF_X1 \mem_reg_wdata[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00295_),
    .Q(mem_reg_wdata[22]),
    .QN(_15297_)
  );
  DFF_X1 \mem_reg_wdata[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00296_),
    .Q(mem_reg_wdata[23]),
    .QN(_15296_)
  );
  DFF_X1 \mem_reg_wdata[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00297_),
    .Q(mem_reg_wdata[24]),
    .QN(_15295_)
  );
  DFF_X1 \mem_reg_wdata[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00298_),
    .Q(mem_reg_wdata[25]),
    .QN(_15294_)
  );
  DFF_X1 \mem_reg_wdata[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00299_),
    .Q(mem_reg_wdata[26]),
    .QN(_15293_)
  );
  DFF_X1 \mem_reg_wdata[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00300_),
    .Q(mem_reg_wdata[27]),
    .QN(_15292_)
  );
  DFF_X1 \mem_reg_wdata[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00301_),
    .Q(mem_reg_wdata[28]),
    .QN(_15291_)
  );
  DFF_X1 \mem_reg_wdata[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00302_),
    .Q(mem_reg_wdata[29]),
    .QN(_15290_)
  );
  DFF_X1 \mem_reg_wdata[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00275_),
    .Q(mem_reg_wdata[2]),
    .QN(_15317_)
  );
  DFF_X1 \mem_reg_wdata[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00303_),
    .Q(mem_reg_wdata[30]),
    .QN(_15289_)
  );
  DFF_X1 \mem_reg_wdata[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00304_),
    .Q(mem_reg_wdata[31]),
    .QN(_15288_)
  );
  DFF_X1 \mem_reg_wdata[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00276_),
    .Q(mem_reg_wdata[3]),
    .QN(_15316_)
  );
  DFF_X1 \mem_reg_wdata[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00277_),
    .Q(mem_reg_wdata[4]),
    .QN(_15315_)
  );
  DFF_X1 \mem_reg_wdata[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00278_),
    .Q(mem_reg_wdata[5]),
    .QN(_15314_)
  );
  DFF_X1 \mem_reg_wdata[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00279_),
    .Q(mem_reg_wdata[6]),
    .QN(_15313_)
  );
  DFF_X1 \mem_reg_wdata[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00280_),
    .Q(mem_reg_wdata[7]),
    .QN(_15312_)
  );
  DFF_X1 \mem_reg_wdata[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00281_),
    .Q(mem_reg_wdata[8]),
    .QN(_15311_)
  );
  DFF_X1 \mem_reg_wdata[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00282_),
    .Q(mem_reg_wdata[9]),
    .QN(_15310_)
  );
  DFF_X1 \mem_reg_xcpt$_DFF_P_  (
    .CK(clock),
    .D(_00007_),
    .Q(mem_reg_xcpt),
    .QN(_take_pc_mem_T)
  );
  DFF_X1 \mem_reg_xcpt_interrupt$_DFF_P_  (
    .CK(clock),
    .D(_00008_),
    .Q(mem_reg_xcpt_interrupt),
    .QN(_15180_)
  );
  DFF_X1 \rf[0][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00751_),
    .Q(\rf[0] [0]),
    .QN(_14863_)
  );
  DFF_X1 \rf[0][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00761_),
    .Q(\rf[0] [10]),
    .QN(_14853_)
  );
  DFF_X1 \rf[0][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00762_),
    .Q(\rf[0] [11]),
    .QN(_14852_)
  );
  DFF_X1 \rf[0][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00763_),
    .Q(\rf[0] [12]),
    .QN(_14851_)
  );
  DFF_X1 \rf[0][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00764_),
    .Q(\rf[0] [13]),
    .QN(_14850_)
  );
  DFF_X1 \rf[0][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00765_),
    .Q(\rf[0] [14]),
    .QN(_14849_)
  );
  DFF_X1 \rf[0][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00766_),
    .Q(\rf[0] [15]),
    .QN(_14848_)
  );
  DFF_X1 \rf[0][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00767_),
    .Q(\rf[0] [16]),
    .QN(_14847_)
  );
  DFF_X1 \rf[0][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00768_),
    .Q(\rf[0] [17]),
    .QN(_14846_)
  );
  DFF_X1 \rf[0][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00769_),
    .Q(\rf[0] [18]),
    .QN(_14845_)
  );
  DFF_X1 \rf[0][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00770_),
    .Q(\rf[0] [19]),
    .QN(_14844_)
  );
  DFF_X1 \rf[0][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00752_),
    .Q(\rf[0] [1]),
    .QN(_14862_)
  );
  DFF_X1 \rf[0][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00771_),
    .Q(\rf[0] [20]),
    .QN(_14843_)
  );
  DFF_X1 \rf[0][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00772_),
    .Q(\rf[0] [21]),
    .QN(_14842_)
  );
  DFF_X1 \rf[0][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00773_),
    .Q(\rf[0] [22]),
    .QN(_14841_)
  );
  DFF_X1 \rf[0][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00774_),
    .Q(\rf[0] [23]),
    .QN(_14840_)
  );
  DFF_X1 \rf[0][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00775_),
    .Q(\rf[0] [24]),
    .QN(_14839_)
  );
  DFF_X1 \rf[0][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00776_),
    .Q(\rf[0] [25]),
    .QN(_14838_)
  );
  DFF_X1 \rf[0][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00777_),
    .Q(\rf[0] [26]),
    .QN(_14837_)
  );
  DFF_X1 \rf[0][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00778_),
    .Q(\rf[0] [27]),
    .QN(_14836_)
  );
  DFF_X1 \rf[0][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00779_),
    .Q(\rf[0] [28]),
    .QN(_14835_)
  );
  DFF_X1 \rf[0][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00780_),
    .Q(\rf[0] [29]),
    .QN(_14834_)
  );
  DFF_X1 \rf[0][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00753_),
    .Q(\rf[0] [2]),
    .QN(_14861_)
  );
  DFF_X1 \rf[0][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00781_),
    .Q(\rf[0] [30]),
    .QN(_14833_)
  );
  DFF_X1 \rf[0][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00625_),
    .Q(\rf[0] [31]),
    .QN(_14988_)
  );
  DFF_X1 \rf[0][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00754_),
    .Q(\rf[0] [3]),
    .QN(_14860_)
  );
  DFF_X1 \rf[0][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00755_),
    .Q(\rf[0] [4]),
    .QN(_14859_)
  );
  DFF_X1 \rf[0][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00756_),
    .Q(\rf[0] [5]),
    .QN(_14858_)
  );
  DFF_X1 \rf[0][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00757_),
    .Q(\rf[0] [6]),
    .QN(_14857_)
  );
  DFF_X1 \rf[0][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00758_),
    .Q(\rf[0] [7]),
    .QN(_14856_)
  );
  DFF_X1 \rf[0][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00759_),
    .Q(\rf[0] [8]),
    .QN(_14855_)
  );
  DFF_X1 \rf[0][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00760_),
    .Q(\rf[0] [9]),
    .QN(_14854_)
  );
  DFF_X1 \rf[10][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00906_),
    .Q(\rf[10] [0]),
    .QN(_14708_)
  );
  DFF_X1 \rf[10][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00916_),
    .Q(\rf[10] [10]),
    .QN(_14698_)
  );
  DFF_X1 \rf[10][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00917_),
    .Q(\rf[10] [11]),
    .QN(_14697_)
  );
  DFF_X1 \rf[10][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00918_),
    .Q(\rf[10] [12]),
    .QN(_14696_)
  );
  DFF_X1 \rf[10][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00919_),
    .Q(\rf[10] [13]),
    .QN(_14695_)
  );
  DFF_X1 \rf[10][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00920_),
    .Q(\rf[10] [14]),
    .QN(_14694_)
  );
  DFF_X1 \rf[10][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00921_),
    .Q(\rf[10] [15]),
    .QN(_14693_)
  );
  DFF_X1 \rf[10][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00922_),
    .Q(\rf[10] [16]),
    .QN(_14692_)
  );
  DFF_X1 \rf[10][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00923_),
    .Q(\rf[10] [17]),
    .QN(_14691_)
  );
  DFF_X1 \rf[10][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00924_),
    .Q(\rf[10] [18]),
    .QN(_14690_)
  );
  DFF_X1 \rf[10][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00925_),
    .Q(\rf[10] [19]),
    .QN(_14689_)
  );
  DFF_X1 \rf[10][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00907_),
    .Q(\rf[10] [1]),
    .QN(_14707_)
  );
  DFF_X1 \rf[10][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00926_),
    .Q(\rf[10] [20]),
    .QN(_14688_)
  );
  DFF_X1 \rf[10][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00927_),
    .Q(\rf[10] [21]),
    .QN(_14687_)
  );
  DFF_X1 \rf[10][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00928_),
    .Q(\rf[10] [22]),
    .QN(_14686_)
  );
  DFF_X1 \rf[10][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00929_),
    .Q(\rf[10] [23]),
    .QN(_14685_)
  );
  DFF_X1 \rf[10][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00930_),
    .Q(\rf[10] [24]),
    .QN(_14684_)
  );
  DFF_X1 \rf[10][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00931_),
    .Q(\rf[10] [25]),
    .QN(_14683_)
  );
  DFF_X1 \rf[10][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00932_),
    .Q(\rf[10] [26]),
    .QN(_14682_)
  );
  DFF_X1 \rf[10][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00933_),
    .Q(\rf[10] [27]),
    .QN(_14681_)
  );
  DFF_X1 \rf[10][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00934_),
    .Q(\rf[10] [28]),
    .QN(_14680_)
  );
  DFF_X1 \rf[10][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00935_),
    .Q(\rf[10] [29]),
    .QN(_14679_)
  );
  DFF_X1 \rf[10][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00908_),
    .Q(\rf[10] [2]),
    .QN(_14706_)
  );
  DFF_X1 \rf[10][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00936_),
    .Q(\rf[10] [30]),
    .QN(_14678_)
  );
  DFF_X1 \rf[10][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00624_),
    .Q(\rf[10] [31]),
    .QN(_14989_)
  );
  DFF_X1 \rf[10][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00909_),
    .Q(\rf[10] [3]),
    .QN(_14705_)
  );
  DFF_X1 \rf[10][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00910_),
    .Q(\rf[10] [4]),
    .QN(_14704_)
  );
  DFF_X1 \rf[10][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00911_),
    .Q(\rf[10] [5]),
    .QN(_14703_)
  );
  DFF_X1 \rf[10][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00912_),
    .Q(\rf[10] [6]),
    .QN(_14702_)
  );
  DFF_X1 \rf[10][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00913_),
    .Q(\rf[10] [7]),
    .QN(_14701_)
  );
  DFF_X1 \rf[10][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00914_),
    .Q(\rf[10] [8]),
    .QN(_14700_)
  );
  DFF_X1 \rf[10][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00915_),
    .Q(\rf[10] [9]),
    .QN(_14699_)
  );
  DFF_X1 \rf[11][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00968_),
    .Q(\rf[11] [0]),
    .QN(_14646_)
  );
  DFF_X1 \rf[11][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00978_),
    .Q(\rf[11] [10]),
    .QN(_14636_)
  );
  DFF_X1 \rf[11][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00979_),
    .Q(\rf[11] [11]),
    .QN(_14635_)
  );
  DFF_X1 \rf[11][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00980_),
    .Q(\rf[11] [12]),
    .QN(_14634_)
  );
  DFF_X1 \rf[11][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00981_),
    .Q(\rf[11] [13]),
    .QN(_14633_)
  );
  DFF_X1 \rf[11][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00982_),
    .Q(\rf[11] [14]),
    .QN(_14632_)
  );
  DFF_X1 \rf[11][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00983_),
    .Q(\rf[11] [15]),
    .QN(_14631_)
  );
  DFF_X1 \rf[11][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00984_),
    .Q(\rf[11] [16]),
    .QN(_14630_)
  );
  DFF_X1 \rf[11][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00985_),
    .Q(\rf[11] [17]),
    .QN(_14629_)
  );
  DFF_X1 \rf[11][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00986_),
    .Q(\rf[11] [18]),
    .QN(_14628_)
  );
  DFF_X1 \rf[11][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00987_),
    .Q(\rf[11] [19]),
    .QN(_14627_)
  );
  DFF_X1 \rf[11][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00969_),
    .Q(\rf[11] [1]),
    .QN(_14645_)
  );
  DFF_X1 \rf[11][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00988_),
    .Q(\rf[11] [20]),
    .QN(_14626_)
  );
  DFF_X1 \rf[11][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00989_),
    .Q(\rf[11] [21]),
    .QN(_14625_)
  );
  DFF_X1 \rf[11][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00990_),
    .Q(\rf[11] [22]),
    .QN(_14624_)
  );
  DFF_X1 \rf[11][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00991_),
    .Q(\rf[11] [23]),
    .QN(_14623_)
  );
  DFF_X1 \rf[11][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00992_),
    .Q(\rf[11] [24]),
    .QN(_14622_)
  );
  DFF_X1 \rf[11][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00993_),
    .Q(\rf[11] [25]),
    .QN(_14621_)
  );
  DFF_X1 \rf[11][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00994_),
    .Q(\rf[11] [26]),
    .QN(_14620_)
  );
  DFF_X1 \rf[11][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00995_),
    .Q(\rf[11] [27]),
    .QN(_14619_)
  );
  DFF_X1 \rf[11][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00996_),
    .Q(\rf[11] [28]),
    .QN(_14618_)
  );
  DFF_X1 \rf[11][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00997_),
    .Q(\rf[11] [29]),
    .QN(_14617_)
  );
  DFF_X1 \rf[11][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00970_),
    .Q(\rf[11] [2]),
    .QN(_14644_)
  );
  DFF_X1 \rf[11][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00998_),
    .Q(\rf[11] [30]),
    .QN(_14616_)
  );
  DFF_X1 \rf[11][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00623_),
    .Q(\rf[11] [31]),
    .QN(_14990_)
  );
  DFF_X1 \rf[11][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00971_),
    .Q(\rf[11] [3]),
    .QN(_14643_)
  );
  DFF_X1 \rf[11][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00972_),
    .Q(\rf[11] [4]),
    .QN(_14642_)
  );
  DFF_X1 \rf[11][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00973_),
    .Q(\rf[11] [5]),
    .QN(_14641_)
  );
  DFF_X1 \rf[11][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00974_),
    .Q(\rf[11] [6]),
    .QN(_14640_)
  );
  DFF_X1 \rf[11][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00975_),
    .Q(\rf[11] [7]),
    .QN(_14639_)
  );
  DFF_X1 \rf[11][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00976_),
    .Q(\rf[11] [8]),
    .QN(_14638_)
  );
  DFF_X1 \rf[11][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00977_),
    .Q(\rf[11] [9]),
    .QN(_14637_)
  );
  DFF_X1 \rf[12][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01030_),
    .Q(\rf[12] [0]),
    .QN(_14584_)
  );
  DFF_X1 \rf[12][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01040_),
    .Q(\rf[12] [10]),
    .QN(_14574_)
  );
  DFF_X1 \rf[12][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01041_),
    .Q(\rf[12] [11]),
    .QN(_14573_)
  );
  DFF_X1 \rf[12][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01042_),
    .Q(\rf[12] [12]),
    .QN(_14572_)
  );
  DFF_X1 \rf[12][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01043_),
    .Q(\rf[12] [13]),
    .QN(_14571_)
  );
  DFF_X1 \rf[12][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01044_),
    .Q(\rf[12] [14]),
    .QN(_14570_)
  );
  DFF_X1 \rf[12][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01045_),
    .Q(\rf[12] [15]),
    .QN(_14569_)
  );
  DFF_X1 \rf[12][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01046_),
    .Q(\rf[12] [16]),
    .QN(_14568_)
  );
  DFF_X1 \rf[12][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01047_),
    .Q(\rf[12] [17]),
    .QN(_14567_)
  );
  DFF_X1 \rf[12][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01048_),
    .Q(\rf[12] [18]),
    .QN(_14566_)
  );
  DFF_X1 \rf[12][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01049_),
    .Q(\rf[12] [19]),
    .QN(_14565_)
  );
  DFF_X1 \rf[12][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01031_),
    .Q(\rf[12] [1]),
    .QN(_14583_)
  );
  DFF_X1 \rf[12][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01050_),
    .Q(\rf[12] [20]),
    .QN(_14564_)
  );
  DFF_X1 \rf[12][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01051_),
    .Q(\rf[12] [21]),
    .QN(_14563_)
  );
  DFF_X1 \rf[12][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01052_),
    .Q(\rf[12] [22]),
    .QN(_14562_)
  );
  DFF_X1 \rf[12][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01053_),
    .Q(\rf[12] [23]),
    .QN(_14561_)
  );
  DFF_X1 \rf[12][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01054_),
    .Q(\rf[12] [24]),
    .QN(_14560_)
  );
  DFF_X1 \rf[12][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01055_),
    .Q(\rf[12] [25]),
    .QN(_14559_)
  );
  DFF_X1 \rf[12][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01056_),
    .Q(\rf[12] [26]),
    .QN(_14558_)
  );
  DFF_X1 \rf[12][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01057_),
    .Q(\rf[12] [27]),
    .QN(_14557_)
  );
  DFF_X1 \rf[12][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01058_),
    .Q(\rf[12] [28]),
    .QN(_14556_)
  );
  DFF_X1 \rf[12][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01059_),
    .Q(\rf[12] [29]),
    .QN(_14555_)
  );
  DFF_X1 \rf[12][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01032_),
    .Q(\rf[12] [2]),
    .QN(_14582_)
  );
  DFF_X1 \rf[12][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01060_),
    .Q(\rf[12] [30]),
    .QN(_14554_)
  );
  DFF_X1 \rf[12][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00622_),
    .Q(\rf[12] [31]),
    .QN(_14991_)
  );
  DFF_X1 \rf[12][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01033_),
    .Q(\rf[12] [3]),
    .QN(_14581_)
  );
  DFF_X1 \rf[12][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01034_),
    .Q(\rf[12] [4]),
    .QN(_14580_)
  );
  DFF_X1 \rf[12][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01035_),
    .Q(\rf[12] [5]),
    .QN(_14579_)
  );
  DFF_X1 \rf[12][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01036_),
    .Q(\rf[12] [6]),
    .QN(_14578_)
  );
  DFF_X1 \rf[12][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01037_),
    .Q(\rf[12] [7]),
    .QN(_14577_)
  );
  DFF_X1 \rf[12][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01038_),
    .Q(\rf[12] [8]),
    .QN(_14576_)
  );
  DFF_X1 \rf[12][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01039_),
    .Q(\rf[12] [9]),
    .QN(_14575_)
  );
  DFF_X1 \rf[13][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01154_),
    .Q(\rf[13] [0]),
    .QN(_14460_)
  );
  DFF_X1 \rf[13][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01164_),
    .Q(\rf[13] [10]),
    .QN(_14450_)
  );
  DFF_X1 \rf[13][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01165_),
    .Q(\rf[13] [11]),
    .QN(_14449_)
  );
  DFF_X1 \rf[13][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01166_),
    .Q(\rf[13] [12]),
    .QN(_14448_)
  );
  DFF_X1 \rf[13][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01167_),
    .Q(\rf[13] [13]),
    .QN(_14447_)
  );
  DFF_X1 \rf[13][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01168_),
    .Q(\rf[13] [14]),
    .QN(_14446_)
  );
  DFF_X1 \rf[13][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01169_),
    .Q(\rf[13] [15]),
    .QN(_14445_)
  );
  DFF_X1 \rf[13][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01170_),
    .Q(\rf[13] [16]),
    .QN(_14444_)
  );
  DFF_X1 \rf[13][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01171_),
    .Q(\rf[13] [17]),
    .QN(_14443_)
  );
  DFF_X1 \rf[13][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01172_),
    .Q(\rf[13] [18]),
    .QN(_14442_)
  );
  DFF_X1 \rf[13][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01173_),
    .Q(\rf[13] [19]),
    .QN(_14441_)
  );
  DFF_X1 \rf[13][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01155_),
    .Q(\rf[13] [1]),
    .QN(_14459_)
  );
  DFF_X1 \rf[13][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01174_),
    .Q(\rf[13] [20]),
    .QN(_14440_)
  );
  DFF_X1 \rf[13][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01175_),
    .Q(\rf[13] [21]),
    .QN(_14439_)
  );
  DFF_X1 \rf[13][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01176_),
    .Q(\rf[13] [22]),
    .QN(_14438_)
  );
  DFF_X1 \rf[13][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01177_),
    .Q(\rf[13] [23]),
    .QN(_14437_)
  );
  DFF_X1 \rf[13][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01178_),
    .Q(\rf[13] [24]),
    .QN(_14436_)
  );
  DFF_X1 \rf[13][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01179_),
    .Q(\rf[13] [25]),
    .QN(_14435_)
  );
  DFF_X1 \rf[13][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01180_),
    .Q(\rf[13] [26]),
    .QN(_14434_)
  );
  DFF_X1 \rf[13][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01181_),
    .Q(\rf[13] [27]),
    .QN(_14433_)
  );
  DFF_X1 \rf[13][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01182_),
    .Q(\rf[13] [28]),
    .QN(_14432_)
  );
  DFF_X1 \rf[13][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01183_),
    .Q(\rf[13] [29]),
    .QN(_14431_)
  );
  DFF_X1 \rf[13][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01156_),
    .Q(\rf[13] [2]),
    .QN(_14458_)
  );
  DFF_X1 \rf[13][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01184_),
    .Q(\rf[13] [30]),
    .QN(_14430_)
  );
  DFF_X1 \rf[13][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00621_),
    .Q(\rf[13] [31]),
    .QN(_14992_)
  );
  DFF_X1 \rf[13][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01157_),
    .Q(\rf[13] [3]),
    .QN(_14457_)
  );
  DFF_X1 \rf[13][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01158_),
    .Q(\rf[13] [4]),
    .QN(_14456_)
  );
  DFF_X1 \rf[13][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01159_),
    .Q(\rf[13] [5]),
    .QN(_14455_)
  );
  DFF_X1 \rf[13][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01160_),
    .Q(\rf[13] [6]),
    .QN(_14454_)
  );
  DFF_X1 \rf[13][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01161_),
    .Q(\rf[13] [7]),
    .QN(_14453_)
  );
  DFF_X1 \rf[13][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01162_),
    .Q(\rf[13] [8]),
    .QN(_14452_)
  );
  DFF_X1 \rf[13][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01163_),
    .Q(\rf[13] [9]),
    .QN(_14451_)
  );
  DFF_X1 \rf[14][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01278_),
    .Q(\rf[14] [0]),
    .QN(_14336_)
  );
  DFF_X1 \rf[14][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01288_),
    .Q(\rf[14] [10]),
    .QN(_14326_)
  );
  DFF_X1 \rf[14][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01289_),
    .Q(\rf[14] [11]),
    .QN(_14325_)
  );
  DFF_X1 \rf[14][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01290_),
    .Q(\rf[14] [12]),
    .QN(_14324_)
  );
  DFF_X1 \rf[14][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01291_),
    .Q(\rf[14] [13]),
    .QN(_14323_)
  );
  DFF_X1 \rf[14][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01292_),
    .Q(\rf[14] [14]),
    .QN(_14322_)
  );
  DFF_X1 \rf[14][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01293_),
    .Q(\rf[14] [15]),
    .QN(_14321_)
  );
  DFF_X1 \rf[14][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01294_),
    .Q(\rf[14] [16]),
    .QN(_14320_)
  );
  DFF_X1 \rf[14][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01295_),
    .Q(\rf[14] [17]),
    .QN(_14319_)
  );
  DFF_X1 \rf[14][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01296_),
    .Q(\rf[14] [18]),
    .QN(_14318_)
  );
  DFF_X1 \rf[14][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01297_),
    .Q(\rf[14] [19]),
    .QN(_14317_)
  );
  DFF_X1 \rf[14][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01279_),
    .Q(\rf[14] [1]),
    .QN(_14335_)
  );
  DFF_X1 \rf[14][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01298_),
    .Q(\rf[14] [20]),
    .QN(_14316_)
  );
  DFF_X1 \rf[14][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01299_),
    .Q(\rf[14] [21]),
    .QN(_14315_)
  );
  DFF_X1 \rf[14][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01300_),
    .Q(\rf[14] [22]),
    .QN(_14314_)
  );
  DFF_X1 \rf[14][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01301_),
    .Q(\rf[14] [23]),
    .QN(_14313_)
  );
  DFF_X1 \rf[14][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01302_),
    .Q(\rf[14] [24]),
    .QN(_14312_)
  );
  DFF_X1 \rf[14][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01303_),
    .Q(\rf[14] [25]),
    .QN(_14311_)
  );
  DFF_X1 \rf[14][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01304_),
    .Q(\rf[14] [26]),
    .QN(_14310_)
  );
  DFF_X1 \rf[14][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01305_),
    .Q(\rf[14] [27]),
    .QN(_14309_)
  );
  DFF_X1 \rf[14][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01306_),
    .Q(\rf[14] [28]),
    .QN(_14308_)
  );
  DFF_X1 \rf[14][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01307_),
    .Q(\rf[14] [29]),
    .QN(_14307_)
  );
  DFF_X1 \rf[14][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01280_),
    .Q(\rf[14] [2]),
    .QN(_14334_)
  );
  DFF_X1 \rf[14][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01308_),
    .Q(\rf[14] [30]),
    .QN(_14306_)
  );
  DFF_X1 \rf[14][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00620_),
    .Q(\rf[14] [31]),
    .QN(_14993_)
  );
  DFF_X1 \rf[14][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01281_),
    .Q(\rf[14] [3]),
    .QN(_14333_)
  );
  DFF_X1 \rf[14][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01282_),
    .Q(\rf[14] [4]),
    .QN(_14332_)
  );
  DFF_X1 \rf[14][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01283_),
    .Q(\rf[14] [5]),
    .QN(_14331_)
  );
  DFF_X1 \rf[14][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01284_),
    .Q(\rf[14] [6]),
    .QN(_14330_)
  );
  DFF_X1 \rf[14][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01285_),
    .Q(\rf[14] [7]),
    .QN(_14329_)
  );
  DFF_X1 \rf[14][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01286_),
    .Q(\rf[14] [8]),
    .QN(_14328_)
  );
  DFF_X1 \rf[14][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01287_),
    .Q(\rf[14] [9]),
    .QN(_14327_)
  );
  DFF_X1 \rf[15][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00782_),
    .Q(\rf[15] [0]),
    .QN(_14832_)
  );
  DFF_X1 \rf[15][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00792_),
    .Q(\rf[15] [10]),
    .QN(_14822_)
  );
  DFF_X1 \rf[15][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00793_),
    .Q(\rf[15] [11]),
    .QN(_14821_)
  );
  DFF_X1 \rf[15][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00794_),
    .Q(\rf[15] [12]),
    .QN(_14820_)
  );
  DFF_X1 \rf[15][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00795_),
    .Q(\rf[15] [13]),
    .QN(_14819_)
  );
  DFF_X1 \rf[15][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00796_),
    .Q(\rf[15] [14]),
    .QN(_14818_)
  );
  DFF_X1 \rf[15][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00797_),
    .Q(\rf[15] [15]),
    .QN(_14817_)
  );
  DFF_X1 \rf[15][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00798_),
    .Q(\rf[15] [16]),
    .QN(_14816_)
  );
  DFF_X1 \rf[15][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00799_),
    .Q(\rf[15] [17]),
    .QN(_14815_)
  );
  DFF_X1 \rf[15][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00800_),
    .Q(\rf[15] [18]),
    .QN(_14814_)
  );
  DFF_X1 \rf[15][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00801_),
    .Q(\rf[15] [19]),
    .QN(_14813_)
  );
  DFF_X1 \rf[15][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00783_),
    .Q(\rf[15] [1]),
    .QN(_14831_)
  );
  DFF_X1 \rf[15][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00802_),
    .Q(\rf[15] [20]),
    .QN(_14812_)
  );
  DFF_X1 \rf[15][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00803_),
    .Q(\rf[15] [21]),
    .QN(_14811_)
  );
  DFF_X1 \rf[15][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00804_),
    .Q(\rf[15] [22]),
    .QN(_14810_)
  );
  DFF_X1 \rf[15][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00805_),
    .Q(\rf[15] [23]),
    .QN(_14809_)
  );
  DFF_X1 \rf[15][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00806_),
    .Q(\rf[15] [24]),
    .QN(_14808_)
  );
  DFF_X1 \rf[15][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00807_),
    .Q(\rf[15] [25]),
    .QN(_14807_)
  );
  DFF_X1 \rf[15][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00808_),
    .Q(\rf[15] [26]),
    .QN(_14806_)
  );
  DFF_X1 \rf[15][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00809_),
    .Q(\rf[15] [27]),
    .QN(_14805_)
  );
  DFF_X1 \rf[15][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00810_),
    .Q(\rf[15] [28]),
    .QN(_14804_)
  );
  DFF_X1 \rf[15][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00811_),
    .Q(\rf[15] [29]),
    .QN(_14803_)
  );
  DFF_X1 \rf[15][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00784_),
    .Q(\rf[15] [2]),
    .QN(_14830_)
  );
  DFF_X1 \rf[15][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00812_),
    .Q(\rf[15] [30]),
    .QN(_14802_)
  );
  DFF_X1 \rf[15][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00619_),
    .Q(\rf[15] [31]),
    .QN(_14994_)
  );
  DFF_X1 \rf[15][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00785_),
    .Q(\rf[15] [3]),
    .QN(_14829_)
  );
  DFF_X1 \rf[15][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00786_),
    .Q(\rf[15] [4]),
    .QN(_14828_)
  );
  DFF_X1 \rf[15][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00787_),
    .Q(\rf[15] [5]),
    .QN(_14827_)
  );
  DFF_X1 \rf[15][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00788_),
    .Q(\rf[15] [6]),
    .QN(_14826_)
  );
  DFF_X1 \rf[15][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00789_),
    .Q(\rf[15] [7]),
    .QN(_14825_)
  );
  DFF_X1 \rf[15][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00790_),
    .Q(\rf[15] [8]),
    .QN(_14824_)
  );
  DFF_X1 \rf[15][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00791_),
    .Q(\rf[15] [9]),
    .QN(_14823_)
  );
  DFF_X1 \rf[16][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00844_),
    .Q(\rf[16] [0]),
    .QN(_14770_)
  );
  DFF_X1 \rf[16][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00854_),
    .Q(\rf[16] [10]),
    .QN(_14760_)
  );
  DFF_X1 \rf[16][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00855_),
    .Q(\rf[16] [11]),
    .QN(_14759_)
  );
  DFF_X1 \rf[16][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00856_),
    .Q(\rf[16] [12]),
    .QN(_14758_)
  );
  DFF_X1 \rf[16][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00857_),
    .Q(\rf[16] [13]),
    .QN(_14757_)
  );
  DFF_X1 \rf[16][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00858_),
    .Q(\rf[16] [14]),
    .QN(_14756_)
  );
  DFF_X1 \rf[16][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00859_),
    .Q(\rf[16] [15]),
    .QN(_14755_)
  );
  DFF_X1 \rf[16][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00860_),
    .Q(\rf[16] [16]),
    .QN(_14754_)
  );
  DFF_X1 \rf[16][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00861_),
    .Q(\rf[16] [17]),
    .QN(_14753_)
  );
  DFF_X1 \rf[16][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00862_),
    .Q(\rf[16] [18]),
    .QN(_14752_)
  );
  DFF_X1 \rf[16][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00863_),
    .Q(\rf[16] [19]),
    .QN(_14751_)
  );
  DFF_X1 \rf[16][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00845_),
    .Q(\rf[16] [1]),
    .QN(_14769_)
  );
  DFF_X1 \rf[16][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00864_),
    .Q(\rf[16] [20]),
    .QN(_14750_)
  );
  DFF_X1 \rf[16][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00865_),
    .Q(\rf[16] [21]),
    .QN(_14749_)
  );
  DFF_X1 \rf[16][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00866_),
    .Q(\rf[16] [22]),
    .QN(_14748_)
  );
  DFF_X1 \rf[16][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00867_),
    .Q(\rf[16] [23]),
    .QN(_14747_)
  );
  DFF_X1 \rf[16][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00868_),
    .Q(\rf[16] [24]),
    .QN(_14746_)
  );
  DFF_X1 \rf[16][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00869_),
    .Q(\rf[16] [25]),
    .QN(_14745_)
  );
  DFF_X1 \rf[16][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00870_),
    .Q(\rf[16] [26]),
    .QN(_14744_)
  );
  DFF_X1 \rf[16][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00871_),
    .Q(\rf[16] [27]),
    .QN(_14743_)
  );
  DFF_X1 \rf[16][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00872_),
    .Q(\rf[16] [28]),
    .QN(_14742_)
  );
  DFF_X1 \rf[16][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00873_),
    .Q(\rf[16] [29]),
    .QN(_14741_)
  );
  DFF_X1 \rf[16][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00846_),
    .Q(\rf[16] [2]),
    .QN(_14768_)
  );
  DFF_X1 \rf[16][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00874_),
    .Q(\rf[16] [30]),
    .QN(_14740_)
  );
  DFF_X1 \rf[16][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00618_),
    .Q(\rf[16] [31]),
    .QN(_14995_)
  );
  DFF_X1 \rf[16][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00847_),
    .Q(\rf[16] [3]),
    .QN(_14767_)
  );
  DFF_X1 \rf[16][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00848_),
    .Q(\rf[16] [4]),
    .QN(_14766_)
  );
  DFF_X1 \rf[16][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00849_),
    .Q(\rf[16] [5]),
    .QN(_14765_)
  );
  DFF_X1 \rf[16][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00850_),
    .Q(\rf[16] [6]),
    .QN(_14764_)
  );
  DFF_X1 \rf[16][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00851_),
    .Q(\rf[16] [7]),
    .QN(_14763_)
  );
  DFF_X1 \rf[16][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00852_),
    .Q(\rf[16] [8]),
    .QN(_14762_)
  );
  DFF_X1 \rf[16][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00853_),
    .Q(\rf[16] [9]),
    .QN(_14761_)
  );
  DFF_X1 \rf[17][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00875_),
    .Q(\rf[17] [0]),
    .QN(_14739_)
  );
  DFF_X1 \rf[17][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00885_),
    .Q(\rf[17] [10]),
    .QN(_14729_)
  );
  DFF_X1 \rf[17][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00886_),
    .Q(\rf[17] [11]),
    .QN(_14728_)
  );
  DFF_X1 \rf[17][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00887_),
    .Q(\rf[17] [12]),
    .QN(_14727_)
  );
  DFF_X1 \rf[17][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00888_),
    .Q(\rf[17] [13]),
    .QN(_14726_)
  );
  DFF_X1 \rf[17][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00889_),
    .Q(\rf[17] [14]),
    .QN(_14725_)
  );
  DFF_X1 \rf[17][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00890_),
    .Q(\rf[17] [15]),
    .QN(_14724_)
  );
  DFF_X1 \rf[17][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00891_),
    .Q(\rf[17] [16]),
    .QN(_14723_)
  );
  DFF_X1 \rf[17][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00892_),
    .Q(\rf[17] [17]),
    .QN(_14722_)
  );
  DFF_X1 \rf[17][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00893_),
    .Q(\rf[17] [18]),
    .QN(_14721_)
  );
  DFF_X1 \rf[17][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00894_),
    .Q(\rf[17] [19]),
    .QN(_14720_)
  );
  DFF_X1 \rf[17][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00876_),
    .Q(\rf[17] [1]),
    .QN(_14738_)
  );
  DFF_X1 \rf[17][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00895_),
    .Q(\rf[17] [20]),
    .QN(_14719_)
  );
  DFF_X1 \rf[17][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00896_),
    .Q(\rf[17] [21]),
    .QN(_14718_)
  );
  DFF_X1 \rf[17][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00897_),
    .Q(\rf[17] [22]),
    .QN(_14717_)
  );
  DFF_X1 \rf[17][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00898_),
    .Q(\rf[17] [23]),
    .QN(_14716_)
  );
  DFF_X1 \rf[17][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00899_),
    .Q(\rf[17] [24]),
    .QN(_14715_)
  );
  DFF_X1 \rf[17][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00900_),
    .Q(\rf[17] [25]),
    .QN(_14714_)
  );
  DFF_X1 \rf[17][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00901_),
    .Q(\rf[17] [26]),
    .QN(_14713_)
  );
  DFF_X1 \rf[17][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00902_),
    .Q(\rf[17] [27]),
    .QN(_14712_)
  );
  DFF_X1 \rf[17][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00903_),
    .Q(\rf[17] [28]),
    .QN(_14711_)
  );
  DFF_X1 \rf[17][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00904_),
    .Q(\rf[17] [29]),
    .QN(_14710_)
  );
  DFF_X1 \rf[17][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00877_),
    .Q(\rf[17] [2]),
    .QN(_14737_)
  );
  DFF_X1 \rf[17][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00905_),
    .Q(\rf[17] [30]),
    .QN(_14709_)
  );
  DFF_X1 \rf[17][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00617_),
    .Q(\rf[17] [31]),
    .QN(_14996_)
  );
  DFF_X1 \rf[17][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00878_),
    .Q(\rf[17] [3]),
    .QN(_14736_)
  );
  DFF_X1 \rf[17][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00879_),
    .Q(\rf[17] [4]),
    .QN(_14735_)
  );
  DFF_X1 \rf[17][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00880_),
    .Q(\rf[17] [5]),
    .QN(_14734_)
  );
  DFF_X1 \rf[17][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00881_),
    .Q(\rf[17] [6]),
    .QN(_14733_)
  );
  DFF_X1 \rf[17][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00882_),
    .Q(\rf[17] [7]),
    .QN(_14732_)
  );
  DFF_X1 \rf[17][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00883_),
    .Q(\rf[17] [8]),
    .QN(_14731_)
  );
  DFF_X1 \rf[17][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00884_),
    .Q(\rf[17] [9]),
    .QN(_14730_)
  );
  DFF_X1 \rf[18][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00937_),
    .Q(\rf[18] [0]),
    .QN(_14677_)
  );
  DFF_X1 \rf[18][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00947_),
    .Q(\rf[18] [10]),
    .QN(_14667_)
  );
  DFF_X1 \rf[18][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00948_),
    .Q(\rf[18] [11]),
    .QN(_14666_)
  );
  DFF_X1 \rf[18][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00949_),
    .Q(\rf[18] [12]),
    .QN(_14665_)
  );
  DFF_X1 \rf[18][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00950_),
    .Q(\rf[18] [13]),
    .QN(_14664_)
  );
  DFF_X1 \rf[18][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00951_),
    .Q(\rf[18] [14]),
    .QN(_14663_)
  );
  DFF_X1 \rf[18][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00952_),
    .Q(\rf[18] [15]),
    .QN(_14662_)
  );
  DFF_X1 \rf[18][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00953_),
    .Q(\rf[18] [16]),
    .QN(_14661_)
  );
  DFF_X1 \rf[18][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00954_),
    .Q(\rf[18] [17]),
    .QN(_14660_)
  );
  DFF_X1 \rf[18][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00955_),
    .Q(\rf[18] [18]),
    .QN(_14659_)
  );
  DFF_X1 \rf[18][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00956_),
    .Q(\rf[18] [19]),
    .QN(_14658_)
  );
  DFF_X1 \rf[18][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00938_),
    .Q(\rf[18] [1]),
    .QN(_14676_)
  );
  DFF_X1 \rf[18][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00957_),
    .Q(\rf[18] [20]),
    .QN(_14657_)
  );
  DFF_X1 \rf[18][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00958_),
    .Q(\rf[18] [21]),
    .QN(_14656_)
  );
  DFF_X1 \rf[18][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00959_),
    .Q(\rf[18] [22]),
    .QN(_14655_)
  );
  DFF_X1 \rf[18][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00960_),
    .Q(\rf[18] [23]),
    .QN(_14654_)
  );
  DFF_X1 \rf[18][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00961_),
    .Q(\rf[18] [24]),
    .QN(_14653_)
  );
  DFF_X1 \rf[18][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00962_),
    .Q(\rf[18] [25]),
    .QN(_14652_)
  );
  DFF_X1 \rf[18][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00963_),
    .Q(\rf[18] [26]),
    .QN(_14651_)
  );
  DFF_X1 \rf[18][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00964_),
    .Q(\rf[18] [27]),
    .QN(_14650_)
  );
  DFF_X1 \rf[18][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00965_),
    .Q(\rf[18] [28]),
    .QN(_14649_)
  );
  DFF_X1 \rf[18][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00966_),
    .Q(\rf[18] [29]),
    .QN(_14648_)
  );
  DFF_X1 \rf[18][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00939_),
    .Q(\rf[18] [2]),
    .QN(_14675_)
  );
  DFF_X1 \rf[18][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00967_),
    .Q(\rf[18] [30]),
    .QN(_14647_)
  );
  DFF_X1 \rf[18][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00616_),
    .Q(\rf[18] [31]),
    .QN(_14997_)
  );
  DFF_X1 \rf[18][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00940_),
    .Q(\rf[18] [3]),
    .QN(_14674_)
  );
  DFF_X1 \rf[18][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00941_),
    .Q(\rf[18] [4]),
    .QN(_14673_)
  );
  DFF_X1 \rf[18][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00942_),
    .Q(\rf[18] [5]),
    .QN(_14672_)
  );
  DFF_X1 \rf[18][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00943_),
    .Q(\rf[18] [6]),
    .QN(_14671_)
  );
  DFF_X1 \rf[18][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00944_),
    .Q(\rf[18] [7]),
    .QN(_14670_)
  );
  DFF_X1 \rf[18][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00945_),
    .Q(\rf[18] [8]),
    .QN(_14669_)
  );
  DFF_X1 \rf[18][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00946_),
    .Q(\rf[18] [9]),
    .QN(_14668_)
  );
  DFF_X1 \rf[19][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00999_),
    .Q(\rf[19] [0]),
    .QN(_14615_)
  );
  DFF_X1 \rf[19][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01009_),
    .Q(\rf[19] [10]),
    .QN(_14605_)
  );
  DFF_X1 \rf[19][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01010_),
    .Q(\rf[19] [11]),
    .QN(_14604_)
  );
  DFF_X1 \rf[19][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01011_),
    .Q(\rf[19] [12]),
    .QN(_14603_)
  );
  DFF_X1 \rf[19][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01012_),
    .Q(\rf[19] [13]),
    .QN(_14602_)
  );
  DFF_X1 \rf[19][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01013_),
    .Q(\rf[19] [14]),
    .QN(_14601_)
  );
  DFF_X1 \rf[19][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01014_),
    .Q(\rf[19] [15]),
    .QN(_14600_)
  );
  DFF_X1 \rf[19][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01015_),
    .Q(\rf[19] [16]),
    .QN(_14599_)
  );
  DFF_X1 \rf[19][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01016_),
    .Q(\rf[19] [17]),
    .QN(_14598_)
  );
  DFF_X1 \rf[19][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01017_),
    .Q(\rf[19] [18]),
    .QN(_14597_)
  );
  DFF_X1 \rf[19][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01018_),
    .Q(\rf[19] [19]),
    .QN(_14596_)
  );
  DFF_X1 \rf[19][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01000_),
    .Q(\rf[19] [1]),
    .QN(_14614_)
  );
  DFF_X1 \rf[19][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01019_),
    .Q(\rf[19] [20]),
    .QN(_14595_)
  );
  DFF_X1 \rf[19][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01020_),
    .Q(\rf[19] [21]),
    .QN(_14594_)
  );
  DFF_X1 \rf[19][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01021_),
    .Q(\rf[19] [22]),
    .QN(_14593_)
  );
  DFF_X1 \rf[19][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01022_),
    .Q(\rf[19] [23]),
    .QN(_14592_)
  );
  DFF_X1 \rf[19][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01023_),
    .Q(\rf[19] [24]),
    .QN(_14591_)
  );
  DFF_X1 \rf[19][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01024_),
    .Q(\rf[19] [25]),
    .QN(_14590_)
  );
  DFF_X1 \rf[19][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01025_),
    .Q(\rf[19] [26]),
    .QN(_14589_)
  );
  DFF_X1 \rf[19][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01026_),
    .Q(\rf[19] [27]),
    .QN(_14588_)
  );
  DFF_X1 \rf[19][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01027_),
    .Q(\rf[19] [28]),
    .QN(_14587_)
  );
  DFF_X1 \rf[19][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01028_),
    .Q(\rf[19] [29]),
    .QN(_14586_)
  );
  DFF_X1 \rf[19][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01001_),
    .Q(\rf[19] [2]),
    .QN(_14613_)
  );
  DFF_X1 \rf[19][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01029_),
    .Q(\rf[19] [30]),
    .QN(_14585_)
  );
  DFF_X1 \rf[19][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00615_),
    .Q(\rf[19] [31]),
    .QN(_14998_)
  );
  DFF_X1 \rf[19][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01002_),
    .Q(\rf[19] [3]),
    .QN(_14612_)
  );
  DFF_X1 \rf[19][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01003_),
    .Q(\rf[19] [4]),
    .QN(_14611_)
  );
  DFF_X1 \rf[19][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01004_),
    .Q(\rf[19] [5]),
    .QN(_14610_)
  );
  DFF_X1 \rf[19][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01005_),
    .Q(\rf[19] [6]),
    .QN(_14609_)
  );
  DFF_X1 \rf[19][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01006_),
    .Q(\rf[19] [7]),
    .QN(_14608_)
  );
  DFF_X1 \rf[19][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01007_),
    .Q(\rf[19] [8]),
    .QN(_14607_)
  );
  DFF_X1 \rf[19][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01008_),
    .Q(\rf[19] [9]),
    .QN(_14606_)
  );
  DFF_X1 \rf[1][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01557_),
    .Q(\rf[1] [0]),
    .QN(_14057_)
  );
  DFF_X1 \rf[1][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01567_),
    .Q(\rf[1] [10]),
    .QN(_14047_)
  );
  DFF_X1 \rf[1][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01568_),
    .Q(\rf[1] [11]),
    .QN(_14046_)
  );
  DFF_X1 \rf[1][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01569_),
    .Q(\rf[1] [12]),
    .QN(_14045_)
  );
  DFF_X1 \rf[1][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01570_),
    .Q(\rf[1] [13]),
    .QN(_14044_)
  );
  DFF_X1 \rf[1][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01571_),
    .Q(\rf[1] [14]),
    .QN(_14043_)
  );
  DFF_X1 \rf[1][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01572_),
    .Q(\rf[1] [15]),
    .QN(_14042_)
  );
  DFF_X1 \rf[1][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01573_),
    .Q(\rf[1] [16]),
    .QN(_14041_)
  );
  DFF_X1 \rf[1][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01574_),
    .Q(\rf[1] [17]),
    .QN(_14040_)
  );
  DFF_X1 \rf[1][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01575_),
    .Q(\rf[1] [18]),
    .QN(_14039_)
  );
  DFF_X1 \rf[1][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01576_),
    .Q(\rf[1] [19]),
    .QN(_14038_)
  );
  DFF_X1 \rf[1][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01558_),
    .Q(\rf[1] [1]),
    .QN(_14056_)
  );
  DFF_X1 \rf[1][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01577_),
    .Q(\rf[1] [20]),
    .QN(_14037_)
  );
  DFF_X1 \rf[1][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01578_),
    .Q(\rf[1] [21]),
    .QN(_14036_)
  );
  DFF_X1 \rf[1][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01579_),
    .Q(\rf[1] [22]),
    .QN(_14035_)
  );
  DFF_X1 \rf[1][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01580_),
    .Q(\rf[1] [23]),
    .QN(_14034_)
  );
  DFF_X1 \rf[1][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01581_),
    .Q(\rf[1] [24]),
    .QN(_14033_)
  );
  DFF_X1 \rf[1][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01582_),
    .Q(\rf[1] [25]),
    .QN(_14032_)
  );
  DFF_X1 \rf[1][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01583_),
    .Q(\rf[1] [26]),
    .QN(_14031_)
  );
  DFF_X1 \rf[1][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01584_),
    .Q(\rf[1] [27]),
    .QN(_14030_)
  );
  DFF_X1 \rf[1][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01585_),
    .Q(\rf[1] [28]),
    .QN(_14029_)
  );
  DFF_X1 \rf[1][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01586_),
    .Q(\rf[1] [29]),
    .QN(_14028_)
  );
  DFF_X1 \rf[1][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01559_),
    .Q(\rf[1] [2]),
    .QN(_14055_)
  );
  DFF_X1 \rf[1][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01587_),
    .Q(\rf[1] [30]),
    .QN(_15562_)
  );
  DFF_X1 \rf[1][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00614_),
    .Q(\rf[1] [31]),
    .QN(_14999_)
  );
  DFF_X1 \rf[1][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01560_),
    .Q(\rf[1] [3]),
    .QN(_14054_)
  );
  DFF_X1 \rf[1][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01561_),
    .Q(\rf[1] [4]),
    .QN(_14053_)
  );
  DFF_X1 \rf[1][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01562_),
    .Q(\rf[1] [5]),
    .QN(_14052_)
  );
  DFF_X1 \rf[1][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01563_),
    .Q(\rf[1] [6]),
    .QN(_14051_)
  );
  DFF_X1 \rf[1][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01564_),
    .Q(\rf[1] [7]),
    .QN(_14050_)
  );
  DFF_X1 \rf[1][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01565_),
    .Q(\rf[1] [8]),
    .QN(_14049_)
  );
  DFF_X1 \rf[1][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01566_),
    .Q(\rf[1] [9]),
    .QN(_14048_)
  );
  DFF_X1 \rf[20][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01061_),
    .Q(\rf[20] [0]),
    .QN(_14553_)
  );
  DFF_X1 \rf[20][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01071_),
    .Q(\rf[20] [10]),
    .QN(_14543_)
  );
  DFF_X1 \rf[20][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01072_),
    .Q(\rf[20] [11]),
    .QN(_14542_)
  );
  DFF_X1 \rf[20][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01073_),
    .Q(\rf[20] [12]),
    .QN(_14541_)
  );
  DFF_X1 \rf[20][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01074_),
    .Q(\rf[20] [13]),
    .QN(_14540_)
  );
  DFF_X1 \rf[20][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01075_),
    .Q(\rf[20] [14]),
    .QN(_14539_)
  );
  DFF_X1 \rf[20][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01076_),
    .Q(\rf[20] [15]),
    .QN(_14538_)
  );
  DFF_X1 \rf[20][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01077_),
    .Q(\rf[20] [16]),
    .QN(_14537_)
  );
  DFF_X1 \rf[20][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01078_),
    .Q(\rf[20] [17]),
    .QN(_14536_)
  );
  DFF_X1 \rf[20][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01079_),
    .Q(\rf[20] [18]),
    .QN(_14535_)
  );
  DFF_X1 \rf[20][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01080_),
    .Q(\rf[20] [19]),
    .QN(_14534_)
  );
  DFF_X1 \rf[20][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01062_),
    .Q(\rf[20] [1]),
    .QN(_14552_)
  );
  DFF_X1 \rf[20][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01081_),
    .Q(\rf[20] [20]),
    .QN(_14533_)
  );
  DFF_X1 \rf[20][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01082_),
    .Q(\rf[20] [21]),
    .QN(_14532_)
  );
  DFF_X1 \rf[20][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01083_),
    .Q(\rf[20] [22]),
    .QN(_14531_)
  );
  DFF_X1 \rf[20][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01084_),
    .Q(\rf[20] [23]),
    .QN(_14530_)
  );
  DFF_X1 \rf[20][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01085_),
    .Q(\rf[20] [24]),
    .QN(_14529_)
  );
  DFF_X1 \rf[20][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01086_),
    .Q(\rf[20] [25]),
    .QN(_14528_)
  );
  DFF_X1 \rf[20][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01087_),
    .Q(\rf[20] [26]),
    .QN(_14527_)
  );
  DFF_X1 \rf[20][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01088_),
    .Q(\rf[20] [27]),
    .QN(_14526_)
  );
  DFF_X1 \rf[20][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01089_),
    .Q(\rf[20] [28]),
    .QN(_14525_)
  );
  DFF_X1 \rf[20][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01090_),
    .Q(\rf[20] [29]),
    .QN(_14524_)
  );
  DFF_X1 \rf[20][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01063_),
    .Q(\rf[20] [2]),
    .QN(_14551_)
  );
  DFF_X1 \rf[20][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01091_),
    .Q(\rf[20] [30]),
    .QN(_14523_)
  );
  DFF_X1 \rf[20][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00613_),
    .Q(\rf[20] [31]),
    .QN(_15000_)
  );
  DFF_X1 \rf[20][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01064_),
    .Q(\rf[20] [3]),
    .QN(_14550_)
  );
  DFF_X1 \rf[20][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01065_),
    .Q(\rf[20] [4]),
    .QN(_14549_)
  );
  DFF_X1 \rf[20][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01066_),
    .Q(\rf[20] [5]),
    .QN(_14548_)
  );
  DFF_X1 \rf[20][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01067_),
    .Q(\rf[20] [6]),
    .QN(_14547_)
  );
  DFF_X1 \rf[20][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01068_),
    .Q(\rf[20] [7]),
    .QN(_14546_)
  );
  DFF_X1 \rf[20][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01069_),
    .Q(\rf[20] [8]),
    .QN(_14545_)
  );
  DFF_X1 \rf[20][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01070_),
    .Q(\rf[20] [9]),
    .QN(_14544_)
  );
  DFF_X1 \rf[21][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01123_),
    .Q(\rf[21] [0]),
    .QN(_14491_)
  );
  DFF_X1 \rf[21][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01133_),
    .Q(\rf[21] [10]),
    .QN(_14481_)
  );
  DFF_X1 \rf[21][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01134_),
    .Q(\rf[21] [11]),
    .QN(_14480_)
  );
  DFF_X1 \rf[21][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01135_),
    .Q(\rf[21] [12]),
    .QN(_14479_)
  );
  DFF_X1 \rf[21][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01136_),
    .Q(\rf[21] [13]),
    .QN(_14478_)
  );
  DFF_X1 \rf[21][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01137_),
    .Q(\rf[21] [14]),
    .QN(_14477_)
  );
  DFF_X1 \rf[21][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01138_),
    .Q(\rf[21] [15]),
    .QN(_14476_)
  );
  DFF_X1 \rf[21][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01139_),
    .Q(\rf[21] [16]),
    .QN(_14475_)
  );
  DFF_X1 \rf[21][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01140_),
    .Q(\rf[21] [17]),
    .QN(_14474_)
  );
  DFF_X1 \rf[21][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01141_),
    .Q(\rf[21] [18]),
    .QN(_14473_)
  );
  DFF_X1 \rf[21][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01142_),
    .Q(\rf[21] [19]),
    .QN(_14472_)
  );
  DFF_X1 \rf[21][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01124_),
    .Q(\rf[21] [1]),
    .QN(_14490_)
  );
  DFF_X1 \rf[21][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01143_),
    .Q(\rf[21] [20]),
    .QN(_14471_)
  );
  DFF_X1 \rf[21][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01144_),
    .Q(\rf[21] [21]),
    .QN(_14470_)
  );
  DFF_X1 \rf[21][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01145_),
    .Q(\rf[21] [22]),
    .QN(_14469_)
  );
  DFF_X1 \rf[21][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01146_),
    .Q(\rf[21] [23]),
    .QN(_14468_)
  );
  DFF_X1 \rf[21][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01147_),
    .Q(\rf[21] [24]),
    .QN(_14467_)
  );
  DFF_X1 \rf[21][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01148_),
    .Q(\rf[21] [25]),
    .QN(_14466_)
  );
  DFF_X1 \rf[21][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01149_),
    .Q(\rf[21] [26]),
    .QN(_14465_)
  );
  DFF_X1 \rf[21][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01150_),
    .Q(\rf[21] [27]),
    .QN(_14464_)
  );
  DFF_X1 \rf[21][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01151_),
    .Q(\rf[21] [28]),
    .QN(_14463_)
  );
  DFF_X1 \rf[21][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01152_),
    .Q(\rf[21] [29]),
    .QN(_14462_)
  );
  DFF_X1 \rf[21][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01125_),
    .Q(\rf[21] [2]),
    .QN(_14489_)
  );
  DFF_X1 \rf[21][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01153_),
    .Q(\rf[21] [30]),
    .QN(_14461_)
  );
  DFF_X1 \rf[21][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00612_),
    .Q(\rf[21] [31]),
    .QN(_15001_)
  );
  DFF_X1 \rf[21][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01126_),
    .Q(\rf[21] [3]),
    .QN(_14488_)
  );
  DFF_X1 \rf[21][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01127_),
    .Q(\rf[21] [4]),
    .QN(_14487_)
  );
  DFF_X1 \rf[21][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01128_),
    .Q(\rf[21] [5]),
    .QN(_14486_)
  );
  DFF_X1 \rf[21][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01129_),
    .Q(\rf[21] [6]),
    .QN(_14485_)
  );
  DFF_X1 \rf[21][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01130_),
    .Q(\rf[21] [7]),
    .QN(_14484_)
  );
  DFF_X1 \rf[21][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01131_),
    .Q(\rf[21] [8]),
    .QN(_14483_)
  );
  DFF_X1 \rf[21][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01132_),
    .Q(\rf[21] [9]),
    .QN(_14482_)
  );
  DFF_X1 \rf[22][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01309_),
    .Q(\rf[22] [0]),
    .QN(_14305_)
  );
  DFF_X1 \rf[22][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01319_),
    .Q(\rf[22] [10]),
    .QN(_14295_)
  );
  DFF_X1 \rf[22][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01320_),
    .Q(\rf[22] [11]),
    .QN(_14294_)
  );
  DFF_X1 \rf[22][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01321_),
    .Q(\rf[22] [12]),
    .QN(_14293_)
  );
  DFF_X1 \rf[22][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01322_),
    .Q(\rf[22] [13]),
    .QN(_14292_)
  );
  DFF_X1 \rf[22][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01323_),
    .Q(\rf[22] [14]),
    .QN(_14291_)
  );
  DFF_X1 \rf[22][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01324_),
    .Q(\rf[22] [15]),
    .QN(_14290_)
  );
  DFF_X1 \rf[22][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01325_),
    .Q(\rf[22] [16]),
    .QN(_14289_)
  );
  DFF_X1 \rf[22][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01326_),
    .Q(\rf[22] [17]),
    .QN(_14288_)
  );
  DFF_X1 \rf[22][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01327_),
    .Q(\rf[22] [18]),
    .QN(_14287_)
  );
  DFF_X1 \rf[22][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01328_),
    .Q(\rf[22] [19]),
    .QN(_14286_)
  );
  DFF_X1 \rf[22][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01310_),
    .Q(\rf[22] [1]),
    .QN(_14304_)
  );
  DFF_X1 \rf[22][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01329_),
    .Q(\rf[22] [20]),
    .QN(_14285_)
  );
  DFF_X1 \rf[22][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01330_),
    .Q(\rf[22] [21]),
    .QN(_14284_)
  );
  DFF_X1 \rf[22][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01331_),
    .Q(\rf[22] [22]),
    .QN(_14283_)
  );
  DFF_X1 \rf[22][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01332_),
    .Q(\rf[22] [23]),
    .QN(_14282_)
  );
  DFF_X1 \rf[22][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01333_),
    .Q(\rf[22] [24]),
    .QN(_14281_)
  );
  DFF_X1 \rf[22][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01334_),
    .Q(\rf[22] [25]),
    .QN(_14280_)
  );
  DFF_X1 \rf[22][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01335_),
    .Q(\rf[22] [26]),
    .QN(_14279_)
  );
  DFF_X1 \rf[22][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01336_),
    .Q(\rf[22] [27]),
    .QN(_14278_)
  );
  DFF_X1 \rf[22][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01337_),
    .Q(\rf[22] [28]),
    .QN(_14277_)
  );
  DFF_X1 \rf[22][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01338_),
    .Q(\rf[22] [29]),
    .QN(_14276_)
  );
  DFF_X1 \rf[22][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01311_),
    .Q(\rf[22] [2]),
    .QN(_14303_)
  );
  DFF_X1 \rf[22][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01339_),
    .Q(\rf[22] [30]),
    .QN(_14275_)
  );
  DFF_X1 \rf[22][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00611_),
    .Q(\rf[22] [31]),
    .QN(_15002_)
  );
  DFF_X1 \rf[22][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01312_),
    .Q(\rf[22] [3]),
    .QN(_14302_)
  );
  DFF_X1 \rf[22][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01313_),
    .Q(\rf[22] [4]),
    .QN(_14301_)
  );
  DFF_X1 \rf[22][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01314_),
    .Q(\rf[22] [5]),
    .QN(_14300_)
  );
  DFF_X1 \rf[22][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01315_),
    .Q(\rf[22] [6]),
    .QN(_14299_)
  );
  DFF_X1 \rf[22][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01316_),
    .Q(\rf[22] [7]),
    .QN(_14298_)
  );
  DFF_X1 \rf[22][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01317_),
    .Q(\rf[22] [8]),
    .QN(_14297_)
  );
  DFF_X1 \rf[22][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01318_),
    .Q(\rf[22] [9]),
    .QN(_14296_)
  );
  DFF_X1 \rf[23][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00657_),
    .Q(\rf[23] [0]),
    .QN(_14956_)
  );
  DFF_X1 \rf[23][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00667_),
    .Q(\rf[23] [10]),
    .QN(_14946_)
  );
  DFF_X1 \rf[23][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00668_),
    .Q(\rf[23] [11]),
    .QN(_14945_)
  );
  DFF_X1 \rf[23][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00669_),
    .Q(\rf[23] [12]),
    .QN(_14944_)
  );
  DFF_X1 \rf[23][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00670_),
    .Q(\rf[23] [13]),
    .QN(_14943_)
  );
  DFF_X1 \rf[23][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00671_),
    .Q(\rf[23] [14]),
    .QN(_14942_)
  );
  DFF_X1 \rf[23][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00672_),
    .Q(\rf[23] [15]),
    .QN(_14941_)
  );
  DFF_X1 \rf[23][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00673_),
    .Q(\rf[23] [16]),
    .QN(_14940_)
  );
  DFF_X1 \rf[23][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00674_),
    .Q(\rf[23] [17]),
    .QN(_14939_)
  );
  DFF_X1 \rf[23][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00675_),
    .Q(\rf[23] [18]),
    .QN(_14938_)
  );
  DFF_X1 \rf[23][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00676_),
    .Q(\rf[23] [19]),
    .QN(_14937_)
  );
  DFF_X1 \rf[23][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00658_),
    .Q(\rf[23] [1]),
    .QN(_14955_)
  );
  DFF_X1 \rf[23][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00677_),
    .Q(\rf[23] [20]),
    .QN(_14936_)
  );
  DFF_X1 \rf[23][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00678_),
    .Q(\rf[23] [21]),
    .QN(_14935_)
  );
  DFF_X1 \rf[23][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00679_),
    .Q(\rf[23] [22]),
    .QN(_14934_)
  );
  DFF_X1 \rf[23][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00680_),
    .Q(\rf[23] [23]),
    .QN(_14933_)
  );
  DFF_X1 \rf[23][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00681_),
    .Q(\rf[23] [24]),
    .QN(_14932_)
  );
  DFF_X1 \rf[23][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00682_),
    .Q(\rf[23] [25]),
    .QN(_14931_)
  );
  DFF_X1 \rf[23][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00683_),
    .Q(\rf[23] [26]),
    .QN(_14930_)
  );
  DFF_X1 \rf[23][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00684_),
    .Q(\rf[23] [27]),
    .QN(_14929_)
  );
  DFF_X1 \rf[23][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00685_),
    .Q(\rf[23] [28]),
    .QN(_14928_)
  );
  DFF_X1 \rf[23][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00686_),
    .Q(\rf[23] [29]),
    .QN(_14927_)
  );
  DFF_X1 \rf[23][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00659_),
    .Q(\rf[23] [2]),
    .QN(_14954_)
  );
  DFF_X1 \rf[23][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00687_),
    .Q(\rf[23] [30]),
    .QN(_14926_)
  );
  DFF_X1 \rf[23][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00610_),
    .Q(\rf[23] [31]),
    .QN(_15003_)
  );
  DFF_X1 \rf[23][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00660_),
    .Q(\rf[23] [3]),
    .QN(_14953_)
  );
  DFF_X1 \rf[23][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00661_),
    .Q(\rf[23] [4]),
    .QN(_14952_)
  );
  DFF_X1 \rf[23][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00662_),
    .Q(\rf[23] [5]),
    .QN(_14951_)
  );
  DFF_X1 \rf[23][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00663_),
    .Q(\rf[23] [6]),
    .QN(_14950_)
  );
  DFF_X1 \rf[23][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00664_),
    .Q(\rf[23] [7]),
    .QN(_14949_)
  );
  DFF_X1 \rf[23][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00665_),
    .Q(\rf[23] [8]),
    .QN(_14948_)
  );
  DFF_X1 \rf[23][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00666_),
    .Q(\rf[23] [9]),
    .QN(_14947_)
  );
  DFF_X1 \rf[24][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01433_),
    .Q(\rf[24] [0]),
    .QN(_14181_)
  );
  DFF_X1 \rf[24][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01443_),
    .Q(\rf[24] [10]),
    .QN(_14171_)
  );
  DFF_X1 \rf[24][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01444_),
    .Q(\rf[24] [11]),
    .QN(_14170_)
  );
  DFF_X1 \rf[24][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01445_),
    .Q(\rf[24] [12]),
    .QN(_14169_)
  );
  DFF_X1 \rf[24][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01446_),
    .Q(\rf[24] [13]),
    .QN(_14168_)
  );
  DFF_X1 \rf[24][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01447_),
    .Q(\rf[24] [14]),
    .QN(_14167_)
  );
  DFF_X1 \rf[24][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01448_),
    .Q(\rf[24] [15]),
    .QN(_14166_)
  );
  DFF_X1 \rf[24][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01449_),
    .Q(\rf[24] [16]),
    .QN(_14165_)
  );
  DFF_X1 \rf[24][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01450_),
    .Q(\rf[24] [17]),
    .QN(_14164_)
  );
  DFF_X1 \rf[24][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01451_),
    .Q(\rf[24] [18]),
    .QN(_14163_)
  );
  DFF_X1 \rf[24][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01452_),
    .Q(\rf[24] [19]),
    .QN(_14162_)
  );
  DFF_X1 \rf[24][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01434_),
    .Q(\rf[24] [1]),
    .QN(_14180_)
  );
  DFF_X1 \rf[24][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01453_),
    .Q(\rf[24] [20]),
    .QN(_14161_)
  );
  DFF_X1 \rf[24][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01454_),
    .Q(\rf[24] [21]),
    .QN(_14160_)
  );
  DFF_X1 \rf[24][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01455_),
    .Q(\rf[24] [22]),
    .QN(_14159_)
  );
  DFF_X1 \rf[24][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01456_),
    .Q(\rf[24] [23]),
    .QN(_14158_)
  );
  DFF_X1 \rf[24][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01457_),
    .Q(\rf[24] [24]),
    .QN(_14157_)
  );
  DFF_X1 \rf[24][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01458_),
    .Q(\rf[24] [25]),
    .QN(_14156_)
  );
  DFF_X1 \rf[24][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01459_),
    .Q(\rf[24] [26]),
    .QN(_14155_)
  );
  DFF_X1 \rf[24][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01460_),
    .Q(\rf[24] [27]),
    .QN(_14154_)
  );
  DFF_X1 \rf[24][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01461_),
    .Q(\rf[24] [28]),
    .QN(_14153_)
  );
  DFF_X1 \rf[24][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01462_),
    .Q(\rf[24] [29]),
    .QN(_14152_)
  );
  DFF_X1 \rf[24][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01435_),
    .Q(\rf[24] [2]),
    .QN(_14179_)
  );
  DFF_X1 \rf[24][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01463_),
    .Q(\rf[24] [30]),
    .QN(_14151_)
  );
  DFF_X1 \rf[24][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00609_),
    .Q(\rf[24] [31]),
    .QN(_15004_)
  );
  DFF_X1 \rf[24][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01436_),
    .Q(\rf[24] [3]),
    .QN(_14178_)
  );
  DFF_X1 \rf[24][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01437_),
    .Q(\rf[24] [4]),
    .QN(_14177_)
  );
  DFF_X1 \rf[24][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01438_),
    .Q(\rf[24] [5]),
    .QN(_14176_)
  );
  DFF_X1 \rf[24][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01439_),
    .Q(\rf[24] [6]),
    .QN(_14175_)
  );
  DFF_X1 \rf[24][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01440_),
    .Q(\rf[24] [7]),
    .QN(_14174_)
  );
  DFF_X1 \rf[24][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01441_),
    .Q(\rf[24] [8]),
    .QN(_14173_)
  );
  DFF_X1 \rf[24][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01442_),
    .Q(\rf[24] [9]),
    .QN(_14172_)
  );
  DFF_X1 \rf[25][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00626_),
    .Q(\rf[25] [0]),
    .QN(_14987_)
  );
  DFF_X1 \rf[25][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00636_),
    .Q(\rf[25] [10]),
    .QN(_14977_)
  );
  DFF_X1 \rf[25][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00637_),
    .Q(\rf[25] [11]),
    .QN(_14976_)
  );
  DFF_X1 \rf[25][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00638_),
    .Q(\rf[25] [12]),
    .QN(_14975_)
  );
  DFF_X1 \rf[25][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00639_),
    .Q(\rf[25] [13]),
    .QN(_14974_)
  );
  DFF_X1 \rf[25][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00640_),
    .Q(\rf[25] [14]),
    .QN(_14973_)
  );
  DFF_X1 \rf[25][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00641_),
    .Q(\rf[25] [15]),
    .QN(_14972_)
  );
  DFF_X1 \rf[25][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00642_),
    .Q(\rf[25] [16]),
    .QN(_14971_)
  );
  DFF_X1 \rf[25][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00643_),
    .Q(\rf[25] [17]),
    .QN(_14970_)
  );
  DFF_X1 \rf[25][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00644_),
    .Q(\rf[25] [18]),
    .QN(_14969_)
  );
  DFF_X1 \rf[25][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00645_),
    .Q(\rf[25] [19]),
    .QN(_14968_)
  );
  DFF_X1 \rf[25][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00627_),
    .Q(\rf[25] [1]),
    .QN(_14986_)
  );
  DFF_X1 \rf[25][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00646_),
    .Q(\rf[25] [20]),
    .QN(_14967_)
  );
  DFF_X1 \rf[25][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00647_),
    .Q(\rf[25] [21]),
    .QN(_14966_)
  );
  DFF_X1 \rf[25][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00648_),
    .Q(\rf[25] [22]),
    .QN(_14965_)
  );
  DFF_X1 \rf[25][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00649_),
    .Q(\rf[25] [23]),
    .QN(_14964_)
  );
  DFF_X1 \rf[25][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00650_),
    .Q(\rf[25] [24]),
    .QN(_14963_)
  );
  DFF_X1 \rf[25][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00651_),
    .Q(\rf[25] [25]),
    .QN(_14962_)
  );
  DFF_X1 \rf[25][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00652_),
    .Q(\rf[25] [26]),
    .QN(_14961_)
  );
  DFF_X1 \rf[25][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00653_),
    .Q(\rf[25] [27]),
    .QN(_14960_)
  );
  DFF_X1 \rf[25][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00654_),
    .Q(\rf[25] [28]),
    .QN(_14959_)
  );
  DFF_X1 \rf[25][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00655_),
    .Q(\rf[25] [29]),
    .QN(_14958_)
  );
  DFF_X1 \rf[25][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00628_),
    .Q(\rf[25] [2]),
    .QN(_14985_)
  );
  DFF_X1 \rf[25][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00656_),
    .Q(\rf[25] [30]),
    .QN(_14957_)
  );
  DFF_X1 \rf[25][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00608_),
    .Q(\rf[25] [31]),
    .QN(_15005_)
  );
  DFF_X1 \rf[25][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00629_),
    .Q(\rf[25] [3]),
    .QN(_14984_)
  );
  DFF_X1 \rf[25][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00630_),
    .Q(\rf[25] [4]),
    .QN(_14983_)
  );
  DFF_X1 \rf[25][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00631_),
    .Q(\rf[25] [5]),
    .QN(_14982_)
  );
  DFF_X1 \rf[25][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00632_),
    .Q(\rf[25] [6]),
    .QN(_14981_)
  );
  DFF_X1 \rf[25][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00633_),
    .Q(\rf[25] [7]),
    .QN(_14980_)
  );
  DFF_X1 \rf[25][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00634_),
    .Q(\rf[25] [8]),
    .QN(_14979_)
  );
  DFF_X1 \rf[25][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00635_),
    .Q(\rf[25] [9]),
    .QN(_14978_)
  );
  DFF_X1 \rf[26][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01340_),
    .Q(\rf[26] [0]),
    .QN(_14274_)
  );
  DFF_X1 \rf[26][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01350_),
    .Q(\rf[26] [10]),
    .QN(_14264_)
  );
  DFF_X1 \rf[26][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01351_),
    .Q(\rf[26] [11]),
    .QN(_14263_)
  );
  DFF_X1 \rf[26][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01352_),
    .Q(\rf[26] [12]),
    .QN(_14262_)
  );
  DFF_X1 \rf[26][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01353_),
    .Q(\rf[26] [13]),
    .QN(_14261_)
  );
  DFF_X1 \rf[26][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01354_),
    .Q(\rf[26] [14]),
    .QN(_14260_)
  );
  DFF_X1 \rf[26][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01355_),
    .Q(\rf[26] [15]),
    .QN(_14259_)
  );
  DFF_X1 \rf[26][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01356_),
    .Q(\rf[26] [16]),
    .QN(_14258_)
  );
  DFF_X1 \rf[26][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01357_),
    .Q(\rf[26] [17]),
    .QN(_14257_)
  );
  DFF_X1 \rf[26][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01358_),
    .Q(\rf[26] [18]),
    .QN(_14256_)
  );
  DFF_X1 \rf[26][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01359_),
    .Q(\rf[26] [19]),
    .QN(_14255_)
  );
  DFF_X1 \rf[26][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01341_),
    .Q(\rf[26] [1]),
    .QN(_14273_)
  );
  DFF_X1 \rf[26][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01360_),
    .Q(\rf[26] [20]),
    .QN(_14254_)
  );
  DFF_X1 \rf[26][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01361_),
    .Q(\rf[26] [21]),
    .QN(_14253_)
  );
  DFF_X1 \rf[26][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01362_),
    .Q(\rf[26] [22]),
    .QN(_14252_)
  );
  DFF_X1 \rf[26][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01363_),
    .Q(\rf[26] [23]),
    .QN(_14251_)
  );
  DFF_X1 \rf[26][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01364_),
    .Q(\rf[26] [24]),
    .QN(_14250_)
  );
  DFF_X1 \rf[26][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01365_),
    .Q(\rf[26] [25]),
    .QN(_14249_)
  );
  DFF_X1 \rf[26][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01366_),
    .Q(\rf[26] [26]),
    .QN(_14248_)
  );
  DFF_X1 \rf[26][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01367_),
    .Q(\rf[26] [27]),
    .QN(_14247_)
  );
  DFF_X1 \rf[26][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01368_),
    .Q(\rf[26] [28]),
    .QN(_14246_)
  );
  DFF_X1 \rf[26][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01369_),
    .Q(\rf[26] [29]),
    .QN(_14245_)
  );
  DFF_X1 \rf[26][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01342_),
    .Q(\rf[26] [2]),
    .QN(_14272_)
  );
  DFF_X1 \rf[26][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01370_),
    .Q(\rf[26] [30]),
    .QN(_14244_)
  );
  DFF_X1 \rf[26][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00607_),
    .Q(\rf[26] [31]),
    .QN(_15006_)
  );
  DFF_X1 \rf[26][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01343_),
    .Q(\rf[26] [3]),
    .QN(_14271_)
  );
  DFF_X1 \rf[26][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01344_),
    .Q(\rf[26] [4]),
    .QN(_14270_)
  );
  DFF_X1 \rf[26][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01345_),
    .Q(\rf[26] [5]),
    .QN(_14269_)
  );
  DFF_X1 \rf[26][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01346_),
    .Q(\rf[26] [6]),
    .QN(_14268_)
  );
  DFF_X1 \rf[26][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01347_),
    .Q(\rf[26] [7]),
    .QN(_14267_)
  );
  DFF_X1 \rf[26][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01348_),
    .Q(\rf[26] [8]),
    .QN(_14266_)
  );
  DFF_X1 \rf[26][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01349_),
    .Q(\rf[26] [9]),
    .QN(_14265_)
  );
  DFF_X1 \rf[27][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01402_),
    .Q(\rf[27] [0]),
    .QN(_14212_)
  );
  DFF_X1 \rf[27][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01412_),
    .Q(\rf[27] [10]),
    .QN(_14202_)
  );
  DFF_X1 \rf[27][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01413_),
    .Q(\rf[27] [11]),
    .QN(_14201_)
  );
  DFF_X1 \rf[27][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01414_),
    .Q(\rf[27] [12]),
    .QN(_14200_)
  );
  DFF_X1 \rf[27][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01415_),
    .Q(\rf[27] [13]),
    .QN(_14199_)
  );
  DFF_X1 \rf[27][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01416_),
    .Q(\rf[27] [14]),
    .QN(_14198_)
  );
  DFF_X1 \rf[27][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01417_),
    .Q(\rf[27] [15]),
    .QN(_14197_)
  );
  DFF_X1 \rf[27][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01418_),
    .Q(\rf[27] [16]),
    .QN(_14196_)
  );
  DFF_X1 \rf[27][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01419_),
    .Q(\rf[27] [17]),
    .QN(_14195_)
  );
  DFF_X1 \rf[27][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01420_),
    .Q(\rf[27] [18]),
    .QN(_14194_)
  );
  DFF_X1 \rf[27][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01421_),
    .Q(\rf[27] [19]),
    .QN(_14193_)
  );
  DFF_X1 \rf[27][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01403_),
    .Q(\rf[27] [1]),
    .QN(_14211_)
  );
  DFF_X1 \rf[27][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01422_),
    .Q(\rf[27] [20]),
    .QN(_14192_)
  );
  DFF_X1 \rf[27][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01423_),
    .Q(\rf[27] [21]),
    .QN(_14191_)
  );
  DFF_X1 \rf[27][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01424_),
    .Q(\rf[27] [22]),
    .QN(_14190_)
  );
  DFF_X1 \rf[27][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01425_),
    .Q(\rf[27] [23]),
    .QN(_14189_)
  );
  DFF_X1 \rf[27][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01426_),
    .Q(\rf[27] [24]),
    .QN(_14188_)
  );
  DFF_X1 \rf[27][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01427_),
    .Q(\rf[27] [25]),
    .QN(_14187_)
  );
  DFF_X1 \rf[27][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01428_),
    .Q(\rf[27] [26]),
    .QN(_14186_)
  );
  DFF_X1 \rf[27][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01429_),
    .Q(\rf[27] [27]),
    .QN(_14185_)
  );
  DFF_X1 \rf[27][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01430_),
    .Q(\rf[27] [28]),
    .QN(_14184_)
  );
  DFF_X1 \rf[27][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01431_),
    .Q(\rf[27] [29]),
    .QN(_14183_)
  );
  DFF_X1 \rf[27][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01404_),
    .Q(\rf[27] [2]),
    .QN(_14210_)
  );
  DFF_X1 \rf[27][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01432_),
    .Q(\rf[27] [30]),
    .QN(_14182_)
  );
  DFF_X1 \rf[27][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00606_),
    .Q(\rf[27] [31]),
    .QN(_15007_)
  );
  DFF_X1 \rf[27][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01405_),
    .Q(\rf[27] [3]),
    .QN(_14209_)
  );
  DFF_X1 \rf[27][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01406_),
    .Q(\rf[27] [4]),
    .QN(_14208_)
  );
  DFF_X1 \rf[27][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01407_),
    .Q(\rf[27] [5]),
    .QN(_14207_)
  );
  DFF_X1 \rf[27][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01408_),
    .Q(\rf[27] [6]),
    .QN(_14206_)
  );
  DFF_X1 \rf[27][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01409_),
    .Q(\rf[27] [7]),
    .QN(_14205_)
  );
  DFF_X1 \rf[27][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01410_),
    .Q(\rf[27] [8]),
    .QN(_14204_)
  );
  DFF_X1 \rf[27][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01411_),
    .Q(\rf[27] [9]),
    .QN(_14203_)
  );
  DFF_X1 \rf[28][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01185_),
    .Q(\rf[28] [0]),
    .QN(_14429_)
  );
  DFF_X1 \rf[28][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01195_),
    .Q(\rf[28] [10]),
    .QN(_14419_)
  );
  DFF_X1 \rf[28][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01196_),
    .Q(\rf[28] [11]),
    .QN(_14418_)
  );
  DFF_X1 \rf[28][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01197_),
    .Q(\rf[28] [12]),
    .QN(_14417_)
  );
  DFF_X1 \rf[28][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01198_),
    .Q(\rf[28] [13]),
    .QN(_14416_)
  );
  DFF_X1 \rf[28][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01199_),
    .Q(\rf[28] [14]),
    .QN(_14415_)
  );
  DFF_X1 \rf[28][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01200_),
    .Q(\rf[28] [15]),
    .QN(_14414_)
  );
  DFF_X1 \rf[28][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01201_),
    .Q(\rf[28] [16]),
    .QN(_14413_)
  );
  DFF_X1 \rf[28][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01202_),
    .Q(\rf[28] [17]),
    .QN(_14412_)
  );
  DFF_X1 \rf[28][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01203_),
    .Q(\rf[28] [18]),
    .QN(_14411_)
  );
  DFF_X1 \rf[28][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01204_),
    .Q(\rf[28] [19]),
    .QN(_14410_)
  );
  DFF_X1 \rf[28][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01186_),
    .Q(\rf[28] [1]),
    .QN(_14428_)
  );
  DFF_X1 \rf[28][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01205_),
    .Q(\rf[28] [20]),
    .QN(_14409_)
  );
  DFF_X1 \rf[28][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01206_),
    .Q(\rf[28] [21]),
    .QN(_14408_)
  );
  DFF_X1 \rf[28][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01207_),
    .Q(\rf[28] [22]),
    .QN(_14407_)
  );
  DFF_X1 \rf[28][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01208_),
    .Q(\rf[28] [23]),
    .QN(_14406_)
  );
  DFF_X1 \rf[28][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01209_),
    .Q(\rf[28] [24]),
    .QN(_14405_)
  );
  DFF_X1 \rf[28][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01210_),
    .Q(\rf[28] [25]),
    .QN(_14404_)
  );
  DFF_X1 \rf[28][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01211_),
    .Q(\rf[28] [26]),
    .QN(_14403_)
  );
  DFF_X1 \rf[28][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01212_),
    .Q(\rf[28] [27]),
    .QN(_14402_)
  );
  DFF_X1 \rf[28][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01213_),
    .Q(\rf[28] [28]),
    .QN(_14401_)
  );
  DFF_X1 \rf[28][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01214_),
    .Q(\rf[28] [29]),
    .QN(_14400_)
  );
  DFF_X1 \rf[28][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01187_),
    .Q(\rf[28] [2]),
    .QN(_14427_)
  );
  DFF_X1 \rf[28][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01215_),
    .Q(\rf[28] [30]),
    .QN(_14399_)
  );
  DFF_X1 \rf[28][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00605_),
    .Q(\rf[28] [31]),
    .QN(_15008_)
  );
  DFF_X1 \rf[28][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01188_),
    .Q(\rf[28] [3]),
    .QN(_14426_)
  );
  DFF_X1 \rf[28][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01189_),
    .Q(\rf[28] [4]),
    .QN(_14425_)
  );
  DFF_X1 \rf[28][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01190_),
    .Q(\rf[28] [5]),
    .QN(_14424_)
  );
  DFF_X1 \rf[28][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01191_),
    .Q(\rf[28] [6]),
    .QN(_14423_)
  );
  DFF_X1 \rf[28][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01192_),
    .Q(\rf[28] [7]),
    .QN(_14422_)
  );
  DFF_X1 \rf[28][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01193_),
    .Q(\rf[28] [8]),
    .QN(_14421_)
  );
  DFF_X1 \rf[28][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01194_),
    .Q(\rf[28] [9]),
    .QN(_14420_)
  );
  DFF_X1 \rf[29][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01216_),
    .Q(\rf[29] [0]),
    .QN(_14398_)
  );
  DFF_X1 \rf[29][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01226_),
    .Q(\rf[29] [10]),
    .QN(_14388_)
  );
  DFF_X1 \rf[29][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01227_),
    .Q(\rf[29] [11]),
    .QN(_14387_)
  );
  DFF_X1 \rf[29][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01228_),
    .Q(\rf[29] [12]),
    .QN(_14386_)
  );
  DFF_X1 \rf[29][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01229_),
    .Q(\rf[29] [13]),
    .QN(_14385_)
  );
  DFF_X1 \rf[29][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01230_),
    .Q(\rf[29] [14]),
    .QN(_14384_)
  );
  DFF_X1 \rf[29][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01231_),
    .Q(\rf[29] [15]),
    .QN(_14383_)
  );
  DFF_X1 \rf[29][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01232_),
    .Q(\rf[29] [16]),
    .QN(_14382_)
  );
  DFF_X1 \rf[29][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01233_),
    .Q(\rf[29] [17]),
    .QN(_14381_)
  );
  DFF_X1 \rf[29][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01234_),
    .Q(\rf[29] [18]),
    .QN(_14380_)
  );
  DFF_X1 \rf[29][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01235_),
    .Q(\rf[29] [19]),
    .QN(_14379_)
  );
  DFF_X1 \rf[29][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01217_),
    .Q(\rf[29] [1]),
    .QN(_14397_)
  );
  DFF_X1 \rf[29][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01236_),
    .Q(\rf[29] [20]),
    .QN(_14378_)
  );
  DFF_X1 \rf[29][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01237_),
    .Q(\rf[29] [21]),
    .QN(_14377_)
  );
  DFF_X1 \rf[29][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01238_),
    .Q(\rf[29] [22]),
    .QN(_14376_)
  );
  DFF_X1 \rf[29][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01239_),
    .Q(\rf[29] [23]),
    .QN(_14375_)
  );
  DFF_X1 \rf[29][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01240_),
    .Q(\rf[29] [24]),
    .QN(_14374_)
  );
  DFF_X1 \rf[29][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01241_),
    .Q(\rf[29] [25]),
    .QN(_14373_)
  );
  DFF_X1 \rf[29][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01242_),
    .Q(\rf[29] [26]),
    .QN(_14372_)
  );
  DFF_X1 \rf[29][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01243_),
    .Q(\rf[29] [27]),
    .QN(_14371_)
  );
  DFF_X1 \rf[29][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01244_),
    .Q(\rf[29] [28]),
    .QN(_14370_)
  );
  DFF_X1 \rf[29][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01245_),
    .Q(\rf[29] [29]),
    .QN(_14369_)
  );
  DFF_X1 \rf[29][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01218_),
    .Q(\rf[29] [2]),
    .QN(_14396_)
  );
  DFF_X1 \rf[29][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01246_),
    .Q(\rf[29] [30]),
    .QN(_14368_)
  );
  DFF_X1 \rf[29][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00604_),
    .Q(\rf[29] [31]),
    .QN(_15009_)
  );
  DFF_X1 \rf[29][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01219_),
    .Q(\rf[29] [3]),
    .QN(_14395_)
  );
  DFF_X1 \rf[29][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01220_),
    .Q(\rf[29] [4]),
    .QN(_14394_)
  );
  DFF_X1 \rf[29][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01221_),
    .Q(\rf[29] [5]),
    .QN(_14393_)
  );
  DFF_X1 \rf[29][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01222_),
    .Q(\rf[29] [6]),
    .QN(_14392_)
  );
  DFF_X1 \rf[29][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01223_),
    .Q(\rf[29] [7]),
    .QN(_14391_)
  );
  DFF_X1 \rf[29][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01224_),
    .Q(\rf[29] [8]),
    .QN(_14390_)
  );
  DFF_X1 \rf[29][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01225_),
    .Q(\rf[29] [9]),
    .QN(_14389_)
  );
  DFF_X1 \rf[2][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01371_),
    .Q(\rf[2] [0]),
    .QN(_14243_)
  );
  DFF_X1 \rf[2][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01381_),
    .Q(\rf[2] [10]),
    .QN(_14233_)
  );
  DFF_X1 \rf[2][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01382_),
    .Q(\rf[2] [11]),
    .QN(_14232_)
  );
  DFF_X1 \rf[2][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01383_),
    .Q(\rf[2] [12]),
    .QN(_14231_)
  );
  DFF_X1 \rf[2][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01384_),
    .Q(\rf[2] [13]),
    .QN(_14230_)
  );
  DFF_X1 \rf[2][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01385_),
    .Q(\rf[2] [14]),
    .QN(_14229_)
  );
  DFF_X1 \rf[2][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01386_),
    .Q(\rf[2] [15]),
    .QN(_14228_)
  );
  DFF_X1 \rf[2][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01387_),
    .Q(\rf[2] [16]),
    .QN(_14227_)
  );
  DFF_X1 \rf[2][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01388_),
    .Q(\rf[2] [17]),
    .QN(_14226_)
  );
  DFF_X1 \rf[2][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01389_),
    .Q(\rf[2] [18]),
    .QN(_14225_)
  );
  DFF_X1 \rf[2][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01390_),
    .Q(\rf[2] [19]),
    .QN(_14224_)
  );
  DFF_X1 \rf[2][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01372_),
    .Q(\rf[2] [1]),
    .QN(_14242_)
  );
  DFF_X1 \rf[2][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01391_),
    .Q(\rf[2] [20]),
    .QN(_14223_)
  );
  DFF_X1 \rf[2][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01392_),
    .Q(\rf[2] [21]),
    .QN(_14222_)
  );
  DFF_X1 \rf[2][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01393_),
    .Q(\rf[2] [22]),
    .QN(_14221_)
  );
  DFF_X1 \rf[2][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01394_),
    .Q(\rf[2] [23]),
    .QN(_14220_)
  );
  DFF_X1 \rf[2][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01395_),
    .Q(\rf[2] [24]),
    .QN(_14219_)
  );
  DFF_X1 \rf[2][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01396_),
    .Q(\rf[2] [25]),
    .QN(_14218_)
  );
  DFF_X1 \rf[2][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01397_),
    .Q(\rf[2] [26]),
    .QN(_14217_)
  );
  DFF_X1 \rf[2][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01398_),
    .Q(\rf[2] [27]),
    .QN(_14216_)
  );
  DFF_X1 \rf[2][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01399_),
    .Q(\rf[2] [28]),
    .QN(_14215_)
  );
  DFF_X1 \rf[2][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01400_),
    .Q(\rf[2] [29]),
    .QN(_14214_)
  );
  DFF_X1 \rf[2][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01373_),
    .Q(\rf[2] [2]),
    .QN(_14241_)
  );
  DFF_X1 \rf[2][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01401_),
    .Q(\rf[2] [30]),
    .QN(_14213_)
  );
  DFF_X1 \rf[2][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00603_),
    .Q(\rf[2] [31]),
    .QN(_15010_)
  );
  DFF_X1 \rf[2][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01374_),
    .Q(\rf[2] [3]),
    .QN(_14240_)
  );
  DFF_X1 \rf[2][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01375_),
    .Q(\rf[2] [4]),
    .QN(_14239_)
  );
  DFF_X1 \rf[2][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01376_),
    .Q(\rf[2] [5]),
    .QN(_14238_)
  );
  DFF_X1 \rf[2][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01377_),
    .Q(\rf[2] [6]),
    .QN(_14237_)
  );
  DFF_X1 \rf[2][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01378_),
    .Q(\rf[2] [7]),
    .QN(_14236_)
  );
  DFF_X1 \rf[2][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01379_),
    .Q(\rf[2] [8]),
    .QN(_14235_)
  );
  DFF_X1 \rf[2][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01380_),
    .Q(\rf[2] [9]),
    .QN(_14234_)
  );
  DFF_X1 \rf[30][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01247_),
    .Q(\rf[30] [0]),
    .QN(_14367_)
  );
  DFF_X1 \rf[30][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01257_),
    .Q(\rf[30] [10]),
    .QN(_14357_)
  );
  DFF_X1 \rf[30][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01258_),
    .Q(\rf[30] [11]),
    .QN(_14356_)
  );
  DFF_X1 \rf[30][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01259_),
    .Q(\rf[30] [12]),
    .QN(_14355_)
  );
  DFF_X1 \rf[30][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01260_),
    .Q(\rf[30] [13]),
    .QN(_14354_)
  );
  DFF_X1 \rf[30][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01261_),
    .Q(\rf[30] [14]),
    .QN(_14353_)
  );
  DFF_X1 \rf[30][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01262_),
    .Q(\rf[30] [15]),
    .QN(_14352_)
  );
  DFF_X1 \rf[30][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01263_),
    .Q(\rf[30] [16]),
    .QN(_14351_)
  );
  DFF_X1 \rf[30][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01264_),
    .Q(\rf[30] [17]),
    .QN(_14350_)
  );
  DFF_X1 \rf[30][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01265_),
    .Q(\rf[30] [18]),
    .QN(_14349_)
  );
  DFF_X1 \rf[30][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01266_),
    .Q(\rf[30] [19]),
    .QN(_14348_)
  );
  DFF_X1 \rf[30][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01248_),
    .Q(\rf[30] [1]),
    .QN(_14366_)
  );
  DFF_X1 \rf[30][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01267_),
    .Q(\rf[30] [20]),
    .QN(_14347_)
  );
  DFF_X1 \rf[30][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01268_),
    .Q(\rf[30] [21]),
    .QN(_14346_)
  );
  DFF_X1 \rf[30][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01269_),
    .Q(\rf[30] [22]),
    .QN(_14345_)
  );
  DFF_X1 \rf[30][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01270_),
    .Q(\rf[30] [23]),
    .QN(_14344_)
  );
  DFF_X1 \rf[30][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01271_),
    .Q(\rf[30] [24]),
    .QN(_14343_)
  );
  DFF_X1 \rf[30][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01272_),
    .Q(\rf[30] [25]),
    .QN(_14342_)
  );
  DFF_X1 \rf[30][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01273_),
    .Q(\rf[30] [26]),
    .QN(_14341_)
  );
  DFF_X1 \rf[30][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01274_),
    .Q(\rf[30] [27]),
    .QN(_14340_)
  );
  DFF_X1 \rf[30][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01275_),
    .Q(\rf[30] [28]),
    .QN(_14339_)
  );
  DFF_X1 \rf[30][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01276_),
    .Q(\rf[30] [29]),
    .QN(_14338_)
  );
  DFF_X1 \rf[30][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01249_),
    .Q(\rf[30] [2]),
    .QN(_14365_)
  );
  DFF_X1 \rf[30][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01277_),
    .Q(\rf[30] [30]),
    .QN(_14337_)
  );
  DFF_X1 \rf[30][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00602_),
    .Q(\rf[30] [31]),
    .QN(_15011_)
  );
  DFF_X1 \rf[30][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01250_),
    .Q(\rf[30] [3]),
    .QN(_14364_)
  );
  DFF_X1 \rf[30][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01251_),
    .Q(\rf[30] [4]),
    .QN(_14363_)
  );
  DFF_X1 \rf[30][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01252_),
    .Q(\rf[30] [5]),
    .QN(_14362_)
  );
  DFF_X1 \rf[30][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01253_),
    .Q(\rf[30] [6]),
    .QN(_14361_)
  );
  DFF_X1 \rf[30][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01254_),
    .Q(\rf[30] [7]),
    .QN(_14360_)
  );
  DFF_X1 \rf[30][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01255_),
    .Q(\rf[30] [8]),
    .QN(_14359_)
  );
  DFF_X1 \rf[30][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01256_),
    .Q(\rf[30] [9]),
    .QN(_14358_)
  );
  DFF_X1 \rf[3][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01526_),
    .Q(\rf[3] [0]),
    .QN(_14088_)
  );
  DFF_X1 \rf[3][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01536_),
    .Q(\rf[3] [10]),
    .QN(_14078_)
  );
  DFF_X1 \rf[3][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01537_),
    .Q(\rf[3] [11]),
    .QN(_14077_)
  );
  DFF_X1 \rf[3][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01538_),
    .Q(\rf[3] [12]),
    .QN(_14076_)
  );
  DFF_X1 \rf[3][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01539_),
    .Q(\rf[3] [13]),
    .QN(_14075_)
  );
  DFF_X1 \rf[3][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01540_),
    .Q(\rf[3] [14]),
    .QN(_14074_)
  );
  DFF_X1 \rf[3][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01541_),
    .Q(\rf[3] [15]),
    .QN(_14073_)
  );
  DFF_X1 \rf[3][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01542_),
    .Q(\rf[3] [16]),
    .QN(_14072_)
  );
  DFF_X1 \rf[3][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01543_),
    .Q(\rf[3] [17]),
    .QN(_14071_)
  );
  DFF_X1 \rf[3][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01544_),
    .Q(\rf[3] [18]),
    .QN(_14070_)
  );
  DFF_X1 \rf[3][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01545_),
    .Q(\rf[3] [19]),
    .QN(_14069_)
  );
  DFF_X1 \rf[3][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01527_),
    .Q(\rf[3] [1]),
    .QN(_14087_)
  );
  DFF_X1 \rf[3][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01546_),
    .Q(\rf[3] [20]),
    .QN(_14068_)
  );
  DFF_X1 \rf[3][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01547_),
    .Q(\rf[3] [21]),
    .QN(_14067_)
  );
  DFF_X1 \rf[3][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01548_),
    .Q(\rf[3] [22]),
    .QN(_14066_)
  );
  DFF_X1 \rf[3][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01549_),
    .Q(\rf[3] [23]),
    .QN(_14065_)
  );
  DFF_X1 \rf[3][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01550_),
    .Q(\rf[3] [24]),
    .QN(_14064_)
  );
  DFF_X1 \rf[3][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01551_),
    .Q(\rf[3] [25]),
    .QN(_14063_)
  );
  DFF_X1 \rf[3][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01552_),
    .Q(\rf[3] [26]),
    .QN(_14062_)
  );
  DFF_X1 \rf[3][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01553_),
    .Q(\rf[3] [27]),
    .QN(_14061_)
  );
  DFF_X1 \rf[3][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01554_),
    .Q(\rf[3] [28]),
    .QN(_14060_)
  );
  DFF_X1 \rf[3][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01555_),
    .Q(\rf[3] [29]),
    .QN(_14059_)
  );
  DFF_X1 \rf[3][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01528_),
    .Q(\rf[3] [2]),
    .QN(_14086_)
  );
  DFF_X1 \rf[3][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01556_),
    .Q(\rf[3] [30]),
    .QN(_14058_)
  );
  DFF_X1 \rf[3][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00601_),
    .Q(\rf[3] [31]),
    .QN(_15012_)
  );
  DFF_X1 \rf[3][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01529_),
    .Q(\rf[3] [3]),
    .QN(_14085_)
  );
  DFF_X1 \rf[3][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01530_),
    .Q(\rf[3] [4]),
    .QN(_14084_)
  );
  DFF_X1 \rf[3][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01531_),
    .Q(\rf[3] [5]),
    .QN(_14083_)
  );
  DFF_X1 \rf[3][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01532_),
    .Q(\rf[3] [6]),
    .QN(_14082_)
  );
  DFF_X1 \rf[3][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01533_),
    .Q(\rf[3] [7]),
    .QN(_14081_)
  );
  DFF_X1 \rf[3][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01534_),
    .Q(\rf[3] [8]),
    .QN(_14080_)
  );
  DFF_X1 \rf[3][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01535_),
    .Q(\rf[3] [9]),
    .QN(_14079_)
  );
  DFF_X1 \rf[4][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00722_),
    .Q(\rf[4] [0]),
    .QN(_14891_)
  );
  DFF_X1 \rf[4][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00732_),
    .Q(\rf[4] [10]),
    .QN(_14881_)
  );
  DFF_X1 \rf[4][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00733_),
    .Q(\rf[4] [11]),
    .QN(_14880_)
  );
  DFF_X1 \rf[4][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00734_),
    .Q(\rf[4] [12]),
    .QN(_14879_)
  );
  DFF_X1 \rf[4][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00735_),
    .Q(\rf[4] [13]),
    .QN(_14878_)
  );
  DFF_X1 \rf[4][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00736_),
    .Q(\rf[4] [14]),
    .QN(_14877_)
  );
  DFF_X1 \rf[4][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00737_),
    .Q(\rf[4] [15]),
    .QN(_14876_)
  );
  DFF_X1 \rf[4][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00738_),
    .Q(\rf[4] [16]),
    .QN(_14875_)
  );
  DFF_X1 \rf[4][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00739_),
    .Q(\rf[4] [17]),
    .QN(_14874_)
  );
  DFF_X1 \rf[4][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00740_),
    .Q(\rf[4] [18]),
    .QN(_14873_)
  );
  DFF_X1 \rf[4][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00741_),
    .Q(\rf[4] [19]),
    .QN(_14872_)
  );
  DFF_X1 \rf[4][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00723_),
    .Q(\rf[4] [1]),
    .QN(_14890_)
  );
  DFF_X1 \rf[4][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00742_),
    .Q(\rf[4] [20]),
    .QN(_14871_)
  );
  DFF_X1 \rf[4][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00743_),
    .Q(\rf[4] [21]),
    .QN(_14870_)
  );
  DFF_X1 \rf[4][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00746_),
    .Q(\rf[4] [22]),
    .QN(_14867_)
  );
  DFF_X1 \rf[4][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00744_),
    .Q(\rf[4] [23]),
    .QN(_14869_)
  );
  DFF_X1 \rf[4][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00745_),
    .Q(\rf[4] [24]),
    .QN(_14868_)
  );
  DFF_X1 \rf[4][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00748_),
    .Q(\rf[4] [25]),
    .QN(_14866_)
  );
  DFF_X1 \rf[4][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00688_),
    .Q(\rf[4] [26]),
    .QN(_14925_)
  );
  DFF_X1 \rf[4][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00749_),
    .Q(\rf[4] [27]),
    .QN(_14865_)
  );
  DFF_X1 \rf[4][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00689_),
    .Q(\rf[4] [28]),
    .QN(_14924_)
  );
  DFF_X1 \rf[4][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00750_),
    .Q(\rf[4] [29]),
    .QN(_14864_)
  );
  DFF_X1 \rf[4][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00724_),
    .Q(\rf[4] [2]),
    .QN(_14889_)
  );
  DFF_X1 \rf[4][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00690_),
    .Q(\rf[4] [30]),
    .QN(_14923_)
  );
  DFF_X1 \rf[4][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00600_),
    .Q(\rf[4] [31]),
    .QN(_15013_)
  );
  DFF_X1 \rf[4][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00725_),
    .Q(\rf[4] [3]),
    .QN(_14888_)
  );
  DFF_X1 \rf[4][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00726_),
    .Q(\rf[4] [4]),
    .QN(_14887_)
  );
  DFF_X1 \rf[4][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00727_),
    .Q(\rf[4] [5]),
    .QN(_14886_)
  );
  DFF_X1 \rf[4][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00728_),
    .Q(\rf[4] [6]),
    .QN(_14885_)
  );
  DFF_X1 \rf[4][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00729_),
    .Q(\rf[4] [7]),
    .QN(_14884_)
  );
  DFF_X1 \rf[4][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00730_),
    .Q(\rf[4] [8]),
    .QN(_14883_)
  );
  DFF_X1 \rf[4][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00731_),
    .Q(\rf[4] [9]),
    .QN(_14882_)
  );
  DFF_X1 \rf[5][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01464_),
    .Q(\rf[5] [0]),
    .QN(_14150_)
  );
  DFF_X1 \rf[5][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01474_),
    .Q(\rf[5] [10]),
    .QN(_14140_)
  );
  DFF_X1 \rf[5][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01475_),
    .Q(\rf[5] [11]),
    .QN(_14139_)
  );
  DFF_X1 \rf[5][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01476_),
    .Q(\rf[5] [12]),
    .QN(_14138_)
  );
  DFF_X1 \rf[5][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01477_),
    .Q(\rf[5] [13]),
    .QN(_14137_)
  );
  DFF_X1 \rf[5][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01478_),
    .Q(\rf[5] [14]),
    .QN(_14136_)
  );
  DFF_X1 \rf[5][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01479_),
    .Q(\rf[5] [15]),
    .QN(_14135_)
  );
  DFF_X1 \rf[5][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01480_),
    .Q(\rf[5] [16]),
    .QN(_14134_)
  );
  DFF_X1 \rf[5][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01481_),
    .Q(\rf[5] [17]),
    .QN(_14133_)
  );
  DFF_X1 \rf[5][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01482_),
    .Q(\rf[5] [18]),
    .QN(_14132_)
  );
  DFF_X1 \rf[5][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01483_),
    .Q(\rf[5] [19]),
    .QN(_14131_)
  );
  DFF_X1 \rf[5][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01465_),
    .Q(\rf[5] [1]),
    .QN(_14149_)
  );
  DFF_X1 \rf[5][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01484_),
    .Q(\rf[5] [20]),
    .QN(_14130_)
  );
  DFF_X1 \rf[5][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01485_),
    .Q(\rf[5] [21]),
    .QN(_14129_)
  );
  DFF_X1 \rf[5][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01486_),
    .Q(\rf[5] [22]),
    .QN(_14128_)
  );
  DFF_X1 \rf[5][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01487_),
    .Q(\rf[5] [23]),
    .QN(_14127_)
  );
  DFF_X1 \rf[5][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01488_),
    .Q(\rf[5] [24]),
    .QN(_14126_)
  );
  DFF_X1 \rf[5][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01489_),
    .Q(\rf[5] [25]),
    .QN(_14125_)
  );
  DFF_X1 \rf[5][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01490_),
    .Q(\rf[5] [26]),
    .QN(_14124_)
  );
  DFF_X1 \rf[5][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01491_),
    .Q(\rf[5] [27]),
    .QN(_14123_)
  );
  DFF_X1 \rf[5][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01492_),
    .Q(\rf[5] [28]),
    .QN(_14122_)
  );
  DFF_X1 \rf[5][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01493_),
    .Q(\rf[5] [29]),
    .QN(_14121_)
  );
  DFF_X1 \rf[5][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01466_),
    .Q(\rf[5] [2]),
    .QN(_14148_)
  );
  DFF_X1 \rf[5][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01494_),
    .Q(\rf[5] [30]),
    .QN(_14120_)
  );
  DFF_X1 \rf[5][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00599_),
    .Q(\rf[5] [31]),
    .QN(_15014_)
  );
  DFF_X1 \rf[5][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01467_),
    .Q(\rf[5] [3]),
    .QN(_14147_)
  );
  DFF_X1 \rf[5][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01468_),
    .Q(\rf[5] [4]),
    .QN(_14146_)
  );
  DFF_X1 \rf[5][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01469_),
    .Q(\rf[5] [5]),
    .QN(_14145_)
  );
  DFF_X1 \rf[5][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01470_),
    .Q(\rf[5] [6]),
    .QN(_14144_)
  );
  DFF_X1 \rf[5][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01471_),
    .Q(\rf[5] [7]),
    .QN(_14143_)
  );
  DFF_X1 \rf[5][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01472_),
    .Q(\rf[5] [8]),
    .QN(_14142_)
  );
  DFF_X1 \rf[5][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01473_),
    .Q(\rf[5] [9]),
    .QN(_14141_)
  );
  DFF_X1 \rf[6][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00691_),
    .Q(\rf[6] [0]),
    .QN(_14922_)
  );
  DFF_X1 \rf[6][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00701_),
    .Q(\rf[6] [10]),
    .QN(_14912_)
  );
  DFF_X1 \rf[6][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00702_),
    .Q(\rf[6] [11]),
    .QN(_14911_)
  );
  DFF_X1 \rf[6][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00703_),
    .Q(\rf[6] [12]),
    .QN(_14910_)
  );
  DFF_X1 \rf[6][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00704_),
    .Q(\rf[6] [13]),
    .QN(_14909_)
  );
  DFF_X1 \rf[6][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00705_),
    .Q(\rf[6] [14]),
    .QN(_14908_)
  );
  DFF_X1 \rf[6][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00706_),
    .Q(\rf[6] [15]),
    .QN(_14907_)
  );
  DFF_X1 \rf[6][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00707_),
    .Q(\rf[6] [16]),
    .QN(_14906_)
  );
  DFF_X1 \rf[6][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00708_),
    .Q(\rf[6] [17]),
    .QN(_14905_)
  );
  DFF_X1 \rf[6][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00709_),
    .Q(\rf[6] [18]),
    .QN(_14904_)
  );
  DFF_X1 \rf[6][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00710_),
    .Q(\rf[6] [19]),
    .QN(_14903_)
  );
  DFF_X1 \rf[6][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00692_),
    .Q(\rf[6] [1]),
    .QN(_14921_)
  );
  DFF_X1 \rf[6][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00711_),
    .Q(\rf[6] [20]),
    .QN(_14902_)
  );
  DFF_X1 \rf[6][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00712_),
    .Q(\rf[6] [21]),
    .QN(_14901_)
  );
  DFF_X1 \rf[6][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00713_),
    .Q(\rf[6] [22]),
    .QN(_14900_)
  );
  DFF_X1 \rf[6][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00714_),
    .Q(\rf[6] [23]),
    .QN(_14899_)
  );
  DFF_X1 \rf[6][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00715_),
    .Q(\rf[6] [24]),
    .QN(_14898_)
  );
  DFF_X1 \rf[6][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00716_),
    .Q(\rf[6] [25]),
    .QN(_14897_)
  );
  DFF_X1 \rf[6][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00717_),
    .Q(\rf[6] [26]),
    .QN(_14896_)
  );
  DFF_X1 \rf[6][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00718_),
    .Q(\rf[6] [27]),
    .QN(_14895_)
  );
  DFF_X1 \rf[6][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00719_),
    .Q(\rf[6] [28]),
    .QN(_14894_)
  );
  DFF_X1 \rf[6][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00720_),
    .Q(\rf[6] [29]),
    .QN(_14893_)
  );
  DFF_X1 \rf[6][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00693_),
    .Q(\rf[6] [2]),
    .QN(_14920_)
  );
  DFF_X1 \rf[6][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00721_),
    .Q(\rf[6] [30]),
    .QN(_14892_)
  );
  DFF_X1 \rf[6][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00598_),
    .Q(\rf[6] [31]),
    .QN(_15015_)
  );
  DFF_X1 \rf[6][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00694_),
    .Q(\rf[6] [3]),
    .QN(_14919_)
  );
  DFF_X1 \rf[6][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00695_),
    .Q(\rf[6] [4]),
    .QN(_14918_)
  );
  DFF_X1 \rf[6][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00696_),
    .Q(\rf[6] [5]),
    .QN(_14917_)
  );
  DFF_X1 \rf[6][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00697_),
    .Q(\rf[6] [6]),
    .QN(_14916_)
  );
  DFF_X1 \rf[6][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00698_),
    .Q(\rf[6] [7]),
    .QN(_14915_)
  );
  DFF_X1 \rf[6][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00699_),
    .Q(\rf[6] [8]),
    .QN(_14914_)
  );
  DFF_X1 \rf[6][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00700_),
    .Q(\rf[6] [9]),
    .QN(_14913_)
  );
  DFF_X1 \rf[7][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01495_),
    .Q(\rf[7] [0]),
    .QN(_14119_)
  );
  DFF_X1 \rf[7][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01505_),
    .Q(\rf[7] [10]),
    .QN(_14109_)
  );
  DFF_X1 \rf[7][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01506_),
    .Q(\rf[7] [11]),
    .QN(_14108_)
  );
  DFF_X1 \rf[7][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01507_),
    .Q(\rf[7] [12]),
    .QN(_14107_)
  );
  DFF_X1 \rf[7][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01508_),
    .Q(\rf[7] [13]),
    .QN(_14106_)
  );
  DFF_X1 \rf[7][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01509_),
    .Q(\rf[7] [14]),
    .QN(_14105_)
  );
  DFF_X1 \rf[7][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01510_),
    .Q(\rf[7] [15]),
    .QN(_14104_)
  );
  DFF_X1 \rf[7][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01511_),
    .Q(\rf[7] [16]),
    .QN(_14103_)
  );
  DFF_X1 \rf[7][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01512_),
    .Q(\rf[7] [17]),
    .QN(_14102_)
  );
  DFF_X1 \rf[7][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01513_),
    .Q(\rf[7] [18]),
    .QN(_14101_)
  );
  DFF_X1 \rf[7][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01514_),
    .Q(\rf[7] [19]),
    .QN(_14100_)
  );
  DFF_X1 \rf[7][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01496_),
    .Q(\rf[7] [1]),
    .QN(_14118_)
  );
  DFF_X1 \rf[7][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01515_),
    .Q(\rf[7] [20]),
    .QN(_14099_)
  );
  DFF_X1 \rf[7][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01516_),
    .Q(\rf[7] [21]),
    .QN(_14098_)
  );
  DFF_X1 \rf[7][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01517_),
    .Q(\rf[7] [22]),
    .QN(_14097_)
  );
  DFF_X1 \rf[7][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01518_),
    .Q(\rf[7] [23]),
    .QN(_14096_)
  );
  DFF_X1 \rf[7][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01519_),
    .Q(\rf[7] [24]),
    .QN(_14095_)
  );
  DFF_X1 \rf[7][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01520_),
    .Q(\rf[7] [25]),
    .QN(_14094_)
  );
  DFF_X1 \rf[7][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01521_),
    .Q(\rf[7] [26]),
    .QN(_14093_)
  );
  DFF_X1 \rf[7][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01522_),
    .Q(\rf[7] [27]),
    .QN(_14092_)
  );
  DFF_X1 \rf[7][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01523_),
    .Q(\rf[7] [28]),
    .QN(_14091_)
  );
  DFF_X1 \rf[7][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01524_),
    .Q(\rf[7] [29]),
    .QN(_14090_)
  );
  DFF_X1 \rf[7][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01497_),
    .Q(\rf[7] [2]),
    .QN(_14117_)
  );
  DFF_X1 \rf[7][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01525_),
    .Q(\rf[7] [30]),
    .QN(_14089_)
  );
  DFF_X1 \rf[7][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00597_),
    .Q(\rf[7] [31]),
    .QN(_15016_)
  );
  DFF_X1 \rf[7][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01498_),
    .Q(\rf[7] [3]),
    .QN(_14116_)
  );
  DFF_X1 \rf[7][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01499_),
    .Q(\rf[7] [4]),
    .QN(_14115_)
  );
  DFF_X1 \rf[7][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01500_),
    .Q(\rf[7] [5]),
    .QN(_14114_)
  );
  DFF_X1 \rf[7][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01501_),
    .Q(\rf[7] [6]),
    .QN(_14113_)
  );
  DFF_X1 \rf[7][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01502_),
    .Q(\rf[7] [7]),
    .QN(_14112_)
  );
  DFF_X1 \rf[7][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01503_),
    .Q(\rf[7] [8]),
    .QN(_14111_)
  );
  DFF_X1 \rf[7][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01504_),
    .Q(\rf[7] [9]),
    .QN(_14110_)
  );
  DFF_X1 \rf[8][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00813_),
    .Q(\rf[8] [0]),
    .QN(_14801_)
  );
  DFF_X1 \rf[8][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00823_),
    .Q(\rf[8] [10]),
    .QN(_14791_)
  );
  DFF_X1 \rf[8][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00824_),
    .Q(\rf[8] [11]),
    .QN(_14790_)
  );
  DFF_X1 \rf[8][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00825_),
    .Q(\rf[8] [12]),
    .QN(_14789_)
  );
  DFF_X1 \rf[8][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00826_),
    .Q(\rf[8] [13]),
    .QN(_14788_)
  );
  DFF_X1 \rf[8][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00827_),
    .Q(\rf[8] [14]),
    .QN(_14787_)
  );
  DFF_X1 \rf[8][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00828_),
    .Q(\rf[8] [15]),
    .QN(_14786_)
  );
  DFF_X1 \rf[8][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00829_),
    .Q(\rf[8] [16]),
    .QN(_14785_)
  );
  DFF_X1 \rf[8][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00830_),
    .Q(\rf[8] [17]),
    .QN(_14784_)
  );
  DFF_X1 \rf[8][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00831_),
    .Q(\rf[8] [18]),
    .QN(_14783_)
  );
  DFF_X1 \rf[8][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00832_),
    .Q(\rf[8] [19]),
    .QN(_14782_)
  );
  DFF_X1 \rf[8][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00814_),
    .Q(\rf[8] [1]),
    .QN(_14800_)
  );
  DFF_X1 \rf[8][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00833_),
    .Q(\rf[8] [20]),
    .QN(_14781_)
  );
  DFF_X1 \rf[8][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00834_),
    .Q(\rf[8] [21]),
    .QN(_14780_)
  );
  DFF_X1 \rf[8][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00835_),
    .Q(\rf[8] [22]),
    .QN(_14779_)
  );
  DFF_X1 \rf[8][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00836_),
    .Q(\rf[8] [23]),
    .QN(_14778_)
  );
  DFF_X1 \rf[8][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00837_),
    .Q(\rf[8] [24]),
    .QN(_14777_)
  );
  DFF_X1 \rf[8][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00838_),
    .Q(\rf[8] [25]),
    .QN(_14776_)
  );
  DFF_X1 \rf[8][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00839_),
    .Q(\rf[8] [26]),
    .QN(_14775_)
  );
  DFF_X1 \rf[8][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00840_),
    .Q(\rf[8] [27]),
    .QN(_14774_)
  );
  DFF_X1 \rf[8][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00841_),
    .Q(\rf[8] [28]),
    .QN(_14773_)
  );
  DFF_X1 \rf[8][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00842_),
    .Q(\rf[8] [29]),
    .QN(_14772_)
  );
  DFF_X1 \rf[8][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00815_),
    .Q(\rf[8] [2]),
    .QN(_14799_)
  );
  DFF_X1 \rf[8][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00843_),
    .Q(\rf[8] [30]),
    .QN(_14771_)
  );
  DFF_X1 \rf[8][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00596_),
    .Q(\rf[8] [31]),
    .QN(_15017_)
  );
  DFF_X1 \rf[8][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00816_),
    .Q(\rf[8] [3]),
    .QN(_14798_)
  );
  DFF_X1 \rf[8][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00817_),
    .Q(\rf[8] [4]),
    .QN(_14797_)
  );
  DFF_X1 \rf[8][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00818_),
    .Q(\rf[8] [5]),
    .QN(_14796_)
  );
  DFF_X1 \rf[8][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00819_),
    .Q(\rf[8] [6]),
    .QN(_14795_)
  );
  DFF_X1 \rf[8][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00820_),
    .Q(\rf[8] [7]),
    .QN(_14794_)
  );
  DFF_X1 \rf[8][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00821_),
    .Q(\rf[8] [8]),
    .QN(_14793_)
  );
  DFF_X1 \rf[8][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00822_),
    .Q(\rf[8] [9]),
    .QN(_14792_)
  );
  DFF_X1 \rf[9][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01092_),
    .Q(\rf[9] [0]),
    .QN(_14522_)
  );
  DFF_X1 \rf[9][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01102_),
    .Q(\rf[9] [10]),
    .QN(_14512_)
  );
  DFF_X1 \rf[9][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01103_),
    .Q(\rf[9] [11]),
    .QN(_14511_)
  );
  DFF_X1 \rf[9][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01104_),
    .Q(\rf[9] [12]),
    .QN(_14510_)
  );
  DFF_X1 \rf[9][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01105_),
    .Q(\rf[9] [13]),
    .QN(_14509_)
  );
  DFF_X1 \rf[9][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01106_),
    .Q(\rf[9] [14]),
    .QN(_14508_)
  );
  DFF_X1 \rf[9][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01107_),
    .Q(\rf[9] [15]),
    .QN(_14507_)
  );
  DFF_X1 \rf[9][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01108_),
    .Q(\rf[9] [16]),
    .QN(_14506_)
  );
  DFF_X1 \rf[9][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01109_),
    .Q(\rf[9] [17]),
    .QN(_14505_)
  );
  DFF_X1 \rf[9][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01110_),
    .Q(\rf[9] [18]),
    .QN(_14504_)
  );
  DFF_X1 \rf[9][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01111_),
    .Q(\rf[9] [19]),
    .QN(_14503_)
  );
  DFF_X1 \rf[9][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01093_),
    .Q(\rf[9] [1]),
    .QN(_14521_)
  );
  DFF_X1 \rf[9][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01112_),
    .Q(\rf[9] [20]),
    .QN(_14502_)
  );
  DFF_X1 \rf[9][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01113_),
    .Q(\rf[9] [21]),
    .QN(_14501_)
  );
  DFF_X1 \rf[9][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01114_),
    .Q(\rf[9] [22]),
    .QN(_14500_)
  );
  DFF_X1 \rf[9][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01115_),
    .Q(\rf[9] [23]),
    .QN(_14499_)
  );
  DFF_X1 \rf[9][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01116_),
    .Q(\rf[9] [24]),
    .QN(_14498_)
  );
  DFF_X1 \rf[9][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01117_),
    .Q(\rf[9] [25]),
    .QN(_14497_)
  );
  DFF_X1 \rf[9][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01118_),
    .Q(\rf[9] [26]),
    .QN(_14496_)
  );
  DFF_X1 \rf[9][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01119_),
    .Q(\rf[9] [27]),
    .QN(_14495_)
  );
  DFF_X1 \rf[9][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01120_),
    .Q(\rf[9] [28]),
    .QN(_14494_)
  );
  DFF_X1 \rf[9][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01121_),
    .Q(\rf[9] [29]),
    .QN(_14493_)
  );
  DFF_X1 \rf[9][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01094_),
    .Q(\rf[9] [2]),
    .QN(_14520_)
  );
  DFF_X1 \rf[9][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01122_),
    .Q(\rf[9] [30]),
    .QN(_14492_)
  );
  DFF_X1 \rf[9][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00595_),
    .Q(\rf[9] [31]),
    .QN(_15018_)
  );
  DFF_X1 \rf[9][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01095_),
    .Q(\rf[9] [3]),
    .QN(_14519_)
  );
  DFF_X1 \rf[9][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01096_),
    .Q(\rf[9] [4]),
    .QN(_14518_)
  );
  DFF_X1 \rf[9][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01097_),
    .Q(\rf[9] [5]),
    .QN(_14517_)
  );
  DFF_X1 \rf[9][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01098_),
    .Q(\rf[9] [6]),
    .QN(_14516_)
  );
  DFF_X1 \rf[9][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01099_),
    .Q(\rf[9] [7]),
    .QN(_14515_)
  );
  DFF_X1 \rf[9][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01100_),
    .Q(\rf[9] [8]),
    .QN(_14514_)
  );
  DFF_X1 \rf[9][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01101_),
    .Q(\rf[9] [9]),
    .QN(_14513_)
  );
  DFF_X1 \wb_ctrl_csr[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00520_),
    .Q(wb_ctrl_csr[0]),
    .QN(_15076_)
  );
  DFF_X1 \wb_ctrl_csr[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00521_),
    .Q(wb_ctrl_csr[1]),
    .QN(_15075_)
  );
  DFF_X1 \wb_ctrl_csr[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00522_),
    .Q(wb_ctrl_csr[2]),
    .QN(_15074_)
  );
  DFF_X1 \wb_ctrl_div$_DFFE_PP_  (
    .CK(clock),
    .D(_00524_),
    .Q(wb_ctrl_div),
    .QN(_15072_)
  );
  DFF_X1 \wb_ctrl_fence_i$_DFFE_PP_  (
    .CK(clock),
    .D(_00519_),
    .Q(wb_ctrl_fence_i),
    .QN(_15077_)
  );
  DFF_X1 \wb_ctrl_mem$_DFFE_PP_  (
    .CK(clock),
    .D(_00525_),
    .Q(wb_ctrl_mem),
    .QN(_15071_)
  );
  DFF_X1 \wb_ctrl_wxd$_DFFE_PP_  (
    .CK(clock),
    .D(_00523_),
    .Q(wb_ctrl_wxd),
    .QN(_15073_)
  );
  DFF_X1 \wb_reg_cause[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00591_),
    .Q(wb_reg_cause[0]),
    .QN(_00016_)
  );
  DFF_X1 \wb_reg_cause[10]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00186_),
    .Q(wb_reg_cause[10]),
    .QN(_15406_)
  );
  DFF_X1 \wb_reg_cause[11]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00187_),
    .Q(wb_reg_cause[11]),
    .QN(_15405_)
  );
  DFF_X1 \wb_reg_cause[12]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00188_),
    .Q(wb_reg_cause[12]),
    .QN(_15404_)
  );
  DFF_X1 \wb_reg_cause[13]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00189_),
    .Q(wb_reg_cause[13]),
    .QN(_15403_)
  );
  DFF_X1 \wb_reg_cause[14]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00190_),
    .Q(wb_reg_cause[14]),
    .QN(_15402_)
  );
  DFF_X1 \wb_reg_cause[15]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00191_),
    .Q(wb_reg_cause[15]),
    .QN(_15401_)
  );
  DFF_X1 \wb_reg_cause[16]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00192_),
    .Q(wb_reg_cause[16]),
    .QN(_15400_)
  );
  DFF_X1 \wb_reg_cause[17]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00193_),
    .Q(wb_reg_cause[17]),
    .QN(_15399_)
  );
  DFF_X1 \wb_reg_cause[18]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00194_),
    .Q(wb_reg_cause[18]),
    .QN(_15398_)
  );
  DFF_X1 \wb_reg_cause[19]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00195_),
    .Q(wb_reg_cause[19]),
    .QN(_15397_)
  );
  DFF_X1 \wb_reg_cause[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00592_),
    .Q(wb_reg_cause[1]),
    .QN(_00015_)
  );
  DFF_X1 \wb_reg_cause[20]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00196_),
    .Q(wb_reg_cause[20]),
    .QN(_15396_)
  );
  DFF_X1 \wb_reg_cause[21]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00197_),
    .Q(wb_reg_cause[21]),
    .QN(_15395_)
  );
  DFF_X1 \wb_reg_cause[22]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00198_),
    .Q(wb_reg_cause[22]),
    .QN(_15394_)
  );
  DFF_X1 \wb_reg_cause[23]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00199_),
    .Q(wb_reg_cause[23]),
    .QN(_15393_)
  );
  DFF_X1 \wb_reg_cause[24]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00200_),
    .Q(wb_reg_cause[24]),
    .QN(_15392_)
  );
  DFF_X1 \wb_reg_cause[25]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00201_),
    .Q(wb_reg_cause[25]),
    .QN(_15391_)
  );
  DFF_X1 \wb_reg_cause[26]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00202_),
    .Q(wb_reg_cause[26]),
    .QN(_15390_)
  );
  DFF_X1 \wb_reg_cause[27]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00203_),
    .Q(wb_reg_cause[27]),
    .QN(_15389_)
  );
  DFF_X1 \wb_reg_cause[28]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00204_),
    .Q(wb_reg_cause[28]),
    .QN(_15388_)
  );
  DFF_X1 \wb_reg_cause[29]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00205_),
    .Q(wb_reg_cause[29]),
    .QN(_15387_)
  );
  DFF_X1 \wb_reg_cause[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00593_),
    .Q(wb_reg_cause[2]),
    .QN(_00014_)
  );
  DFF_X1 \wb_reg_cause[30]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00206_),
    .Q(wb_reg_cause[30]),
    .QN(_15386_)
  );
  DFF_X1 \wb_reg_cause[31]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00207_),
    .Q(wb_reg_cause[31]),
    .QN(_15554_)
  );
  DFF_X1 \wb_reg_cause[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00594_),
    .Q(wb_reg_cause[3]),
    .QN(_00013_)
  );
  DFF_X1 \wb_reg_cause[4]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00180_),
    .Q(wb_reg_cause[4]),
    .QN(_00030_)
  );
  DFF_X1 \wb_reg_cause[5]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00181_),
    .Q(wb_reg_cause[5]),
    .QN(_15411_)
  );
  DFF_X1 \wb_reg_cause[6]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00182_),
    .Q(wb_reg_cause[6]),
    .QN(_15410_)
  );
  DFF_X1 \wb_reg_cause[7]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00183_),
    .Q(wb_reg_cause[7]),
    .QN(_15409_)
  );
  DFF_X1 \wb_reg_cause[8]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00184_),
    .Q(wb_reg_cause[8]),
    .QN(_15408_)
  );
  DFF_X1 \wb_reg_cause[9]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00185_),
    .Q(wb_reg_cause[9]),
    .QN(_15407_)
  );
  DFF_X1 \wb_reg_flush_pipe$_DFF_P_  (
    .CK(clock),
    .D(_00009_),
    .Q(wb_reg_flush_pipe),
    .QN(_15555_)
  );
  DFF_X1 \wb_reg_inst[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00529_),
    .Q(wb_reg_inst[10]),
    .QN(_15068_)
  );
  DFF_X1 \wb_reg_inst[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00530_),
    .Q(wb_reg_inst[11]),
    .QN(_15067_)
  );
  DFF_X1 \wb_reg_inst[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00531_),
    .Q(wb_reg_inst[16]),
    .QN(_15066_)
  );
  DFF_X1 \wb_reg_inst[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00532_),
    .Q(wb_reg_inst[17]),
    .QN(_15065_)
  );
  DFF_X1 \wb_reg_inst[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00533_),
    .Q(wb_reg_inst[18]),
    .QN(_15064_)
  );
  DFF_X1 \wb_reg_inst[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00534_),
    .Q(wb_reg_inst[19]),
    .QN(_15063_)
  );
  DFF_X1 \wb_reg_inst[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00535_),
    .Q(wb_reg_inst[20]),
    .QN(_15062_)
  );
  DFF_X1 \wb_reg_inst[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00536_),
    .Q(wb_reg_inst[21]),
    .QN(_15061_)
  );
  DFF_X1 \wb_reg_inst[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00537_),
    .Q(wb_reg_inst[22]),
    .QN(_15060_)
  );
  DFF_X1 \wb_reg_inst[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00538_),
    .Q(wb_reg_inst[23]),
    .QN(_15059_)
  );
  DFF_X1 \wb_reg_inst[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00539_),
    .Q(wb_reg_inst[24]),
    .QN(_15058_)
  );
  DFF_X1 \wb_reg_inst[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00540_),
    .Q(wb_reg_inst[25]),
    .QN(_15057_)
  );
  DFF_X1 \wb_reg_inst[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00541_),
    .Q(wb_reg_inst[26]),
    .QN(_15056_)
  );
  DFF_X1 \wb_reg_inst[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00542_),
    .Q(wb_reg_inst[27]),
    .QN(_15055_)
  );
  DFF_X1 \wb_reg_inst[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00543_),
    .Q(wb_reg_inst[28]),
    .QN(_15054_)
  );
  DFF_X1 \wb_reg_inst[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00544_),
    .Q(wb_reg_inst[29]),
    .QN(_15053_)
  );
  DFF_X1 \wb_reg_inst[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00545_),
    .Q(wb_reg_inst[30]),
    .QN(_15052_)
  );
  DFF_X1 \wb_reg_inst[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00546_),
    .Q(wb_reg_inst[31]),
    .QN(_15051_)
  );
  DFF_X1 \wb_reg_inst[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00526_),
    .Q(wb_reg_inst[7]),
    .QN(_00029_)
  );
  DFF_X1 \wb_reg_inst[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00527_),
    .Q(wb_reg_inst[8]),
    .QN(_15070_)
  );
  DFF_X1 \wb_reg_inst[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00528_),
    .Q(wb_reg_inst[9]),
    .QN(_15069_)
  );
  DFF_X1 \wb_reg_pc[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00208_),
    .Q(wb_reg_pc[0]),
    .QN(_15384_)
  );
  DFF_X1 \wb_reg_pc[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00218_),
    .Q(wb_reg_pc[10]),
    .QN(_15374_)
  );
  DFF_X1 \wb_reg_pc[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00219_),
    .Q(wb_reg_pc[11]),
    .QN(_15373_)
  );
  DFF_X1 \wb_reg_pc[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00220_),
    .Q(wb_reg_pc[12]),
    .QN(_15372_)
  );
  DFF_X1 \wb_reg_pc[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00221_),
    .Q(wb_reg_pc[13]),
    .QN(_15371_)
  );
  DFF_X1 \wb_reg_pc[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00222_),
    .Q(wb_reg_pc[14]),
    .QN(_15370_)
  );
  DFF_X1 \wb_reg_pc[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00223_),
    .Q(wb_reg_pc[15]),
    .QN(_15369_)
  );
  DFF_X1 \wb_reg_pc[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00224_),
    .Q(wb_reg_pc[16]),
    .QN(_15368_)
  );
  DFF_X1 \wb_reg_pc[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00225_),
    .Q(wb_reg_pc[17]),
    .QN(_15367_)
  );
  DFF_X1 \wb_reg_pc[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00226_),
    .Q(wb_reg_pc[18]),
    .QN(_15366_)
  );
  DFF_X1 \wb_reg_pc[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00227_),
    .Q(wb_reg_pc[19]),
    .QN(_15365_)
  );
  DFF_X1 \wb_reg_pc[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00209_),
    .Q(wb_reg_pc[1]),
    .QN(_15383_)
  );
  DFF_X1 \wb_reg_pc[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00228_),
    .Q(wb_reg_pc[20]),
    .QN(_15364_)
  );
  DFF_X1 \wb_reg_pc[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00229_),
    .Q(wb_reg_pc[21]),
    .QN(_15363_)
  );
  DFF_X1 \wb_reg_pc[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00230_),
    .Q(wb_reg_pc[22]),
    .QN(_15362_)
  );
  DFF_X1 \wb_reg_pc[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00231_),
    .Q(wb_reg_pc[23]),
    .QN(_15361_)
  );
  DFF_X1 \wb_reg_pc[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00232_),
    .Q(wb_reg_pc[24]),
    .QN(_15360_)
  );
  DFF_X1 \wb_reg_pc[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00233_),
    .Q(wb_reg_pc[25]),
    .QN(_15359_)
  );
  DFF_X1 \wb_reg_pc[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00234_),
    .Q(wb_reg_pc[26]),
    .QN(_15358_)
  );
  DFF_X1 \wb_reg_pc[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00235_),
    .Q(wb_reg_pc[27]),
    .QN(_15357_)
  );
  DFF_X1 \wb_reg_pc[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00236_),
    .Q(wb_reg_pc[28]),
    .QN(_15356_)
  );
  DFF_X1 \wb_reg_pc[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00237_),
    .Q(wb_reg_pc[29]),
    .QN(_15355_)
  );
  DFF_X1 \wb_reg_pc[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00210_),
    .Q(wb_reg_pc[2]),
    .QN(_15382_)
  );
  DFF_X1 \wb_reg_pc[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00238_),
    .Q(wb_reg_pc[30]),
    .QN(_15354_)
  );
  DFF_X1 \wb_reg_pc[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00239_),
    .Q(wb_reg_pc[31]),
    .QN(_15353_)
  );
  DFF_X1 \wb_reg_pc[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00211_),
    .Q(wb_reg_pc[3]),
    .QN(_15381_)
  );
  DFF_X1 \wb_reg_pc[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00212_),
    .Q(wb_reg_pc[4]),
    .QN(_15380_)
  );
  DFF_X1 \wb_reg_pc[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00213_),
    .Q(wb_reg_pc[5]),
    .QN(_15379_)
  );
  DFF_X1 \wb_reg_pc[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00214_),
    .Q(wb_reg_pc[6]),
    .QN(_15378_)
  );
  DFF_X1 \wb_reg_pc[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00215_),
    .Q(wb_reg_pc[7]),
    .QN(_15377_)
  );
  DFF_X1 \wb_reg_pc[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00216_),
    .Q(wb_reg_pc[8]),
    .QN(_15376_)
  );
  DFF_X1 \wb_reg_pc[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00217_),
    .Q(wb_reg_pc[9]),
    .QN(_15375_)
  );
  DFF_X1 \wb_reg_raw_inst[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00101_),
    .Q(wb_reg_raw_inst[0]),
    .QN(_15489_)
  );
  DFF_X1 \wb_reg_raw_inst[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00111_),
    .Q(wb_reg_raw_inst[10]),
    .QN(_15479_)
  );
  DFF_X1 \wb_reg_raw_inst[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00112_),
    .Q(wb_reg_raw_inst[11]),
    .QN(_15478_)
  );
  DFF_X1 \wb_reg_raw_inst[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00113_),
    .Q(wb_reg_raw_inst[12]),
    .QN(_15477_)
  );
  DFF_X1 \wb_reg_raw_inst[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00114_),
    .Q(wb_reg_raw_inst[13]),
    .QN(_15476_)
  );
  DFF_X1 \wb_reg_raw_inst[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00115_),
    .Q(wb_reg_raw_inst[14]),
    .QN(_15475_)
  );
  DFF_X1 \wb_reg_raw_inst[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00116_),
    .Q(wb_reg_raw_inst[15]),
    .QN(_15474_)
  );
  DFF_X1 \wb_reg_raw_inst[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00102_),
    .Q(wb_reg_raw_inst[1]),
    .QN(_15488_)
  );
  DFF_X1 \wb_reg_raw_inst[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00103_),
    .Q(wb_reg_raw_inst[2]),
    .QN(_15487_)
  );
  DFF_X1 \wb_reg_raw_inst[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00104_),
    .Q(wb_reg_raw_inst[3]),
    .QN(_15486_)
  );
  DFF_X1 \wb_reg_raw_inst[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00105_),
    .Q(wb_reg_raw_inst[4]),
    .QN(_15485_)
  );
  DFF_X1 \wb_reg_raw_inst[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00106_),
    .Q(wb_reg_raw_inst[5]),
    .QN(_15484_)
  );
  DFF_X1 \wb_reg_raw_inst[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00107_),
    .Q(wb_reg_raw_inst[6]),
    .QN(_15483_)
  );
  DFF_X1 \wb_reg_raw_inst[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00108_),
    .Q(wb_reg_raw_inst[7]),
    .QN(_15482_)
  );
  DFF_X1 \wb_reg_raw_inst[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00109_),
    .Q(wb_reg_raw_inst[8]),
    .QN(_15481_)
  );
  DFF_X1 \wb_reg_raw_inst[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00110_),
    .Q(wb_reg_raw_inst[9]),
    .QN(_15480_)
  );
  DFF_X1 \wb_reg_replay$_DFF_P_  (
    .CK(clock),
    .D(_00010_),
    .Q(wb_reg_replay),
    .QN(_15556_)
  );
  DFF_X1 \wb_reg_valid$_DFF_P_  (
    .CK(clock),
    .D(_wb_reg_valid_T),
    .Q(wb_reg_valid),
    .QN(_15385_)
  );
  DFF_X1 \wb_reg_wdata[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00117_),
    .Q(wb_reg_wdata[0]),
    .QN(_15473_)
  );
  DFF_X1 \wb_reg_wdata[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00127_),
    .Q(wb_reg_wdata[10]),
    .QN(_15463_)
  );
  DFF_X1 \wb_reg_wdata[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00128_),
    .Q(wb_reg_wdata[11]),
    .QN(_15462_)
  );
  DFF_X1 \wb_reg_wdata[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00129_),
    .Q(wb_reg_wdata[12]),
    .QN(_15461_)
  );
  DFF_X1 \wb_reg_wdata[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00130_),
    .Q(wb_reg_wdata[13]),
    .QN(_15460_)
  );
  DFF_X1 \wb_reg_wdata[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00131_),
    .Q(wb_reg_wdata[14]),
    .QN(_15459_)
  );
  DFF_X1 \wb_reg_wdata[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00132_),
    .Q(wb_reg_wdata[15]),
    .QN(_15458_)
  );
  DFF_X1 \wb_reg_wdata[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00133_),
    .Q(wb_reg_wdata[16]),
    .QN(_15457_)
  );
  DFF_X1 \wb_reg_wdata[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00134_),
    .Q(wb_reg_wdata[17]),
    .QN(_15456_)
  );
  DFF_X1 \wb_reg_wdata[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00135_),
    .Q(wb_reg_wdata[18]),
    .QN(_15455_)
  );
  DFF_X1 \wb_reg_wdata[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00136_),
    .Q(wb_reg_wdata[19]),
    .QN(_15454_)
  );
  DFF_X1 \wb_reg_wdata[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00118_),
    .Q(wb_reg_wdata[1]),
    .QN(_15472_)
  );
  DFF_X1 \wb_reg_wdata[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00137_),
    .Q(wb_reg_wdata[20]),
    .QN(_15453_)
  );
  DFF_X1 \wb_reg_wdata[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00138_),
    .Q(wb_reg_wdata[21]),
    .QN(_15452_)
  );
  DFF_X1 \wb_reg_wdata[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00139_),
    .Q(wb_reg_wdata[22]),
    .QN(_15451_)
  );
  DFF_X1 \wb_reg_wdata[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00140_),
    .Q(wb_reg_wdata[23]),
    .QN(_15450_)
  );
  DFF_X1 \wb_reg_wdata[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00141_),
    .Q(wb_reg_wdata[24]),
    .QN(_15449_)
  );
  DFF_X1 \wb_reg_wdata[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00142_),
    .Q(wb_reg_wdata[25]),
    .QN(_15448_)
  );
  DFF_X1 \wb_reg_wdata[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00143_),
    .Q(wb_reg_wdata[26]),
    .QN(_15447_)
  );
  DFF_X1 \wb_reg_wdata[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00144_),
    .Q(wb_reg_wdata[27]),
    .QN(_15446_)
  );
  DFF_X1 \wb_reg_wdata[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00145_),
    .Q(wb_reg_wdata[28]),
    .QN(_15445_)
  );
  DFF_X1 \wb_reg_wdata[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00146_),
    .Q(wb_reg_wdata[29]),
    .QN(_15444_)
  );
  DFF_X1 \wb_reg_wdata[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00119_),
    .Q(wb_reg_wdata[2]),
    .QN(_15471_)
  );
  DFF_X1 \wb_reg_wdata[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00147_),
    .Q(wb_reg_wdata[30]),
    .QN(_15443_)
  );
  DFF_X1 \wb_reg_wdata[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00148_),
    .Q(wb_reg_wdata[31]),
    .QN(_15442_)
  );
  DFF_X1 \wb_reg_wdata[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00120_),
    .Q(wb_reg_wdata[3]),
    .QN(_15470_)
  );
  DFF_X1 \wb_reg_wdata[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00121_),
    .Q(wb_reg_wdata[4]),
    .QN(_15469_)
  );
  DFF_X1 \wb_reg_wdata[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00122_),
    .Q(wb_reg_wdata[5]),
    .QN(_15468_)
  );
  DFF_X1 \wb_reg_wdata[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00123_),
    .Q(wb_reg_wdata[6]),
    .QN(_15467_)
  );
  DFF_X1 \wb_reg_wdata[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00124_),
    .Q(wb_reg_wdata[7]),
    .QN(_15466_)
  );
  DFF_X1 \wb_reg_wdata[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00125_),
    .Q(wb_reg_wdata[8]),
    .QN(_15465_)
  );
  DFF_X1 \wb_reg_wdata[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00126_),
    .Q(wb_reg_wdata[9]),
    .QN(_15464_)
  );
  DFF_X1 \wb_reg_xcpt$_DFF_P_  (
    .CK(clock),
    .D(_00011_),
    .Q(wb_reg_xcpt),
    .QN(tval_dmem_addr)
  );
  assign _15563_[1] = ex_reg_mem_size[1];
  assign _15564_[0] = ex_reg_mem_size[0];
  assign PlusArgTimeout_clock = clock;
  assign PlusArgTimeout_io_count = csr_io_time;
  assign PlusArgTimeout_reset = reset;
  assign { _T_11[4:2], _T_11[0] } = { 3'h0, ibuf_io_inst_0_bits_xcpt1_ae_inst };
  assign { _T_113[2], _T_113[0] } = 2'h2;
  assign _T_114[2] = 1'h1;
  assign _T_115[2] = 1'h1;
  assign _T_116 = { 3'h1, _T_115[1:0] };
  assign { _T_118[4], _T_118[2] } = 2'h1;
  assign { _T_119[4], _T_119[2] } = 2'h1;
  assign _T_12[4:2] = { ibuf_io_inst_0_bits_xcpt1_gf_inst, 1'h0, ibuf_io_inst_0_bits_xcpt1_gf_inst };
  assign _T_13[3] = ibuf_io_inst_0_bits_xcpt1_pf_inst;
  assign _T_143[0] = 1'h0;
  assign _T_35 = { ibuf_io_inst_0_bits_xcpt1_pf_inst, ibuf_io_inst_0_bits_xcpt1_gf_inst, ibuf_io_inst_0_bits_xcpt1_ae_inst };
  assign _T_37 = { 2'h0, ibuf_io_inst_0_bits_xcpt0_ae_inst };
  assign _T_40 = 1'h0;
  assign _T_41 = 1'h0;
  assign _T_42 = 1'h0;
  assign _T_74[2] = _T_74[3];
  assign _T_93 = _T_118[3];
  assign _bypass_src_T[1] = 1'h1;
  assign _bypass_src_T_2[1] = 1'h1;
  assign _csr_io_rw_cmd_T[1:0] = 2'h0;
  assign _csr_io_rw_cmd_T_1 = { wb_reg_valid, 2'h3 };
  assign _ctrl_stalld_T_15 = 1'h0;
  assign _ex_imm_b11_T_5 = ex_reg_inst[20];
  assign _ex_imm_b11_T_8 = ex_reg_inst[7];
  assign _ex_imm_b19_12_T_4 = ex_reg_inst[19:12];
  assign _ex_imm_b30_20_T_2 = ex_reg_inst[30:20];
  assign _ex_imm_sign_T_2 = ex_reg_inst[31];
  assign { _ex_op2_T_1[3], _ex_op2_T_1[1:0] } = { 1'h0, ex_reg_rvc, 1'h0 };
  assign _ex_rs_T_13 = { ex_reg_rs_msb_1, ex_reg_rs_lsb_1 };
  assign _ex_rs_T_6 = { ex_reg_rs_msb_0, ex_reg_rs_lsb_0 };
  assign _id_ctrl_decoder_decoded_T[7:6] = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1] };
  assign _id_ctrl_decoder_decoded_T_10[8:1] = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], csr_io_decode_0_inst[3], _id_ctrl_decoder_decoded_T[3:0] };
  assign _id_ctrl_decoder_decoded_T_100 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:3], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], csr_io_decode_0_inst[13], csr_io_decode_0_inst[14] };
  assign _id_ctrl_decoder_decoded_T_102 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], csr_io_decode_0_inst[13], csr_io_decode_0_inst[14] };
  assign _id_ctrl_decoder_decoded_T_104 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], _id_ctrl_decoder_decoded_T[2:1], csr_io_decode_0_inst[12], csr_io_decode_0_inst[13], csr_io_decode_0_inst[14] };
  assign _id_ctrl_decoder_decoded_T_106[13:6] = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[25] };
  assign _id_ctrl_decoder_decoded_T_108 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[12], csr_io_decode_0_inst[25], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign _id_ctrl_decoder_decoded_T_110 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[13], csr_io_decode_0_inst[25], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign { _id_ctrl_decoder_decoded_T_112[13:7], _id_ctrl_decoder_decoded_T_112[5:0] } = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], csr_io_decode_0_inst[3], _id_ctrl_decoder_decoded_T[3], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0], csr_io_decode_0_inst[27], _id_ctrl_decoder_decoded_T_106[2:0] };
  assign { _id_ctrl_decoder_decoded_T_114[16:10], _id_ctrl_decoder_decoded_T_114[4:0] } = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], csr_io_decode_0_inst[3], _id_ctrl_decoder_decoded_T[3], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T_106[4], csr_io_decode_0_inst[28], _id_ctrl_decoder_decoded_T_106[2:0] };
  assign _id_ctrl_decoder_decoded_T_116 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], csr_io_decode_0_inst[3], _id_ctrl_decoder_decoded_T[3], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T_112[6], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_114[9:5], _id_ctrl_decoder_decoded_T_106[4], csr_io_decode_0_inst[28], _id_ctrl_decoder_decoded_T_106[2:0] };
  assign { _id_ctrl_decoder_decoded_T_118[27:24], _id_ctrl_decoder_decoded_T_118[18:16], _id_ctrl_decoder_decoded_T_118[10:6], _id_ctrl_decoder_decoded_T_118[4:0] } = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0], csr_io_decode_0_inst[20], _id_ctrl_decoder_decoded_T_114[8], csr_io_decode_0_inst[22], _id_ctrl_decoder_decoded_T_114[6:5], _id_ctrl_decoder_decoded_T_106[5:4], csr_io_decode_0_inst[28], _id_ctrl_decoder_decoded_T_106[1:0] };
  assign _id_ctrl_decoder_decoded_T_12 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], _id_ctrl_decoder_decoded_T[4], csr_io_decode_0_inst[4], _id_ctrl_decoder_decoded_T[1] };
  assign _id_ctrl_decoder_decoded_T_120 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], _id_ctrl_decoder_decoded_T_118[23:19], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[15:11], csr_io_decode_0_inst[20], _id_ctrl_decoder_decoded_T_114[8], csr_io_decode_0_inst[22], _id_ctrl_decoder_decoded_T_114[6:5], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:4], csr_io_decode_0_inst[28], _id_ctrl_decoder_decoded_T_106[1:0] };
  assign _id_ctrl_decoder_decoded_T_122 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], csr_io_decode_0_inst[3], _id_ctrl_decoder_decoded_T[3], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T_112[6], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0], csr_io_decode_0_inst[27], csr_io_decode_0_inst[28], _id_ctrl_decoder_decoded_T_106[2:0] };
  assign _id_ctrl_decoder_decoded_T_124 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], csr_io_decode_0_inst[3], _id_ctrl_decoder_decoded_T[3], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T_112[6], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_106[4:3], csr_io_decode_0_inst[29] };
  assign _id_ctrl_decoder_decoded_T_126 = { csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], _id_ctrl_decoder_decoded_T_118[23:19], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[15:11], _id_ctrl_decoder_decoded_T_114[9], csr_io_decode_0_inst[21], _id_ctrl_decoder_decoded_T_114[7:5], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:4], csr_io_decode_0_inst[28], csr_io_decode_0_inst[29], _id_ctrl_decoder_decoded_T_106[1:0] };
  assign _id_ctrl_decoder_decoded_T_128 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], _id_ctrl_decoder_decoded_T_118[23:19], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[15:11], _id_ctrl_decoder_decoded_T_114[9], csr_io_decode_0_inst[21], _id_ctrl_decoder_decoded_T_114[7:5], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:4], csr_io_decode_0_inst[28], csr_io_decode_0_inst[29], _id_ctrl_decoder_decoded_T_106[1:0] };
  assign _id_ctrl_decoder_decoded_T_130 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:2], csr_io_decode_0_inst[30], _id_ctrl_decoder_decoded_T_106[0] };
  assign _id_ctrl_decoder_decoded_T_132 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], csr_io_decode_0_inst[3], _id_ctrl_decoder_decoded_T[3], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T_112[6], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_106[4:3], csr_io_decode_0_inst[30] };
  assign _id_ctrl_decoder_decoded_T_134 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[12], _id_ctrl_decoder_decoded_T[0], csr_io_decode_0_inst[14], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:2], csr_io_decode_0_inst[30], _id_ctrl_decoder_decoded_T_106[0] };
  assign _id_ctrl_decoder_decoded_T_136 = { csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], _id_ctrl_decoder_decoded_T_118[23:19], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[15:11], _id_ctrl_decoder_decoded_T_114[9], csr_io_decode_0_inst[21], _id_ctrl_decoder_decoded_T_114[7:6], csr_io_decode_0_inst[24], csr_io_decode_0_inst[25], _id_ctrl_decoder_decoded_T_106[5], csr_io_decode_0_inst[27], csr_io_decode_0_inst[28], csr_io_decode_0_inst[29], csr_io_decode_0_inst[30], _id_ctrl_decoder_decoded_T_106[0] };
  assign _id_ctrl_decoder_decoded_T_138 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], _id_ctrl_decoder_decoded_T_118[23:19], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[15:11], _id_ctrl_decoder_decoded_T_114[9], csr_io_decode_0_inst[21], _id_ctrl_decoder_decoded_T_114[7:6], csr_io_decode_0_inst[24], csr_io_decode_0_inst[25], _id_ctrl_decoder_decoded_T_106[5], csr_io_decode_0_inst[27], csr_io_decode_0_inst[28], csr_io_decode_0_inst[29], csr_io_decode_0_inst[30], _id_ctrl_decoder_decoded_T_106[0] };
  assign _id_ctrl_decoder_decoded_T_14 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], _id_ctrl_decoder_decoded_T[4], csr_io_decode_0_inst[4], _id_ctrl_decoder_decoded_T[2:1] };
  assign _id_ctrl_decoder_decoded_T_140 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], csr_io_decode_0_inst[3], _id_ctrl_decoder_decoded_T[3], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T_112[6], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_106[4:3], csr_io_decode_0_inst[31] };
  assign _id_ctrl_decoder_decoded_T_16 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:3], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T_10[0] };
  assign _id_ctrl_decoder_decoded_T_18 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:3], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0] };
  assign _id_ctrl_decoder_decoded_T_2 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], _id_ctrl_decoder_decoded_T[2:1], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0] };
  assign _id_ctrl_decoder_decoded_T_20 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:3], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1:0], _id_ctrl_decoder_decoded_T_10[0] };
  assign _id_ctrl_decoder_decoded_T_22 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:2], _id_ctrl_decoder_decoded_T_106[0] };
  assign _id_ctrl_decoder_decoded_T_24 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign _id_ctrl_decoder_decoded_T_26 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:3], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], _id_ctrl_decoder_decoded_T[0] };
  assign _id_ctrl_decoder_decoded_T_28 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:3], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0] };
  assign _id_ctrl_decoder_decoded_T_30 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[4:3], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0] };
  assign _id_ctrl_decoder_decoded_T_32 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], _id_ctrl_decoder_decoded_T[4:3], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0] };
  assign _id_ctrl_decoder_decoded_T_34 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], csr_io_decode_0_inst[3], _id_ctrl_decoder_decoded_T[3], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6] };
  assign _id_ctrl_decoder_decoded_T_36 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], _id_ctrl_decoder_decoded_T_118[23:19], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[15:11], _id_ctrl_decoder_decoded_T_114[8:5], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign _id_ctrl_decoder_decoded_T_38 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], _id_ctrl_decoder_decoded_T_118[23:19], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[15:11], _id_ctrl_decoder_decoded_T_114[8:5], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign _id_ctrl_decoder_decoded_T_4 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:3], _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T_10[0] };
  assign _id_ctrl_decoder_decoded_T_40 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], csr_io_decode_0_inst[3], _id_ctrl_decoder_decoded_T[3:1], csr_io_decode_0_inst[12], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0] };
  assign _id_ctrl_decoder_decoded_T_42 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[12], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign _id_ctrl_decoder_decoded_T_44 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], _id_ctrl_decoder_decoded_T[2:1], csr_io_decode_0_inst[12], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign _id_ctrl_decoder_decoded_T_46 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], csr_io_decode_0_inst[12], _id_ctrl_decoder_decoded_T[0] };
  assign _id_ctrl_decoder_decoded_T_48 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:3], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], csr_io_decode_0_inst[12], _id_ctrl_decoder_decoded_T[0] };
  assign _id_ctrl_decoder_decoded_T_50 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], csr_io_decode_0_inst[12], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0] };
  assign _id_ctrl_decoder_decoded_T_52 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], csr_io_decode_0_inst[12] };
  assign _id_ctrl_decoder_decoded_T_54 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], _id_ctrl_decoder_decoded_T[2:1], csr_io_decode_0_inst[13] };
  assign _id_ctrl_decoder_decoded_T_56 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], _id_ctrl_decoder_decoded_T[2:1], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0] };
  assign _id_ctrl_decoder_decoded_T_58 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], csr_io_decode_0_inst[3], _id_ctrl_decoder_decoded_T[3], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T_112[6], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_106[4:3] };
  assign _id_ctrl_decoder_decoded_T_6 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], _id_ctrl_decoder_decoded_T[2:1], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T_10[0] };
  assign _id_ctrl_decoder_decoded_T_60 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign _id_ctrl_decoder_decoded_T_62 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign _id_ctrl_decoder_decoded_T_64 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], csr_io_decode_0_inst[13] };
  assign _id_ctrl_decoder_decoded_T_66 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0] };
  assign _id_ctrl_decoder_decoded_T_68 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], _id_ctrl_decoder_decoded_T[2:1], csr_io_decode_0_inst[12], csr_io_decode_0_inst[13] };
  assign _id_ctrl_decoder_decoded_T_70 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[12], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign _id_ctrl_decoder_decoded_T_72 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], _id_ctrl_decoder_decoded_T[2:1], _id_ctrl_decoder_decoded_T_112[6], csr_io_decode_0_inst[14] };
  assign _id_ctrl_decoder_decoded_T_74 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[14], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign _id_ctrl_decoder_decoded_T_76 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:3], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], csr_io_decode_0_inst[14] };
  assign _id_ctrl_decoder_decoded_T_78 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[12], _id_ctrl_decoder_decoded_T[0], csr_io_decode_0_inst[14], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:2], _id_ctrl_decoder_decoded_T_106[0] };
  assign _id_ctrl_decoder_decoded_T_8 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:3], _id_ctrl_decoder_decoded_T[1:0], _id_ctrl_decoder_decoded_T_10[0] };
  assign _id_ctrl_decoder_decoded_T_80 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], _id_ctrl_decoder_decoded_T[2:1], csr_io_decode_0_inst[12], _id_ctrl_decoder_decoded_T[0], csr_io_decode_0_inst[14], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:2], _id_ctrl_decoder_decoded_T_106[0] };
  assign _id_ctrl_decoder_decoded_T_82 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[12], _id_ctrl_decoder_decoded_T[0], csr_io_decode_0_inst[14], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign _id_ctrl_decoder_decoded_T_84 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[12], _id_ctrl_decoder_decoded_T[0], csr_io_decode_0_inst[14], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:2], _id_ctrl_decoder_decoded_T_106[0] };
  assign _id_ctrl_decoder_decoded_T_86 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[12], csr_io_decode_0_inst[14], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign _id_ctrl_decoder_decoded_T_88 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], csr_io_decode_0_inst[12], csr_io_decode_0_inst[14] };
  assign _id_ctrl_decoder_decoded_T_90 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:3], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], csr_io_decode_0_inst[12], csr_io_decode_0_inst[14] };
  assign _id_ctrl_decoder_decoded_T_92 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], csr_io_decode_0_inst[12], csr_io_decode_0_inst[14] };
  assign _id_ctrl_decoder_decoded_T_94 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], _id_ctrl_decoder_decoded_T[2:1], csr_io_decode_0_inst[13], csr_io_decode_0_inst[14] };
  assign _id_ctrl_decoder_decoded_T_96 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[13], csr_io_decode_0_inst[14], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign _id_ctrl_decoder_decoded_T_98 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], csr_io_decode_0_inst[13], csr_io_decode_0_inst[14] };
  assign _id_illegal_insn_T_11 = 1'h0;
  assign _id_illegal_insn_T_15 = 1'h0;
  assign _id_illegal_insn_T_33 = 1'h0;
  assign _io_fpu_time_T = csr_io_time;
  assign _mem_br_target_T_3 = { mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[7], mem_reg_inst[30:25], mem_reg_inst[11:8], 1'h0 };
  assign _mem_br_target_T_5 = { mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[19:12], mem_reg_inst[20], mem_reg_inst[30:21], 1'h0 };
  assign { _mem_br_target_T_6[3], _mem_br_target_T_6[1:0] } = { 1'h0, mem_reg_rvc, 1'h0 };
  assign { _mem_br_target_T_7[30:20], _mem_br_target_T_7[0] } = { _mem_br_target_T_7[31], _mem_br_target_T_7[31], _mem_br_target_T_7[31], _mem_br_target_T_7[31], _mem_br_target_T_7[31], _mem_br_target_T_7[31], _mem_br_target_T_7[31], _mem_br_target_T_7[31], _mem_br_target_T_7[31], _mem_br_target_T_7[31], _mem_br_target_T_7[31], 1'h0 };
  assign { _mem_br_target_T_8[30:20], _mem_br_target_T_8[0] } = { _mem_br_target_T_8[31], _mem_br_target_T_8[31], _mem_br_target_T_8[31], _mem_br_target_T_8[31], _mem_br_target_T_8[31], _mem_br_target_T_8[31], _mem_br_target_T_8[31], _mem_br_target_T_8[31], _mem_br_target_T_8[31], _mem_br_target_T_8[31], _mem_br_target_T_8[31], 1'h0 };
  assign _mem_reg_load_T_1 = 1'h0;
  assign _mem_reg_rs2_T_3 = { _ex_op2_T[7:0], _ex_op2_T[7:0], _ex_op2_T[7:0], _ex_op2_T[7:0] };
  assign _mem_reg_rs2_T_6 = { _ex_op2_T[15:0], _ex_op2_T[15:0] };
  assign _mem_reg_rs2_T_7[15:0] = _ex_op2_T[15:0];
  assign _mem_reg_wdata_T = alu_io_out;
  assign _wb_reg_replay_T = io_imem_req_bits_speculative;
  assign alu_io_fn = ex_ctrl_alu_fn;
  assign bpu_io_ea = mem_reg_wdata;
  assign coreMonitorBundle_inst = csr_io_trace_0_insn;
  assign coreMonitorBundle_pc = csr_io_trace_0_iaddr;
  assign csr_clock = clock;
  assign csr_io_bp_0_address = bpu_io_bp_0_address;
  assign csr_io_bp_0_control_action = bpu_io_bp_0_control_action;
  assign csr_io_bp_0_control_r = bpu_io_bp_0_control_r;
  assign csr_io_bp_0_control_tmatch = bpu_io_bp_0_control_tmatch;
  assign csr_io_bp_0_control_w = bpu_io_bp_0_control_w;
  assign csr_io_bp_0_control_x = bpu_io_bp_0_control_x;
  assign csr_io_customCSRs_0_value[1] = io_ptw_customCSRs_csrs_0_value[1];
  assign csr_io_gva = 1'h0;
  assign csr_io_hartid = io_hartid;
  assign csr_io_inst_0 = { _csr_io_inst_0_T_3, wb_reg_raw_inst[15:0] };
  assign csr_io_interrupts_debug = io_interrupts_debug;
  assign csr_io_interrupts_meip = io_interrupts_meip;
  assign csr_io_interrupts_msip = io_interrupts_msip;
  assign csr_io_interrupts_mtip = io_interrupts_mtip;
  assign csr_io_pc = wb_reg_pc;
  assign csr_io_rw_addr = wb_reg_inst[31:20];
  assign csr_io_rw_cmd[1:0] = wb_ctrl_csr[1:0];
  assign csr_io_rw_wdata = wb_reg_wdata;
  assign csr_io_status_debug = bpu_io_status_debug;
  assign csr_io_ungated_clock = clock;
  assign csr_reset = reset;
  assign div_clock = clock;
  assign div_io_req_bits_fn = ex_ctrl_alu_fn;
  assign div_io_req_bits_in1 = _ex_op1_T;
  assign div_io_req_bits_in2 = _ex_op2_T;
  assign div_io_req_bits_tag = ex_reg_inst[11:7];
  assign div_reset = reset;
  assign dmem_resp_waddr = io_dmem_resp_bits_tag[5:1];
  assign ex_ctrl_fp = 1'h0;
  assign ex_ctrl_mem_cmd[4] = 1'h0;
  assign ex_ctrl_mul = 1'h0;
  assign ex_ctrl_rfs1 = 1'h0;
  assign ex_ctrl_rfs2 = 1'h0;
  assign ex_ctrl_rocc = 1'h0;
  assign ex_ctrl_wfd = 1'h0;
  assign ex_dcache_tag = { ex_reg_inst[11:7], 1'h0 };
  assign ex_rs_1 = _ex_op2_T;
  assign ex_waddr = ex_reg_inst[11:7];
  assign ibuf_clock = clock;
  assign ibuf_io_imem_bits_data = io_imem_resp_bits_data;
  assign ibuf_io_imem_bits_pc = io_imem_resp_bits_pc;
  assign ibuf_io_imem_bits_replay = io_imem_resp_bits_replay;
  assign ibuf_io_imem_bits_xcpt_ae_inst = io_imem_resp_bits_xcpt_ae_inst;
  assign ibuf_io_imem_valid = io_imem_resp_valid;
  assign ibuf_io_inst_0_bits_inst_bits = csr_io_decode_0_inst;
  assign ibuf_io_pc = bpu_io_pc;
  assign ibuf_reset = reset;
  assign id_amo_aq = csr_io_decode_0_inst[26];
  assign id_amo_rl = csr_io_decode_0_inst[25];
  assign id_ctrl_decoder_1 = 1'h0;
  assign id_ctrl_decoder_15[4] = 1'h0;
  assign id_ctrl_decoder_16 = 1'h0;
  assign id_ctrl_decoder_17 = 1'h0;
  assign id_ctrl_decoder_19 = 1'h0;
  assign id_ctrl_decoder_2 = 1'h0;
  assign id_ctrl_decoder_20 = 1'h0;
  assign id_ctrl_decoder_27 = 1'h0;
  assign id_ctrl_decoder_8 = 1'h0;
  assign id_ctrl_decoder_decoded_andMatrixInput_0 = csr_io_decode_0_inst[0];
  assign id_ctrl_decoder_decoded_andMatrixInput_1 = csr_io_decode_0_inst[1];
  assign id_ctrl_decoder_decoded_andMatrixInput_10 = _id_ctrl_decoder_decoded_T_118[5];
  assign id_ctrl_decoder_decoded_andMatrixInput_10_20 = csr_io_decode_0_inst[27];
  assign id_ctrl_decoder_decoded_andMatrixInput_11 = _id_ctrl_decoder_decoded_T_106[5];
  assign id_ctrl_decoder_decoded_andMatrixInput_11_1 = _id_ctrl_decoder_decoded_T_106[1];
  assign id_ctrl_decoder_decoded_andMatrixInput_12 = _id_ctrl_decoder_decoded_T_106[4];
  assign id_ctrl_decoder_decoded_andMatrixInput_12_2 = _id_ctrl_decoder_decoded_T_118[15];
  assign id_ctrl_decoder_decoded_andMatrixInput_12_25 = csr_io_decode_0_inst[29];
  assign id_ctrl_decoder_decoded_andMatrixInput_12_33 = csr_io_decode_0_inst[31];
  assign id_ctrl_decoder_decoded_andMatrixInput_13 = _id_ctrl_decoder_decoded_T_106[3];
  assign id_ctrl_decoder_decoded_andMatrixInput_13_1 = _id_ctrl_decoder_decoded_T_118[14];
  assign id_ctrl_decoder_decoded_andMatrixInput_13_19 = csr_io_decode_0_inst[28];
  assign id_ctrl_decoder_decoded_andMatrixInput_14 = _id_ctrl_decoder_decoded_T_106[2];
  assign id_ctrl_decoder_decoded_andMatrixInput_14_1 = _id_ctrl_decoder_decoded_T_118[13];
  assign id_ctrl_decoder_decoded_andMatrixInput_15 = _id_ctrl_decoder_decoded_T_106[0];
  assign id_ctrl_decoder_decoded_andMatrixInput_15_1 = _id_ctrl_decoder_decoded_T_118[12];
  assign id_ctrl_decoder_decoded_andMatrixInput_15_14 = csr_io_decode_0_inst[30];
  assign id_ctrl_decoder_decoded_andMatrixInput_16 = _id_ctrl_decoder_decoded_T_118[11];
  assign id_ctrl_decoder_decoded_andMatrixInput_17 = _id_ctrl_decoder_decoded_T_114[8];
  assign id_ctrl_decoder_decoded_andMatrixInput_17_3 = csr_io_decode_0_inst[20];
  assign id_ctrl_decoder_decoded_andMatrixInput_17_5 = csr_io_decode_0_inst[21];
  assign id_ctrl_decoder_decoded_andMatrixInput_18 = _id_ctrl_decoder_decoded_T_114[7];
  assign id_ctrl_decoder_decoded_andMatrixInput_19 = _id_ctrl_decoder_decoded_T_114[6];
  assign id_ctrl_decoder_decoded_andMatrixInput_19_3 = csr_io_decode_0_inst[22];
  assign id_ctrl_decoder_decoded_andMatrixInput_2 = _id_ctrl_decoder_decoded_T[5];
  assign id_ctrl_decoder_decoded_andMatrixInput_20 = _id_ctrl_decoder_decoded_T_114[5];
  assign id_ctrl_decoder_decoded_andMatrixInput_20_6 = csr_io_decode_0_inst[24];
  assign id_ctrl_decoder_decoded_andMatrixInput_2_5 = csr_io_decode_0_inst[2];
  assign id_ctrl_decoder_decoded_andMatrixInput_3 = _id_ctrl_decoder_decoded_T[4];
  assign id_ctrl_decoder_decoded_andMatrixInput_3_5 = csr_io_decode_0_inst[3];
  assign id_ctrl_decoder_decoded_andMatrixInput_4 = _id_ctrl_decoder_decoded_T[3];
  assign id_ctrl_decoder_decoded_andMatrixInput_4_18 = _id_ctrl_decoder_decoded_T_118[23];
  assign id_ctrl_decoder_decoded_andMatrixInput_4_6 = csr_io_decode_0_inst[4];
  assign id_ctrl_decoder_decoded_andMatrixInput_5 = _id_ctrl_decoder_decoded_T[2];
  assign id_ctrl_decoder_decoded_andMatrixInput_5_18 = _id_ctrl_decoder_decoded_T_118[22];
  assign id_ctrl_decoder_decoded_andMatrixInput_5_8 = csr_io_decode_0_inst[5];
  assign id_ctrl_decoder_decoded_andMatrixInput_6 = _id_ctrl_decoder_decoded_T[1];
  assign id_ctrl_decoder_decoded_andMatrixInput_6_1 = _id_ctrl_decoder_decoded_T_112[6];
  assign id_ctrl_decoder_decoded_andMatrixInput_6_12 = csr_io_decode_0_inst[6];
  assign id_ctrl_decoder_decoded_andMatrixInput_6_17 = _id_ctrl_decoder_decoded_T_118[21];
  assign id_ctrl_decoder_decoded_andMatrixInput_7 = _id_ctrl_decoder_decoded_T[0];
  assign id_ctrl_decoder_decoded_andMatrixInput_7_15 = _id_ctrl_decoder_decoded_T_118[20];
  assign id_ctrl_decoder_decoded_andMatrixInput_7_17 = csr_io_decode_0_inst[12];
  assign id_ctrl_decoder_decoded_andMatrixInput_7_2 = _id_ctrl_decoder_decoded_T_10[0];
  assign id_ctrl_decoder_decoded_andMatrixInput_7_24 = csr_io_decode_0_inst[13];
  assign id_ctrl_decoder_decoded_andMatrixInput_7_50 = csr_io_decode_0_inst[25];
  assign id_ctrl_decoder_decoded_andMatrixInput_7_54 = _id_ctrl_decoder_decoded_T_114[9];
  assign id_ctrl_decoder_decoded_andMatrixInput_8_22 = csr_io_decode_0_inst[14];
  assign id_ctrl_decoder_decoded_andMatrixInput_8_8 = _id_ctrl_decoder_decoded_T_118[19];
  assign id_ctrl_decoder_decoded_hi_58 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], csr_io_decode_0_inst[3], _id_ctrl_decoder_decoded_T[3], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T_112[6], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0] };
  assign id_ctrl_decoder_decoded_hi_lo_17 = { _id_ctrl_decoder_decoded_T_118[20:19], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[15:14] };
  assign id_ctrl_decoder_decoded_hi_lo_18 = { _id_ctrl_decoder_decoded_T_118[22:19], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[15] };
  assign id_ctrl_decoder_decoded_hi_lo_62 = { _id_ctrl_decoder_decoded_T_118[19], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[15:13] };
  assign id_ctrl_decoder_decoded_invInputs[31:2] = { _id_ctrl_decoder_decoded_T_106[0], _id_ctrl_decoder_decoded_T_106[1], _id_ctrl_decoder_decoded_T_106[2], _id_ctrl_decoder_decoded_T_106[3], _id_ctrl_decoder_decoded_T_106[4], _id_ctrl_decoder_decoded_T_106[5], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_114[5], _id_ctrl_decoder_decoded_T_114[6], _id_ctrl_decoder_decoded_T_114[7], _id_ctrl_decoder_decoded_T_114[8], _id_ctrl_decoder_decoded_T_114[9], _id_ctrl_decoder_decoded_T_118[11], _id_ctrl_decoder_decoded_T_118[12], _id_ctrl_decoder_decoded_T_118[13], _id_ctrl_decoder_decoded_T_118[14], _id_ctrl_decoder_decoded_T_118[15], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T_118[19], _id_ctrl_decoder_decoded_T_118[20], _id_ctrl_decoder_decoded_T_118[21], _id_ctrl_decoder_decoded_T_118[22], _id_ctrl_decoder_decoded_T_118[23], _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T[2], _id_ctrl_decoder_decoded_T[3], _id_ctrl_decoder_decoded_T[4], _id_ctrl_decoder_decoded_T[5] };
  assign { id_ctrl_decoder_decoded_invMatrixOutputs[39:38], id_ctrl_decoder_decoded_invMatrixOutputs[32], id_ctrl_decoder_decoded_invMatrixOutputs[18], id_ctrl_decoder_decoded_invMatrixOutputs[13:9], id_ctrl_decoder_decoded_invMatrixOutputs[0] } = 10'h000;
  assign id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_lo[2] = 1'h0;
  assign { id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi[8], id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi[3:0] } = 5'h00;
  assign { id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo[9], id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo[0] } = 2'h0;
  assign id_ctrl_decoder_decoded_lo_11 = { _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:2], _id_ctrl_decoder_decoded_T_106[0] };
  assign id_ctrl_decoder_decoded_lo_12 = _id_ctrl_decoder_decoded_T_106[5:0];
  assign id_ctrl_decoder_decoded_lo_18 = { _id_ctrl_decoder_decoded_T_118[13:11], _id_ctrl_decoder_decoded_T_114[8:5], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign id_ctrl_decoder_decoded_lo_19 = { _id_ctrl_decoder_decoded_T_118[14:11], _id_ctrl_decoder_decoded_T_114[8:5], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign id_ctrl_decoder_decoded_lo_22 = { _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign id_ctrl_decoder_decoded_lo_29 = { _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T_112[6], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_106[4:3] };
  assign id_ctrl_decoder_decoded_lo_31 = { _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign id_ctrl_decoder_decoded_lo_35 = { csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign id_ctrl_decoder_decoded_lo_37 = { csr_io_decode_0_inst[14], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign id_ctrl_decoder_decoded_lo_39 = { csr_io_decode_0_inst[14], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:2], _id_ctrl_decoder_decoded_T_106[0] };
  assign id_ctrl_decoder_decoded_lo_40 = { _id_ctrl_decoder_decoded_T[0], csr_io_decode_0_inst[14], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:2], _id_ctrl_decoder_decoded_T_106[0] };
  assign id_ctrl_decoder_decoded_lo_41 = { csr_io_decode_0_inst[14], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign id_ctrl_decoder_decoded_lo_53 = { csr_io_decode_0_inst[25], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign id_ctrl_decoder_decoded_lo_56 = { _id_ctrl_decoder_decoded_T_112[6], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0], csr_io_decode_0_inst[27], _id_ctrl_decoder_decoded_T_106[2:0] };
  assign id_ctrl_decoder_decoded_lo_57 = { _id_ctrl_decoder_decoded_T_114[7:5], _id_ctrl_decoder_decoded_T_106[4], csr_io_decode_0_inst[28], _id_ctrl_decoder_decoded_T_106[2:0] };
  assign id_ctrl_decoder_decoded_lo_58 = { _id_ctrl_decoder_decoded_T_114[9:5], _id_ctrl_decoder_decoded_T_106[4], csr_io_decode_0_inst[28], _id_ctrl_decoder_decoded_T_106[2:0] };
  assign id_ctrl_decoder_decoded_lo_59 = { _id_ctrl_decoder_decoded_T_118[13:11], csr_io_decode_0_inst[20], _id_ctrl_decoder_decoded_T_114[8], csr_io_decode_0_inst[22], _id_ctrl_decoder_decoded_T_114[6:5], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:4], csr_io_decode_0_inst[28], _id_ctrl_decoder_decoded_T_106[1:0] };
  assign id_ctrl_decoder_decoded_lo_60 = { _id_ctrl_decoder_decoded_T_118[14:11], csr_io_decode_0_inst[20], _id_ctrl_decoder_decoded_T_114[8], csr_io_decode_0_inst[22], _id_ctrl_decoder_decoded_T_114[6:5], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:4], csr_io_decode_0_inst[28], _id_ctrl_decoder_decoded_T_106[1:0] };
  assign id_ctrl_decoder_decoded_lo_61 = { csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0], csr_io_decode_0_inst[27], csr_io_decode_0_inst[28], _id_ctrl_decoder_decoded_T_106[2:0] };
  assign id_ctrl_decoder_decoded_lo_62 = { _id_ctrl_decoder_decoded_T_112[6], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_106[4:3], csr_io_decode_0_inst[29] };
  assign id_ctrl_decoder_decoded_lo_63 = { _id_ctrl_decoder_decoded_T_118[12:11], _id_ctrl_decoder_decoded_T_114[9], csr_io_decode_0_inst[21], _id_ctrl_decoder_decoded_T_114[7:5], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:4], csr_io_decode_0_inst[28], csr_io_decode_0_inst[29], _id_ctrl_decoder_decoded_T_106[1:0] };
  assign id_ctrl_decoder_decoded_lo_64 = { _id_ctrl_decoder_decoded_T_118[14:11], _id_ctrl_decoder_decoded_T_114[9], csr_io_decode_0_inst[21], _id_ctrl_decoder_decoded_T_114[7:5], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:4], csr_io_decode_0_inst[28], csr_io_decode_0_inst[29], _id_ctrl_decoder_decoded_T_106[1:0] };
  assign id_ctrl_decoder_decoded_lo_65 = { _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:2], csr_io_decode_0_inst[30], _id_ctrl_decoder_decoded_T_106[0] };
  assign id_ctrl_decoder_decoded_lo_66 = { _id_ctrl_decoder_decoded_T_112[6], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_106[4:3], csr_io_decode_0_inst[30] };
  assign id_ctrl_decoder_decoded_lo_67 = { csr_io_decode_0_inst[14], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:2], csr_io_decode_0_inst[30], _id_ctrl_decoder_decoded_T_106[0] };
  assign id_ctrl_decoder_decoded_lo_68 = { _id_ctrl_decoder_decoded_T_118[12:11], _id_ctrl_decoder_decoded_T_114[9], csr_io_decode_0_inst[21], _id_ctrl_decoder_decoded_T_114[7:6], csr_io_decode_0_inst[24], csr_io_decode_0_inst[25], _id_ctrl_decoder_decoded_T_106[5], csr_io_decode_0_inst[27], csr_io_decode_0_inst[28], csr_io_decode_0_inst[29], csr_io_decode_0_inst[30], _id_ctrl_decoder_decoded_T_106[0] };
  assign id_ctrl_decoder_decoded_lo_69 = { _id_ctrl_decoder_decoded_T_118[14:11], _id_ctrl_decoder_decoded_T_114[9], csr_io_decode_0_inst[21], _id_ctrl_decoder_decoded_T_114[7:6], csr_io_decode_0_inst[24], csr_io_decode_0_inst[25], _id_ctrl_decoder_decoded_T_106[5], csr_io_decode_0_inst[27], csr_io_decode_0_inst[28], csr_io_decode_0_inst[29], csr_io_decode_0_inst[30], _id_ctrl_decoder_decoded_T_106[0] };
  assign id_ctrl_decoder_decoded_lo_70 = { _id_ctrl_decoder_decoded_T_112[6], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_106[4:3], csr_io_decode_0_inst[31] };
  assign id_ctrl_decoder_decoded_lo_lo_15 = { _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign id_ctrl_decoder_decoded_lo_lo_56 = { _id_ctrl_decoder_decoded_T_114[5], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:4], csr_io_decode_0_inst[28], _id_ctrl_decoder_decoded_T_106[1:0] };
  assign id_ctrl_decoder_decoded_lo_lo_60 = { _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:4], csr_io_decode_0_inst[28], csr_io_decode_0_inst[29], _id_ctrl_decoder_decoded_T_106[1:0] };
  assign id_ctrl_decoder_decoded_lo_lo_61 = { _id_ctrl_decoder_decoded_T_114[5], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:4], csr_io_decode_0_inst[28], csr_io_decode_0_inst[29], _id_ctrl_decoder_decoded_T_106[1:0] };
  assign id_ctrl_decoder_decoded_lo_lo_65 = { csr_io_decode_0_inst[25], _id_ctrl_decoder_decoded_T_106[5], csr_io_decode_0_inst[27], csr_io_decode_0_inst[28], csr_io_decode_0_inst[29], csr_io_decode_0_inst[30], _id_ctrl_decoder_decoded_T_106[0] };
  assign id_ctrl_decoder_decoded_lo_lo_66 = { csr_io_decode_0_inst[24], csr_io_decode_0_inst[25], _id_ctrl_decoder_decoded_T_106[5], csr_io_decode_0_inst[27], csr_io_decode_0_inst[28], csr_io_decode_0_inst[29], csr_io_decode_0_inst[30], _id_ctrl_decoder_decoded_T_106[0] };
  assign { id_ctrl_decoder_decoded_orMatrixOutputs[39:38], id_ctrl_decoder_decoded_orMatrixOutputs[32], id_ctrl_decoder_decoded_orMatrixOutputs[18], id_ctrl_decoder_decoded_orMatrixOutputs[13:9], id_ctrl_decoder_decoded_orMatrixOutputs[0] } = 10'h000;
  assign id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_6[2] = 1'h0;
  assign { id_ctrl_decoder_decoded_orMatrixOutputs_lo_17[18], id_ctrl_decoder_decoded_orMatrixOutputs_lo_17[13:9], id_ctrl_decoder_decoded_orMatrixOutputs_lo_17[0] } = 7'h00;
  assign { id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_10[9], id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_10[0] } = 2'h0;
  assign id_ctrl_decoder_decoded_plaInput = csr_io_decode_0_inst;
  assign id_fence_succ = csr_io_decode_0_inst[23:20];
  assign id_raddr1 = ibuf_io_inst_0_bits_inst_rs1;
  assign id_raddr2 = ibuf_io_inst_0_bits_inst_rs2;
  assign id_waddr = ibuf_io_inst_0_bits_inst_rd;
  assign inst[15:0] = ibuf_io_inst_0_bits_raw[15:0];
  assign io_dmem_req_bits_addr = alu_io_adder_out;
  assign io_dmem_req_bits_cmd = { 1'h0, ex_ctrl_mem_cmd[3:0] };
  assign io_dmem_req_bits_dv = 1'h0;
  assign io_dmem_req_bits_size = ex_reg_mem_size;
  assign io_dmem_req_bits_tag = { 1'h0, ex_reg_inst[11:7], 1'h0 };
  assign io_dmem_s1_data_data = mem_reg_rs2;
  assign io_imem_might_request = imem_might_request_reg;
  assign io_imem_req_valid = ibuf_io_kill;
  assign io_imem_resp_ready = ibuf_io_imem_ready;
  assign { io_ptw_customCSRs_csrs_0_value[31:2], io_ptw_customCSRs_csrs_0_value[0] } = { csr_io_customCSRs_0_value[31:2], csr_io_customCSRs_0_value[0] };
  assign io_ptw_pmp_0_addr = csr_io_pmp_0_addr;
  assign io_ptw_pmp_0_cfg_a = csr_io_pmp_0_cfg_a;
  assign io_ptw_pmp_0_cfg_l = csr_io_pmp_0_cfg_l;
  assign io_ptw_pmp_0_cfg_r = csr_io_pmp_0_cfg_r;
  assign io_ptw_pmp_0_cfg_w = csr_io_pmp_0_cfg_w;
  assign io_ptw_pmp_0_cfg_x = csr_io_pmp_0_cfg_x;
  assign io_ptw_pmp_0_mask = csr_io_pmp_0_mask;
  assign io_ptw_pmp_1_addr = csr_io_pmp_1_addr;
  assign io_ptw_pmp_1_cfg_a = csr_io_pmp_1_cfg_a;
  assign io_ptw_pmp_1_cfg_l = csr_io_pmp_1_cfg_l;
  assign io_ptw_pmp_1_cfg_r = csr_io_pmp_1_cfg_r;
  assign io_ptw_pmp_1_cfg_w = csr_io_pmp_1_cfg_w;
  assign io_ptw_pmp_1_cfg_x = csr_io_pmp_1_cfg_x;
  assign io_ptw_pmp_1_mask = csr_io_pmp_1_mask;
  assign io_ptw_pmp_2_addr = csr_io_pmp_2_addr;
  assign io_ptw_pmp_2_cfg_a = csr_io_pmp_2_cfg_a;
  assign io_ptw_pmp_2_cfg_l = csr_io_pmp_2_cfg_l;
  assign io_ptw_pmp_2_cfg_r = csr_io_pmp_2_cfg_r;
  assign io_ptw_pmp_2_cfg_w = csr_io_pmp_2_cfg_w;
  assign io_ptw_pmp_2_cfg_x = csr_io_pmp_2_cfg_x;
  assign io_ptw_pmp_2_mask = csr_io_pmp_2_mask;
  assign io_ptw_pmp_3_addr = csr_io_pmp_3_addr;
  assign io_ptw_pmp_3_cfg_a = csr_io_pmp_3_cfg_a;
  assign io_ptw_pmp_3_cfg_l = csr_io_pmp_3_cfg_l;
  assign io_ptw_pmp_3_cfg_r = csr_io_pmp_3_cfg_r;
  assign io_ptw_pmp_3_cfg_w = csr_io_pmp_3_cfg_w;
  assign io_ptw_pmp_3_cfg_x = csr_io_pmp_3_cfg_x;
  assign io_ptw_pmp_3_mask = csr_io_pmp_3_mask;
  assign io_ptw_pmp_4_addr = csr_io_pmp_4_addr;
  assign io_ptw_pmp_4_cfg_a = csr_io_pmp_4_cfg_a;
  assign io_ptw_pmp_4_cfg_l = csr_io_pmp_4_cfg_l;
  assign io_ptw_pmp_4_cfg_r = csr_io_pmp_4_cfg_r;
  assign io_ptw_pmp_4_cfg_w = csr_io_pmp_4_cfg_w;
  assign io_ptw_pmp_4_cfg_x = csr_io_pmp_4_cfg_x;
  assign io_ptw_pmp_4_mask = csr_io_pmp_4_mask;
  assign io_ptw_pmp_5_addr = csr_io_pmp_5_addr;
  assign io_ptw_pmp_5_cfg_a = csr_io_pmp_5_cfg_a;
  assign io_ptw_pmp_5_cfg_l = csr_io_pmp_5_cfg_l;
  assign io_ptw_pmp_5_cfg_r = csr_io_pmp_5_cfg_r;
  assign io_ptw_pmp_5_cfg_w = csr_io_pmp_5_cfg_w;
  assign io_ptw_pmp_5_cfg_x = csr_io_pmp_5_cfg_x;
  assign io_ptw_pmp_5_mask = csr_io_pmp_5_mask;
  assign io_ptw_pmp_6_addr = csr_io_pmp_6_addr;
  assign io_ptw_pmp_6_cfg_a = csr_io_pmp_6_cfg_a;
  assign io_ptw_pmp_6_cfg_l = csr_io_pmp_6_cfg_l;
  assign io_ptw_pmp_6_cfg_r = csr_io_pmp_6_cfg_r;
  assign io_ptw_pmp_6_cfg_w = csr_io_pmp_6_cfg_w;
  assign io_ptw_pmp_6_cfg_x = csr_io_pmp_6_cfg_x;
  assign io_ptw_pmp_6_mask = csr_io_pmp_6_mask;
  assign io_ptw_pmp_7_addr = csr_io_pmp_7_addr;
  assign io_ptw_pmp_7_cfg_a = csr_io_pmp_7_cfg_a;
  assign io_ptw_pmp_7_cfg_l = csr_io_pmp_7_cfg_l;
  assign io_ptw_pmp_7_cfg_r = csr_io_pmp_7_cfg_r;
  assign io_ptw_pmp_7_cfg_w = csr_io_pmp_7_cfg_w;
  assign io_ptw_pmp_7_cfg_x = csr_io_pmp_7_cfg_x;
  assign io_ptw_pmp_7_mask = csr_io_pmp_7_mask;
  assign io_ptw_status_debug = bpu_io_status_debug;
  assign io_rocc_cmd_valid = 1'h0;
  assign io_wfi = csr_io_status_wfi;
  assign ll_wdata = div_io_resp_bits_data;
  assign mem_br_target[0] = mem_reg_pc[0];
  assign mem_br_target_b10_5 = mem_reg_inst[30:25];
  assign mem_br_target_b4_1 = mem_reg_inst[11:8];
  assign mem_br_target_hi_hi_hi = mem_reg_inst[31];
  assign mem_br_target_hi_hi_lo = { mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31] };
  assign mem_br_target_hi_lo_hi = { mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31] };
  assign mem_br_target_hi_lo_hi_1 = mem_reg_inst[19:12];
  assign mem_br_target_hi_lo_lo = mem_reg_inst[7];
  assign mem_br_target_hi_lo_lo_1 = mem_reg_inst[20];
  assign mem_br_target_sign = mem_reg_inst[31];
  assign mem_ctrl_fp = 1'h0;
  assign mem_ctrl_mul = 1'h0;
  assign mem_ctrl_rocc = 1'h0;
  assign mem_ldst_cause[1] = 1'h1;
  assign mem_npc[0] = 1'h0;
  assign mem_reg_hls_or_dv = 1'h0;
  assign mem_waddr = mem_reg_inst[11:7];
  assign r = { _r[31:1], 1'h0 };
  assign replay_wb_rocc = 1'h0;
  assign rf_MPORT_mask = 1'h1;
  assign rf_id_rs_MPORT_1_en = 1'h1;
  assign rf_id_rs_MPORT_en = 1'h1;
  assign size = ex_reg_mem_size;
  assign take_pc_mem_wb = ibuf_io_kill;
  assign wb_ctrl_rocc = 1'h0;
  assign wb_reg_hls_or_dv = 1'h0;
  assign wb_valid = csr_io_retire;
  assign wb_waddr = wb_reg_inst[11:7];
  assign wb_xcpt = csr_io_exception;
endmodule
