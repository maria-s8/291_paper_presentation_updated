module \$paramod$1e0019554db24e403a85d4260c10a25441229a90\plusarg_reader (out);
  output [31:0] out;
  wire [31:0] out;
  assign out = 32'd0;
endmodule
module ALU(io_fn, io_in2, io_in1, io_out, io_adder_out, io_cmp_out);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire [31:0] _GEN_0;
  wire [31:0] _GEN_1;
  wire [31:0] _GEN_10;
  wire [31:0] _GEN_11;
  wire [31:0] _GEN_2;
  wire [31:0] _GEN_3;
  wire [31:0] _GEN_4;
  wire [31:0] _GEN_5;
  wire [31:0] _GEN_6;
  wire [31:0] _GEN_7;
  wire [31:0] _GEN_8;
  wire [31:0] _GEN_9;
  wire _shift_logic_T_1;
  wire [31:0] _shin_T_10;
  wire [31:0] _shin_T_11;
  wire [31:0] _shin_T_16;
  wire [31:0] _shin_T_18;
  wire [31:0] _shin_T_20;
  wire [31:0] _shin_T_21;
  wire [31:0] _shin_T_26;
  wire [31:0] _shin_T_28;
  wire [31:0] _shin_T_30;
  wire [31:0] _shin_T_31;
  wire [31:0] _shin_T_36;
  wire [31:0] _shin_T_38;
  wire [31:0] _shin_T_40;
  wire [31:0] _shin_T_41;
  wire [31:0] _shin_T_46;
  wire [31:0] _shin_T_48;
  wire [31:0] _shin_T_50;
  wire [31:0] _shin_T_51;
  wire [31:0] _shin_T_6;
  wire [31:0] _shin_T_8;
  wire [31:0] _shout_l_T_13;
  wire [31:0] _shout_l_T_15;
  wire [31:0] _shout_l_T_17;
  wire [31:0] _shout_l_T_18;
  wire [31:0] _shout_l_T_23;
  wire [31:0] _shout_l_T_25;
  wire [31:0] _shout_l_T_27;
  wire [31:0] _shout_l_T_28;
  wire [31:0] _shout_l_T_3;
  wire [31:0] _shout_l_T_33;
  wire [31:0] _shout_l_T_35;
  wire [31:0] _shout_l_T_37;
  wire [31:0] _shout_l_T_38;
  wire [31:0] _shout_l_T_43;
  wire [31:0] _shout_l_T_45;
  wire [31:0] _shout_l_T_47;
  wire [31:0] _shout_l_T_5;
  wire [31:0] _shout_l_T_7;
  wire [31:0] _shout_l_T_8;
  wire [32:0] _shout_r_T_5;
  output [31:0] io_adder_out;
  wire [31:0] io_adder_out;
  output io_cmp_out;
  wire io_cmp_out;
  input [3:0] io_fn;
  wire [3:0] io_fn;
  input [31:0] io_in1;
  wire [31:0] io_in1;
  input [31:0] io_in2;
  wire [31:0] io_in2;
  output [31:0] io_out;
  wire [31:0] io_out;
  wire [4:0] shamt;
  wire [31:0] shout_l;
  wire [31:0] shout_r;
  INV_X1 _0784_ (
    .A(io_fn[2]),
    .ZN(_0000_)
  );
  INV_X1 _0785_ (
    .A(io_fn[0]),
    .ZN(_0001_)
  );
  INV_X1 _0786_ (
    .A(io_fn[3]),
    .ZN(_0002_)
  );
  INV_X1 _0787_ (
    .A(io_fn[1]),
    .ZN(_0003_)
  );
  INV_X1 _0788_ (
    .A(io_in2[0]),
    .ZN(_0004_)
  );
  INV_X1 _0789_ (
    .A(io_in2[1]),
    .ZN(_0005_)
  );
  INV_X1 _0790_ (
    .A(io_in2[31]),
    .ZN(_0006_)
  );
  INV_X1 _0791_ (
    .A(io_in1[31]),
    .ZN(_0007_)
  );
  XOR2_X1 _0792_ (
    .A(io_fn[3]),
    .B(io_in2[22]),
    .Z(_0008_)
  );
  AND2_X1 _0793_ (
    .A1(io_in1[22]),
    .A2(_0008_),
    .ZN(_0009_)
  );
  XOR2_X1 _0794_ (
    .A(io_in1[22]),
    .B(_0008_),
    .Z(_0010_)
  );
  XOR2_X1 _0795_ (
    .A(io_fn[3]),
    .B(io_in2[21]),
    .Z(_0011_)
  );
  AND2_X1 _0796_ (
    .A1(io_in1[21]),
    .A2(_0011_),
    .ZN(_0012_)
  );
  OR2_X1 _0797_ (
    .A1(io_in1[21]),
    .A2(_0011_),
    .ZN(_0013_)
  );
  XOR2_X1 _0798_ (
    .A(io_fn[3]),
    .B(io_in2[20]),
    .Z(_0014_)
  );
  AND2_X1 _0799_ (
    .A1(io_in1[20]),
    .A2(_0014_),
    .ZN(_0015_)
  );
  XOR2_X1 _0800_ (
    .A(io_in1[20]),
    .B(_0014_),
    .Z(_0016_)
  );
  XOR2_X1 _0801_ (
    .A(io_fn[3]),
    .B(io_in2[19]),
    .Z(_0017_)
  );
  AND2_X1 _0802_ (
    .A1(io_in1[19]),
    .A2(_0017_),
    .ZN(_0018_)
  );
  XOR2_X1 _0803_ (
    .A(io_in1[19]),
    .B(_0017_),
    .Z(_0019_)
  );
  XOR2_X1 _0804_ (
    .A(io_fn[3]),
    .B(io_in2[18]),
    .Z(_0020_)
  );
  AND2_X1 _0805_ (
    .A1(io_in1[18]),
    .A2(_0020_),
    .ZN(_0021_)
  );
  XOR2_X1 _0806_ (
    .A(io_in1[18]),
    .B(_0020_),
    .Z(_0022_)
  );
  XOR2_X1 _0807_ (
    .A(io_fn[3]),
    .B(io_in2[17]),
    .Z(_0023_)
  );
  AND2_X1 _0808_ (
    .A1(io_in1[17]),
    .A2(_0023_),
    .ZN(_0024_)
  );
  XOR2_X1 _0809_ (
    .A(io_fn[3]),
    .B(io_in2[16]),
    .Z(_0025_)
  );
  AND2_X1 _0810_ (
    .A1(io_in1[16]),
    .A2(_0025_),
    .ZN(_0026_)
  );
  XOR2_X1 _0811_ (
    .A(io_fn[3]),
    .B(io_in2[15]),
    .Z(_0027_)
  );
  OR2_X1 _0812_ (
    .A1(io_in1[15]),
    .A2(_0027_),
    .ZN(_0028_)
  );
  AND2_X1 _0813_ (
    .A1(io_in1[15]),
    .A2(_0027_),
    .ZN(_0029_)
  );
  XOR2_X1 _0814_ (
    .A(io_in1[15]),
    .B(_0027_),
    .Z(_0030_)
  );
  XOR2_X1 _0815_ (
    .A(io_fn[3]),
    .B(io_in2[14]),
    .Z(_0031_)
  );
  AND2_X1 _0816_ (
    .A1(io_in1[14]),
    .A2(_0031_),
    .ZN(_0032_)
  );
  XOR2_X1 _0817_ (
    .A(io_in1[14]),
    .B(_0031_),
    .Z(_0033_)
  );
  XOR2_X1 _0818_ (
    .A(io_fn[3]),
    .B(io_in2[13]),
    .Z(_0034_)
  );
  AND2_X1 _0819_ (
    .A1(io_in1[13]),
    .A2(_0034_),
    .ZN(_0035_)
  );
  OR2_X1 _0820_ (
    .A1(io_in1[13]),
    .A2(_0034_),
    .ZN(_0036_)
  );
  XOR2_X1 _0821_ (
    .A(io_in1[13]),
    .B(_0034_),
    .Z(_0037_)
  );
  XOR2_X1 _0822_ (
    .A(io_fn[3]),
    .B(io_in2[12]),
    .Z(_0038_)
  );
  AND2_X1 _0823_ (
    .A1(io_in1[12]),
    .A2(_0038_),
    .ZN(_0039_)
  );
  XOR2_X1 _0824_ (
    .A(io_in1[12]),
    .B(_0038_),
    .Z(_0040_)
  );
  XOR2_X1 _0825_ (
    .A(io_fn[3]),
    .B(io_in2[11]),
    .Z(_0041_)
  );
  AND2_X1 _0826_ (
    .A1(io_in1[11]),
    .A2(_0041_),
    .ZN(_0042_)
  );
  OR2_X1 _0827_ (
    .A1(io_in1[11]),
    .A2(_0041_),
    .ZN(_0043_)
  );
  XOR2_X1 _0828_ (
    .A(io_in1[11]),
    .B(_0041_),
    .Z(_0044_)
  );
  XOR2_X1 _0829_ (
    .A(io_fn[3]),
    .B(io_in2[10]),
    .Z(_0045_)
  );
  AND2_X1 _0830_ (
    .A1(io_in1[10]),
    .A2(_0045_),
    .ZN(_0046_)
  );
  XOR2_X1 _0831_ (
    .A(io_in1[10]),
    .B(_0045_),
    .Z(_0047_)
  );
  XOR2_X1 _0832_ (
    .A(io_fn[3]),
    .B(io_in2[9]),
    .Z(_0048_)
  );
  AND2_X1 _0833_ (
    .A1(io_in1[9]),
    .A2(_0048_),
    .ZN(_0049_)
  );
  XOR2_X1 _0834_ (
    .A(io_in1[9]),
    .B(_0048_),
    .Z(_0050_)
  );
  XOR2_X1 _0835_ (
    .A(io_fn[3]),
    .B(io_in2[8]),
    .Z(_0051_)
  );
  AND2_X1 _0836_ (
    .A1(io_in1[8]),
    .A2(_0051_),
    .ZN(_0052_)
  );
  XOR2_X1 _0837_ (
    .A(io_fn[3]),
    .B(io_in2[7]),
    .Z(_0053_)
  );
  AND2_X1 _0838_ (
    .A1(io_in1[7]),
    .A2(_0053_),
    .ZN(_0054_)
  );
  XOR2_X1 _0839_ (
    .A(io_in1[7]),
    .B(_0053_),
    .Z(_0055_)
  );
  XOR2_X1 _0840_ (
    .A(io_fn[3]),
    .B(io_in2[6]),
    .Z(_0056_)
  );
  AND2_X1 _0841_ (
    .A1(io_in1[6]),
    .A2(_0056_),
    .ZN(_0057_)
  );
  XOR2_X1 _0842_ (
    .A(io_in1[6]),
    .B(_0056_),
    .Z(_0058_)
  );
  XOR2_X1 _0843_ (
    .A(io_fn[3]),
    .B(io_in2[5]),
    .Z(_0059_)
  );
  AND2_X1 _0844_ (
    .A1(io_in1[5]),
    .A2(_0059_),
    .ZN(_0060_)
  );
  XOR2_X1 _0845_ (
    .A(io_fn[3]),
    .B(io_in2[4]),
    .Z(_0061_)
  );
  AND2_X1 _0846_ (
    .A1(io_in1[4]),
    .A2(_0061_),
    .ZN(_0062_)
  );
  XOR2_X1 _0847_ (
    .A(io_fn[3]),
    .B(io_in2[3]),
    .Z(_0063_)
  );
  AND2_X1 _0848_ (
    .A1(io_in1[3]),
    .A2(_0063_),
    .ZN(_0064_)
  );
  XOR2_X1 _0849_ (
    .A(io_fn[3]),
    .B(io_in2[2]),
    .Z(_0065_)
  );
  AND2_X1 _0850_ (
    .A1(io_in1[2]),
    .A2(_0065_),
    .ZN(_0066_)
  );
  OR2_X1 _0851_ (
    .A1(io_fn[3]),
    .A2(_0005_),
    .ZN(_0067_)
  );
  XOR2_X1 _0852_ (
    .A(io_fn[3]),
    .B(io_in2[1]),
    .Z(_0068_)
  );
  AND2_X1 _0853_ (
    .A1(io_in1[1]),
    .A2(_0068_),
    .ZN(_0069_)
  );
  OR2_X1 _0854_ (
    .A1(io_fn[3]),
    .A2(_0004_),
    .ZN(_0070_)
  );
  XOR2_X1 _0855_ (
    .A(io_fn[3]),
    .B(io_in2[0]),
    .Z(_0071_)
  );
  AND2_X1 _0856_ (
    .A1(io_in1[0]),
    .A2(_0071_),
    .ZN(_0072_)
  );
  XOR2_X1 _0857_ (
    .A(io_in1[1]),
    .B(_0068_),
    .Z(_0073_)
  );
  INV_X1 _0858_ (
    .A(_0073_),
    .ZN(_0074_)
  );
  AND2_X1 _0859_ (
    .A1(_0072_),
    .A2(_0073_),
    .ZN(_0075_)
  );
  OR2_X1 _0860_ (
    .A1(_0069_),
    .A2(_0075_),
    .ZN(_0076_)
  );
  XOR2_X1 _0861_ (
    .A(io_in1[2]),
    .B(_0065_),
    .Z(_0077_)
  );
  AND2_X1 _0862_ (
    .A1(_0076_),
    .A2(_0077_),
    .ZN(_0078_)
  );
  OR2_X1 _0863_ (
    .A1(_0066_),
    .A2(_0078_),
    .ZN(_0079_)
  );
  XOR2_X1 _0864_ (
    .A(io_in1[3]),
    .B(_0063_),
    .Z(_0080_)
  );
  AND2_X1 _0865_ (
    .A1(_0079_),
    .A2(_0080_),
    .ZN(_0081_)
  );
  OR2_X1 _0866_ (
    .A1(_0064_),
    .A2(_0081_),
    .ZN(_0082_)
  );
  XOR2_X1 _0867_ (
    .A(io_in1[4]),
    .B(_0061_),
    .Z(_0083_)
  );
  AND2_X1 _0868_ (
    .A1(_0082_),
    .A2(_0083_),
    .ZN(_0084_)
  );
  OR2_X1 _0869_ (
    .A1(_0062_),
    .A2(_0084_),
    .ZN(_0085_)
  );
  XOR2_X1 _0870_ (
    .A(io_in1[5]),
    .B(_0059_),
    .Z(_0086_)
  );
  AND2_X1 _0871_ (
    .A1(_0085_),
    .A2(_0086_),
    .ZN(_0087_)
  );
  OR2_X1 _0872_ (
    .A1(_0060_),
    .A2(_0087_),
    .ZN(_0088_)
  );
  AND2_X1 _0873_ (
    .A1(_0058_),
    .A2(_0088_),
    .ZN(_0089_)
  );
  OR2_X1 _0874_ (
    .A1(_0057_),
    .A2(_0089_),
    .ZN(_0090_)
  );
  AND2_X1 _0875_ (
    .A1(_0055_),
    .A2(_0090_),
    .ZN(_0091_)
  );
  OR2_X1 _0876_ (
    .A1(_0054_),
    .A2(_0091_),
    .ZN(_0092_)
  );
  XOR2_X1 _0877_ (
    .A(io_in1[8]),
    .B(_0051_),
    .Z(_0093_)
  );
  AND2_X1 _0878_ (
    .A1(_0092_),
    .A2(_0093_),
    .ZN(_0094_)
  );
  OR2_X1 _0879_ (
    .A1(_0052_),
    .A2(_0094_),
    .ZN(_0095_)
  );
  AND2_X1 _0880_ (
    .A1(_0050_),
    .A2(_0095_),
    .ZN(_0096_)
  );
  OR2_X1 _0881_ (
    .A1(_0049_),
    .A2(_0096_),
    .ZN(_0097_)
  );
  AND2_X1 _0882_ (
    .A1(_0047_),
    .A2(_0097_),
    .ZN(_0098_)
  );
  AND2_X1 _0883_ (
    .A1(_0044_),
    .A2(_0098_),
    .ZN(_0099_)
  );
  AND2_X1 _0884_ (
    .A1(_0043_),
    .A2(_0046_),
    .ZN(_0100_)
  );
  OR2_X1 _0885_ (
    .A1(_0042_),
    .A2(_0100_),
    .ZN(_0101_)
  );
  OR2_X1 _0886_ (
    .A1(_0099_),
    .A2(_0101_),
    .ZN(_0102_)
  );
  AND2_X1 _0887_ (
    .A1(_0040_),
    .A2(_0102_),
    .ZN(_0103_)
  );
  AND2_X1 _0888_ (
    .A1(_0037_),
    .A2(_0103_),
    .ZN(_0104_)
  );
  OR2_X1 _0889_ (
    .A1(_0035_),
    .A2(_0039_),
    .ZN(_0105_)
  );
  AND2_X1 _0890_ (
    .A1(_0036_),
    .A2(_0105_),
    .ZN(_0106_)
  );
  OR2_X1 _0891_ (
    .A1(_0104_),
    .A2(_0106_),
    .ZN(_0107_)
  );
  AND2_X1 _0892_ (
    .A1(_0033_),
    .A2(_0107_),
    .ZN(_0108_)
  );
  AND2_X1 _0893_ (
    .A1(_0030_),
    .A2(_0108_),
    .ZN(_0109_)
  );
  OR2_X1 _0894_ (
    .A1(_0029_),
    .A2(_0032_),
    .ZN(_0110_)
  );
  AND2_X1 _0895_ (
    .A1(_0028_),
    .A2(_0110_),
    .ZN(_0111_)
  );
  OR2_X1 _0896_ (
    .A1(_0109_),
    .A2(_0111_),
    .ZN(_0112_)
  );
  XOR2_X1 _0897_ (
    .A(io_in1[16]),
    .B(_0025_),
    .Z(_0113_)
  );
  AND2_X1 _0898_ (
    .A1(_0112_),
    .A2(_0113_),
    .ZN(_0114_)
  );
  OR2_X1 _0899_ (
    .A1(_0026_),
    .A2(_0114_),
    .ZN(_0115_)
  );
  XOR2_X1 _0900_ (
    .A(io_in1[17]),
    .B(_0023_),
    .Z(_0116_)
  );
  AND2_X1 _0901_ (
    .A1(_0115_),
    .A2(_0116_),
    .ZN(_0117_)
  );
  OR2_X1 _0902_ (
    .A1(_0024_),
    .A2(_0117_),
    .ZN(_0118_)
  );
  AND2_X1 _0903_ (
    .A1(_0022_),
    .A2(_0118_),
    .ZN(_0119_)
  );
  OR2_X1 _0904_ (
    .A1(_0021_),
    .A2(_0119_),
    .ZN(_0120_)
  );
  AND2_X1 _0905_ (
    .A1(_0019_),
    .A2(_0120_),
    .ZN(_0121_)
  );
  OR2_X1 _0906_ (
    .A1(_0018_),
    .A2(_0121_),
    .ZN(_0122_)
  );
  AND2_X1 _0907_ (
    .A1(_0016_),
    .A2(_0122_),
    .ZN(_0123_)
  );
  OR2_X1 _0908_ (
    .A1(_0015_),
    .A2(_0123_),
    .ZN(_0124_)
  );
  AND2_X1 _0909_ (
    .A1(_0013_),
    .A2(_0124_),
    .ZN(_0125_)
  );
  OR2_X1 _0910_ (
    .A1(_0012_),
    .A2(_0125_),
    .ZN(_0126_)
  );
  AND2_X1 _0911_ (
    .A1(_0010_),
    .A2(_0126_),
    .ZN(_0127_)
  );
  XOR2_X1 _0912_ (
    .A(_0010_),
    .B(_0126_),
    .Z(_0128_)
  );
  XOR2_X1 _0913_ (
    .A(_0016_),
    .B(_0122_),
    .Z(_0129_)
  );
  XOR2_X1 _0914_ (
    .A(_0115_),
    .B(_0116_),
    .Z(_0130_)
  );
  XOR2_X1 _0915_ (
    .A(_0112_),
    .B(_0113_),
    .Z(_0131_)
  );
  XOR2_X1 _0916_ (
    .A(_0033_),
    .B(_0107_),
    .Z(_0132_)
  );
  XOR2_X1 _0917_ (
    .A(_0092_),
    .B(_0093_),
    .Z(_0133_)
  );
  XOR2_X1 _0918_ (
    .A(io_in1[0]),
    .B(_0071_),
    .Z(_0134_)
  );
  AND2_X1 _0919_ (
    .A1(io_fn[3]),
    .A2(_0134_),
    .ZN(_0135_)
  );
  AND2_X1 _0920_ (
    .A1(_0073_),
    .A2(_0135_),
    .ZN(_0136_)
  );
  XOR2_X1 _0921_ (
    .A(_0076_),
    .B(_0077_),
    .Z(_0137_)
  );
  AND2_X1 _0922_ (
    .A1(_0136_),
    .A2(_0137_),
    .ZN(_0138_)
  );
  XOR2_X1 _0923_ (
    .A(_0079_),
    .B(_0080_),
    .Z(_0139_)
  );
  AND2_X1 _0924_ (
    .A1(_0138_),
    .A2(_0139_),
    .ZN(_0140_)
  );
  XOR2_X1 _0925_ (
    .A(_0082_),
    .B(_0083_),
    .Z(_0141_)
  );
  AND2_X1 _0926_ (
    .A1(_0140_),
    .A2(_0141_),
    .ZN(_0142_)
  );
  XOR2_X1 _0927_ (
    .A(_0085_),
    .B(_0086_),
    .Z(_0143_)
  );
  AND2_X1 _0928_ (
    .A1(_0142_),
    .A2(_0143_),
    .ZN(_0144_)
  );
  XOR2_X1 _0929_ (
    .A(_0058_),
    .B(_0088_),
    .Z(_0145_)
  );
  AND2_X1 _0930_ (
    .A1(_0144_),
    .A2(_0145_),
    .ZN(_0146_)
  );
  XOR2_X1 _0931_ (
    .A(_0055_),
    .B(_0090_),
    .Z(_0147_)
  );
  AND2_X1 _0932_ (
    .A1(_0146_),
    .A2(_0147_),
    .ZN(_0148_)
  );
  AND2_X1 _0933_ (
    .A1(_0133_),
    .A2(_0148_),
    .ZN(_0149_)
  );
  XOR2_X1 _0934_ (
    .A(_0050_),
    .B(_0095_),
    .Z(_0150_)
  );
  AND2_X1 _0935_ (
    .A1(_0149_),
    .A2(_0150_),
    .ZN(_0151_)
  );
  XOR2_X1 _0936_ (
    .A(_0047_),
    .B(_0097_),
    .Z(_0152_)
  );
  AND2_X1 _0937_ (
    .A1(_0151_),
    .A2(_0152_),
    .ZN(_0153_)
  );
  OR2_X1 _0938_ (
    .A1(_0046_),
    .A2(_0098_),
    .ZN(_0154_)
  );
  XOR2_X1 _0939_ (
    .A(_0044_),
    .B(_0154_),
    .Z(_0155_)
  );
  AND2_X1 _0940_ (
    .A1(_0153_),
    .A2(_0155_),
    .ZN(_0156_)
  );
  XOR2_X1 _0941_ (
    .A(_0040_),
    .B(_0102_),
    .Z(_0157_)
  );
  AND2_X1 _0942_ (
    .A1(_0156_),
    .A2(_0157_),
    .ZN(_0158_)
  );
  OR2_X1 _0943_ (
    .A1(_0039_),
    .A2(_0103_),
    .ZN(_0159_)
  );
  XOR2_X1 _0944_ (
    .A(_0037_),
    .B(_0159_),
    .Z(_0160_)
  );
  AND2_X1 _0945_ (
    .A1(_0158_),
    .A2(_0160_),
    .ZN(_0161_)
  );
  AND2_X1 _0946_ (
    .A1(_0132_),
    .A2(_0161_),
    .ZN(_0162_)
  );
  OR2_X1 _0947_ (
    .A1(_0032_),
    .A2(_0108_),
    .ZN(_0163_)
  );
  XOR2_X1 _0948_ (
    .A(_0030_),
    .B(_0163_),
    .Z(_0164_)
  );
  AND2_X1 _0949_ (
    .A1(_0162_),
    .A2(_0164_),
    .ZN(_0165_)
  );
  AND2_X1 _0950_ (
    .A1(_0131_),
    .A2(_0165_),
    .ZN(_0166_)
  );
  AND2_X1 _0951_ (
    .A1(_0130_),
    .A2(_0166_),
    .ZN(_0167_)
  );
  XOR2_X1 _0952_ (
    .A(_0022_),
    .B(_0118_),
    .Z(_0168_)
  );
  AND2_X1 _0953_ (
    .A1(_0167_),
    .A2(_0168_),
    .ZN(_0169_)
  );
  XOR2_X1 _0954_ (
    .A(_0019_),
    .B(_0120_),
    .Z(_0170_)
  );
  AND2_X1 _0955_ (
    .A1(_0169_),
    .A2(_0170_),
    .ZN(_0171_)
  );
  AND2_X1 _0956_ (
    .A1(_0129_),
    .A2(_0171_),
    .ZN(_0172_)
  );
  XOR2_X1 _0957_ (
    .A(io_in1[21]),
    .B(_0011_),
    .Z(_0173_)
  );
  XOR2_X1 _0958_ (
    .A(_0124_),
    .B(_0173_),
    .Z(_0174_)
  );
  AND2_X1 _0959_ (
    .A1(_0172_),
    .A2(_0174_),
    .ZN(_0175_)
  );
  AND2_X1 _0960_ (
    .A1(_0128_),
    .A2(_0175_),
    .ZN(_0176_)
  );
  XOR2_X1 _0961_ (
    .A(io_fn[3]),
    .B(io_in2[23]),
    .Z(_0177_)
  );
  AND2_X1 _0962_ (
    .A1(io_in1[23]),
    .A2(_0177_),
    .ZN(_0178_)
  );
  OR2_X1 _0963_ (
    .A1(io_in1[23]),
    .A2(_0177_),
    .ZN(_0179_)
  );
  XOR2_X1 _0964_ (
    .A(io_in1[23]),
    .B(_0177_),
    .Z(_0180_)
  );
  OR2_X1 _0965_ (
    .A1(_0009_),
    .A2(_0127_),
    .ZN(_0181_)
  );
  XOR2_X1 _0966_ (
    .A(_0180_),
    .B(_0181_),
    .Z(_0182_)
  );
  AND2_X1 _0967_ (
    .A1(_0176_),
    .A2(_0182_),
    .ZN(_0183_)
  );
  XOR2_X1 _0968_ (
    .A(io_fn[3]),
    .B(io_in2[24]),
    .Z(_0184_)
  );
  AND2_X1 _0969_ (
    .A1(io_in1[24]),
    .A2(_0184_),
    .ZN(_0185_)
  );
  XOR2_X1 _0970_ (
    .A(io_in1[24]),
    .B(_0184_),
    .Z(_0186_)
  );
  AND2_X1 _0971_ (
    .A1(_0179_),
    .A2(_0181_),
    .ZN(_0187_)
  );
  OR2_X1 _0972_ (
    .A1(_0178_),
    .A2(_0187_),
    .ZN(_0188_)
  );
  AND2_X1 _0973_ (
    .A1(_0186_),
    .A2(_0188_),
    .ZN(_0189_)
  );
  XOR2_X1 _0974_ (
    .A(_0186_),
    .B(_0188_),
    .Z(_0190_)
  );
  AND2_X1 _0975_ (
    .A1(_0183_),
    .A2(_0190_),
    .ZN(_0191_)
  );
  XOR2_X1 _0976_ (
    .A(io_fn[3]),
    .B(io_in2[25]),
    .Z(_0192_)
  );
  AND2_X1 _0977_ (
    .A1(io_in1[25]),
    .A2(_0192_),
    .ZN(_0193_)
  );
  XOR2_X1 _0978_ (
    .A(io_in1[25]),
    .B(_0192_),
    .Z(_0194_)
  );
  OR2_X1 _0979_ (
    .A1(_0185_),
    .A2(_0189_),
    .ZN(_0195_)
  );
  AND2_X1 _0980_ (
    .A1(_0194_),
    .A2(_0195_),
    .ZN(_0196_)
  );
  XOR2_X1 _0981_ (
    .A(_0194_),
    .B(_0195_),
    .Z(_0197_)
  );
  AND2_X1 _0982_ (
    .A1(_0191_),
    .A2(_0197_),
    .ZN(_0198_)
  );
  XOR2_X1 _0983_ (
    .A(io_fn[3]),
    .B(io_in2[26]),
    .Z(_0199_)
  );
  AND2_X1 _0984_ (
    .A1(io_in1[26]),
    .A2(_0199_),
    .ZN(_0200_)
  );
  XOR2_X1 _0985_ (
    .A(io_in1[26]),
    .B(_0199_),
    .Z(_0201_)
  );
  OR2_X1 _0986_ (
    .A1(_0193_),
    .A2(_0196_),
    .ZN(_0202_)
  );
  AND2_X1 _0987_ (
    .A1(_0201_),
    .A2(_0202_),
    .ZN(_0203_)
  );
  XOR2_X1 _0988_ (
    .A(_0201_),
    .B(_0202_),
    .Z(_0204_)
  );
  AND2_X1 _0989_ (
    .A1(_0198_),
    .A2(_0204_),
    .ZN(_0205_)
  );
  XOR2_X1 _0990_ (
    .A(io_fn[3]),
    .B(io_in2[27]),
    .Z(_0206_)
  );
  AND2_X1 _0991_ (
    .A1(io_in1[27]),
    .A2(_0206_),
    .ZN(_0207_)
  );
  XOR2_X1 _0992_ (
    .A(io_in1[27]),
    .B(_0206_),
    .Z(_0208_)
  );
  OR2_X1 _0993_ (
    .A1(_0200_),
    .A2(_0203_),
    .ZN(_0209_)
  );
  AND2_X1 _0994_ (
    .A1(_0208_),
    .A2(_0209_),
    .ZN(_0210_)
  );
  XOR2_X1 _0995_ (
    .A(_0208_),
    .B(_0209_),
    .Z(_0211_)
  );
  AND2_X1 _0996_ (
    .A1(_0205_),
    .A2(_0211_),
    .ZN(_0212_)
  );
  OR2_X1 _0997_ (
    .A1(_0207_),
    .A2(_0210_),
    .ZN(_0213_)
  );
  XOR2_X1 _0998_ (
    .A(io_fn[3]),
    .B(io_in2[28]),
    .Z(_0214_)
  );
  AND2_X1 _0999_ (
    .A1(io_in1[28]),
    .A2(_0214_),
    .ZN(_0215_)
  );
  XOR2_X1 _1000_ (
    .A(io_in1[28]),
    .B(_0214_),
    .Z(_0216_)
  );
  AND2_X1 _1001_ (
    .A1(_0213_),
    .A2(_0216_),
    .ZN(_0217_)
  );
  XOR2_X1 _1002_ (
    .A(_0213_),
    .B(_0216_),
    .Z(_0218_)
  );
  AND2_X1 _1003_ (
    .A1(_0212_),
    .A2(_0218_),
    .ZN(_0219_)
  );
  XOR2_X1 _1004_ (
    .A(io_fn[3]),
    .B(io_in2[29]),
    .Z(_0220_)
  );
  AND2_X1 _1005_ (
    .A1(io_in1[29]),
    .A2(_0220_),
    .ZN(_0221_)
  );
  XOR2_X1 _1006_ (
    .A(io_in1[29]),
    .B(_0220_),
    .Z(_0222_)
  );
  OR2_X1 _1007_ (
    .A1(_0215_),
    .A2(_0217_),
    .ZN(_0223_)
  );
  AND2_X1 _1008_ (
    .A1(_0222_),
    .A2(_0223_),
    .ZN(_0224_)
  );
  XOR2_X1 _1009_ (
    .A(_0222_),
    .B(_0223_),
    .Z(_0225_)
  );
  AND2_X1 _1010_ (
    .A1(_0219_),
    .A2(_0225_),
    .ZN(_0226_)
  );
  OR2_X1 _1011_ (
    .A1(_0221_),
    .A2(_0224_),
    .ZN(_0227_)
  );
  XOR2_X1 _1012_ (
    .A(io_fn[3]),
    .B(io_in2[30]),
    .Z(_0228_)
  );
  AND2_X1 _1013_ (
    .A1(io_in1[30]),
    .A2(_0228_),
    .ZN(_0229_)
  );
  XOR2_X1 _1014_ (
    .A(io_in1[30]),
    .B(_0228_),
    .Z(_0230_)
  );
  AND2_X1 _1015_ (
    .A1(_0227_),
    .A2(_0230_),
    .ZN(_0231_)
  );
  XOR2_X1 _1016_ (
    .A(_0227_),
    .B(_0230_),
    .Z(_0232_)
  );
  AND2_X1 _1017_ (
    .A1(_0226_),
    .A2(_0232_),
    .ZN(_0233_)
  );
  OR2_X1 _1018_ (
    .A1(_0229_),
    .A2(_0231_),
    .ZN(_0234_)
  );
  AND2_X1 _1019_ (
    .A1(io_in2[31]),
    .A2(_0007_),
    .ZN(_0235_)
  );
  AND2_X1 _1020_ (
    .A1(_0006_),
    .A2(io_in1[31]),
    .ZN(_0236_)
  );
  OR2_X1 _1021_ (
    .A1(_0235_),
    .A2(_0236_),
    .ZN(_0237_)
  );
  INV_X1 _1022_ (
    .A(_0237_),
    .ZN(_0238_)
  );
  AND2_X1 _1023_ (
    .A1(io_fn[3]),
    .A2(_0238_),
    .ZN(_0239_)
  );
  XOR2_X1 _1024_ (
    .A(io_fn[3]),
    .B(_0237_),
    .Z(_0240_)
  );
  XOR2_X1 _1025_ (
    .A(_0234_),
    .B(_0240_),
    .Z(_0241_)
  );
  XOR2_X1 _1026_ (
    .A(_0233_),
    .B(_0241_),
    .Z(io_adder_out[31])
  );
  OR2_X1 _1027_ (
    .A1(io_fn[3]),
    .A2(_0134_),
    .ZN(_0242_)
  );
  XOR2_X1 _1028_ (
    .A(io_in2[0]),
    .B(io_in1[0]),
    .Z(io_adder_out[0])
  );
  AND2_X1 _1029_ (
    .A1(_0239_),
    .A2(io_adder_out[31]),
    .ZN(_0243_)
  );
  AND2_X1 _1030_ (
    .A1(io_fn[3]),
    .A2(io_fn[1]),
    .ZN(_0244_)
  );
  AND2_X1 _1031_ (
    .A1(_0235_),
    .A2(_0244_),
    .ZN(_0245_)
  );
  AND2_X1 _1032_ (
    .A1(io_fn[3]),
    .A2(_0003_),
    .ZN(_0246_)
  );
  AND2_X1 _1033_ (
    .A1(_0236_),
    .A2(_0246_),
    .ZN(_0247_)
  );
  OR2_X1 _1034_ (
    .A1(_0245_),
    .A2(_0247_),
    .ZN(_0248_)
  );
  OR2_X1 _1035_ (
    .A1(_0243_),
    .A2(_0248_),
    .ZN(_0249_)
  );
  AND2_X1 _1036_ (
    .A1(io_fn[2]),
    .A2(_0249_),
    .ZN(_0250_)
  );
  AND2_X1 _1037_ (
    .A1(_0000_),
    .A2(_0244_),
    .ZN(_0251_)
  );
  AND2_X1 _1038_ (
    .A1(io_fn[2]),
    .A2(_0002_),
    .ZN(_0252_)
  );
  AND2_X1 _1039_ (
    .A1(_0003_),
    .A2(_0252_),
    .ZN(_0253_)
  );
  OR2_X1 _1040_ (
    .A1(_0251_),
    .A2(_0253_),
    .ZN(_0254_)
  );
  AND2_X1 _1041_ (
    .A1(io_fn[0]),
    .A2(_0254_),
    .ZN(_0255_)
  );
  INV_X1 _1042_ (
    .A(_0255_),
    .ZN(_0256_)
  );
  MUX2_X1 _1043_ (
    .A(io_in1[30]),
    .B(io_in1[1]),
    .S(_0255_),
    .Z(_0257_)
  );
  OR2_X1 _1044_ (
    .A1(_0004_),
    .A2(_0257_),
    .ZN(_0258_)
  );
  AND2_X1 _1045_ (
    .A1(io_in1[31]),
    .A2(_0256_),
    .ZN(_0259_)
  );
  AND2_X1 _1046_ (
    .A1(io_in1[0]),
    .A2(_0255_),
    .ZN(_0260_)
  );
  OR2_X1 _1047_ (
    .A1(io_in2[0]),
    .A2(_0260_),
    .ZN(_0261_)
  );
  OR2_X1 _1048_ (
    .A1(_0259_),
    .A2(_0261_),
    .ZN(_0262_)
  );
  AND2_X1 _1049_ (
    .A1(_0258_),
    .A2(_0262_),
    .ZN(_0263_)
  );
  MUX2_X1 _1050_ (
    .A(io_in1[29]),
    .B(io_in1[2]),
    .S(_0255_),
    .Z(_0264_)
  );
  MUX2_X1 _1051_ (
    .A(io_in1[28]),
    .B(io_in1[3]),
    .S(_0255_),
    .Z(_0265_)
  );
  MUX2_X1 _1052_ (
    .A(_0264_),
    .B(_0265_),
    .S(io_in2[0]),
    .Z(_0266_)
  );
  MUX2_X1 _1053_ (
    .A(_0263_),
    .B(_0266_),
    .S(io_in2[1]),
    .Z(_0267_)
  );
  MUX2_X1 _1054_ (
    .A(io_in1[27]),
    .B(io_in1[4]),
    .S(_0255_),
    .Z(_0268_)
  );
  MUX2_X1 _1055_ (
    .A(io_in1[26]),
    .B(io_in1[5]),
    .S(_0255_),
    .Z(_0269_)
  );
  MUX2_X1 _1056_ (
    .A(_0268_),
    .B(_0269_),
    .S(io_in2[0]),
    .Z(_0270_)
  );
  MUX2_X1 _1057_ (
    .A(io_in1[25]),
    .B(io_in1[6]),
    .S(_0255_),
    .Z(_0271_)
  );
  MUX2_X1 _1058_ (
    .A(io_in1[24]),
    .B(io_in1[7]),
    .S(_0255_),
    .Z(_0272_)
  );
  MUX2_X1 _1059_ (
    .A(_0271_),
    .B(_0272_),
    .S(io_in2[0]),
    .Z(_0273_)
  );
  MUX2_X1 _1060_ (
    .A(_0270_),
    .B(_0273_),
    .S(io_in2[1]),
    .Z(_0274_)
  );
  MUX2_X1 _1061_ (
    .A(_0267_),
    .B(_0274_),
    .S(io_in2[2]),
    .Z(_0275_)
  );
  MUX2_X1 _1062_ (
    .A(io_in1[23]),
    .B(io_in1[8]),
    .S(_0255_),
    .Z(_0276_)
  );
  MUX2_X1 _1063_ (
    .A(io_in1[22]),
    .B(io_in1[9]),
    .S(_0255_),
    .Z(_0277_)
  );
  MUX2_X1 _1064_ (
    .A(_0276_),
    .B(_0277_),
    .S(io_in2[0]),
    .Z(_0278_)
  );
  MUX2_X1 _1065_ (
    .A(io_in1[21]),
    .B(io_in1[10]),
    .S(_0255_),
    .Z(_0279_)
  );
  MUX2_X1 _1066_ (
    .A(io_in1[20]),
    .B(io_in1[11]),
    .S(_0255_),
    .Z(_0280_)
  );
  MUX2_X1 _1067_ (
    .A(_0279_),
    .B(_0280_),
    .S(io_in2[0]),
    .Z(_0281_)
  );
  MUX2_X1 _1068_ (
    .A(_0278_),
    .B(_0281_),
    .S(io_in2[1]),
    .Z(_0282_)
  );
  MUX2_X1 _1069_ (
    .A(io_in1[19]),
    .B(io_in1[12]),
    .S(_0255_),
    .Z(_0283_)
  );
  MUX2_X1 _1070_ (
    .A(io_in1[18]),
    .B(io_in1[13]),
    .S(_0255_),
    .Z(_0284_)
  );
  MUX2_X1 _1071_ (
    .A(_0283_),
    .B(_0284_),
    .S(io_in2[0]),
    .Z(_0285_)
  );
  MUX2_X1 _1072_ (
    .A(io_in1[17]),
    .B(io_in1[14]),
    .S(_0255_),
    .Z(_0286_)
  );
  MUX2_X1 _1073_ (
    .A(io_in1[16]),
    .B(io_in1[15]),
    .S(_0255_),
    .Z(_0287_)
  );
  MUX2_X1 _1074_ (
    .A(_0286_),
    .B(_0287_),
    .S(io_in2[0]),
    .Z(_0288_)
  );
  MUX2_X1 _1075_ (
    .A(_0285_),
    .B(_0288_),
    .S(io_in2[1]),
    .Z(_0289_)
  );
  MUX2_X1 _1076_ (
    .A(_0282_),
    .B(_0289_),
    .S(io_in2[2]),
    .Z(_0290_)
  );
  MUX2_X1 _1077_ (
    .A(_0275_),
    .B(_0290_),
    .S(io_in2[3]),
    .Z(_0291_)
  );
  MUX2_X1 _1078_ (
    .A(io_in1[15]),
    .B(io_in1[16]),
    .S(_0255_),
    .Z(_0292_)
  );
  MUX2_X1 _1079_ (
    .A(io_in1[14]),
    .B(io_in1[17]),
    .S(_0255_),
    .Z(_0293_)
  );
  MUX2_X1 _1080_ (
    .A(_0292_),
    .B(_0293_),
    .S(io_in2[0]),
    .Z(_0294_)
  );
  MUX2_X1 _1081_ (
    .A(io_in1[13]),
    .B(io_in1[18]),
    .S(_0255_),
    .Z(_0295_)
  );
  MUX2_X1 _1082_ (
    .A(io_in1[12]),
    .B(io_in1[19]),
    .S(_0255_),
    .Z(_0296_)
  );
  MUX2_X1 _1083_ (
    .A(_0295_),
    .B(_0296_),
    .S(io_in2[0]),
    .Z(_0297_)
  );
  MUX2_X1 _1084_ (
    .A(_0294_),
    .B(_0297_),
    .S(io_in2[1]),
    .Z(_0298_)
  );
  MUX2_X1 _1085_ (
    .A(io_in1[11]),
    .B(io_in1[20]),
    .S(_0255_),
    .Z(_0299_)
  );
  MUX2_X1 _1086_ (
    .A(io_in1[10]),
    .B(io_in1[21]),
    .S(_0255_),
    .Z(_0300_)
  );
  MUX2_X1 _1087_ (
    .A(_0299_),
    .B(_0300_),
    .S(io_in2[0]),
    .Z(_0301_)
  );
  MUX2_X1 _1088_ (
    .A(io_in1[9]),
    .B(io_in1[22]),
    .S(_0255_),
    .Z(_0302_)
  );
  MUX2_X1 _1089_ (
    .A(io_in1[8]),
    .B(io_in1[23]),
    .S(_0255_),
    .Z(_0303_)
  );
  MUX2_X1 _1090_ (
    .A(_0302_),
    .B(_0303_),
    .S(io_in2[0]),
    .Z(_0304_)
  );
  MUX2_X1 _1091_ (
    .A(_0301_),
    .B(_0304_),
    .S(io_in2[1]),
    .Z(_0305_)
  );
  MUX2_X1 _1092_ (
    .A(_0298_),
    .B(_0305_),
    .S(io_in2[2]),
    .Z(_0306_)
  );
  MUX2_X1 _1093_ (
    .A(io_in1[7]),
    .B(io_in1[24]),
    .S(_0255_),
    .Z(_0307_)
  );
  MUX2_X1 _1094_ (
    .A(io_in1[6]),
    .B(io_in1[25]),
    .S(_0255_),
    .Z(_0308_)
  );
  MUX2_X1 _1095_ (
    .A(_0307_),
    .B(_0308_),
    .S(io_in2[0]),
    .Z(_0309_)
  );
  MUX2_X1 _1096_ (
    .A(io_in1[5]),
    .B(io_in1[26]),
    .S(_0255_),
    .Z(_0310_)
  );
  MUX2_X1 _1097_ (
    .A(io_in1[4]),
    .B(io_in1[27]),
    .S(_0255_),
    .Z(_0311_)
  );
  MUX2_X1 _1098_ (
    .A(_0310_),
    .B(_0311_),
    .S(io_in2[0]),
    .Z(_0312_)
  );
  MUX2_X1 _1099_ (
    .A(_0309_),
    .B(_0312_),
    .S(io_in2[1]),
    .Z(_0313_)
  );
  MUX2_X1 _1100_ (
    .A(io_in1[3]),
    .B(io_in1[28]),
    .S(_0255_),
    .Z(_0314_)
  );
  MUX2_X1 _1101_ (
    .A(io_in1[2]),
    .B(io_in1[29]),
    .S(_0255_),
    .Z(_0315_)
  );
  MUX2_X1 _1102_ (
    .A(_0314_),
    .B(_0315_),
    .S(io_in2[0]),
    .Z(_0316_)
  );
  MUX2_X1 _1103_ (
    .A(io_in1[1]),
    .B(io_in1[30]),
    .S(_0255_),
    .Z(_0317_)
  );
  MUX2_X1 _1104_ (
    .A(io_in1[0]),
    .B(io_in1[31]),
    .S(_0255_),
    .Z(_0318_)
  );
  MUX2_X1 _1105_ (
    .A(_0317_),
    .B(_0318_),
    .S(io_in2[0]),
    .Z(_0319_)
  );
  MUX2_X1 _1106_ (
    .A(_0316_),
    .B(_0319_),
    .S(io_in2[1]),
    .Z(_0320_)
  );
  MUX2_X1 _1107_ (
    .A(_0313_),
    .B(_0320_),
    .S(io_in2[2]),
    .Z(_0321_)
  );
  MUX2_X1 _1108_ (
    .A(_0306_),
    .B(_0321_),
    .S(io_in2[3]),
    .Z(_0322_)
  );
  MUX2_X1 _1109_ (
    .A(_0291_),
    .B(_0322_),
    .S(io_in2[4]),
    .Z(_0323_)
  );
  AND2_X1 _1110_ (
    .A1(_0255_),
    .A2(_0323_),
    .ZN(_0324_)
  );
  AND2_X1 _1111_ (
    .A1(_0070_),
    .A2(_0318_),
    .ZN(_0325_)
  );
  AND2_X1 _1112_ (
    .A1(_0067_),
    .A2(_0325_),
    .ZN(_0326_)
  );
  AND2_X1 _1113_ (
    .A1(io_fn[3]),
    .A2(_0318_),
    .ZN(_0327_)
  );
  MUX2_X1 _1114_ (
    .A(_0326_),
    .B(_0327_),
    .S(io_in2[2]),
    .Z(_0328_)
  );
  MUX2_X1 _1115_ (
    .A(_0328_),
    .B(_0327_),
    .S(io_in2[3]),
    .Z(_0329_)
  );
  MUX2_X1 _1116_ (
    .A(_0329_),
    .B(_0327_),
    .S(io_in2[4]),
    .Z(_0330_)
  );
  AND2_X1 _1117_ (
    .A1(_0000_),
    .A2(_0002_),
    .ZN(_0331_)
  );
  AND2_X1 _1118_ (
    .A1(_0003_),
    .A2(_0331_),
    .ZN(_0332_)
  );
  AND2_X1 _1119_ (
    .A1(io_fn[0]),
    .A2(_0332_),
    .ZN(_0333_)
  );
  AND2_X1 _1120_ (
    .A1(_0330_),
    .A2(_0333_),
    .ZN(_0334_)
  );
  OR2_X1 _1121_ (
    .A1(_0251_),
    .A2(_0332_),
    .ZN(_0335_)
  );
  AND2_X1 _1122_ (
    .A1(_0001_),
    .A2(_0335_),
    .ZN(_0336_)
  );
  AND2_X1 _1123_ (
    .A1(io_adder_out[0]),
    .A2(_0336_),
    .ZN(_0337_)
  );
  AND2_X1 _1124_ (
    .A1(io_fn[1]),
    .A2(_0252_),
    .ZN(_0338_)
  );
  AND2_X1 _1125_ (
    .A1(io_in2[0]),
    .A2(io_in1[0]),
    .ZN(_0339_)
  );
  AND2_X1 _1126_ (
    .A1(_0338_),
    .A2(_0339_),
    .ZN(_0340_)
  );
  AND2_X1 _1127_ (
    .A1(_0001_),
    .A2(_0252_),
    .ZN(_0341_)
  );
  AND2_X1 _1128_ (
    .A1(_0134_),
    .A2(_0341_),
    .ZN(_0342_)
  );
  OR2_X1 _1129_ (
    .A1(_0340_),
    .A2(_0342_),
    .ZN(_0343_)
  );
  OR2_X1 _1130_ (
    .A1(_0337_),
    .A2(_0343_),
    .ZN(_0344_)
  );
  OR2_X1 _1131_ (
    .A1(_0334_),
    .A2(_0344_),
    .ZN(_0345_)
  );
  OR2_X1 _1132_ (
    .A1(_0324_),
    .A2(_0345_),
    .ZN(_0346_)
  );
  OR2_X1 _1133_ (
    .A1(_0250_),
    .A2(_0346_),
    .ZN(io_out[0])
  );
  XOR2_X1 _1134_ (
    .A(_0072_),
    .B(_0073_),
    .Z(_0347_)
  );
  MUX2_X1 _1135_ (
    .A(_0347_),
    .B(_0074_),
    .S(_0135_),
    .Z(io_adder_out[1])
  );
  MUX2_X1 _1136_ (
    .A(_0319_),
    .B(_0327_),
    .S(io_in2[1]),
    .Z(_0348_)
  );
  MUX2_X1 _1137_ (
    .A(_0348_),
    .B(_0327_),
    .S(io_in2[2]),
    .Z(_0349_)
  );
  MUX2_X1 _1138_ (
    .A(_0349_),
    .B(_0327_),
    .S(io_in2[3]),
    .Z(_0350_)
  );
  MUX2_X1 _1139_ (
    .A(_0350_),
    .B(_0327_),
    .S(io_in2[4]),
    .Z(_0351_)
  );
  AND2_X1 _1140_ (
    .A1(_0333_),
    .A2(_0351_),
    .ZN(_0352_)
  );
  MUX2_X1 _1141_ (
    .A(_0257_),
    .B(_0264_),
    .S(io_in2[0]),
    .Z(_0353_)
  );
  MUX2_X1 _1142_ (
    .A(_0265_),
    .B(_0268_),
    .S(io_in2[0]),
    .Z(_0354_)
  );
  MUX2_X1 _1143_ (
    .A(_0353_),
    .B(_0354_),
    .S(io_in2[1]),
    .Z(_0355_)
  );
  MUX2_X1 _1144_ (
    .A(_0269_),
    .B(_0271_),
    .S(io_in2[0]),
    .Z(_0356_)
  );
  MUX2_X1 _1145_ (
    .A(_0272_),
    .B(_0276_),
    .S(io_in2[0]),
    .Z(_0357_)
  );
  MUX2_X1 _1146_ (
    .A(_0356_),
    .B(_0357_),
    .S(io_in2[1]),
    .Z(_0358_)
  );
  MUX2_X1 _1147_ (
    .A(_0355_),
    .B(_0358_),
    .S(io_in2[2]),
    .Z(_0359_)
  );
  MUX2_X1 _1148_ (
    .A(_0277_),
    .B(_0279_),
    .S(io_in2[0]),
    .Z(_0360_)
  );
  MUX2_X1 _1149_ (
    .A(_0280_),
    .B(_0283_),
    .S(io_in2[0]),
    .Z(_0361_)
  );
  MUX2_X1 _1150_ (
    .A(_0360_),
    .B(_0361_),
    .S(io_in2[1]),
    .Z(_0362_)
  );
  MUX2_X1 _1151_ (
    .A(_0284_),
    .B(_0286_),
    .S(io_in2[0]),
    .Z(_0363_)
  );
  MUX2_X1 _1152_ (
    .A(_0287_),
    .B(_0292_),
    .S(io_in2[0]),
    .Z(_0364_)
  );
  MUX2_X1 _1153_ (
    .A(_0363_),
    .B(_0364_),
    .S(io_in2[1]),
    .Z(_0365_)
  );
  MUX2_X1 _1154_ (
    .A(_0362_),
    .B(_0365_),
    .S(io_in2[2]),
    .Z(_0366_)
  );
  MUX2_X1 _1155_ (
    .A(_0359_),
    .B(_0366_),
    .S(io_in2[3]),
    .Z(_0367_)
  );
  MUX2_X1 _1156_ (
    .A(_0293_),
    .B(_0295_),
    .S(io_in2[0]),
    .Z(_0368_)
  );
  MUX2_X1 _1157_ (
    .A(_0296_),
    .B(_0299_),
    .S(io_in2[0]),
    .Z(_0369_)
  );
  MUX2_X1 _1158_ (
    .A(_0368_),
    .B(_0369_),
    .S(io_in2[1]),
    .Z(_0370_)
  );
  MUX2_X1 _1159_ (
    .A(_0300_),
    .B(_0302_),
    .S(io_in2[0]),
    .Z(_0371_)
  );
  MUX2_X1 _1160_ (
    .A(_0303_),
    .B(_0307_),
    .S(io_in2[0]),
    .Z(_0372_)
  );
  MUX2_X1 _1161_ (
    .A(_0371_),
    .B(_0372_),
    .S(io_in2[1]),
    .Z(_0373_)
  );
  MUX2_X1 _1162_ (
    .A(_0370_),
    .B(_0373_),
    .S(io_in2[2]),
    .Z(_0374_)
  );
  MUX2_X1 _1163_ (
    .A(_0308_),
    .B(_0310_),
    .S(io_in2[0]),
    .Z(_0375_)
  );
  MUX2_X1 _1164_ (
    .A(_0311_),
    .B(_0314_),
    .S(io_in2[0]),
    .Z(_0376_)
  );
  MUX2_X1 _1165_ (
    .A(_0375_),
    .B(_0376_),
    .S(io_in2[1]),
    .Z(_0377_)
  );
  MUX2_X1 _1166_ (
    .A(_0315_),
    .B(_0317_),
    .S(io_in2[0]),
    .Z(_0378_)
  );
  MUX2_X1 _1167_ (
    .A(_0325_),
    .B(_0378_),
    .S(_0005_),
    .Z(_0379_)
  );
  MUX2_X1 _1168_ (
    .A(_0377_),
    .B(_0379_),
    .S(io_in2[2]),
    .Z(_0380_)
  );
  MUX2_X1 _1169_ (
    .A(_0374_),
    .B(_0380_),
    .S(io_in2[3]),
    .Z(_0381_)
  );
  MUX2_X1 _1170_ (
    .A(_0367_),
    .B(_0381_),
    .S(io_in2[4]),
    .Z(_0382_)
  );
  AND2_X1 _1171_ (
    .A1(_0255_),
    .A2(_0382_),
    .ZN(_0383_)
  );
  AND2_X1 _1172_ (
    .A1(_0336_),
    .A2(io_adder_out[1]),
    .ZN(_0384_)
  );
  AND2_X1 _1173_ (
    .A1(_0073_),
    .A2(_0341_),
    .ZN(_0385_)
  );
  AND2_X1 _1174_ (
    .A1(io_in2[1]),
    .A2(io_in1[1]),
    .ZN(_0386_)
  );
  AND2_X1 _1175_ (
    .A1(_0338_),
    .A2(_0386_),
    .ZN(_0387_)
  );
  OR2_X1 _1176_ (
    .A1(_0385_),
    .A2(_0387_),
    .ZN(_0388_)
  );
  OR2_X1 _1177_ (
    .A1(_0384_),
    .A2(_0388_),
    .ZN(_0389_)
  );
  OR2_X1 _1178_ (
    .A1(_0383_),
    .A2(_0389_),
    .ZN(_0390_)
  );
  OR2_X1 _1179_ (
    .A1(_0352_),
    .A2(_0390_),
    .ZN(io_out[1])
  );
  XOR2_X1 _1180_ (
    .A(_0136_),
    .B(_0137_),
    .Z(io_adder_out[2])
  );
  MUX2_X1 _1181_ (
    .A(_0379_),
    .B(_0327_),
    .S(io_in2[2]),
    .Z(_0391_)
  );
  MUX2_X1 _1182_ (
    .A(_0391_),
    .B(_0327_),
    .S(io_in2[3]),
    .Z(_0392_)
  );
  MUX2_X1 _1183_ (
    .A(_0392_),
    .B(_0327_),
    .S(io_in2[4]),
    .Z(_0393_)
  );
  AND2_X1 _1184_ (
    .A1(_0333_),
    .A2(_0393_),
    .ZN(_0394_)
  );
  MUX2_X1 _1185_ (
    .A(_0266_),
    .B(_0270_),
    .S(io_in2[1]),
    .Z(_0395_)
  );
  MUX2_X1 _1186_ (
    .A(_0273_),
    .B(_0278_),
    .S(io_in2[1]),
    .Z(_0396_)
  );
  MUX2_X1 _1187_ (
    .A(_0395_),
    .B(_0396_),
    .S(io_in2[2]),
    .Z(_0397_)
  );
  MUX2_X1 _1188_ (
    .A(_0281_),
    .B(_0285_),
    .S(io_in2[1]),
    .Z(_0398_)
  );
  MUX2_X1 _1189_ (
    .A(_0288_),
    .B(_0294_),
    .S(io_in2[1]),
    .Z(_0399_)
  );
  MUX2_X1 _1190_ (
    .A(_0398_),
    .B(_0399_),
    .S(io_in2[2]),
    .Z(_0400_)
  );
  MUX2_X1 _1191_ (
    .A(_0397_),
    .B(_0400_),
    .S(io_in2[3]),
    .Z(_0401_)
  );
  MUX2_X1 _1192_ (
    .A(_0297_),
    .B(_0301_),
    .S(io_in2[1]),
    .Z(_0402_)
  );
  MUX2_X1 _1193_ (
    .A(_0304_),
    .B(_0309_),
    .S(io_in2[1]),
    .Z(_0403_)
  );
  MUX2_X1 _1194_ (
    .A(_0402_),
    .B(_0403_),
    .S(io_in2[2]),
    .Z(_0404_)
  );
  MUX2_X1 _1195_ (
    .A(_0312_),
    .B(_0316_),
    .S(io_in2[1]),
    .Z(_0405_)
  );
  MUX2_X1 _1196_ (
    .A(_0405_),
    .B(_0348_),
    .S(io_in2[2]),
    .Z(_0406_)
  );
  MUX2_X1 _1197_ (
    .A(_0404_),
    .B(_0406_),
    .S(io_in2[3]),
    .Z(_0407_)
  );
  MUX2_X1 _1198_ (
    .A(_0401_),
    .B(_0407_),
    .S(io_in2[4]),
    .Z(_0408_)
  );
  AND2_X1 _1199_ (
    .A1(_0255_),
    .A2(_0408_),
    .ZN(_0409_)
  );
  AND2_X1 _1200_ (
    .A1(_0336_),
    .A2(io_adder_out[2]),
    .ZN(_0410_)
  );
  AND2_X1 _1201_ (
    .A1(_0077_),
    .A2(_0341_),
    .ZN(_0411_)
  );
  AND2_X1 _1202_ (
    .A1(io_in2[2]),
    .A2(io_in1[2]),
    .ZN(_0412_)
  );
  AND2_X1 _1203_ (
    .A1(_0338_),
    .A2(_0412_),
    .ZN(_0413_)
  );
  OR2_X1 _1204_ (
    .A1(_0411_),
    .A2(_0413_),
    .ZN(_0414_)
  );
  OR2_X1 _1205_ (
    .A1(_0410_),
    .A2(_0414_),
    .ZN(_0415_)
  );
  OR2_X1 _1206_ (
    .A1(_0409_),
    .A2(_0415_),
    .ZN(_0416_)
  );
  OR2_X1 _1207_ (
    .A1(_0394_),
    .A2(_0416_),
    .ZN(io_out[2])
  );
  XOR2_X1 _1208_ (
    .A(_0138_),
    .B(_0139_),
    .Z(io_adder_out[3])
  );
  MUX2_X1 _1209_ (
    .A(_0320_),
    .B(_0327_),
    .S(io_in2[2]),
    .Z(_0417_)
  );
  MUX2_X1 _1210_ (
    .A(_0417_),
    .B(_0327_),
    .S(io_in2[3]),
    .Z(_0418_)
  );
  MUX2_X1 _1211_ (
    .A(_0418_),
    .B(_0327_),
    .S(io_in2[4]),
    .Z(_0419_)
  );
  AND2_X1 _1212_ (
    .A1(_0333_),
    .A2(_0419_),
    .ZN(_0420_)
  );
  MUX2_X1 _1213_ (
    .A(_0354_),
    .B(_0356_),
    .S(io_in2[1]),
    .Z(_0421_)
  );
  MUX2_X1 _1214_ (
    .A(_0357_),
    .B(_0360_),
    .S(io_in2[1]),
    .Z(_0422_)
  );
  MUX2_X1 _1215_ (
    .A(_0421_),
    .B(_0422_),
    .S(io_in2[2]),
    .Z(_0423_)
  );
  MUX2_X1 _1216_ (
    .A(_0361_),
    .B(_0363_),
    .S(io_in2[1]),
    .Z(_0424_)
  );
  MUX2_X1 _1217_ (
    .A(_0364_),
    .B(_0368_),
    .S(io_in2[1]),
    .Z(_0425_)
  );
  MUX2_X1 _1218_ (
    .A(_0424_),
    .B(_0425_),
    .S(io_in2[2]),
    .Z(_0426_)
  );
  MUX2_X1 _1219_ (
    .A(_0423_),
    .B(_0426_),
    .S(io_in2[3]),
    .Z(_0427_)
  );
  MUX2_X1 _1220_ (
    .A(_0369_),
    .B(_0371_),
    .S(io_in2[1]),
    .Z(_0428_)
  );
  MUX2_X1 _1221_ (
    .A(_0372_),
    .B(_0375_),
    .S(io_in2[1]),
    .Z(_0429_)
  );
  MUX2_X1 _1222_ (
    .A(_0428_),
    .B(_0429_),
    .S(io_in2[2]),
    .Z(_0430_)
  );
  MUX2_X1 _1223_ (
    .A(_0376_),
    .B(_0378_),
    .S(io_in2[1]),
    .Z(_0431_)
  );
  MUX2_X1 _1224_ (
    .A(_0431_),
    .B(_0326_),
    .S(io_in2[2]),
    .Z(_0432_)
  );
  MUX2_X1 _1225_ (
    .A(_0430_),
    .B(_0432_),
    .S(io_in2[3]),
    .Z(_0433_)
  );
  MUX2_X1 _1226_ (
    .A(_0427_),
    .B(_0433_),
    .S(io_in2[4]),
    .Z(_0434_)
  );
  AND2_X1 _1227_ (
    .A1(_0255_),
    .A2(_0434_),
    .ZN(_0435_)
  );
  AND2_X1 _1228_ (
    .A1(_0336_),
    .A2(io_adder_out[3]),
    .ZN(_0436_)
  );
  AND2_X1 _1229_ (
    .A1(_0080_),
    .A2(_0341_),
    .ZN(_0437_)
  );
  AND2_X1 _1230_ (
    .A1(io_in2[3]),
    .A2(io_in1[3]),
    .ZN(_0438_)
  );
  AND2_X1 _1231_ (
    .A1(_0338_),
    .A2(_0438_),
    .ZN(_0439_)
  );
  OR2_X1 _1232_ (
    .A1(_0437_),
    .A2(_0439_),
    .ZN(_0440_)
  );
  OR2_X1 _1233_ (
    .A1(_0436_),
    .A2(_0440_),
    .ZN(_0441_)
  );
  OR2_X1 _1234_ (
    .A1(_0435_),
    .A2(_0441_),
    .ZN(_0442_)
  );
  OR2_X1 _1235_ (
    .A1(_0420_),
    .A2(_0442_),
    .ZN(io_out[3])
  );
  XOR2_X1 _1236_ (
    .A(_0140_),
    .B(_0141_),
    .Z(io_adder_out[4])
  );
  MUX2_X1 _1237_ (
    .A(_0432_),
    .B(_0327_),
    .S(io_in2[3]),
    .Z(_0443_)
  );
  MUX2_X1 _1238_ (
    .A(_0443_),
    .B(_0327_),
    .S(io_in2[4]),
    .Z(_0444_)
  );
  AND2_X1 _1239_ (
    .A1(_0333_),
    .A2(_0444_),
    .ZN(_0445_)
  );
  MUX2_X1 _1240_ (
    .A(_0274_),
    .B(_0282_),
    .S(io_in2[2]),
    .Z(_0446_)
  );
  MUX2_X1 _1241_ (
    .A(_0289_),
    .B(_0298_),
    .S(io_in2[2]),
    .Z(_0447_)
  );
  MUX2_X1 _1242_ (
    .A(_0446_),
    .B(_0447_),
    .S(io_in2[3]),
    .Z(_0448_)
  );
  MUX2_X1 _1243_ (
    .A(_0305_),
    .B(_0313_),
    .S(io_in2[2]),
    .Z(_0449_)
  );
  MUX2_X1 _1244_ (
    .A(_0449_),
    .B(_0417_),
    .S(io_in2[3]),
    .Z(_0450_)
  );
  MUX2_X1 _1245_ (
    .A(_0448_),
    .B(_0450_),
    .S(io_in2[4]),
    .Z(_0451_)
  );
  AND2_X1 _1246_ (
    .A1(_0255_),
    .A2(_0451_),
    .ZN(_0452_)
  );
  AND2_X1 _1247_ (
    .A1(_0336_),
    .A2(io_adder_out[4]),
    .ZN(_0453_)
  );
  AND2_X1 _1248_ (
    .A1(_0083_),
    .A2(_0341_),
    .ZN(_0454_)
  );
  AND2_X1 _1249_ (
    .A1(io_in2[4]),
    .A2(io_in1[4]),
    .ZN(_0455_)
  );
  AND2_X1 _1250_ (
    .A1(_0338_),
    .A2(_0455_),
    .ZN(_0456_)
  );
  OR2_X1 _1251_ (
    .A1(_0454_),
    .A2(_0456_),
    .ZN(_0457_)
  );
  OR2_X1 _1252_ (
    .A1(_0453_),
    .A2(_0457_),
    .ZN(_0458_)
  );
  OR2_X1 _1253_ (
    .A1(_0452_),
    .A2(_0458_),
    .ZN(_0459_)
  );
  OR2_X1 _1254_ (
    .A1(_0445_),
    .A2(_0459_),
    .ZN(io_out[4])
  );
  XOR2_X1 _1255_ (
    .A(_0142_),
    .B(_0143_),
    .Z(io_adder_out[5])
  );
  MUX2_X1 _1256_ (
    .A(_0406_),
    .B(_0327_),
    .S(io_in2[3]),
    .Z(_0460_)
  );
  MUX2_X1 _1257_ (
    .A(_0460_),
    .B(_0327_),
    .S(io_in2[4]),
    .Z(_0461_)
  );
  AND2_X1 _1258_ (
    .A1(_0333_),
    .A2(_0461_),
    .ZN(_0462_)
  );
  AND2_X1 _1259_ (
    .A1(io_in2[5]),
    .A2(io_in1[5]),
    .ZN(_0463_)
  );
  AND2_X1 _1260_ (
    .A1(_0338_),
    .A2(_0463_),
    .ZN(_0464_)
  );
  AND2_X1 _1261_ (
    .A1(_0086_),
    .A2(_0341_),
    .ZN(_0465_)
  );
  OR2_X1 _1262_ (
    .A1(_0464_),
    .A2(_0465_),
    .ZN(_0466_)
  );
  OR2_X1 _1263_ (
    .A1(_0462_),
    .A2(_0466_),
    .ZN(_0467_)
  );
  AND2_X1 _1264_ (
    .A1(_0336_),
    .A2(io_adder_out[5]),
    .ZN(_0468_)
  );
  MUX2_X1 _1265_ (
    .A(_0358_),
    .B(_0362_),
    .S(io_in2[2]),
    .Z(_0469_)
  );
  MUX2_X1 _1266_ (
    .A(_0365_),
    .B(_0370_),
    .S(io_in2[2]),
    .Z(_0470_)
  );
  MUX2_X1 _1267_ (
    .A(_0469_),
    .B(_0470_),
    .S(io_in2[3]),
    .Z(_0471_)
  );
  MUX2_X1 _1268_ (
    .A(_0373_),
    .B(_0377_),
    .S(io_in2[2]),
    .Z(_0472_)
  );
  MUX2_X1 _1269_ (
    .A(_0472_),
    .B(_0391_),
    .S(io_in2[3]),
    .Z(_0473_)
  );
  MUX2_X1 _1270_ (
    .A(_0471_),
    .B(_0473_),
    .S(io_in2[4]),
    .Z(_0474_)
  );
  AND2_X1 _1271_ (
    .A1(_0255_),
    .A2(_0474_),
    .ZN(_0475_)
  );
  OR2_X1 _1272_ (
    .A1(_0468_),
    .A2(_0475_),
    .ZN(_0476_)
  );
  OR2_X1 _1273_ (
    .A1(_0467_),
    .A2(_0476_),
    .ZN(io_out[5])
  );
  XOR2_X1 _1274_ (
    .A(_0144_),
    .B(_0145_),
    .Z(io_adder_out[6])
  );
  AND2_X1 _1275_ (
    .A1(_0336_),
    .A2(io_adder_out[6]),
    .ZN(_0477_)
  );
  MUX2_X1 _1276_ (
    .A(_0396_),
    .B(_0398_),
    .S(io_in2[2]),
    .Z(_0478_)
  );
  MUX2_X1 _1277_ (
    .A(_0399_),
    .B(_0402_),
    .S(io_in2[2]),
    .Z(_0479_)
  );
  MUX2_X1 _1278_ (
    .A(_0478_),
    .B(_0479_),
    .S(io_in2[3]),
    .Z(_0480_)
  );
  MUX2_X1 _1279_ (
    .A(_0403_),
    .B(_0405_),
    .S(io_in2[2]),
    .Z(_0481_)
  );
  MUX2_X1 _1280_ (
    .A(_0481_),
    .B(_0349_),
    .S(io_in2[3]),
    .Z(_0482_)
  );
  MUX2_X1 _1281_ (
    .A(_0480_),
    .B(_0482_),
    .S(io_in2[4]),
    .Z(_0483_)
  );
  AND2_X1 _1282_ (
    .A1(_0255_),
    .A2(_0483_),
    .ZN(_0484_)
  );
  MUX2_X1 _1283_ (
    .A(_0380_),
    .B(_0327_),
    .S(io_in2[3]),
    .Z(_0485_)
  );
  MUX2_X1 _1284_ (
    .A(_0485_),
    .B(_0327_),
    .S(io_in2[4]),
    .Z(_0486_)
  );
  AND2_X1 _1285_ (
    .A1(_0333_),
    .A2(_0486_),
    .ZN(_0487_)
  );
  AND2_X1 _1286_ (
    .A1(io_in2[6]),
    .A2(io_in1[6]),
    .ZN(_0488_)
  );
  AND2_X1 _1287_ (
    .A1(_0338_),
    .A2(_0488_),
    .ZN(_0489_)
  );
  AND2_X1 _1288_ (
    .A1(_0058_),
    .A2(_0341_),
    .ZN(_0490_)
  );
  OR2_X1 _1289_ (
    .A1(_0489_),
    .A2(_0490_),
    .ZN(_0491_)
  );
  OR2_X1 _1290_ (
    .A1(_0487_),
    .A2(_0491_),
    .ZN(_0492_)
  );
  OR2_X1 _1291_ (
    .A1(_0484_),
    .A2(_0492_),
    .ZN(_0493_)
  );
  OR2_X1 _1292_ (
    .A1(_0477_),
    .A2(_0493_),
    .ZN(io_out[6])
  );
  XOR2_X1 _1293_ (
    .A(_0146_),
    .B(_0147_),
    .Z(io_adder_out[7])
  );
  AND2_X1 _1294_ (
    .A1(_0336_),
    .A2(io_adder_out[7]),
    .ZN(_0494_)
  );
  MUX2_X1 _1295_ (
    .A(_0422_),
    .B(_0424_),
    .S(io_in2[2]),
    .Z(_0495_)
  );
  MUX2_X1 _1296_ (
    .A(_0425_),
    .B(_0428_),
    .S(io_in2[2]),
    .Z(_0496_)
  );
  MUX2_X1 _1297_ (
    .A(_0495_),
    .B(_0496_),
    .S(io_in2[3]),
    .Z(_0497_)
  );
  MUX2_X1 _1298_ (
    .A(_0429_),
    .B(_0431_),
    .S(io_in2[2]),
    .Z(_0498_)
  );
  MUX2_X1 _1299_ (
    .A(_0498_),
    .B(_0328_),
    .S(io_in2[3]),
    .Z(_0499_)
  );
  MUX2_X1 _1300_ (
    .A(_0497_),
    .B(_0499_),
    .S(io_in2[4]),
    .Z(_0500_)
  );
  AND2_X1 _1301_ (
    .A1(_0255_),
    .A2(_0500_),
    .ZN(_0501_)
  );
  MUX2_X1 _1302_ (
    .A(_0321_),
    .B(_0327_),
    .S(io_in2[3]),
    .Z(_0502_)
  );
  MUX2_X1 _1303_ (
    .A(_0502_),
    .B(_0327_),
    .S(io_in2[4]),
    .Z(_0503_)
  );
  AND2_X1 _1304_ (
    .A1(_0333_),
    .A2(_0503_),
    .ZN(_0504_)
  );
  AND2_X1 _1305_ (
    .A1(_0055_),
    .A2(_0341_),
    .ZN(_0505_)
  );
  AND2_X1 _1306_ (
    .A1(io_in2[7]),
    .A2(io_in1[7]),
    .ZN(_0506_)
  );
  AND2_X1 _1307_ (
    .A1(_0338_),
    .A2(_0506_),
    .ZN(_0507_)
  );
  OR2_X1 _1308_ (
    .A1(_0505_),
    .A2(_0507_),
    .ZN(_0508_)
  );
  OR2_X1 _1309_ (
    .A1(_0504_),
    .A2(_0508_),
    .ZN(_0509_)
  );
  OR2_X1 _1310_ (
    .A1(_0501_),
    .A2(_0509_),
    .ZN(_0510_)
  );
  OR2_X1 _1311_ (
    .A1(_0494_),
    .A2(_0510_),
    .ZN(io_out[7])
  );
  XOR2_X1 _1312_ (
    .A(_0133_),
    .B(_0148_),
    .Z(io_adder_out[8])
  );
  AND2_X1 _1313_ (
    .A1(_0336_),
    .A2(io_adder_out[8]),
    .ZN(_0511_)
  );
  MUX2_X1 _1314_ (
    .A(_0499_),
    .B(_0327_),
    .S(io_in2[4]),
    .Z(_0512_)
  );
  AND2_X1 _1315_ (
    .A1(_0333_),
    .A2(_0512_),
    .ZN(_0513_)
  );
  MUX2_X1 _1316_ (
    .A(_0290_),
    .B(_0306_),
    .S(io_in2[3]),
    .Z(_0514_)
  );
  MUX2_X1 _1317_ (
    .A(_0514_),
    .B(_0502_),
    .S(io_in2[4]),
    .Z(_0515_)
  );
  AND2_X1 _1318_ (
    .A1(_0255_),
    .A2(_0515_),
    .ZN(_0516_)
  );
  AND2_X1 _1319_ (
    .A1(_0093_),
    .A2(_0341_),
    .ZN(_0517_)
  );
  AND2_X1 _1320_ (
    .A1(io_in2[8]),
    .A2(io_in1[8]),
    .ZN(_0518_)
  );
  AND2_X1 _1321_ (
    .A1(_0338_),
    .A2(_0518_),
    .ZN(_0519_)
  );
  OR2_X1 _1322_ (
    .A1(_0513_),
    .A2(_0517_),
    .ZN(_0520_)
  );
  OR2_X1 _1323_ (
    .A1(_0516_),
    .A2(_0519_),
    .ZN(_0521_)
  );
  OR2_X1 _1324_ (
    .A1(_0520_),
    .A2(_0521_),
    .ZN(_0522_)
  );
  OR2_X1 _1325_ (
    .A1(_0511_),
    .A2(_0522_),
    .ZN(io_out[8])
  );
  XOR2_X1 _1326_ (
    .A(_0149_),
    .B(_0150_),
    .Z(io_adder_out[9])
  );
  AND2_X1 _1327_ (
    .A1(_0336_),
    .A2(io_adder_out[9]),
    .ZN(_0523_)
  );
  MUX2_X1 _1328_ (
    .A(_0482_),
    .B(_0327_),
    .S(io_in2[4]),
    .Z(_0524_)
  );
  AND2_X1 _1329_ (
    .A1(_0333_),
    .A2(_0524_),
    .ZN(_0525_)
  );
  MUX2_X1 _1330_ (
    .A(_0366_),
    .B(_0374_),
    .S(io_in2[3]),
    .Z(_0526_)
  );
  MUX2_X1 _1331_ (
    .A(_0526_),
    .B(_0485_),
    .S(io_in2[4]),
    .Z(_0527_)
  );
  AND2_X1 _1332_ (
    .A1(_0255_),
    .A2(_0527_),
    .ZN(_0528_)
  );
  AND2_X1 _1333_ (
    .A1(_0050_),
    .A2(_0341_),
    .ZN(_0529_)
  );
  AND2_X1 _1334_ (
    .A1(io_in2[9]),
    .A2(io_in1[9]),
    .ZN(_0530_)
  );
  AND2_X1 _1335_ (
    .A1(_0338_),
    .A2(_0530_),
    .ZN(_0531_)
  );
  OR2_X1 _1336_ (
    .A1(_0529_),
    .A2(_0531_),
    .ZN(_0532_)
  );
  OR2_X1 _1337_ (
    .A1(_0528_),
    .A2(_0532_),
    .ZN(_0533_)
  );
  OR2_X1 _1338_ (
    .A1(_0525_),
    .A2(_0533_),
    .ZN(_0534_)
  );
  OR2_X1 _1339_ (
    .A1(_0523_),
    .A2(_0534_),
    .ZN(io_out[9])
  );
  XOR2_X1 _1340_ (
    .A(_0151_),
    .B(_0152_),
    .Z(io_adder_out[10])
  );
  AND2_X1 _1341_ (
    .A1(_0336_),
    .A2(io_adder_out[10]),
    .ZN(_0535_)
  );
  MUX2_X1 _1342_ (
    .A(_0400_),
    .B(_0404_),
    .S(io_in2[3]),
    .Z(_0536_)
  );
  MUX2_X1 _1343_ (
    .A(_0536_),
    .B(_0460_),
    .S(io_in2[4]),
    .Z(_0537_)
  );
  AND2_X1 _1344_ (
    .A1(_0255_),
    .A2(_0537_),
    .ZN(_0538_)
  );
  MUX2_X1 _1345_ (
    .A(_0473_),
    .B(_0327_),
    .S(io_in2[4]),
    .Z(_0539_)
  );
  AND2_X1 _1346_ (
    .A1(_0333_),
    .A2(_0539_),
    .ZN(_0540_)
  );
  AND2_X1 _1347_ (
    .A1(io_in2[10]),
    .A2(io_in1[10]),
    .ZN(_0541_)
  );
  AND2_X1 _1348_ (
    .A1(_0338_),
    .A2(_0541_),
    .ZN(_0542_)
  );
  AND2_X1 _1349_ (
    .A1(_0047_),
    .A2(_0341_),
    .ZN(_0543_)
  );
  OR2_X1 _1350_ (
    .A1(_0542_),
    .A2(_0543_),
    .ZN(_0544_)
  );
  OR2_X1 _1351_ (
    .A1(_0540_),
    .A2(_0544_),
    .ZN(_0545_)
  );
  OR2_X1 _1352_ (
    .A1(_0538_),
    .A2(_0545_),
    .ZN(_0546_)
  );
  OR2_X1 _1353_ (
    .A1(_0535_),
    .A2(_0546_),
    .ZN(io_out[10])
  );
  XOR2_X1 _1354_ (
    .A(_0153_),
    .B(_0155_),
    .Z(io_adder_out[11])
  );
  AND2_X1 _1355_ (
    .A1(_0336_),
    .A2(io_adder_out[11]),
    .ZN(_0547_)
  );
  MUX2_X1 _1356_ (
    .A(_0426_),
    .B(_0430_),
    .S(io_in2[3]),
    .Z(_0548_)
  );
  MUX2_X1 _1357_ (
    .A(_0548_),
    .B(_0443_),
    .S(io_in2[4]),
    .Z(_0549_)
  );
  AND2_X1 _1358_ (
    .A1(_0255_),
    .A2(_0549_),
    .ZN(_0550_)
  );
  AND2_X1 _1359_ (
    .A1(_0044_),
    .A2(_0341_),
    .ZN(_0551_)
  );
  AND2_X1 _1360_ (
    .A1(io_in2[11]),
    .A2(io_in1[11]),
    .ZN(_0552_)
  );
  AND2_X1 _1361_ (
    .A1(_0338_),
    .A2(_0552_),
    .ZN(_0553_)
  );
  OR2_X1 _1362_ (
    .A1(_0551_),
    .A2(_0553_),
    .ZN(_0554_)
  );
  OR2_X1 _1363_ (
    .A1(_0550_),
    .A2(_0554_),
    .ZN(_0555_)
  );
  MUX2_X1 _1364_ (
    .A(_0450_),
    .B(_0327_),
    .S(io_in2[4]),
    .Z(_0556_)
  );
  AND2_X1 _1365_ (
    .A1(_0333_),
    .A2(_0556_),
    .ZN(_0557_)
  );
  OR2_X1 _1366_ (
    .A1(_0555_),
    .A2(_0557_),
    .ZN(_0558_)
  );
  OR2_X1 _1367_ (
    .A1(_0547_),
    .A2(_0558_),
    .ZN(io_out[11])
  );
  XOR2_X1 _1368_ (
    .A(_0156_),
    .B(_0157_),
    .Z(io_adder_out[12])
  );
  AND2_X1 _1369_ (
    .A1(_0336_),
    .A2(io_adder_out[12]),
    .ZN(_0559_)
  );
  MUX2_X1 _1370_ (
    .A(_0447_),
    .B(_0449_),
    .S(io_in2[3]),
    .Z(_0560_)
  );
  MUX2_X1 _1371_ (
    .A(_0560_),
    .B(_0418_),
    .S(io_in2[4]),
    .Z(_0561_)
  );
  AND2_X1 _1372_ (
    .A1(_0255_),
    .A2(_0561_),
    .ZN(_0562_)
  );
  MUX2_X1 _1373_ (
    .A(_0433_),
    .B(_0327_),
    .S(io_in2[4]),
    .Z(_0563_)
  );
  AND2_X1 _1374_ (
    .A1(_0333_),
    .A2(_0563_),
    .ZN(_0564_)
  );
  AND2_X1 _1375_ (
    .A1(io_in2[12]),
    .A2(io_in1[12]),
    .ZN(_0565_)
  );
  AND2_X1 _1376_ (
    .A1(_0338_),
    .A2(_0565_),
    .ZN(_0566_)
  );
  AND2_X1 _1377_ (
    .A1(_0040_),
    .A2(_0341_),
    .ZN(_0567_)
  );
  OR2_X1 _1378_ (
    .A1(_0566_),
    .A2(_0567_),
    .ZN(_0568_)
  );
  OR2_X1 _1379_ (
    .A1(_0564_),
    .A2(_0568_),
    .ZN(_0569_)
  );
  OR2_X1 _1380_ (
    .A1(_0562_),
    .A2(_0569_),
    .ZN(_0570_)
  );
  OR2_X1 _1381_ (
    .A1(_0559_),
    .A2(_0570_),
    .ZN(io_out[12])
  );
  XOR2_X1 _1382_ (
    .A(_0158_),
    .B(_0160_),
    .Z(io_adder_out[13])
  );
  AND2_X1 _1383_ (
    .A1(_0336_),
    .A2(io_adder_out[13]),
    .ZN(_0571_)
  );
  MUX2_X1 _1384_ (
    .A(_0470_),
    .B(_0472_),
    .S(io_in2[3]),
    .Z(_0572_)
  );
  MUX2_X1 _1385_ (
    .A(_0572_),
    .B(_0392_),
    .S(io_in2[4]),
    .Z(_0573_)
  );
  AND2_X1 _1386_ (
    .A1(_0255_),
    .A2(_0573_),
    .ZN(_0574_)
  );
  AND2_X1 _1387_ (
    .A1(_0037_),
    .A2(_0341_),
    .ZN(_0575_)
  );
  AND2_X1 _1388_ (
    .A1(io_in2[13]),
    .A2(io_in1[13]),
    .ZN(_0576_)
  );
  AND2_X1 _1389_ (
    .A1(_0338_),
    .A2(_0576_),
    .ZN(_0577_)
  );
  OR2_X1 _1390_ (
    .A1(_0575_),
    .A2(_0577_),
    .ZN(_0578_)
  );
  OR2_X1 _1391_ (
    .A1(_0574_),
    .A2(_0578_),
    .ZN(_0579_)
  );
  MUX2_X1 _1392_ (
    .A(_0407_),
    .B(_0327_),
    .S(io_in2[4]),
    .Z(_0580_)
  );
  AND2_X1 _1393_ (
    .A1(_0333_),
    .A2(_0580_),
    .ZN(_0581_)
  );
  OR2_X1 _1394_ (
    .A1(_0579_),
    .A2(_0581_),
    .ZN(_0582_)
  );
  OR2_X1 _1395_ (
    .A1(_0571_),
    .A2(_0582_),
    .ZN(io_out[13])
  );
  XOR2_X1 _1396_ (
    .A(_0132_),
    .B(_0161_),
    .Z(io_adder_out[14])
  );
  AND2_X1 _1397_ (
    .A1(_0336_),
    .A2(io_adder_out[14]),
    .ZN(_0583_)
  );
  MUX2_X1 _1398_ (
    .A(_0479_),
    .B(_0481_),
    .S(io_in2[3]),
    .Z(_0584_)
  );
  MUX2_X1 _1399_ (
    .A(_0584_),
    .B(_0350_),
    .S(io_in2[4]),
    .Z(_0585_)
  );
  AND2_X1 _1400_ (
    .A1(_0255_),
    .A2(_0585_),
    .ZN(_0586_)
  );
  AND2_X1 _1401_ (
    .A1(_0033_),
    .A2(_0341_),
    .ZN(_0587_)
  );
  AND2_X1 _1402_ (
    .A1(io_in2[14]),
    .A2(io_in1[14]),
    .ZN(_0588_)
  );
  AND2_X1 _1403_ (
    .A1(_0338_),
    .A2(_0588_),
    .ZN(_0589_)
  );
  OR2_X1 _1404_ (
    .A1(_0587_),
    .A2(_0589_),
    .ZN(_0590_)
  );
  OR2_X1 _1405_ (
    .A1(_0586_),
    .A2(_0590_),
    .ZN(_0591_)
  );
  MUX2_X1 _1406_ (
    .A(_0381_),
    .B(_0327_),
    .S(io_in2[4]),
    .Z(_0592_)
  );
  AND2_X1 _1407_ (
    .A1(_0333_),
    .A2(_0592_),
    .ZN(_0593_)
  );
  OR2_X1 _1408_ (
    .A1(_0591_),
    .A2(_0593_),
    .ZN(_0594_)
  );
  OR2_X1 _1409_ (
    .A1(_0583_),
    .A2(_0594_),
    .ZN(io_out[14])
  );
  XOR2_X1 _1410_ (
    .A(_0162_),
    .B(_0164_),
    .Z(io_adder_out[15])
  );
  AND2_X1 _1411_ (
    .A1(_0336_),
    .A2(io_adder_out[15]),
    .ZN(_0595_)
  );
  MUX2_X1 _1412_ (
    .A(_0496_),
    .B(_0498_),
    .S(io_in2[3]),
    .Z(_0596_)
  );
  MUX2_X1 _1413_ (
    .A(_0596_),
    .B(_0329_),
    .S(io_in2[4]),
    .Z(_0597_)
  );
  AND2_X1 _1414_ (
    .A1(_0255_),
    .A2(_0597_),
    .ZN(_0598_)
  );
  MUX2_X1 _1415_ (
    .A(_0322_),
    .B(_0327_),
    .S(io_in2[4]),
    .Z(_0599_)
  );
  AND2_X1 _1416_ (
    .A1(_0333_),
    .A2(_0599_),
    .ZN(_0600_)
  );
  AND2_X1 _1417_ (
    .A1(_0030_),
    .A2(_0341_),
    .ZN(_0601_)
  );
  AND2_X1 _1418_ (
    .A1(io_in2[15]),
    .A2(io_in1[15]),
    .ZN(_0602_)
  );
  AND2_X1 _1419_ (
    .A1(_0338_),
    .A2(_0602_),
    .ZN(_0603_)
  );
  OR2_X1 _1420_ (
    .A1(_0600_),
    .A2(_0601_),
    .ZN(_0604_)
  );
  OR2_X1 _1421_ (
    .A1(_0598_),
    .A2(_0603_),
    .ZN(_0605_)
  );
  OR2_X1 _1422_ (
    .A1(_0604_),
    .A2(_0605_),
    .ZN(_0606_)
  );
  OR2_X1 _1423_ (
    .A1(_0595_),
    .A2(_0606_),
    .ZN(io_out[15])
  );
  XOR2_X1 _1424_ (
    .A(_0131_),
    .B(_0165_),
    .Z(io_adder_out[16])
  );
  AND2_X1 _1425_ (
    .A1(_0336_),
    .A2(io_adder_out[16]),
    .ZN(_0607_)
  );
  AND2_X1 _1426_ (
    .A1(_0255_),
    .A2(_0599_),
    .ZN(_0608_)
  );
  AND2_X1 _1427_ (
    .A1(_0113_),
    .A2(_0341_),
    .ZN(_0609_)
  );
  AND2_X1 _1428_ (
    .A1(io_in2[16]),
    .A2(io_in1[16]),
    .ZN(_0610_)
  );
  AND2_X1 _1429_ (
    .A1(_0338_),
    .A2(_0610_),
    .ZN(_0611_)
  );
  OR2_X1 _1430_ (
    .A1(_0609_),
    .A2(_0611_),
    .ZN(_0612_)
  );
  OR2_X1 _1431_ (
    .A1(_0608_),
    .A2(_0612_),
    .ZN(_0613_)
  );
  AND2_X1 _1432_ (
    .A1(_0333_),
    .A2(_0597_),
    .ZN(_0614_)
  );
  OR2_X1 _1433_ (
    .A1(_0613_),
    .A2(_0614_),
    .ZN(_0615_)
  );
  OR2_X1 _1434_ (
    .A1(_0607_),
    .A2(_0615_),
    .ZN(io_out[16])
  );
  XOR2_X1 _1435_ (
    .A(_0130_),
    .B(_0166_),
    .Z(io_adder_out[17])
  );
  AND2_X1 _1436_ (
    .A1(_0336_),
    .A2(io_adder_out[17]),
    .ZN(_0616_)
  );
  AND2_X1 _1437_ (
    .A1(_0333_),
    .A2(_0585_),
    .ZN(_0617_)
  );
  AND2_X1 _1438_ (
    .A1(_0255_),
    .A2(_0592_),
    .ZN(_0618_)
  );
  AND2_X1 _1439_ (
    .A1(io_in2[17]),
    .A2(io_in1[17]),
    .ZN(_0619_)
  );
  AND2_X1 _1440_ (
    .A1(_0338_),
    .A2(_0619_),
    .ZN(_0620_)
  );
  AND2_X1 _1441_ (
    .A1(_0116_),
    .A2(_0341_),
    .ZN(_0621_)
  );
  OR2_X1 _1442_ (
    .A1(_0620_),
    .A2(_0621_),
    .ZN(_0622_)
  );
  OR2_X1 _1443_ (
    .A1(_0618_),
    .A2(_0622_),
    .ZN(_0623_)
  );
  OR2_X1 _1444_ (
    .A1(_0617_),
    .A2(_0623_),
    .ZN(_0624_)
  );
  OR2_X1 _1445_ (
    .A1(_0616_),
    .A2(_0624_),
    .ZN(io_out[17])
  );
  XOR2_X1 _1446_ (
    .A(_0167_),
    .B(_0168_),
    .Z(io_adder_out[18])
  );
  AND2_X1 _1447_ (
    .A1(_0336_),
    .A2(io_adder_out[18]),
    .ZN(_0625_)
  );
  AND2_X1 _1448_ (
    .A1(_0255_),
    .A2(_0580_),
    .ZN(_0626_)
  );
  AND2_X1 _1449_ (
    .A1(_0022_),
    .A2(_0341_),
    .ZN(_0627_)
  );
  AND2_X1 _1450_ (
    .A1(io_in2[18]),
    .A2(io_in1[18]),
    .ZN(_0628_)
  );
  AND2_X1 _1451_ (
    .A1(_0338_),
    .A2(_0628_),
    .ZN(_0629_)
  );
  OR2_X1 _1452_ (
    .A1(_0627_),
    .A2(_0629_),
    .ZN(_0630_)
  );
  OR2_X1 _1453_ (
    .A1(_0626_),
    .A2(_0630_),
    .ZN(_0631_)
  );
  AND2_X1 _1454_ (
    .A1(_0333_),
    .A2(_0573_),
    .ZN(_0632_)
  );
  OR2_X1 _1455_ (
    .A1(_0631_),
    .A2(_0632_),
    .ZN(_0633_)
  );
  OR2_X1 _1456_ (
    .A1(_0625_),
    .A2(_0633_),
    .ZN(io_out[18])
  );
  XOR2_X1 _1457_ (
    .A(_0169_),
    .B(_0170_),
    .Z(io_adder_out[19])
  );
  AND2_X1 _1458_ (
    .A1(_0336_),
    .A2(io_adder_out[19]),
    .ZN(_0634_)
  );
  AND2_X1 _1459_ (
    .A1(_0255_),
    .A2(_0563_),
    .ZN(_0635_)
  );
  AND2_X1 _1460_ (
    .A1(_0019_),
    .A2(_0341_),
    .ZN(_0636_)
  );
  AND2_X1 _1461_ (
    .A1(io_in2[19]),
    .A2(io_in1[19]),
    .ZN(_0637_)
  );
  AND2_X1 _1462_ (
    .A1(_0338_),
    .A2(_0637_),
    .ZN(_0638_)
  );
  OR2_X1 _1463_ (
    .A1(_0636_),
    .A2(_0638_),
    .ZN(_0639_)
  );
  OR2_X1 _1464_ (
    .A1(_0635_),
    .A2(_0639_),
    .ZN(_0640_)
  );
  AND2_X1 _1465_ (
    .A1(_0333_),
    .A2(_0561_),
    .ZN(_0641_)
  );
  OR2_X1 _1466_ (
    .A1(_0640_),
    .A2(_0641_),
    .ZN(_0642_)
  );
  OR2_X1 _1467_ (
    .A1(_0634_),
    .A2(_0642_),
    .ZN(io_out[19])
  );
  XOR2_X1 _1468_ (
    .A(_0129_),
    .B(_0171_),
    .Z(io_adder_out[20])
  );
  AND2_X1 _1469_ (
    .A1(_0336_),
    .A2(io_adder_out[20]),
    .ZN(_0643_)
  );
  AND2_X1 _1470_ (
    .A1(_0255_),
    .A2(_0556_),
    .ZN(_0644_)
  );
  AND2_X1 _1471_ (
    .A1(_0016_),
    .A2(_0341_),
    .ZN(_0645_)
  );
  AND2_X1 _1472_ (
    .A1(io_in2[20]),
    .A2(io_in1[20]),
    .ZN(_0646_)
  );
  AND2_X1 _1473_ (
    .A1(_0338_),
    .A2(_0646_),
    .ZN(_0647_)
  );
  OR2_X1 _1474_ (
    .A1(_0645_),
    .A2(_0647_),
    .ZN(_0648_)
  );
  OR2_X1 _1475_ (
    .A1(_0644_),
    .A2(_0648_),
    .ZN(_0649_)
  );
  AND2_X1 _1476_ (
    .A1(_0333_),
    .A2(_0549_),
    .ZN(_0650_)
  );
  OR2_X1 _1477_ (
    .A1(_0649_),
    .A2(_0650_),
    .ZN(_0651_)
  );
  OR2_X1 _1478_ (
    .A1(_0643_),
    .A2(_0651_),
    .ZN(io_out[20])
  );
  XOR2_X1 _1479_ (
    .A(_0172_),
    .B(_0174_),
    .Z(io_adder_out[21])
  );
  AND2_X1 _1480_ (
    .A1(_0336_),
    .A2(io_adder_out[21]),
    .ZN(_0652_)
  );
  AND2_X1 _1481_ (
    .A1(_0255_),
    .A2(_0539_),
    .ZN(_0653_)
  );
  AND2_X1 _1482_ (
    .A1(_0173_),
    .A2(_0341_),
    .ZN(_0654_)
  );
  AND2_X1 _1483_ (
    .A1(io_in2[21]),
    .A2(io_in1[21]),
    .ZN(_0655_)
  );
  AND2_X1 _1484_ (
    .A1(_0338_),
    .A2(_0655_),
    .ZN(_0656_)
  );
  OR2_X1 _1485_ (
    .A1(_0654_),
    .A2(_0656_),
    .ZN(_0657_)
  );
  OR2_X1 _1486_ (
    .A1(_0653_),
    .A2(_0657_),
    .ZN(_0658_)
  );
  AND2_X1 _1487_ (
    .A1(_0333_),
    .A2(_0537_),
    .ZN(_0659_)
  );
  OR2_X1 _1488_ (
    .A1(_0658_),
    .A2(_0659_),
    .ZN(_0660_)
  );
  OR2_X1 _1489_ (
    .A1(_0652_),
    .A2(_0660_),
    .ZN(io_out[21])
  );
  XOR2_X1 _1490_ (
    .A(_0128_),
    .B(_0175_),
    .Z(io_adder_out[22])
  );
  AND2_X1 _1491_ (
    .A1(_0336_),
    .A2(io_adder_out[22]),
    .ZN(_0661_)
  );
  AND2_X1 _1492_ (
    .A1(_0255_),
    .A2(_0524_),
    .ZN(_0662_)
  );
  AND2_X1 _1493_ (
    .A1(_0333_),
    .A2(_0527_),
    .ZN(_0663_)
  );
  AND2_X1 _1494_ (
    .A1(io_in2[22]),
    .A2(io_in1[22]),
    .ZN(_0664_)
  );
  AND2_X1 _1495_ (
    .A1(_0338_),
    .A2(_0664_),
    .ZN(_0665_)
  );
  AND2_X1 _1496_ (
    .A1(_0010_),
    .A2(_0341_),
    .ZN(_0666_)
  );
  OR2_X1 _1497_ (
    .A1(_0665_),
    .A2(_0666_),
    .ZN(_0667_)
  );
  OR2_X1 _1498_ (
    .A1(_0663_),
    .A2(_0667_),
    .ZN(_0668_)
  );
  OR2_X1 _1499_ (
    .A1(_0662_),
    .A2(_0668_),
    .ZN(_0669_)
  );
  OR2_X1 _1500_ (
    .A1(_0661_),
    .A2(_0669_),
    .ZN(io_out[22])
  );
  XOR2_X1 _1501_ (
    .A(_0176_),
    .B(_0182_),
    .Z(io_adder_out[23])
  );
  AND2_X1 _1502_ (
    .A1(_0336_),
    .A2(io_adder_out[23]),
    .ZN(_0670_)
  );
  AND2_X1 _1503_ (
    .A1(_0255_),
    .A2(_0512_),
    .ZN(_0671_)
  );
  AND2_X1 _1504_ (
    .A1(_0333_),
    .A2(_0515_),
    .ZN(_0672_)
  );
  AND2_X1 _1505_ (
    .A1(_0180_),
    .A2(_0341_),
    .ZN(_0673_)
  );
  AND2_X1 _1506_ (
    .A1(io_in2[23]),
    .A2(io_in1[23]),
    .ZN(_0674_)
  );
  AND2_X1 _1507_ (
    .A1(_0338_),
    .A2(_0674_),
    .ZN(_0675_)
  );
  OR2_X1 _1508_ (
    .A1(_0673_),
    .A2(_0675_),
    .ZN(_0676_)
  );
  OR2_X1 _1509_ (
    .A1(_0672_),
    .A2(_0676_),
    .ZN(_0677_)
  );
  OR2_X1 _1510_ (
    .A1(_0671_),
    .A2(_0677_),
    .ZN(_0678_)
  );
  OR2_X1 _1511_ (
    .A1(_0670_),
    .A2(_0678_),
    .ZN(io_out[23])
  );
  XOR2_X1 _1512_ (
    .A(_0183_),
    .B(_0190_),
    .Z(io_adder_out[24])
  );
  AND2_X1 _1513_ (
    .A1(_0336_),
    .A2(io_adder_out[24]),
    .ZN(_0679_)
  );
  AND2_X1 _1514_ (
    .A1(_0255_),
    .A2(_0503_),
    .ZN(_0680_)
  );
  AND2_X1 _1515_ (
    .A1(_0186_),
    .A2(_0341_),
    .ZN(_0681_)
  );
  AND2_X1 _1516_ (
    .A1(io_in2[24]),
    .A2(io_in1[24]),
    .ZN(_0682_)
  );
  AND2_X1 _1517_ (
    .A1(_0338_),
    .A2(_0682_),
    .ZN(_0683_)
  );
  OR2_X1 _1518_ (
    .A1(_0681_),
    .A2(_0683_),
    .ZN(_0684_)
  );
  OR2_X1 _1519_ (
    .A1(_0680_),
    .A2(_0684_),
    .ZN(_0685_)
  );
  AND2_X1 _1520_ (
    .A1(_0333_),
    .A2(_0500_),
    .ZN(_0686_)
  );
  OR2_X1 _1521_ (
    .A1(_0685_),
    .A2(_0686_),
    .ZN(_0687_)
  );
  OR2_X1 _1522_ (
    .A1(_0679_),
    .A2(_0687_),
    .ZN(io_out[24])
  );
  XOR2_X1 _1523_ (
    .A(_0191_),
    .B(_0197_),
    .Z(io_adder_out[25])
  );
  AND2_X1 _1524_ (
    .A1(_0336_),
    .A2(io_adder_out[25]),
    .ZN(_0688_)
  );
  AND2_X1 _1525_ (
    .A1(_0255_),
    .A2(_0486_),
    .ZN(_0689_)
  );
  AND2_X1 _1526_ (
    .A1(_0194_),
    .A2(_0341_),
    .ZN(_0690_)
  );
  AND2_X1 _1527_ (
    .A1(io_in2[25]),
    .A2(io_in1[25]),
    .ZN(_0691_)
  );
  AND2_X1 _1528_ (
    .A1(_0338_),
    .A2(_0691_),
    .ZN(_0692_)
  );
  OR2_X1 _1529_ (
    .A1(_0690_),
    .A2(_0692_),
    .ZN(_0693_)
  );
  OR2_X1 _1530_ (
    .A1(_0689_),
    .A2(_0693_),
    .ZN(_0694_)
  );
  AND2_X1 _1531_ (
    .A1(_0333_),
    .A2(_0483_),
    .ZN(_0695_)
  );
  OR2_X1 _1532_ (
    .A1(_0694_),
    .A2(_0695_),
    .ZN(_0696_)
  );
  OR2_X1 _1533_ (
    .A1(_0688_),
    .A2(_0696_),
    .ZN(io_out[25])
  );
  XOR2_X1 _1534_ (
    .A(_0198_),
    .B(_0204_),
    .Z(io_adder_out[26])
  );
  AND2_X1 _1535_ (
    .A1(_0336_),
    .A2(io_adder_out[26]),
    .ZN(_0697_)
  );
  AND2_X1 _1536_ (
    .A1(_0255_),
    .A2(_0461_),
    .ZN(_0698_)
  );
  AND2_X1 _1537_ (
    .A1(_0333_),
    .A2(_0474_),
    .ZN(_0699_)
  );
  AND2_X1 _1538_ (
    .A1(_0201_),
    .A2(_0341_),
    .ZN(_0700_)
  );
  AND2_X1 _1539_ (
    .A1(io_in2[26]),
    .A2(io_in1[26]),
    .ZN(_0701_)
  );
  AND2_X1 _1540_ (
    .A1(_0338_),
    .A2(_0701_),
    .ZN(_0702_)
  );
  OR2_X1 _1541_ (
    .A1(_0700_),
    .A2(_0702_),
    .ZN(_0703_)
  );
  OR2_X1 _1542_ (
    .A1(_0699_),
    .A2(_0703_),
    .ZN(_0704_)
  );
  OR2_X1 _1543_ (
    .A1(_0698_),
    .A2(_0704_),
    .ZN(_0705_)
  );
  OR2_X1 _1544_ (
    .A1(_0697_),
    .A2(_0705_),
    .ZN(io_out[26])
  );
  XOR2_X1 _1545_ (
    .A(_0205_),
    .B(_0211_),
    .Z(io_adder_out[27])
  );
  AND2_X1 _1546_ (
    .A1(_0336_),
    .A2(io_adder_out[27]),
    .ZN(_0706_)
  );
  AND2_X1 _1547_ (
    .A1(_0255_),
    .A2(_0444_),
    .ZN(_0707_)
  );
  AND2_X1 _1548_ (
    .A1(_0208_),
    .A2(_0341_),
    .ZN(_0708_)
  );
  AND2_X1 _1549_ (
    .A1(io_in2[27]),
    .A2(io_in1[27]),
    .ZN(_0709_)
  );
  AND2_X1 _1550_ (
    .A1(_0338_),
    .A2(_0709_),
    .ZN(_0710_)
  );
  OR2_X1 _1551_ (
    .A1(_0708_),
    .A2(_0710_),
    .ZN(_0711_)
  );
  OR2_X1 _1552_ (
    .A1(_0707_),
    .A2(_0711_),
    .ZN(_0712_)
  );
  AND2_X1 _1553_ (
    .A1(_0333_),
    .A2(_0451_),
    .ZN(_0713_)
  );
  OR2_X1 _1554_ (
    .A1(_0712_),
    .A2(_0713_),
    .ZN(_0714_)
  );
  OR2_X1 _1555_ (
    .A1(_0706_),
    .A2(_0714_),
    .ZN(io_out[27])
  );
  XOR2_X1 _1556_ (
    .A(_0212_),
    .B(_0218_),
    .Z(io_adder_out[28])
  );
  AND2_X1 _1557_ (
    .A1(_0336_),
    .A2(io_adder_out[28]),
    .ZN(_0715_)
  );
  AND2_X1 _1558_ (
    .A1(_0255_),
    .A2(_0419_),
    .ZN(_0716_)
  );
  AND2_X1 _1559_ (
    .A1(_0216_),
    .A2(_0341_),
    .ZN(_0717_)
  );
  AND2_X1 _1560_ (
    .A1(io_in2[28]),
    .A2(io_in1[28]),
    .ZN(_0718_)
  );
  AND2_X1 _1561_ (
    .A1(_0338_),
    .A2(_0718_),
    .ZN(_0719_)
  );
  OR2_X1 _1562_ (
    .A1(_0717_),
    .A2(_0719_),
    .ZN(_0720_)
  );
  OR2_X1 _1563_ (
    .A1(_0716_),
    .A2(_0720_),
    .ZN(_0721_)
  );
  AND2_X1 _1564_ (
    .A1(_0333_),
    .A2(_0434_),
    .ZN(_0722_)
  );
  OR2_X1 _1565_ (
    .A1(_0721_),
    .A2(_0722_),
    .ZN(_0723_)
  );
  OR2_X1 _1566_ (
    .A1(_0715_),
    .A2(_0723_),
    .ZN(io_out[28])
  );
  XOR2_X1 _1567_ (
    .A(_0219_),
    .B(_0225_),
    .Z(io_adder_out[29])
  );
  AND2_X1 _1568_ (
    .A1(_0336_),
    .A2(io_adder_out[29]),
    .ZN(_0724_)
  );
  AND2_X1 _1569_ (
    .A1(_0333_),
    .A2(_0408_),
    .ZN(_0725_)
  );
  AND2_X1 _1570_ (
    .A1(_0255_),
    .A2(_0393_),
    .ZN(_0726_)
  );
  AND2_X1 _1571_ (
    .A1(_0222_),
    .A2(_0341_),
    .ZN(_0727_)
  );
  AND2_X1 _1572_ (
    .A1(io_in2[29]),
    .A2(io_in1[29]),
    .ZN(_0728_)
  );
  AND2_X1 _1573_ (
    .A1(_0338_),
    .A2(_0728_),
    .ZN(_0729_)
  );
  OR2_X1 _1574_ (
    .A1(_0727_),
    .A2(_0729_),
    .ZN(_0730_)
  );
  OR2_X1 _1575_ (
    .A1(_0726_),
    .A2(_0730_),
    .ZN(_0731_)
  );
  OR2_X1 _1576_ (
    .A1(_0725_),
    .A2(_0731_),
    .ZN(_0732_)
  );
  OR2_X1 _1577_ (
    .A1(_0724_),
    .A2(_0732_),
    .ZN(io_out[29])
  );
  XOR2_X1 _1578_ (
    .A(_0226_),
    .B(_0232_),
    .Z(io_adder_out[30])
  );
  AND2_X1 _1579_ (
    .A1(_0336_),
    .A2(io_adder_out[30]),
    .ZN(_0733_)
  );
  AND2_X1 _1580_ (
    .A1(_0333_),
    .A2(_0382_),
    .ZN(_0734_)
  );
  AND2_X1 _1581_ (
    .A1(_0255_),
    .A2(_0351_),
    .ZN(_0735_)
  );
  AND2_X1 _1582_ (
    .A1(_0230_),
    .A2(_0341_),
    .ZN(_0736_)
  );
  AND2_X1 _1583_ (
    .A1(io_in2[30]),
    .A2(io_in1[30]),
    .ZN(_0737_)
  );
  AND2_X1 _1584_ (
    .A1(_0338_),
    .A2(_0737_),
    .ZN(_0738_)
  );
  OR2_X1 _1585_ (
    .A1(_0736_),
    .A2(_0738_),
    .ZN(_0739_)
  );
  OR2_X1 _1586_ (
    .A1(_0735_),
    .A2(_0739_),
    .ZN(_0740_)
  );
  OR2_X1 _1587_ (
    .A1(_0734_),
    .A2(_0740_),
    .ZN(_0741_)
  );
  OR2_X1 _1588_ (
    .A1(_0733_),
    .A2(_0741_),
    .ZN(io_out[30])
  );
  AND2_X1 _1589_ (
    .A1(io_adder_out[31]),
    .A2(_0336_),
    .ZN(_0742_)
  );
  AND2_X1 _1590_ (
    .A1(_0323_),
    .A2(_0333_),
    .ZN(_0743_)
  );
  AND2_X1 _1591_ (
    .A1(_0255_),
    .A2(_0330_),
    .ZN(_0744_)
  );
  AND2_X1 _1592_ (
    .A1(_0237_),
    .A2(_0341_),
    .ZN(_0745_)
  );
  AND2_X1 _1593_ (
    .A1(io_in2[31]),
    .A2(io_in1[31]),
    .ZN(_0746_)
  );
  AND2_X1 _1594_ (
    .A1(_0338_),
    .A2(_0746_),
    .ZN(_0747_)
  );
  OR2_X1 _1595_ (
    .A1(_0745_),
    .A2(_0747_),
    .ZN(_0748_)
  );
  OR2_X1 _1596_ (
    .A1(_0744_),
    .A2(_0748_),
    .ZN(_0749_)
  );
  OR2_X1 _1597_ (
    .A1(_0743_),
    .A2(_0749_),
    .ZN(_0750_)
  );
  OR2_X1 _1598_ (
    .A1(_0742_),
    .A2(_0750_),
    .ZN(io_out[31])
  );
  OR2_X1 _1599_ (
    .A1(_0222_),
    .A2(_0230_),
    .ZN(_0751_)
  );
  OR2_X1 _1600_ (
    .A1(_0240_),
    .A2(_0751_),
    .ZN(_0752_)
  );
  OR2_X1 _1601_ (
    .A1(_0194_),
    .A2(_0201_),
    .ZN(_0753_)
  );
  OR2_X1 _1602_ (
    .A1(_0208_),
    .A2(_0216_),
    .ZN(_0754_)
  );
  OR2_X1 _1603_ (
    .A1(_0753_),
    .A2(_0754_),
    .ZN(_0755_)
  );
  OR2_X1 _1604_ (
    .A1(_0116_),
    .A2(_0173_),
    .ZN(_0756_)
  );
  OR2_X1 _1605_ (
    .A1(_0180_),
    .A2(_0186_),
    .ZN(_0757_)
  );
  OR2_X1 _1606_ (
    .A1(_0756_),
    .A2(_0757_),
    .ZN(_0758_)
  );
  OR2_X1 _1607_ (
    .A1(_0755_),
    .A2(_0758_),
    .ZN(_0759_)
  );
  OR2_X1 _1608_ (
    .A1(_0752_),
    .A2(_0759_),
    .ZN(_0760_)
  );
  OR2_X1 _1609_ (
    .A1(_0010_),
    .A2(_0016_),
    .ZN(_0761_)
  );
  OR2_X1 _1610_ (
    .A1(_0019_),
    .A2(_0022_),
    .ZN(_0762_)
  );
  OR2_X1 _1611_ (
    .A1(_0761_),
    .A2(_0762_),
    .ZN(_0763_)
  );
  OR2_X1 _1612_ (
    .A1(_0242_),
    .A2(_0763_),
    .ZN(_0764_)
  );
  OR2_X1 _1613_ (
    .A1(_0044_),
    .A2(_0047_),
    .ZN(_0765_)
  );
  OR2_X1 _1614_ (
    .A1(_0050_),
    .A2(_0055_),
    .ZN(_0766_)
  );
  OR2_X1 _1615_ (
    .A1(_0765_),
    .A2(_0766_),
    .ZN(_0767_)
  );
  OR2_X1 _1616_ (
    .A1(_0030_),
    .A2(_0033_),
    .ZN(_0768_)
  );
  OR2_X1 _1617_ (
    .A1(_0037_),
    .A2(_0040_),
    .ZN(_0769_)
  );
  OR2_X1 _1618_ (
    .A1(_0768_),
    .A2(_0769_),
    .ZN(_0770_)
  );
  OR2_X1 _1619_ (
    .A1(_0767_),
    .A2(_0770_),
    .ZN(_0771_)
  );
  OR2_X1 _1620_ (
    .A1(_0083_),
    .A2(_0086_),
    .ZN(_0772_)
  );
  OR2_X1 _1621_ (
    .A1(_0093_),
    .A2(_0113_),
    .ZN(_0773_)
  );
  OR2_X1 _1622_ (
    .A1(_0772_),
    .A2(_0773_),
    .ZN(_0774_)
  );
  OR2_X1 _1623_ (
    .A1(_0058_),
    .A2(_0073_),
    .ZN(_0775_)
  );
  OR2_X1 _1624_ (
    .A1(_0077_),
    .A2(_0080_),
    .ZN(_0776_)
  );
  OR2_X1 _1625_ (
    .A1(_0775_),
    .A2(_0776_),
    .ZN(_0777_)
  );
  OR2_X1 _1626_ (
    .A1(_0774_),
    .A2(_0777_),
    .ZN(_0778_)
  );
  OR2_X1 _1627_ (
    .A1(_0771_),
    .A2(_0778_),
    .ZN(_0779_)
  );
  OR2_X1 _1628_ (
    .A1(_0764_),
    .A2(_0779_),
    .ZN(_0780_)
  );
  OR2_X1 _1629_ (
    .A1(_0760_),
    .A2(_0780_),
    .ZN(_0781_)
  );
  INV_X1 _1630_ (
    .A(_0781_),
    .ZN(_0782_)
  );
  OR2_X1 _1631_ (
    .A1(_0249_),
    .A2(_0782_),
    .ZN(_0783_)
  );
  XOR2_X1 _1632_ (
    .A(io_fn[0]),
    .B(_0783_),
    .Z(io_cmp_out)
  );
  assign _GEN_0 = { 31'h00000000, io_fn[3] };
  assign _GEN_1 = { 16'h0000, io_in1[31:16] };
  assign _GEN_10[31] = 1'h0;
  assign _GEN_11[31:1] = 31'h00000000;
  assign _GEN_2 = { 8'h00, io_in1[15:0], io_in1[31:24] };
  assign _GEN_3 = { 4'h0, io_in1[7:0], io_in1[15:8], io_in1[23:16], io_in1[31:28] };
  assign _GEN_4 = { 2'h0, io_in1[3:0], io_in1[7:4], io_in1[11:8], io_in1[15:12], io_in1[19:16], io_in1[23:20], io_in1[27:24], io_in1[31:30] };
  assign _GEN_5 = { 1'h0, io_in1[1:0], io_in1[3:2], io_in1[5:4], io_in1[7:6], io_in1[9:8], io_in1[11:10], io_in1[13:12], io_in1[15:14], io_in1[17:16], io_in1[19:18], io_in1[21:20], io_in1[23:22], io_in1[25:24], io_in1[27:26], io_in1[29:28], io_in1[31] };
  assign { _GEN_6[31:15], _GEN_6[13:0] } = { 16'h0000, _GEN_10[0], _GEN_10[2:1], _GEN_10[4:3], _GEN_10[6:5], _GEN_10[8:7], _GEN_10[10:9], _GEN_10[12:11], _GEN_10[14:13] };
  assign _GEN_7 = { 8'h00, _GEN_10[16:15], _GEN_10[18:17], _GEN_10[20:19], _GEN_10[22:21], _GEN_10[24:23], _GEN_10[26:25], _GEN_10[28:27], _GEN_10[30:29], _GEN_10[0], _GEN_6[14], _GEN_10[2:1], _GEN_10[4:3], _GEN_10[6:5] };
  assign _GEN_8 = { 4'h0, _GEN_10[24:23], _GEN_10[26:25], _GEN_10[28:27], _GEN_10[30:29], _GEN_10[16:15], _GEN_10[18:17], _GEN_10[20:19], _GEN_10[22:21], _GEN_10[8:7], _GEN_10[10:9], _GEN_10[12:11], _GEN_10[14:13], _GEN_10[0], _GEN_6[14], _GEN_10[2:1] };
  assign _GEN_9 = { 2'h0, _GEN_10[28:27], _GEN_10[30:29], _GEN_10[24:23], _GEN_10[26:25], _GEN_10[20:19], _GEN_10[22:21], _GEN_10[16:15], _GEN_10[18:17], _GEN_10[12:11], _GEN_10[14:13], _GEN_10[8:7], _GEN_10[10:9], _GEN_10[4:3], _GEN_10[6:5], _GEN_10[0], _GEN_6[14] };
  assign _shift_logic_T_1 = _GEN_11[0];
  assign _shin_T_10 = { io_in1[15:0], 16'h0000 };
  assign _shin_T_11 = { io_in1[15:0], io_in1[31:16] };
  assign _shin_T_16 = { 8'h00, io_in1[15:8], 8'h00, io_in1[31:24] };
  assign _shin_T_18 = { io_in1[7:0], io_in1[31:16], 8'h00 };
  assign _shin_T_20 = { io_in1[7:0], 8'h00, io_in1[23:16], 8'h00 };
  assign _shin_T_21 = { io_in1[7:0], io_in1[15:8], io_in1[23:16], io_in1[31:24] };
  assign _shin_T_26 = { 4'h0, io_in1[7:4], 4'h0, io_in1[15:12], 4'h0, io_in1[23:20], 4'h0, io_in1[31:28] };
  assign _shin_T_28 = { io_in1[3:0], io_in1[15:8], io_in1[23:16], io_in1[31:24], 4'h0 };
  assign _shin_T_30 = { io_in1[3:0], 4'h0, io_in1[11:8], 4'h0, io_in1[19:16], 4'h0, io_in1[27:24], 4'h0 };
  assign _shin_T_31 = { io_in1[3:0], io_in1[7:4], io_in1[11:8], io_in1[15:12], io_in1[19:16], io_in1[23:20], io_in1[27:24], io_in1[31:28] };
  assign _shin_T_36 = { 2'h0, io_in1[3:2], 2'h0, io_in1[7:6], 2'h0, io_in1[11:10], 2'h0, io_in1[15:14], 2'h0, io_in1[19:18], 2'h0, io_in1[23:22], 2'h0, io_in1[27:26], 2'h0, io_in1[31:30] };
  assign _shin_T_38 = { io_in1[1:0], io_in1[7:4], io_in1[11:8], io_in1[15:12], io_in1[19:16], io_in1[23:20], io_in1[27:24], io_in1[31:28], 2'h0 };
  assign _shin_T_40 = { io_in1[1:0], 2'h0, io_in1[5:4], 2'h0, io_in1[9:8], 2'h0, io_in1[13:12], 2'h0, io_in1[17:16], 2'h0, io_in1[21:20], 2'h0, io_in1[25:24], 2'h0, io_in1[29:28], 2'h0 };
  assign _shin_T_41 = { io_in1[1:0], io_in1[3:2], io_in1[5:4], io_in1[7:6], io_in1[9:8], io_in1[11:10], io_in1[13:12], io_in1[15:14], io_in1[17:16], io_in1[19:18], io_in1[21:20], io_in1[23:22], io_in1[25:24], io_in1[27:26], io_in1[29:28], io_in1[31:30] };
  assign _shin_T_46 = { 1'h0, io_in1[1], 1'h0, io_in1[3], 1'h0, io_in1[5], 1'h0, io_in1[7], 1'h0, io_in1[9], 1'h0, io_in1[11], 1'h0, io_in1[13], 1'h0, io_in1[15], 1'h0, io_in1[17], 1'h0, io_in1[19], 1'h0, io_in1[21], 1'h0, io_in1[23], 1'h0, io_in1[25], 1'h0, io_in1[27], 1'h0, io_in1[29], 1'h0, io_in1[31] };
  assign _shin_T_48 = { io_in1[0], io_in1[3:2], io_in1[5:4], io_in1[7:6], io_in1[9:8], io_in1[11:10], io_in1[13:12], io_in1[15:14], io_in1[17:16], io_in1[19:18], io_in1[21:20], io_in1[23:22], io_in1[25:24], io_in1[27:26], io_in1[29:28], io_in1[31:30], 1'h0 };
  assign _shin_T_50 = { io_in1[0], 1'h0, io_in1[2], 1'h0, io_in1[4], 1'h0, io_in1[6], 1'h0, io_in1[8], 1'h0, io_in1[10], 1'h0, io_in1[12], 1'h0, io_in1[14], 1'h0, io_in1[16], 1'h0, io_in1[18], 1'h0, io_in1[20], 1'h0, io_in1[22], 1'h0, io_in1[24], 1'h0, io_in1[26], 1'h0, io_in1[28], 1'h0, io_in1[30], 1'h0 };
  assign _shin_T_51 = { io_in1[0], io_in1[1], io_in1[2], io_in1[3], io_in1[4], io_in1[5], io_in1[6], io_in1[7], io_in1[8], io_in1[9], io_in1[10], io_in1[11], io_in1[12], io_in1[13], io_in1[14], io_in1[15], io_in1[16], io_in1[17], io_in1[18], io_in1[19], io_in1[20], io_in1[21], io_in1[22], io_in1[23], io_in1[24], io_in1[25], io_in1[26], io_in1[27], io_in1[28], io_in1[29], io_in1[30], io_in1[31] };
  assign _shin_T_6 = { 16'h0000, io_in1[31:16] };
  assign _shin_T_8 = { io_in1[15:0], 16'h0000 };
  assign _shout_l_T_13 = { 8'h00, _GEN_10[16:15], _GEN_10[18:17], _GEN_10[20:19], _GEN_10[22:21], 8'h00, _GEN_10[0], _GEN_6[14], _GEN_10[2:1], _GEN_10[4:3], _GEN_10[6:5] };
  assign _shout_l_T_15 = { _GEN_10[24:23], _GEN_10[26:25], _GEN_10[28:27], _GEN_10[30:29], _GEN_10[0], _GEN_6[14], _GEN_10[2:1], _GEN_10[4:3], _GEN_10[6:5], _GEN_10[8:7], _GEN_10[10:9], _GEN_10[12:11], _GEN_10[14:13], 8'h00 };
  assign _shout_l_T_17 = { _GEN_10[24:23], _GEN_10[26:25], _GEN_10[28:27], _GEN_10[30:29], 8'h00, _GEN_10[8:7], _GEN_10[10:9], _GEN_10[12:11], _GEN_10[14:13], 8'h00 };
  assign _shout_l_T_18 = { _GEN_10[24:23], _GEN_10[26:25], _GEN_10[28:27], _GEN_10[30:29], _GEN_10[16:15], _GEN_10[18:17], _GEN_10[20:19], _GEN_10[22:21], _GEN_10[8:7], _GEN_10[10:9], _GEN_10[12:11], _GEN_10[14:13], _GEN_10[0], _GEN_6[14], _GEN_10[2:1], _GEN_10[4:3], _GEN_10[6:5] };
  assign _shout_l_T_23 = { 4'h0, _GEN_10[24:23], _GEN_10[26:25], 4'h0, _GEN_10[16:15], _GEN_10[18:17], 4'h0, _GEN_10[8:7], _GEN_10[10:9], 4'h0, _GEN_10[0], _GEN_6[14], _GEN_10[2:1] };
  assign _shout_l_T_25 = { _GEN_10[28:27], _GEN_10[30:29], _GEN_10[16:15], _GEN_10[18:17], _GEN_10[20:19], _GEN_10[22:21], _GEN_10[8:7], _GEN_10[10:9], _GEN_10[12:11], _GEN_10[14:13], _GEN_10[0], _GEN_6[14], _GEN_10[2:1], _GEN_10[4:3], _GEN_10[6:5], 4'h0 };
  assign _shout_l_T_27 = { _GEN_10[28:27], _GEN_10[30:29], 4'h0, _GEN_10[20:19], _GEN_10[22:21], 4'h0, _GEN_10[12:11], _GEN_10[14:13], 4'h0, _GEN_10[4:3], _GEN_10[6:5], 4'h0 };
  assign _shout_l_T_28 = { _GEN_10[28:27], _GEN_10[30:29], _GEN_10[24:23], _GEN_10[26:25], _GEN_10[20:19], _GEN_10[22:21], _GEN_10[16:15], _GEN_10[18:17], _GEN_10[12:11], _GEN_10[14:13], _GEN_10[8:7], _GEN_10[10:9], _GEN_10[4:3], _GEN_10[6:5], _GEN_10[0], _GEN_6[14], _GEN_10[2:1] };
  assign _shout_l_T_3 = { 16'h0000, _GEN_10[0], _GEN_6[14], _GEN_10[2:1], _GEN_10[4:3], _GEN_10[6:5], _GEN_10[8:7], _GEN_10[10:9], _GEN_10[12:11], _GEN_10[14:13] };
  assign _shout_l_T_33 = { 2'h0, _GEN_10[28:27], 2'h0, _GEN_10[24:23], 2'h0, _GEN_10[20:19], 2'h0, _GEN_10[16:15], 2'h0, _GEN_10[12:11], 2'h0, _GEN_10[8:7], 2'h0, _GEN_10[4:3], 2'h0, _GEN_10[0], _GEN_6[14] };
  assign _shout_l_T_35 = { _GEN_10[30:29], _GEN_10[24:23], _GEN_10[26:25], _GEN_10[20:19], _GEN_10[22:21], _GEN_10[16:15], _GEN_10[18:17], _GEN_10[12:11], _GEN_10[14:13], _GEN_10[8:7], _GEN_10[10:9], _GEN_10[4:3], _GEN_10[6:5], _GEN_10[0], _GEN_6[14], _GEN_10[2:1], 2'h0 };
  assign _shout_l_T_37 = { _GEN_10[30:29], 2'h0, _GEN_10[26:25], 2'h0, _GEN_10[22:21], 2'h0, _GEN_10[18:17], 2'h0, _GEN_10[14:13], 2'h0, _GEN_10[10:9], 2'h0, _GEN_10[6:5], 2'h0, _GEN_10[2:1], 2'h0 };
  assign _shout_l_T_38 = { _GEN_10[30:0], _GEN_6[14] };
  assign _shout_l_T_43 = { 1'h0, _GEN_10[30], 1'h0, _GEN_10[28], 1'h0, _GEN_10[26], 1'h0, _GEN_10[24], 1'h0, _GEN_10[22], 1'h0, _GEN_10[20], 1'h0, _GEN_10[18], 1'h0, _GEN_10[16], 1'h0, _GEN_10[14], 1'h0, _GEN_10[12], 1'h0, _GEN_10[10], 1'h0, _GEN_10[8], 1'h0, _GEN_10[6], 1'h0, _GEN_10[4], 1'h0, _GEN_10[2], 1'h0, _GEN_10[0] };
  assign _shout_l_T_45 = { _GEN_10[29:0], _GEN_6[14], 1'h0 };
  assign _shout_l_T_47 = { _GEN_10[29], 1'h0, _GEN_10[27], 1'h0, _GEN_10[25], 1'h0, _GEN_10[23], 1'h0, _GEN_10[21], 1'h0, _GEN_10[19], 1'h0, _GEN_10[17], 1'h0, _GEN_10[15], 1'h0, _GEN_10[13], 1'h0, _GEN_10[11], 1'h0, _GEN_10[9], 1'h0, _GEN_10[7], 1'h0, _GEN_10[5], 1'h0, _GEN_10[3], 1'h0, _GEN_10[1], 1'h0, _GEN_6[14], 1'h0 };
  assign _shout_l_T_5 = { _GEN_10[16:15], _GEN_10[18:17], _GEN_10[20:19], _GEN_10[22:21], _GEN_10[24:23], _GEN_10[26:25], _GEN_10[28:27], _GEN_10[30:29], 16'h0000 };
  assign _shout_l_T_7 = { _GEN_10[16:15], _GEN_10[18:17], _GEN_10[20:19], _GEN_10[22:21], _GEN_10[24:23], _GEN_10[26:25], _GEN_10[28:27], _GEN_10[30:29], 16'h0000 };
  assign _shout_l_T_8 = { _GEN_10[16:15], _GEN_10[18:17], _GEN_10[20:19], _GEN_10[22:21], _GEN_10[24:23], _GEN_10[26:25], _GEN_10[28:27], _GEN_10[30:29], _GEN_10[0], _GEN_6[14], _GEN_10[2:1], _GEN_10[4:3], _GEN_10[6:5], _GEN_10[8:7], _GEN_10[10:9], _GEN_10[12:11], _GEN_10[14:13] };
  assign _shout_r_T_5[31:0] = { _GEN_10[0], _GEN_6[14], _GEN_10[2:1], _GEN_10[4:3], _GEN_10[6:5], _GEN_10[8:7], _GEN_10[10:9], _GEN_10[12:11], _GEN_10[14:13], _GEN_10[16:15], _GEN_10[18:17], _GEN_10[20:19], _GEN_10[22:21], _GEN_10[24:23], _GEN_10[26:25], _GEN_10[28:27], _GEN_10[30:29] };
  assign shamt = io_in2[4:0];
  assign shout_l = { _GEN_10[29], _GEN_10[30], _GEN_10[27], _GEN_10[28], _GEN_10[25], _GEN_10[26], _GEN_10[23], _GEN_10[24], _GEN_10[21], _GEN_10[22], _GEN_10[19], _GEN_10[20], _GEN_10[17], _GEN_10[18], _GEN_10[15], _GEN_10[16], _GEN_10[13], _GEN_10[14], _GEN_10[11], _GEN_10[12], _GEN_10[9], _GEN_10[10], _GEN_10[7], _GEN_10[8], _GEN_10[5], _GEN_10[6], _GEN_10[3], _GEN_10[4], _GEN_10[1], _GEN_10[2], _GEN_6[14], _GEN_10[0] };
  assign shout_r = { _GEN_10[0], _GEN_6[14], _GEN_10[2:1], _GEN_10[4:3], _GEN_10[6:5], _GEN_10[8:7], _GEN_10[10:9], _GEN_10[12:11], _GEN_10[14:13], _GEN_10[16:15], _GEN_10[18:17], _GEN_10[20:19], _GEN_10[22:21], _GEN_10[24:23], _GEN_10[26:25], _GEN_10[28:27], _GEN_10[30:29] };
endmodule
module BreakpointUnit(io_status_debug, io_bp_0_control_action, io_bp_0_control_tmatch, io_bp_0_control_x, io_bp_0_control_w, io_bp_0_control_r, io_bp_0_address, io_pc, io_ea, io_xcpt_if, io_xcpt_ld, io_xcpt_st, io_debug_if, io_debug_ld, io_debug_st);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire [31:0] _GEN_11;
  wire _r_T_10;
  wire _r_T_12;
  wire [3:0] _r_T_13;
  wire _r_T_8;
  input [31:0] io_bp_0_address;
  wire [31:0] io_bp_0_address;
  input io_bp_0_control_action;
  wire io_bp_0_control_action;
  input io_bp_0_control_r;
  wire io_bp_0_control_r;
  input [1:0] io_bp_0_control_tmatch;
  wire [1:0] io_bp_0_control_tmatch;
  input io_bp_0_control_w;
  wire io_bp_0_control_w;
  input io_bp_0_control_x;
  wire io_bp_0_control_x;
  output io_debug_if;
  wire io_debug_if;
  output io_debug_ld;
  wire io_debug_ld;
  output io_debug_st;
  wire io_debug_st;
  input [31:0] io_ea;
  wire [31:0] io_ea;
  input [31:0] io_pc;
  wire [31:0] io_pc;
  input io_status_debug;
  wire io_status_debug;
  output io_xcpt_if;
  wire io_xcpt_if;
  output io_xcpt_ld;
  wire io_xcpt_ld;
  output io_xcpt_st;
  wire io_xcpt_st;
  INV_X1 _0506_ (
    .A(io_bp_0_control_tmatch[1]),
    .ZN(_0000_)
  );
  INV_X1 _0507_ (
    .A(io_status_debug),
    .ZN(_0001_)
  );
  INV_X1 _0508_ (
    .A(io_ea[5]),
    .ZN(_0002_)
  );
  INV_X1 _0509_ (
    .A(io_ea[6]),
    .ZN(_0003_)
  );
  INV_X1 _0510_ (
    .A(io_ea[7]),
    .ZN(_0004_)
  );
  INV_X1 _0511_ (
    .A(io_ea[8]),
    .ZN(_0005_)
  );
  INV_X1 _0512_ (
    .A(io_ea[9]),
    .ZN(_0006_)
  );
  INV_X1 _0513_ (
    .A(io_ea[10]),
    .ZN(_0007_)
  );
  INV_X1 _0514_ (
    .A(io_ea[11]),
    .ZN(_0008_)
  );
  INV_X1 _0515_ (
    .A(io_ea[12]),
    .ZN(_0009_)
  );
  INV_X1 _0516_ (
    .A(io_ea[13]),
    .ZN(_0010_)
  );
  INV_X1 _0517_ (
    .A(io_ea[16]),
    .ZN(_0011_)
  );
  INV_X1 _0518_ (
    .A(io_ea[17]),
    .ZN(_0012_)
  );
  INV_X1 _0519_ (
    .A(io_ea[18]),
    .ZN(_0013_)
  );
  INV_X1 _0520_ (
    .A(io_ea[19]),
    .ZN(_0014_)
  );
  INV_X1 _0521_ (
    .A(io_ea[20]),
    .ZN(_0015_)
  );
  INV_X1 _0522_ (
    .A(io_ea[21]),
    .ZN(_0016_)
  );
  INV_X1 _0523_ (
    .A(io_ea[22]),
    .ZN(_0017_)
  );
  INV_X1 _0524_ (
    .A(io_ea[23]),
    .ZN(_0018_)
  );
  INV_X1 _0525_ (
    .A(io_ea[24]),
    .ZN(_0019_)
  );
  INV_X1 _0526_ (
    .A(io_ea[25]),
    .ZN(_0020_)
  );
  INV_X1 _0527_ (
    .A(io_ea[28]),
    .ZN(_0021_)
  );
  INV_X1 _0528_ (
    .A(io_ea[29]),
    .ZN(_0022_)
  );
  INV_X1 _0529_ (
    .A(io_ea[30]),
    .ZN(_0023_)
  );
  INV_X1 _0530_ (
    .A(io_ea[31]),
    .ZN(_0024_)
  );
  INV_X1 _0531_ (
    .A(io_pc[0]),
    .ZN(_0025_)
  );
  INV_X1 _0532_ (
    .A(io_pc[1]),
    .ZN(_0026_)
  );
  INV_X1 _0533_ (
    .A(io_pc[2]),
    .ZN(_0027_)
  );
  INV_X1 _0534_ (
    .A(io_pc[3]),
    .ZN(_0028_)
  );
  INV_X1 _0535_ (
    .A(io_pc[4]),
    .ZN(_0029_)
  );
  INV_X1 _0536_ (
    .A(io_pc[5]),
    .ZN(_0030_)
  );
  INV_X1 _0537_ (
    .A(io_pc[6]),
    .ZN(_0031_)
  );
  INV_X1 _0538_ (
    .A(io_pc[7]),
    .ZN(_0032_)
  );
  INV_X1 _0539_ (
    .A(io_pc[8]),
    .ZN(_0033_)
  );
  INV_X1 _0540_ (
    .A(io_pc[9]),
    .ZN(_0034_)
  );
  INV_X1 _0541_ (
    .A(io_pc[10]),
    .ZN(_0035_)
  );
  INV_X1 _0542_ (
    .A(io_pc[11]),
    .ZN(_0036_)
  );
  INV_X1 _0543_ (
    .A(io_pc[12]),
    .ZN(_0037_)
  );
  INV_X1 _0544_ (
    .A(io_pc[13]),
    .ZN(_0038_)
  );
  INV_X1 _0545_ (
    .A(io_pc[14]),
    .ZN(_0039_)
  );
  INV_X1 _0546_ (
    .A(io_pc[15]),
    .ZN(_0040_)
  );
  INV_X1 _0547_ (
    .A(io_pc[16]),
    .ZN(_0041_)
  );
  INV_X1 _0548_ (
    .A(io_pc[17]),
    .ZN(_0042_)
  );
  INV_X1 _0549_ (
    .A(io_pc[18]),
    .ZN(_0043_)
  );
  INV_X1 _0550_ (
    .A(io_pc[19]),
    .ZN(_0044_)
  );
  INV_X1 _0551_ (
    .A(io_pc[20]),
    .ZN(_0045_)
  );
  INV_X1 _0552_ (
    .A(io_pc[21]),
    .ZN(_0046_)
  );
  INV_X1 _0553_ (
    .A(io_pc[22]),
    .ZN(_0047_)
  );
  INV_X1 _0554_ (
    .A(io_pc[23]),
    .ZN(_0048_)
  );
  INV_X1 _0555_ (
    .A(io_pc[24]),
    .ZN(_0049_)
  );
  INV_X1 _0556_ (
    .A(io_pc[25]),
    .ZN(_0050_)
  );
  INV_X1 _0557_ (
    .A(io_pc[26]),
    .ZN(_0051_)
  );
  INV_X1 _0558_ (
    .A(io_pc[27]),
    .ZN(_0052_)
  );
  INV_X1 _0559_ (
    .A(io_pc[28]),
    .ZN(_0053_)
  );
  INV_X1 _0560_ (
    .A(io_pc[29]),
    .ZN(_0054_)
  );
  INV_X1 _0561_ (
    .A(io_pc[30]),
    .ZN(_0055_)
  );
  INV_X1 _0562_ (
    .A(io_pc[31]),
    .ZN(_0056_)
  );
  INV_X1 _0563_ (
    .A(io_bp_0_control_action),
    .ZN(_0057_)
  );
  INV_X1 _0564_ (
    .A(io_bp_0_address[0]),
    .ZN(_0058_)
  );
  INV_X1 _0565_ (
    .A(io_bp_0_address[1]),
    .ZN(_0059_)
  );
  INV_X1 _0566_ (
    .A(io_bp_0_address[2]),
    .ZN(_0060_)
  );
  INV_X1 _0567_ (
    .A(io_bp_0_address[3]),
    .ZN(_0061_)
  );
  INV_X1 _0568_ (
    .A(io_bp_0_address[4]),
    .ZN(_0062_)
  );
  INV_X1 _0569_ (
    .A(io_bp_0_address[5]),
    .ZN(_0063_)
  );
  INV_X1 _0570_ (
    .A(io_bp_0_address[6]),
    .ZN(_0064_)
  );
  INV_X1 _0571_ (
    .A(io_bp_0_address[7]),
    .ZN(_0065_)
  );
  INV_X1 _0572_ (
    .A(io_bp_0_address[8]),
    .ZN(_0066_)
  );
  INV_X1 _0573_ (
    .A(io_bp_0_address[9]),
    .ZN(_0067_)
  );
  INV_X1 _0574_ (
    .A(io_bp_0_address[12]),
    .ZN(_0068_)
  );
  INV_X1 _0575_ (
    .A(io_bp_0_address[13]),
    .ZN(_0069_)
  );
  INV_X1 _0576_ (
    .A(io_bp_0_address[14]),
    .ZN(_0070_)
  );
  INV_X1 _0577_ (
    .A(io_bp_0_address[15]),
    .ZN(_0071_)
  );
  INV_X1 _0578_ (
    .A(io_bp_0_address[16]),
    .ZN(_0072_)
  );
  INV_X1 _0579_ (
    .A(io_bp_0_address[17]),
    .ZN(_0073_)
  );
  INV_X1 _0580_ (
    .A(io_bp_0_address[20]),
    .ZN(_0074_)
  );
  INV_X1 _0581_ (
    .A(io_bp_0_address[21]),
    .ZN(_0075_)
  );
  INV_X1 _0582_ (
    .A(io_bp_0_address[22]),
    .ZN(_0076_)
  );
  INV_X1 _0583_ (
    .A(io_bp_0_address[23]),
    .ZN(_0077_)
  );
  INV_X1 _0584_ (
    .A(io_bp_0_address[24]),
    .ZN(_0078_)
  );
  INV_X1 _0585_ (
    .A(io_bp_0_address[25]),
    .ZN(_0079_)
  );
  INV_X1 _0586_ (
    .A(io_bp_0_address[26]),
    .ZN(_0080_)
  );
  INV_X1 _0587_ (
    .A(io_bp_0_address[27]),
    .ZN(_0081_)
  );
  INV_X1 _0588_ (
    .A(io_bp_0_address[28]),
    .ZN(_0082_)
  );
  INV_X1 _0589_ (
    .A(io_bp_0_address[29]),
    .ZN(_0083_)
  );
  INV_X1 _0590_ (
    .A(io_bp_0_address[30]),
    .ZN(_0084_)
  );
  INV_X1 _0591_ (
    .A(io_bp_0_address[31]),
    .ZN(_0085_)
  );
  INV_X1 _0592_ (
    .A(io_bp_0_control_tmatch[0]),
    .ZN(_0086_)
  );
  AND2_X1 _0593_ (
    .A1(io_pc[31]),
    .A2(_0085_),
    .ZN(_0087_)
  );
  OR2_X1 _0594_ (
    .A1(_0056_),
    .A2(io_bp_0_address[31]),
    .ZN(_0088_)
  );
  AND2_X1 _0595_ (
    .A1(io_pc[30]),
    .A2(_0084_),
    .ZN(_0089_)
  );
  OR2_X1 _0596_ (
    .A1(_0055_),
    .A2(io_bp_0_address[30]),
    .ZN(_0090_)
  );
  AND2_X1 _0597_ (
    .A1(_0088_),
    .A2(_0090_),
    .ZN(_0091_)
  );
  OR2_X1 _0598_ (
    .A1(_0087_),
    .A2(_0089_),
    .ZN(_0092_)
  );
  AND2_X1 _0599_ (
    .A1(_0055_),
    .A2(io_bp_0_address[30]),
    .ZN(_0093_)
  );
  AND2_X1 _0600_ (
    .A1(_0056_),
    .A2(io_bp_0_address[31]),
    .ZN(_0094_)
  );
  AND2_X1 _0601_ (
    .A1(_0054_),
    .A2(io_bp_0_address[29]),
    .ZN(_0095_)
  );
  OR2_X1 _0602_ (
    .A1(_0053_),
    .A2(io_bp_0_address[28]),
    .ZN(_0096_)
  );
  OR2_X1 _0603_ (
    .A1(_0054_),
    .A2(io_bp_0_address[29]),
    .ZN(_0097_)
  );
  OR2_X1 _0604_ (
    .A1(_0093_),
    .A2(_0094_),
    .ZN(_0098_)
  );
  OR2_X1 _0605_ (
    .A1(_0092_),
    .A2(_0098_),
    .ZN(_0099_)
  );
  XOR2_X1 _0606_ (
    .A(io_pc[28]),
    .B(io_bp_0_address[28]),
    .Z(_0100_)
  );
  XOR2_X1 _0607_ (
    .A(io_pc[29]),
    .B(io_bp_0_address[29]),
    .Z(_0101_)
  );
  OR2_X1 _0608_ (
    .A1(_0100_),
    .A2(_0101_),
    .ZN(_0102_)
  );
  OR2_X1 _0609_ (
    .A1(_0099_),
    .A2(_0102_),
    .ZN(_0103_)
  );
  AND2_X1 _0610_ (
    .A1(io_pc[17]),
    .A2(_0073_),
    .ZN(_0104_)
  );
  OR2_X1 _0611_ (
    .A1(_0042_),
    .A2(io_bp_0_address[17]),
    .ZN(_0105_)
  );
  AND2_X1 _0612_ (
    .A1(_0041_),
    .A2(io_bp_0_address[16]),
    .ZN(_0106_)
  );
  OR2_X1 _0613_ (
    .A1(_0104_),
    .A2(_0106_),
    .ZN(_0107_)
  );
  AND2_X1 _0614_ (
    .A1(io_pc[16]),
    .A2(_0072_),
    .ZN(_0108_)
  );
  OR2_X1 _0615_ (
    .A1(_0041_),
    .A2(io_bp_0_address[16]),
    .ZN(_0109_)
  );
  AND2_X1 _0616_ (
    .A1(_0045_),
    .A2(io_bp_0_address[20]),
    .ZN(_0110_)
  );
  AND2_X1 _0617_ (
    .A1(_0046_),
    .A2(io_bp_0_address[21]),
    .ZN(_0111_)
  );
  AND2_X1 _0618_ (
    .A1(_0047_),
    .A2(io_bp_0_address[22]),
    .ZN(_0112_)
  );
  OR2_X1 _0619_ (
    .A1(_0111_),
    .A2(_0112_),
    .ZN(_0113_)
  );
  OR2_X1 _0620_ (
    .A1(_0048_),
    .A2(io_bp_0_address[23]),
    .ZN(_0114_)
  );
  OR2_X1 _0621_ (
    .A1(_0047_),
    .A2(io_bp_0_address[22]),
    .ZN(_0115_)
  );
  AND2_X1 _0622_ (
    .A1(_0114_),
    .A2(_0115_),
    .ZN(_0116_)
  );
  OR2_X1 _0623_ (
    .A1(_0044_),
    .A2(io_bp_0_address[19]),
    .ZN(_0117_)
  );
  AND2_X1 _0624_ (
    .A1(_0044_),
    .A2(io_bp_0_address[19]),
    .ZN(_0118_)
  );
  XOR2_X1 _0625_ (
    .A(io_pc[19]),
    .B(io_bp_0_address[19]),
    .Z(_0119_)
  );
  OR2_X1 _0626_ (
    .A1(_0043_),
    .A2(io_bp_0_address[18]),
    .ZN(_0120_)
  );
  XOR2_X1 _0627_ (
    .A(io_pc[18]),
    .B(io_bp_0_address[18]),
    .Z(_0121_)
  );
  OR2_X1 _0628_ (
    .A1(_0119_),
    .A2(_0121_),
    .ZN(_0122_)
  );
  AND2_X1 _0629_ (
    .A1(_0048_),
    .A2(io_bp_0_address[23]),
    .ZN(_0123_)
  );
  AND2_X1 _0630_ (
    .A1(io_pc[21]),
    .A2(_0075_),
    .ZN(_0124_)
  );
  OR2_X1 _0631_ (
    .A1(_0046_),
    .A2(io_bp_0_address[21]),
    .ZN(_0125_)
  );
  AND2_X1 _0632_ (
    .A1(_0042_),
    .A2(io_bp_0_address[17]),
    .ZN(_0126_)
  );
  OR2_X1 _0633_ (
    .A1(_0045_),
    .A2(io_bp_0_address[20]),
    .ZN(_0127_)
  );
  OR2_X1 _0634_ (
    .A1(_0107_),
    .A2(_0122_),
    .ZN(_0128_)
  );
  XOR2_X1 _0635_ (
    .A(io_pc[23]),
    .B(io_bp_0_address[23]),
    .Z(_0129_)
  );
  XOR2_X1 _0636_ (
    .A(io_pc[22]),
    .B(io_bp_0_address[22]),
    .Z(_0130_)
  );
  OR2_X1 _0637_ (
    .A1(_0129_),
    .A2(_0130_),
    .ZN(_0131_)
  );
  OR2_X1 _0638_ (
    .A1(_0111_),
    .A2(_0131_),
    .ZN(_0132_)
  );
  OR2_X1 _0639_ (
    .A1(_0108_),
    .A2(_0126_),
    .ZN(_0133_)
  );
  XOR2_X1 _0640_ (
    .A(io_pc[20]),
    .B(io_bp_0_address[20]),
    .Z(_0134_)
  );
  OR2_X1 _0641_ (
    .A1(_0124_),
    .A2(_0134_),
    .ZN(_0135_)
  );
  OR2_X1 _0642_ (
    .A1(_0133_),
    .A2(_0135_),
    .ZN(_0136_)
  );
  OR2_X1 _0643_ (
    .A1(_0132_),
    .A2(_0136_),
    .ZN(_0137_)
  );
  OR2_X1 _0644_ (
    .A1(_0128_),
    .A2(_0137_),
    .ZN(_0138_)
  );
  OR2_X1 _0645_ (
    .A1(_0052_),
    .A2(io_bp_0_address[27]),
    .ZN(_0139_)
  );
  AND2_X1 _0646_ (
    .A1(_0052_),
    .A2(io_bp_0_address[27]),
    .ZN(_0140_)
  );
  XOR2_X1 _0647_ (
    .A(io_pc[27]),
    .B(io_bp_0_address[27]),
    .Z(_0141_)
  );
  OR2_X1 _0648_ (
    .A1(_0051_),
    .A2(io_bp_0_address[26]),
    .ZN(_0142_)
  );
  XOR2_X1 _0649_ (
    .A(io_pc[26]),
    .B(io_bp_0_address[26]),
    .Z(_0143_)
  );
  OR2_X1 _0650_ (
    .A1(_0141_),
    .A2(_0143_),
    .ZN(_0144_)
  );
  AND2_X1 _0651_ (
    .A1(_0050_),
    .A2(io_bp_0_address[25]),
    .ZN(_0145_)
  );
  AND2_X1 _0652_ (
    .A1(_0049_),
    .A2(io_bp_0_address[24]),
    .ZN(_0146_)
  );
  OR2_X1 _0653_ (
    .A1(_0145_),
    .A2(_0146_),
    .ZN(_0147_)
  );
  AND2_X1 _0654_ (
    .A1(io_pc[25]),
    .A2(_0079_),
    .ZN(_0148_)
  );
  OR2_X1 _0655_ (
    .A1(_0050_),
    .A2(io_bp_0_address[25]),
    .ZN(_0149_)
  );
  AND2_X1 _0656_ (
    .A1(io_pc[24]),
    .A2(_0078_),
    .ZN(_0150_)
  );
  OR2_X1 _0657_ (
    .A1(_0049_),
    .A2(io_bp_0_address[24]),
    .ZN(_0151_)
  );
  AND2_X1 _0658_ (
    .A1(_0149_),
    .A2(_0151_),
    .ZN(_0152_)
  );
  OR2_X1 _0659_ (
    .A1(_0148_),
    .A2(_0150_),
    .ZN(_0153_)
  );
  OR2_X1 _0660_ (
    .A1(_0147_),
    .A2(_0153_),
    .ZN(_0154_)
  );
  OR2_X1 _0661_ (
    .A1(_0144_),
    .A2(_0154_),
    .ZN(_0155_)
  );
  OR2_X1 _0662_ (
    .A1(_0103_),
    .A2(_0155_),
    .ZN(_0156_)
  );
  OR2_X1 _0663_ (
    .A1(_0138_),
    .A2(_0156_),
    .ZN(_0157_)
  );
  AND2_X1 _0664_ (
    .A1(io_pc[5]),
    .A2(_0063_),
    .ZN(_0158_)
  );
  OR2_X1 _0665_ (
    .A1(_0030_),
    .A2(io_bp_0_address[5]),
    .ZN(_0159_)
  );
  AND2_X1 _0666_ (
    .A1(io_pc[6]),
    .A2(_0064_),
    .ZN(_0160_)
  );
  OR2_X1 _0667_ (
    .A1(_0031_),
    .A2(io_bp_0_address[6]),
    .ZN(_0161_)
  );
  AND2_X1 _0668_ (
    .A1(_0159_),
    .A2(_0161_),
    .ZN(_0162_)
  );
  OR2_X1 _0669_ (
    .A1(_0158_),
    .A2(_0160_),
    .ZN(_0163_)
  );
  AND2_X1 _0670_ (
    .A1(_0032_),
    .A2(io_bp_0_address[7]),
    .ZN(_0164_)
  );
  AND2_X1 _0671_ (
    .A1(_0031_),
    .A2(io_bp_0_address[6]),
    .ZN(_0165_)
  );
  OR2_X1 _0672_ (
    .A1(_0164_),
    .A2(_0165_),
    .ZN(_0166_)
  );
  AND2_X1 _0673_ (
    .A1(_0030_),
    .A2(io_bp_0_address[5]),
    .ZN(_0167_)
  );
  AND2_X1 _0674_ (
    .A1(_0029_),
    .A2(io_bp_0_address[4]),
    .ZN(_0168_)
  );
  OR2_X1 _0675_ (
    .A1(_0167_),
    .A2(_0168_),
    .ZN(_0169_)
  );
  OR2_X1 _0676_ (
    .A1(_0166_),
    .A2(_0169_),
    .ZN(_0170_)
  );
  OR2_X1 _0677_ (
    .A1(_0163_),
    .A2(_0170_),
    .ZN(_0171_)
  );
  AND2_X1 _0678_ (
    .A1(_0025_),
    .A2(io_bp_0_address[0]),
    .ZN(_0172_)
  );
  XOR2_X1 _0679_ (
    .A(io_pc[0]),
    .B(io_bp_0_address[0]),
    .Z(_0173_)
  );
  AND2_X1 _0680_ (
    .A1(_0086_),
    .A2(_0173_),
    .ZN(_0174_)
  );
  AND2_X1 _0681_ (
    .A1(io_pc[4]),
    .A2(_0062_),
    .ZN(_0175_)
  );
  OR2_X1 _0682_ (
    .A1(_0029_),
    .A2(io_bp_0_address[4]),
    .ZN(_0176_)
  );
  AND2_X1 _0683_ (
    .A1(io_pc[7]),
    .A2(_0065_),
    .ZN(_0177_)
  );
  OR2_X1 _0684_ (
    .A1(_0032_),
    .A2(io_bp_0_address[7]),
    .ZN(_0178_)
  );
  OR2_X1 _0685_ (
    .A1(io_bp_0_control_tmatch[1]),
    .A2(_0177_),
    .ZN(_0179_)
  );
  OR2_X1 _0686_ (
    .A1(_0175_),
    .A2(_0179_),
    .ZN(_0180_)
  );
  OR2_X1 _0687_ (
    .A1(_0174_),
    .A2(_0180_),
    .ZN(_0181_)
  );
  OR2_X1 _0688_ (
    .A1(_0171_),
    .A2(_0181_),
    .ZN(_0182_)
  );
  OR2_X1 _0689_ (
    .A1(_0036_),
    .A2(io_bp_0_address[11]),
    .ZN(_0183_)
  );
  OR2_X1 _0690_ (
    .A1(_0035_),
    .A2(io_bp_0_address[10]),
    .ZN(_0184_)
  );
  AND2_X1 _0691_ (
    .A1(_0183_),
    .A2(_0184_),
    .ZN(_0185_)
  );
  AND2_X1 _0692_ (
    .A1(_0036_),
    .A2(io_bp_0_address[11]),
    .ZN(_0186_)
  );
  XOR2_X1 _0693_ (
    .A(io_pc[11]),
    .B(io_bp_0_address[11]),
    .Z(_0187_)
  );
  XOR2_X1 _0694_ (
    .A(io_pc[10]),
    .B(io_bp_0_address[10]),
    .Z(_0188_)
  );
  OR2_X1 _0695_ (
    .A1(_0187_),
    .A2(_0188_),
    .ZN(_0189_)
  );
  AND2_X1 _0696_ (
    .A1(_0034_),
    .A2(io_bp_0_address[9]),
    .ZN(_0190_)
  );
  AND2_X1 _0697_ (
    .A1(_0033_),
    .A2(io_bp_0_address[8]),
    .ZN(_0191_)
  );
  OR2_X1 _0698_ (
    .A1(_0190_),
    .A2(_0191_),
    .ZN(_0192_)
  );
  AND2_X1 _0699_ (
    .A1(io_pc[9]),
    .A2(_0067_),
    .ZN(_0193_)
  );
  OR2_X1 _0700_ (
    .A1(_0034_),
    .A2(io_bp_0_address[9]),
    .ZN(_0194_)
  );
  AND2_X1 _0701_ (
    .A1(io_pc[8]),
    .A2(_0066_),
    .ZN(_0195_)
  );
  OR2_X1 _0702_ (
    .A1(_0033_),
    .A2(io_bp_0_address[8]),
    .ZN(_0196_)
  );
  AND2_X1 _0703_ (
    .A1(_0194_),
    .A2(_0196_),
    .ZN(_0197_)
  );
  OR2_X1 _0704_ (
    .A1(_0193_),
    .A2(_0195_),
    .ZN(_0198_)
  );
  OR2_X1 _0705_ (
    .A1(_0192_),
    .A2(_0198_),
    .ZN(_0199_)
  );
  OR2_X1 _0706_ (
    .A1(_0189_),
    .A2(_0199_),
    .ZN(_0200_)
  );
  AND2_X1 _0707_ (
    .A1(io_bp_0_address[0]),
    .A2(io_bp_0_control_tmatch[0]),
    .ZN(_0201_)
  );
  INV_X1 _0708_ (
    .A(_0201_),
    .ZN(_0202_)
  );
  AND2_X1 _0709_ (
    .A1(io_bp_0_address[1]),
    .A2(_0201_),
    .ZN(_0203_)
  );
  INV_X1 _0710_ (
    .A(_0203_),
    .ZN(_0204_)
  );
  AND2_X1 _0711_ (
    .A1(io_bp_0_address[2]),
    .A2(_0203_),
    .ZN(_0205_)
  );
  INV_X1 _0712_ (
    .A(_0205_),
    .ZN(_0206_)
  );
  AND2_X1 _0713_ (
    .A1(_0028_),
    .A2(io_bp_0_address[3]),
    .ZN(_0207_)
  );
  OR2_X1 _0714_ (
    .A1(_0028_),
    .A2(io_bp_0_address[3]),
    .ZN(_0208_)
  );
  XOR2_X1 _0715_ (
    .A(io_pc[3]),
    .B(io_bp_0_address[3]),
    .Z(_0209_)
  );
  AND2_X1 _0716_ (
    .A1(_0206_),
    .A2(_0209_),
    .ZN(_0210_)
  );
  OR2_X1 _0717_ (
    .A1(_0200_),
    .A2(_0210_),
    .ZN(_0211_)
  );
  OR2_X1 _0718_ (
    .A1(_0182_),
    .A2(_0211_),
    .ZN(_0212_)
  );
  AND2_X1 _0719_ (
    .A1(_0040_),
    .A2(io_bp_0_address[15]),
    .ZN(_0213_)
  );
  OR2_X1 _0720_ (
    .A1(_0039_),
    .A2(io_bp_0_address[14]),
    .ZN(_0214_)
  );
  AND2_X1 _0721_ (
    .A1(_0038_),
    .A2(io_bp_0_address[13]),
    .ZN(_0215_)
  );
  OR2_X1 _0722_ (
    .A1(_0040_),
    .A2(io_bp_0_address[15]),
    .ZN(_0216_)
  );
  XOR2_X1 _0723_ (
    .A(io_pc[14]),
    .B(io_bp_0_address[14]),
    .Z(_0217_)
  );
  XOR2_X1 _0724_ (
    .A(io_pc[15]),
    .B(io_bp_0_address[15]),
    .Z(_0218_)
  );
  OR2_X1 _0725_ (
    .A1(_0217_),
    .A2(_0218_),
    .ZN(_0219_)
  );
  OR2_X1 _0726_ (
    .A1(_0215_),
    .A2(_0219_),
    .ZN(_0220_)
  );
  AND2_X1 _0727_ (
    .A1(io_pc[13]),
    .A2(_0069_),
    .ZN(_0221_)
  );
  OR2_X1 _0728_ (
    .A1(_0038_),
    .A2(io_bp_0_address[13]),
    .ZN(_0222_)
  );
  OR2_X1 _0729_ (
    .A1(_0037_),
    .A2(io_bp_0_address[12]),
    .ZN(_0223_)
  );
  AND2_X1 _0730_ (
    .A1(_0222_),
    .A2(_0223_),
    .ZN(_0224_)
  );
  XOR2_X1 _0731_ (
    .A(io_pc[12]),
    .B(io_bp_0_address[12]),
    .Z(_0225_)
  );
  OR2_X1 _0732_ (
    .A1(_0221_),
    .A2(_0225_),
    .ZN(_0226_)
  );
  OR2_X1 _0733_ (
    .A1(_0220_),
    .A2(_0226_),
    .ZN(_0227_)
  );
  OR2_X1 _0734_ (
    .A1(_0026_),
    .A2(io_bp_0_address[1]),
    .ZN(_0228_)
  );
  AND2_X1 _0735_ (
    .A1(_0026_),
    .A2(io_bp_0_address[1]),
    .ZN(_0229_)
  );
  XOR2_X1 _0736_ (
    .A(io_pc[1]),
    .B(io_bp_0_address[1]),
    .Z(_0230_)
  );
  AND2_X1 _0737_ (
    .A1(_0202_),
    .A2(_0230_),
    .ZN(_0231_)
  );
  AND2_X1 _0738_ (
    .A1(_0027_),
    .A2(io_bp_0_address[2]),
    .ZN(_0232_)
  );
  OR2_X1 _0739_ (
    .A1(_0027_),
    .A2(io_bp_0_address[2]),
    .ZN(_0233_)
  );
  XOR2_X1 _0740_ (
    .A(io_pc[2]),
    .B(io_bp_0_address[2]),
    .Z(_0234_)
  );
  OR2_X1 _0741_ (
    .A1(_0231_),
    .A2(_0234_),
    .ZN(_0235_)
  );
  AND2_X1 _0742_ (
    .A1(_0204_),
    .A2(_0235_),
    .ZN(_0236_)
  );
  OR2_X1 _0743_ (
    .A1(_0227_),
    .A2(_0236_),
    .ZN(_0237_)
  );
  OR2_X1 _0744_ (
    .A1(_0212_),
    .A2(_0237_),
    .ZN(_0238_)
  );
  OR2_X1 _0745_ (
    .A1(_0157_),
    .A2(_0238_),
    .ZN(_0239_)
  );
  INV_X1 _0746_ (
    .A(_0239_),
    .ZN(_0240_)
  );
  AND2_X1 _0747_ (
    .A1(_0172_),
    .A2(_0228_),
    .ZN(_0241_)
  );
  OR2_X1 _0748_ (
    .A1(_0229_),
    .A2(_0232_),
    .ZN(_0242_)
  );
  OR2_X1 _0749_ (
    .A1(_0241_),
    .A2(_0242_),
    .ZN(_0243_)
  );
  AND2_X1 _0750_ (
    .A1(_0208_),
    .A2(_0233_),
    .ZN(_0244_)
  );
  AND2_X1 _0751_ (
    .A1(_0243_),
    .A2(_0244_),
    .ZN(_0245_)
  );
  OR2_X1 _0752_ (
    .A1(_0207_),
    .A2(_0245_),
    .ZN(_0246_)
  );
  AND2_X1 _0753_ (
    .A1(_0176_),
    .A2(_0246_),
    .ZN(_0247_)
  );
  OR2_X1 _0754_ (
    .A1(_0169_),
    .A2(_0247_),
    .ZN(_0248_)
  );
  AND2_X1 _0755_ (
    .A1(_0162_),
    .A2(_0248_),
    .ZN(_0249_)
  );
  OR2_X1 _0756_ (
    .A1(_0166_),
    .A2(_0249_),
    .ZN(_0250_)
  );
  AND2_X1 _0757_ (
    .A1(_0178_),
    .A2(_0250_),
    .ZN(_0251_)
  );
  OR2_X1 _0758_ (
    .A1(_0200_),
    .A2(_0251_),
    .ZN(_0252_)
  );
  OR2_X1 _0759_ (
    .A1(_0185_),
    .A2(_0186_),
    .ZN(_0253_)
  );
  OR2_X1 _0760_ (
    .A1(_0190_),
    .A2(_0197_),
    .ZN(_0254_)
  );
  OR2_X1 _0761_ (
    .A1(_0189_),
    .A2(_0254_),
    .ZN(_0255_)
  );
  AND2_X1 _0762_ (
    .A1(_0253_),
    .A2(_0255_),
    .ZN(_0256_)
  );
  AND2_X1 _0763_ (
    .A1(_0252_),
    .A2(_0256_),
    .ZN(_0257_)
  );
  OR2_X1 _0764_ (
    .A1(_0227_),
    .A2(_0257_),
    .ZN(_0258_)
  );
  OR2_X1 _0765_ (
    .A1(_0220_),
    .A2(_0224_),
    .ZN(_0259_)
  );
  OR2_X1 _0766_ (
    .A1(_0213_),
    .A2(_0214_),
    .ZN(_0260_)
  );
  AND2_X1 _0767_ (
    .A1(_0216_),
    .A2(_0260_),
    .ZN(_0261_)
  );
  AND2_X1 _0768_ (
    .A1(_0259_),
    .A2(_0261_),
    .ZN(_0262_)
  );
  AND2_X1 _0769_ (
    .A1(_0258_),
    .A2(_0262_),
    .ZN(_0263_)
  );
  OR2_X1 _0770_ (
    .A1(_0157_),
    .A2(_0263_),
    .ZN(_0264_)
  );
  AND2_X1 _0771_ (
    .A1(_0139_),
    .A2(_0142_),
    .ZN(_0265_)
  );
  OR2_X1 _0772_ (
    .A1(_0140_),
    .A2(_0265_),
    .ZN(_0266_)
  );
  OR2_X1 _0773_ (
    .A1(_0145_),
    .A2(_0152_),
    .ZN(_0267_)
  );
  OR2_X1 _0774_ (
    .A1(_0144_),
    .A2(_0267_),
    .ZN(_0268_)
  );
  AND2_X1 _0775_ (
    .A1(_0266_),
    .A2(_0268_),
    .ZN(_0269_)
  );
  OR2_X1 _0776_ (
    .A1(_0109_),
    .A2(_0126_),
    .ZN(_0270_)
  );
  AND2_X1 _0777_ (
    .A1(_0105_),
    .A2(_0270_),
    .ZN(_0271_)
  );
  OR2_X1 _0778_ (
    .A1(_0122_),
    .A2(_0271_),
    .ZN(_0272_)
  );
  OR2_X1 _0779_ (
    .A1(_0118_),
    .A2(_0120_),
    .ZN(_0273_)
  );
  AND2_X1 _0780_ (
    .A1(_0117_),
    .A2(_0127_),
    .ZN(_0274_)
  );
  AND2_X1 _0781_ (
    .A1(_0273_),
    .A2(_0274_),
    .ZN(_0275_)
  );
  AND2_X1 _0782_ (
    .A1(_0272_),
    .A2(_0275_),
    .ZN(_0276_)
  );
  OR2_X1 _0783_ (
    .A1(_0110_),
    .A2(_0276_),
    .ZN(_0277_)
  );
  AND2_X1 _0784_ (
    .A1(_0125_),
    .A2(_0277_),
    .ZN(_0278_)
  );
  OR2_X1 _0785_ (
    .A1(_0113_),
    .A2(_0278_),
    .ZN(_0279_)
  );
  AND2_X1 _0786_ (
    .A1(_0116_),
    .A2(_0279_),
    .ZN(_0280_)
  );
  OR2_X1 _0787_ (
    .A1(_0095_),
    .A2(_0096_),
    .ZN(_0281_)
  );
  AND2_X1 _0788_ (
    .A1(_0097_),
    .A2(_0281_),
    .ZN(_0282_)
  );
  OR2_X1 _0789_ (
    .A1(_0099_),
    .A2(_0282_),
    .ZN(_0283_)
  );
  OR2_X1 _0790_ (
    .A1(_0091_),
    .A2(_0094_),
    .ZN(_0284_)
  );
  OR2_X1 _0791_ (
    .A1(_0103_),
    .A2(_0269_),
    .ZN(_0285_)
  );
  AND2_X1 _0792_ (
    .A1(_0283_),
    .A2(_0285_),
    .ZN(_0286_)
  );
  OR2_X1 _0793_ (
    .A1(_0123_),
    .A2(_0156_),
    .ZN(_0287_)
  );
  OR2_X1 _0794_ (
    .A1(_0280_),
    .A2(_0287_),
    .ZN(_0288_)
  );
  AND2_X1 _0795_ (
    .A1(_0284_),
    .A2(_0288_),
    .ZN(_0289_)
  );
  AND2_X1 _0796_ (
    .A1(_0286_),
    .A2(_0289_),
    .ZN(_0290_)
  );
  AND2_X1 _0797_ (
    .A1(_0264_),
    .A2(_0290_),
    .ZN(_0291_)
  );
  XOR2_X1 _0798_ (
    .A(_0086_),
    .B(_0291_),
    .Z(_0292_)
  );
  AND2_X1 _0799_ (
    .A1(io_bp_0_control_tmatch[1]),
    .A2(_0292_),
    .ZN(_0293_)
  );
  OR2_X1 _0800_ (
    .A1(_0240_),
    .A2(_0293_),
    .ZN(_0294_)
  );
  AND2_X1 _0801_ (
    .A1(_0001_),
    .A2(io_bp_0_control_x),
    .ZN(_0295_)
  );
  AND2_X1 _0802_ (
    .A1(_0294_),
    .A2(_0295_),
    .ZN(_0296_)
  );
  AND2_X1 _0803_ (
    .A1(_0057_),
    .A2(_0296_),
    .ZN(io_xcpt_if)
  );
  AND2_X1 _0804_ (
    .A1(io_ea[31]),
    .A2(_0085_),
    .ZN(_0297_)
  );
  OR2_X1 _0805_ (
    .A1(_0024_),
    .A2(io_bp_0_address[31]),
    .ZN(_0298_)
  );
  AND2_X1 _0806_ (
    .A1(io_ea[28]),
    .A2(_0082_),
    .ZN(_0299_)
  );
  OR2_X1 _0807_ (
    .A1(_0021_),
    .A2(io_bp_0_address[28]),
    .ZN(_0300_)
  );
  AND2_X1 _0808_ (
    .A1(_0298_),
    .A2(_0300_),
    .ZN(_0301_)
  );
  AND2_X1 _0809_ (
    .A1(io_ea[30]),
    .A2(_0084_),
    .ZN(_0302_)
  );
  OR2_X1 _0810_ (
    .A1(_0023_),
    .A2(io_bp_0_address[30]),
    .ZN(_0303_)
  );
  OR2_X1 _0811_ (
    .A1(io_ea[25]),
    .A2(_0079_),
    .ZN(_0304_)
  );
  AND2_X1 _0812_ (
    .A1(_0303_),
    .A2(_0304_),
    .ZN(_0305_)
  );
  AND2_X1 _0813_ (
    .A1(_0301_),
    .A2(_0305_),
    .ZN(_0306_)
  );
  OR2_X1 _0814_ (
    .A1(io_ea[31]),
    .A2(_0085_),
    .ZN(_0307_)
  );
  OR2_X1 _0815_ (
    .A1(io_ea[30]),
    .A2(_0084_),
    .ZN(_0308_)
  );
  AND2_X1 _0816_ (
    .A1(_0307_),
    .A2(_0308_),
    .ZN(_0309_)
  );
  OR2_X1 _0817_ (
    .A1(io_ea[29]),
    .A2(_0083_),
    .ZN(_0310_)
  );
  OR2_X1 _0818_ (
    .A1(io_ea[28]),
    .A2(_0082_),
    .ZN(_0311_)
  );
  AND2_X1 _0819_ (
    .A1(_0310_),
    .A2(_0311_),
    .ZN(_0312_)
  );
  AND2_X1 _0820_ (
    .A1(_0309_),
    .A2(_0312_),
    .ZN(_0313_)
  );
  AND2_X1 _0821_ (
    .A1(_0306_),
    .A2(_0313_),
    .ZN(_0314_)
  );
  AND2_X1 _0822_ (
    .A1(io_ea[27]),
    .A2(_0081_),
    .ZN(_0315_)
  );
  OR2_X1 _0823_ (
    .A1(io_ea[27]),
    .A2(_0081_),
    .ZN(_0316_)
  );
  XOR2_X1 _0824_ (
    .A(io_ea[27]),
    .B(io_bp_0_address[27]),
    .Z(_0317_)
  );
  AND2_X1 _0825_ (
    .A1(io_ea[26]),
    .A2(_0080_),
    .ZN(_0318_)
  );
  XOR2_X1 _0826_ (
    .A(io_ea[26]),
    .B(io_bp_0_address[26]),
    .Z(_0319_)
  );
  OR2_X1 _0827_ (
    .A1(_0317_),
    .A2(_0319_),
    .ZN(_0320_)
  );
  INV_X1 _0828_ (
    .A(_0320_),
    .ZN(_0321_)
  );
  OR2_X1 _0829_ (
    .A1(io_ea[24]),
    .A2(_0078_),
    .ZN(_0322_)
  );
  AND2_X1 _0830_ (
    .A1(io_ea[25]),
    .A2(_0079_),
    .ZN(_0323_)
  );
  OR2_X1 _0831_ (
    .A1(_0020_),
    .A2(io_bp_0_address[25]),
    .ZN(_0324_)
  );
  AND2_X1 _0832_ (
    .A1(_0322_),
    .A2(_0324_),
    .ZN(_0325_)
  );
  AND2_X1 _0833_ (
    .A1(io_ea[29]),
    .A2(_0083_),
    .ZN(_0326_)
  );
  OR2_X1 _0834_ (
    .A1(_0022_),
    .A2(io_bp_0_address[29]),
    .ZN(_0327_)
  );
  AND2_X1 _0835_ (
    .A1(io_ea[24]),
    .A2(_0078_),
    .ZN(_0328_)
  );
  OR2_X1 _0836_ (
    .A1(_0019_),
    .A2(io_bp_0_address[24]),
    .ZN(_0329_)
  );
  AND2_X1 _0837_ (
    .A1(_0327_),
    .A2(_0329_),
    .ZN(_0330_)
  );
  AND2_X1 _0838_ (
    .A1(_0325_),
    .A2(_0330_),
    .ZN(_0331_)
  );
  AND2_X1 _0839_ (
    .A1(_0321_),
    .A2(_0331_),
    .ZN(_0332_)
  );
  AND2_X1 _0840_ (
    .A1(_0314_),
    .A2(_0332_),
    .ZN(_0333_)
  );
  OR2_X1 _0841_ (
    .A1(io_ea[22]),
    .A2(_0076_),
    .ZN(_0334_)
  );
  OR2_X1 _0842_ (
    .A1(io_ea[21]),
    .A2(_0075_),
    .ZN(_0335_)
  );
  AND2_X1 _0843_ (
    .A1(_0334_),
    .A2(_0335_),
    .ZN(_0336_)
  );
  AND2_X1 _0844_ (
    .A1(io_ea[21]),
    .A2(_0075_),
    .ZN(_0337_)
  );
  OR2_X1 _0845_ (
    .A1(_0016_),
    .A2(io_bp_0_address[21]),
    .ZN(_0338_)
  );
  AND2_X1 _0846_ (
    .A1(io_ea[23]),
    .A2(_0077_),
    .ZN(_0339_)
  );
  OR2_X1 _0847_ (
    .A1(_0018_),
    .A2(io_bp_0_address[23]),
    .ZN(_0340_)
  );
  AND2_X1 _0848_ (
    .A1(io_ea[22]),
    .A2(_0076_),
    .ZN(_0341_)
  );
  OR2_X1 _0849_ (
    .A1(_0017_),
    .A2(io_bp_0_address[22]),
    .ZN(_0342_)
  );
  AND2_X1 _0850_ (
    .A1(_0340_),
    .A2(_0342_),
    .ZN(_0343_)
  );
  OR2_X1 _0851_ (
    .A1(_0339_),
    .A2(_0341_),
    .ZN(_0344_)
  );
  OR2_X1 _0852_ (
    .A1(_0012_),
    .A2(io_bp_0_address[17]),
    .ZN(_0345_)
  );
  OR2_X1 _0853_ (
    .A1(_0011_),
    .A2(io_bp_0_address[16]),
    .ZN(_0346_)
  );
  AND2_X1 _0854_ (
    .A1(_0345_),
    .A2(_0346_),
    .ZN(_0347_)
  );
  OR2_X1 _0855_ (
    .A1(_0014_),
    .A2(io_bp_0_address[19]),
    .ZN(_0348_)
  );
  OR2_X1 _0856_ (
    .A1(_0013_),
    .A2(io_bp_0_address[18]),
    .ZN(_0349_)
  );
  AND2_X1 _0857_ (
    .A1(_0348_),
    .A2(_0349_),
    .ZN(_0350_)
  );
  AND2_X1 _0858_ (
    .A1(_0014_),
    .A2(io_bp_0_address[19]),
    .ZN(_0351_)
  );
  XOR2_X1 _0859_ (
    .A(io_ea[19]),
    .B(io_bp_0_address[19]),
    .Z(_0352_)
  );
  XOR2_X1 _0860_ (
    .A(io_ea[18]),
    .B(io_bp_0_address[18]),
    .Z(_0353_)
  );
  OR2_X1 _0861_ (
    .A1(_0352_),
    .A2(_0353_),
    .ZN(_0354_)
  );
  OR2_X1 _0862_ (
    .A1(io_ea[23]),
    .A2(_0077_),
    .ZN(_0355_)
  );
  OR2_X1 _0863_ (
    .A1(_0015_),
    .A2(io_bp_0_address[20]),
    .ZN(_0356_)
  );
  AND2_X1 _0864_ (
    .A1(_0355_),
    .A2(_0356_),
    .ZN(_0357_)
  );
  OR2_X1 _0865_ (
    .A1(io_ea[20]),
    .A2(_0074_),
    .ZN(_0358_)
  );
  AND2_X1 _0866_ (
    .A1(_0012_),
    .A2(io_bp_0_address[17]),
    .ZN(_0359_)
  );
  AND2_X1 _0867_ (
    .A1(_0338_),
    .A2(_0358_),
    .ZN(_0360_)
  );
  AND2_X1 _0868_ (
    .A1(_0357_),
    .A2(_0360_),
    .ZN(_0361_)
  );
  AND2_X1 _0869_ (
    .A1(_0336_),
    .A2(_0361_),
    .ZN(_0362_)
  );
  AND2_X1 _0870_ (
    .A1(_0343_),
    .A2(_0362_),
    .ZN(_0363_)
  );
  XOR2_X1 _0871_ (
    .A(io_ea[17]),
    .B(io_bp_0_address[17]),
    .Z(_0364_)
  );
  XOR2_X1 _0872_ (
    .A(io_ea[16]),
    .B(io_bp_0_address[16]),
    .Z(_0365_)
  );
  OR2_X1 _0873_ (
    .A1(_0354_),
    .A2(_0365_),
    .ZN(_0366_)
  );
  OR2_X1 _0874_ (
    .A1(_0364_),
    .A2(_0366_),
    .ZN(_0367_)
  );
  INV_X1 _0875_ (
    .A(_0367_),
    .ZN(_0368_)
  );
  AND2_X1 _0876_ (
    .A1(_0363_),
    .A2(_0368_),
    .ZN(_0369_)
  );
  AND2_X1 _0877_ (
    .A1(_0333_),
    .A2(_0369_),
    .ZN(_0370_)
  );
  AND2_X1 _0878_ (
    .A1(io_ea[14]),
    .A2(_0070_),
    .ZN(_0371_)
  );
  AND2_X1 _0879_ (
    .A1(_0006_),
    .A2(io_bp_0_address[9]),
    .ZN(_0372_)
  );
  OR2_X1 _0880_ (
    .A1(io_ea[13]),
    .A2(_0069_),
    .ZN(_0373_)
  );
  OR2_X1 _0881_ (
    .A1(_0009_),
    .A2(io_bp_0_address[12]),
    .ZN(_0374_)
  );
  OR2_X1 _0882_ (
    .A1(io_ea[15]),
    .A2(_0071_),
    .ZN(_0375_)
  );
  OR2_X1 _0883_ (
    .A1(io_ea[14]),
    .A2(_0070_),
    .ZN(_0376_)
  );
  AND2_X1 _0884_ (
    .A1(_0375_),
    .A2(_0376_),
    .ZN(_0377_)
  );
  AND2_X1 _0885_ (
    .A1(io_ea[15]),
    .A2(_0071_),
    .ZN(_0378_)
  );
  AND2_X1 _0886_ (
    .A1(io_ea[13]),
    .A2(_0069_),
    .ZN(_0379_)
  );
  OR2_X1 _0887_ (
    .A1(_0010_),
    .A2(io_bp_0_address[13]),
    .ZN(_0380_)
  );
  OR2_X1 _0888_ (
    .A1(_0008_),
    .A2(io_bp_0_address[11]),
    .ZN(_0381_)
  );
  AND2_X1 _0889_ (
    .A1(_0008_),
    .A2(io_bp_0_address[11]),
    .ZN(_0382_)
  );
  XOR2_X1 _0890_ (
    .A(io_ea[11]),
    .B(io_bp_0_address[11]),
    .Z(_0383_)
  );
  OR2_X1 _0891_ (
    .A1(_0007_),
    .A2(io_bp_0_address[10]),
    .ZN(_0384_)
  );
  XOR2_X1 _0892_ (
    .A(io_ea[10]),
    .B(io_bp_0_address[10]),
    .Z(_0385_)
  );
  OR2_X1 _0893_ (
    .A1(_0383_),
    .A2(_0385_),
    .ZN(_0386_)
  );
  AND2_X1 _0894_ (
    .A1(_0005_),
    .A2(io_bp_0_address[8]),
    .ZN(_0387_)
  );
  OR2_X1 _0895_ (
    .A1(_0006_),
    .A2(io_bp_0_address[9]),
    .ZN(_0388_)
  );
  OR2_X1 _0896_ (
    .A1(io_ea[12]),
    .A2(_0068_),
    .ZN(_0389_)
  );
  OR2_X1 _0897_ (
    .A1(_0005_),
    .A2(io_bp_0_address[8]),
    .ZN(_0390_)
  );
  OR2_X1 _0898_ (
    .A1(_0371_),
    .A2(_0387_),
    .ZN(_0391_)
  );
  XOR2_X1 _0899_ (
    .A(io_ea[9]),
    .B(io_bp_0_address[9]),
    .Z(_0392_)
  );
  OR2_X1 _0900_ (
    .A1(_0391_),
    .A2(_0392_),
    .ZN(_0393_)
  );
  OR2_X1 _0901_ (
    .A1(_0378_),
    .A2(_0393_),
    .ZN(_0394_)
  );
  XOR2_X1 _0902_ (
    .A(io_ea[12]),
    .B(io_bp_0_address[12]),
    .Z(_0395_)
  );
  OR2_X1 _0903_ (
    .A1(_0386_),
    .A2(_0395_),
    .ZN(_0396_)
  );
  OR2_X1 _0904_ (
    .A1(_0394_),
    .A2(_0396_),
    .ZN(_0397_)
  );
  INV_X1 _0905_ (
    .A(_0397_),
    .ZN(_0398_)
  );
  AND2_X1 _0906_ (
    .A1(_0380_),
    .A2(_0390_),
    .ZN(_0399_)
  );
  AND2_X1 _0907_ (
    .A1(_0373_),
    .A2(_0377_),
    .ZN(_0400_)
  );
  AND2_X1 _0908_ (
    .A1(_0399_),
    .A2(_0400_),
    .ZN(_0401_)
  );
  AND2_X1 _0909_ (
    .A1(_0398_),
    .A2(_0401_),
    .ZN(_0402_)
  );
  AND2_X1 _0910_ (
    .A1(io_ea[7]),
    .A2(_0065_),
    .ZN(_0403_)
  );
  OR2_X1 _0911_ (
    .A1(_0004_),
    .A2(io_bp_0_address[7]),
    .ZN(_0404_)
  );
  OR2_X1 _0912_ (
    .A1(io_ea[7]),
    .A2(_0065_),
    .ZN(_0405_)
  );
  OR2_X1 _0913_ (
    .A1(io_ea[6]),
    .A2(_0064_),
    .ZN(_0406_)
  );
  AND2_X1 _0914_ (
    .A1(_0405_),
    .A2(_0406_),
    .ZN(_0407_)
  );
  AND2_X1 _0915_ (
    .A1(io_ea[6]),
    .A2(_0064_),
    .ZN(_0408_)
  );
  OR2_X1 _0916_ (
    .A1(_0003_),
    .A2(io_bp_0_address[6]),
    .ZN(_0409_)
  );
  AND2_X1 _0917_ (
    .A1(io_ea[5]),
    .A2(_0063_),
    .ZN(_0410_)
  );
  OR2_X1 _0918_ (
    .A1(_0002_),
    .A2(io_bp_0_address[5]),
    .ZN(_0411_)
  );
  OR2_X1 _0919_ (
    .A1(_0408_),
    .A2(_0410_),
    .ZN(_0412_)
  );
  AND2_X1 _0920_ (
    .A1(io_ea[4]),
    .A2(_0062_),
    .ZN(_0413_)
  );
  OR2_X1 _0921_ (
    .A1(io_ea[3]),
    .A2(_0061_),
    .ZN(_0414_)
  );
  AND2_X1 _0922_ (
    .A1(io_ea[1]),
    .A2(_0059_),
    .ZN(_0415_)
  );
  OR2_X1 _0923_ (
    .A1(io_ea[0]),
    .A2(_0058_),
    .ZN(_0416_)
  );
  OR2_X1 _0924_ (
    .A1(_0415_),
    .A2(_0416_),
    .ZN(_0417_)
  );
  OR2_X1 _0925_ (
    .A1(io_ea[2]),
    .A2(_0060_),
    .ZN(_0418_)
  );
  OR2_X1 _0926_ (
    .A1(io_ea[1]),
    .A2(_0059_),
    .ZN(_0419_)
  );
  AND2_X1 _0927_ (
    .A1(_0418_),
    .A2(_0419_),
    .ZN(_0420_)
  );
  AND2_X1 _0928_ (
    .A1(_0417_),
    .A2(_0420_),
    .ZN(_0421_)
  );
  AND2_X1 _0929_ (
    .A1(io_ea[3]),
    .A2(_0061_),
    .ZN(_0422_)
  );
  AND2_X1 _0930_ (
    .A1(io_ea[2]),
    .A2(_0060_),
    .ZN(_0423_)
  );
  OR2_X1 _0931_ (
    .A1(_0422_),
    .A2(_0423_),
    .ZN(_0424_)
  );
  OR2_X1 _0932_ (
    .A1(_0421_),
    .A2(_0424_),
    .ZN(_0425_)
  );
  AND2_X1 _0933_ (
    .A1(_0414_),
    .A2(_0425_),
    .ZN(_0426_)
  );
  OR2_X1 _0934_ (
    .A1(_0413_),
    .A2(_0426_),
    .ZN(_0427_)
  );
  OR2_X1 _0935_ (
    .A1(io_ea[5]),
    .A2(_0063_),
    .ZN(_0428_)
  );
  OR2_X1 _0936_ (
    .A1(io_ea[4]),
    .A2(_0062_),
    .ZN(_0429_)
  );
  AND2_X1 _0937_ (
    .A1(_0428_),
    .A2(_0429_),
    .ZN(_0430_)
  );
  AND2_X1 _0938_ (
    .A1(_0427_),
    .A2(_0430_),
    .ZN(_0431_)
  );
  OR2_X1 _0939_ (
    .A1(_0412_),
    .A2(_0431_),
    .ZN(_0432_)
  );
  AND2_X1 _0940_ (
    .A1(_0407_),
    .A2(_0432_),
    .ZN(_0433_)
  );
  OR2_X1 _0941_ (
    .A1(_0403_),
    .A2(_0433_),
    .ZN(_0434_)
  );
  AND2_X1 _0942_ (
    .A1(_0402_),
    .A2(_0434_),
    .ZN(_0435_)
  );
  OR2_X1 _0943_ (
    .A1(_0372_),
    .A2(_0390_),
    .ZN(_0436_)
  );
  AND2_X1 _0944_ (
    .A1(_0388_),
    .A2(_0436_),
    .ZN(_0437_)
  );
  OR2_X1 _0945_ (
    .A1(_0386_),
    .A2(_0437_),
    .ZN(_0438_)
  );
  OR2_X1 _0946_ (
    .A1(_0382_),
    .A2(_0384_),
    .ZN(_0439_)
  );
  AND2_X1 _0947_ (
    .A1(_0381_),
    .A2(_0439_),
    .ZN(_0440_)
  );
  AND2_X1 _0948_ (
    .A1(_0374_),
    .A2(_0440_),
    .ZN(_0441_)
  );
  AND2_X1 _0949_ (
    .A1(_0438_),
    .A2(_0441_),
    .ZN(_0442_)
  );
  INV_X1 _0950_ (
    .A(_0442_),
    .ZN(_0443_)
  );
  AND2_X1 _0951_ (
    .A1(_0373_),
    .A2(_0389_),
    .ZN(_0444_)
  );
  AND2_X1 _0952_ (
    .A1(_0443_),
    .A2(_0444_),
    .ZN(_0445_)
  );
  OR2_X1 _0953_ (
    .A1(_0371_),
    .A2(_0379_),
    .ZN(_0446_)
  );
  OR2_X1 _0954_ (
    .A1(_0445_),
    .A2(_0446_),
    .ZN(_0447_)
  );
  AND2_X1 _0955_ (
    .A1(_0377_),
    .A2(_0447_),
    .ZN(_0448_)
  );
  OR2_X1 _0956_ (
    .A1(_0378_),
    .A2(_0448_),
    .ZN(_0449_)
  );
  OR2_X1 _0957_ (
    .A1(_0435_),
    .A2(_0449_),
    .ZN(_0450_)
  );
  AND2_X1 _0958_ (
    .A1(_0370_),
    .A2(_0450_),
    .ZN(_0451_)
  );
  OR2_X1 _0959_ (
    .A1(_0347_),
    .A2(_0359_),
    .ZN(_0452_)
  );
  OR2_X1 _0960_ (
    .A1(_0354_),
    .A2(_0452_),
    .ZN(_0453_)
  );
  OR2_X1 _0961_ (
    .A1(_0350_),
    .A2(_0351_),
    .ZN(_0454_)
  );
  AND2_X1 _0962_ (
    .A1(_0356_),
    .A2(_0454_),
    .ZN(_0455_)
  );
  AND2_X1 _0963_ (
    .A1(_0453_),
    .A2(_0455_),
    .ZN(_0456_)
  );
  INV_X1 _0964_ (
    .A(_0456_),
    .ZN(_0457_)
  );
  AND2_X1 _0965_ (
    .A1(_0358_),
    .A2(_0457_),
    .ZN(_0458_)
  );
  OR2_X1 _0966_ (
    .A1(_0337_),
    .A2(_0458_),
    .ZN(_0459_)
  );
  AND2_X1 _0967_ (
    .A1(_0336_),
    .A2(_0459_),
    .ZN(_0460_)
  );
  OR2_X1 _0968_ (
    .A1(_0344_),
    .A2(_0460_),
    .ZN(_0461_)
  );
  AND2_X1 _0969_ (
    .A1(_0333_),
    .A2(_0355_),
    .ZN(_0462_)
  );
  AND2_X1 _0970_ (
    .A1(_0461_),
    .A2(_0462_),
    .ZN(_0463_)
  );
  AND2_X1 _0971_ (
    .A1(_0304_),
    .A2(_0328_),
    .ZN(_0464_)
  );
  OR2_X1 _0972_ (
    .A1(_0323_),
    .A2(_0464_),
    .ZN(_0465_)
  );
  AND2_X1 _0973_ (
    .A1(_0321_),
    .A2(_0465_),
    .ZN(_0466_)
  );
  AND2_X1 _0974_ (
    .A1(_0316_),
    .A2(_0318_),
    .ZN(_0467_)
  );
  OR2_X1 _0975_ (
    .A1(_0299_),
    .A2(_0315_),
    .ZN(_0468_)
  );
  OR2_X1 _0976_ (
    .A1(_0467_),
    .A2(_0468_),
    .ZN(_0469_)
  );
  OR2_X1 _0977_ (
    .A1(_0466_),
    .A2(_0469_),
    .ZN(_0470_)
  );
  AND2_X1 _0978_ (
    .A1(_0312_),
    .A2(_0470_),
    .ZN(_0471_)
  );
  OR2_X1 _0979_ (
    .A1(_0302_),
    .A2(_0326_),
    .ZN(_0472_)
  );
  OR2_X1 _0980_ (
    .A1(_0471_),
    .A2(_0472_),
    .ZN(_0473_)
  );
  AND2_X1 _0981_ (
    .A1(_0309_),
    .A2(_0473_),
    .ZN(_0474_)
  );
  OR2_X1 _0982_ (
    .A1(_0297_),
    .A2(_0474_),
    .ZN(_0475_)
  );
  OR2_X1 _0983_ (
    .A1(_0463_),
    .A2(_0475_),
    .ZN(_0476_)
  );
  OR2_X1 _0984_ (
    .A1(_0451_),
    .A2(_0476_),
    .ZN(_0477_)
  );
  XOR2_X1 _0985_ (
    .A(io_bp_0_control_tmatch[0]),
    .B(_0477_),
    .Z(_0478_)
  );
  AND2_X1 _0986_ (
    .A1(io_bp_0_control_tmatch[1]),
    .A2(_0478_),
    .ZN(_0479_)
  );
  XOR2_X1 _0987_ (
    .A(io_ea[3]),
    .B(_0061_),
    .Z(_0480_)
  );
  OR2_X1 _0988_ (
    .A1(_0205_),
    .A2(_0480_),
    .ZN(_0481_)
  );
  XOR2_X1 _0989_ (
    .A(io_ea[0]),
    .B(_0058_),
    .Z(_0482_)
  );
  OR2_X1 _0990_ (
    .A1(io_bp_0_control_tmatch[0]),
    .A2(_0482_),
    .ZN(_0483_)
  );
  AND2_X1 _0991_ (
    .A1(_0000_),
    .A2(_0428_),
    .ZN(_0484_)
  );
  AND2_X1 _0992_ (
    .A1(_0411_),
    .A2(_0484_),
    .ZN(_0485_)
  );
  AND2_X1 _0993_ (
    .A1(_0483_),
    .A2(_0485_),
    .ZN(_0486_)
  );
  AND2_X1 _0994_ (
    .A1(_0404_),
    .A2(_0409_),
    .ZN(_0487_)
  );
  AND2_X1 _0995_ (
    .A1(_0407_),
    .A2(_0487_),
    .ZN(_0488_)
  );
  XOR2_X1 _0996_ (
    .A(io_ea[4]),
    .B(_0062_),
    .Z(_0489_)
  );
  AND2_X1 _0997_ (
    .A1(_0488_),
    .A2(_0489_),
    .ZN(_0490_)
  );
  AND2_X1 _0998_ (
    .A1(_0481_),
    .A2(_0490_),
    .ZN(_0491_)
  );
  AND2_X1 _0999_ (
    .A1(_0486_),
    .A2(_0491_),
    .ZN(_0492_)
  );
  XOR2_X1 _1000_ (
    .A(io_ea[1]),
    .B(_0059_),
    .Z(_0493_)
  );
  OR2_X1 _1001_ (
    .A1(_0201_),
    .A2(_0493_),
    .ZN(_0494_)
  );
  XOR2_X1 _1002_ (
    .A(io_ea[2]),
    .B(_0060_),
    .Z(_0495_)
  );
  AND2_X1 _1003_ (
    .A1(_0494_),
    .A2(_0495_),
    .ZN(_0496_)
  );
  OR2_X1 _1004_ (
    .A1(_0203_),
    .A2(_0496_),
    .ZN(_0497_)
  );
  AND2_X1 _1005_ (
    .A1(_0492_),
    .A2(_0497_),
    .ZN(_0498_)
  );
  AND2_X1 _1006_ (
    .A1(_0402_),
    .A2(_0498_),
    .ZN(_0499_)
  );
  AND2_X1 _1007_ (
    .A1(_0370_),
    .A2(_0499_),
    .ZN(_0500_)
  );
  OR2_X1 _1008_ (
    .A1(_0479_),
    .A2(_0500_),
    .ZN(_0501_)
  );
  AND2_X1 _1009_ (
    .A1(_0001_),
    .A2(io_bp_0_control_r),
    .ZN(_0502_)
  );
  AND2_X1 _1010_ (
    .A1(_0501_),
    .A2(_0502_),
    .ZN(_0503_)
  );
  AND2_X1 _1011_ (
    .A1(_0057_),
    .A2(_0503_),
    .ZN(io_xcpt_ld)
  );
  AND2_X1 _1012_ (
    .A1(_0001_),
    .A2(io_bp_0_control_w),
    .ZN(_0504_)
  );
  AND2_X1 _1013_ (
    .A1(_0501_),
    .A2(_0504_),
    .ZN(_0505_)
  );
  AND2_X1 _1014_ (
    .A1(_0057_),
    .A2(_0505_),
    .ZN(io_xcpt_st)
  );
  AND2_X1 _1015_ (
    .A1(io_bp_0_control_action),
    .A2(_0296_),
    .ZN(io_debug_if)
  );
  AND2_X1 _1016_ (
    .A1(io_bp_0_control_action),
    .A2(_0503_),
    .ZN(io_debug_ld)
  );
  AND2_X1 _1017_ (
    .A1(io_bp_0_control_action),
    .A2(_0505_),
    .ZN(io_debug_st)
  );
  assign { _GEN_11[31:4], _GEN_11[0] } = { 28'h0000000, io_bp_0_control_tmatch[0] };
  assign _r_T_10 = _GEN_11[2];
  assign _r_T_12 = _GEN_11[3];
  assign _r_T_13 = { _GEN_11[3:1], io_bp_0_control_tmatch[0] };
  assign _r_T_8 = _GEN_11[1];
endmodule
module CSRFile(clock, reset, io_ungated_clock, io_interrupts_debug, io_interrupts_mtip, io_interrupts_msip, io_interrupts_meip, io_hartid, io_rw_addr, io_rw_cmd, io_rw_rdata, io_rw_wdata, io_decode_0_inst, io_decode_0_fp_illegal, io_decode_0_fp_csr, io_decode_0_rocc_illegal, io_decode_0_read_illegal, io_decode_0_write_illegal, io_decode_0_write_flush, io_decode_0_system_illegal, io_csr_stall
, io_eret, io_singleStep, io_status_debug, io_status_cease, io_status_wfi, io_status_isa, io_status_dprv, io_status_dv, io_status_prv, io_status_v, io_status_sd, io_status_zero2, io_status_mpv, io_status_gva, io_status_mbe, io_status_sbe, io_status_sxl, io_status_uxl, io_status_sd_rv32, io_status_zero1, io_status_tsr
, io_status_tw, io_status_tvm, io_status_mxr, io_status_sum, io_status_mprv, io_status_xs, io_status_fs, io_status_mpp, io_status_vs, io_status_spp, io_status_mpie, io_status_ube, io_status_spie, io_status_upie, io_status_mie, io_status_hie, io_status_sie, io_status_uie, io_evec, io_exception, io_retire
, io_cause, io_pc, io_tval, io_gva, io_time, io_interrupt, io_interrupt_cause, io_bp_0_control_action, io_bp_0_control_tmatch, io_bp_0_control_x, io_bp_0_control_w, io_bp_0_control_r, io_bp_0_address, io_pmp_0_cfg_l, io_pmp_0_cfg_a, io_pmp_0_cfg_x, io_pmp_0_cfg_w, io_pmp_0_cfg_r, io_pmp_0_addr, io_pmp_0_mask, io_pmp_1_cfg_l
, io_pmp_1_cfg_a, io_pmp_1_cfg_x, io_pmp_1_cfg_w, io_pmp_1_cfg_r, io_pmp_1_addr, io_pmp_1_mask, io_pmp_2_cfg_l, io_pmp_2_cfg_a, io_pmp_2_cfg_x, io_pmp_2_cfg_w, io_pmp_2_cfg_r, io_pmp_2_addr, io_pmp_2_mask, io_pmp_3_cfg_l, io_pmp_3_cfg_a, io_pmp_3_cfg_x, io_pmp_3_cfg_w, io_pmp_3_cfg_r, io_pmp_3_addr, io_pmp_3_mask, io_pmp_4_cfg_l
, io_pmp_4_cfg_a, io_pmp_4_cfg_x, io_pmp_4_cfg_w, io_pmp_4_cfg_r, io_pmp_4_addr, io_pmp_4_mask, io_pmp_5_cfg_l, io_pmp_5_cfg_a, io_pmp_5_cfg_x, io_pmp_5_cfg_w, io_pmp_5_cfg_r, io_pmp_5_addr, io_pmp_5_mask, io_pmp_6_cfg_l, io_pmp_6_cfg_a, io_pmp_6_cfg_x, io_pmp_6_cfg_w, io_pmp_6_cfg_r, io_pmp_6_addr, io_pmp_6_mask, io_pmp_7_cfg_l
, io_pmp_7_cfg_a, io_pmp_7_cfg_x, io_pmp_7_cfg_w, io_pmp_7_cfg_r, io_pmp_7_addr, io_pmp_7_mask, io_inhibit_cycle, io_inst_0, io_trace_0_valid, io_trace_0_iaddr, io_trace_0_insn, io_trace_0_exception, io_customCSRs_0_value);
  wire [31:0] _0000_;
  wire [31:0] _0001_;
  wire [31:0] _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire _1340_;
  wire _1341_;
  wire _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  wire _1351_;
  wire _1352_;
  wire _1353_;
  wire _1354_;
  wire _1355_;
  wire _1356_;
  wire _1357_;
  wire _1358_;
  wire _1359_;
  wire _1360_;
  wire _1361_;
  wire _1362_;
  wire _1363_;
  wire _1364_;
  wire _1365_;
  wire _1366_;
  wire _1367_;
  wire _1368_;
  wire _1369_;
  wire _1370_;
  wire _1371_;
  wire _1372_;
  wire _1373_;
  wire _1374_;
  wire _1375_;
  wire _1376_;
  wire _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire _1382_;
  wire _1383_;
  wire _1384_;
  wire _1385_;
  wire _1386_;
  wire _1387_;
  wire _1388_;
  wire _1389_;
  wire _1390_;
  wire _1391_;
  wire _1392_;
  wire _1393_;
  wire _1394_;
  wire _1395_;
  wire _1396_;
  wire _1397_;
  wire _1398_;
  wire _1399_;
  wire _1400_;
  wire _1401_;
  wire _1402_;
  wire _1403_;
  wire _1404_;
  wire _1405_;
  wire _1406_;
  wire _1407_;
  wire _1408_;
  wire _1409_;
  wire _1410_;
  wire _1411_;
  wire _1412_;
  wire _1413_;
  wire _1414_;
  wire _1415_;
  wire _1416_;
  wire _1417_;
  wire _1418_;
  wire _1419_;
  wire _1420_;
  wire _1421_;
  wire _1422_;
  wire _1423_;
  wire _1424_;
  wire _1425_;
  wire _1426_;
  wire _1427_;
  wire _1428_;
  wire _1429_;
  wire _1430_;
  wire _1431_;
  wire _1432_;
  wire _1433_;
  wire _1434_;
  wire _1435_;
  wire _1436_;
  wire _1437_;
  wire _1438_;
  wire _1439_;
  wire _1440_;
  wire _1441_;
  wire _1442_;
  wire _1443_;
  wire _1444_;
  wire _1445_;
  wire _1446_;
  wire _1447_;
  wire _1448_;
  wire _1449_;
  wire _1450_;
  wire _1451_;
  wire _1452_;
  wire _1453_;
  wire _1454_;
  wire _1455_;
  wire _1456_;
  wire _1457_;
  wire _1458_;
  wire _1459_;
  wire _1460_;
  wire _1461_;
  wire _1462_;
  wire _1463_;
  wire _1464_;
  wire _1465_;
  wire _1466_;
  wire _1467_;
  wire _1468_;
  wire _1469_;
  wire _1470_;
  wire _1471_;
  wire _1472_;
  wire _1473_;
  wire _1474_;
  wire _1475_;
  wire _1476_;
  wire _1477_;
  wire _1478_;
  wire _1479_;
  wire _1480_;
  wire _1481_;
  wire _1482_;
  wire _1483_;
  wire _1484_;
  wire _1485_;
  wire _1486_;
  wire _1487_;
  wire _1488_;
  wire _1489_;
  wire _1490_;
  wire _1491_;
  wire _1492_;
  wire _1493_;
  wire _1494_;
  wire _1495_;
  wire _1496_;
  wire _1497_;
  wire _1498_;
  wire _1499_;
  wire _1500_;
  wire _1501_;
  wire _1502_;
  wire _1503_;
  wire _1504_;
  wire _1505_;
  wire _1506_;
  wire _1507_;
  wire _1508_;
  wire _1509_;
  wire _1510_;
  wire _1511_;
  wire _1512_;
  wire _1513_;
  wire _1514_;
  wire _1515_;
  wire _1516_;
  wire _1517_;
  wire _1518_;
  wire _1519_;
  wire _1520_;
  wire _1521_;
  wire _1522_;
  wire _1523_;
  wire _1524_;
  wire _1525_;
  wire _1526_;
  wire _1527_;
  wire _1528_;
  wire _1529_;
  wire _1530_;
  wire _1531_;
  wire _1532_;
  wire _1533_;
  wire _1534_;
  wire _1535_;
  wire _1536_;
  wire _1537_;
  wire _1538_;
  wire _1539_;
  wire _1540_;
  wire _1541_;
  wire _1542_;
  wire _1543_;
  wire _1544_;
  wire _1545_;
  wire _1546_;
  wire _1547_;
  wire _1548_;
  wire _1549_;
  wire _1550_;
  wire _1551_;
  wire _1552_;
  wire _1553_;
  wire _1554_;
  wire _1555_;
  wire _1556_;
  wire _1557_;
  wire _1558_;
  wire _1559_;
  wire _1560_;
  wire _1561_;
  wire _1562_;
  wire _1563_;
  wire _1564_;
  wire _1565_;
  wire _1566_;
  wire _1567_;
  wire _1568_;
  wire _1569_;
  wire _1570_;
  wire _1571_;
  wire _1572_;
  wire _1573_;
  wire _1574_;
  wire _1575_;
  wire _1576_;
  wire _1577_;
  wire _1578_;
  wire _1579_;
  wire _1580_;
  wire _1581_;
  wire _1582_;
  wire _1583_;
  wire _1584_;
  wire _1585_;
  wire _1586_;
  wire _1587_;
  wire _1588_;
  wire _1589_;
  wire _1590_;
  wire _1591_;
  wire _1592_;
  wire _1593_;
  wire _1594_;
  wire _1595_;
  wire _1596_;
  wire _1597_;
  wire _1598_;
  wire _1599_;
  wire _1600_;
  wire _1601_;
  wire _1602_;
  wire _1603_;
  wire _1604_;
  wire _1605_;
  wire _1606_;
  wire _1607_;
  wire _1608_;
  wire _1609_;
  wire _1610_;
  wire _1611_;
  wire _1612_;
  wire _1613_;
  wire _1614_;
  wire _1615_;
  wire _1616_;
  wire _1617_;
  wire _1618_;
  wire _1619_;
  wire _1620_;
  wire _1621_;
  wire _1622_;
  wire _1623_;
  wire _1624_;
  wire _1625_;
  wire _1626_;
  wire _1627_;
  wire _1628_;
  wire _1629_;
  wire _1630_;
  wire _1631_;
  wire _1632_;
  wire _1633_;
  wire _1634_;
  wire _1635_;
  wire _1636_;
  wire _1637_;
  wire _1638_;
  wire _1639_;
  wire _1640_;
  wire _1641_;
  wire _1642_;
  wire _1643_;
  wire _1644_;
  wire _1645_;
  wire _1646_;
  wire _1647_;
  wire _1648_;
  wire _1649_;
  wire _1650_;
  wire _1651_;
  wire _1652_;
  wire _1653_;
  wire _1654_;
  wire _1655_;
  wire _1656_;
  wire _1657_;
  wire _1658_;
  wire _1659_;
  wire _1660_;
  wire _1661_;
  wire _1662_;
  wire _1663_;
  wire _1664_;
  wire _1665_;
  wire _1666_;
  wire _1667_;
  wire _1668_;
  wire _1669_;
  wire _1670_;
  wire _1671_;
  wire _1672_;
  wire _1673_;
  wire _1674_;
  wire _1675_;
  wire _1676_;
  wire _1677_;
  wire _1678_;
  wire _1679_;
  wire _1680_;
  wire _1681_;
  wire _1682_;
  wire _1683_;
  wire _1684_;
  wire _1685_;
  wire _1686_;
  wire _1687_;
  wire _1688_;
  wire _1689_;
  wire _1690_;
  wire _1691_;
  wire _1692_;
  wire _1693_;
  wire _1694_;
  wire _1695_;
  wire _1696_;
  wire _1697_;
  wire _1698_;
  wire _1699_;
  wire _1700_;
  wire _1701_;
  wire _1702_;
  wire _1703_;
  wire _1704_;
  wire _1705_;
  wire _1706_;
  wire _1707_;
  wire _1708_;
  wire _1709_;
  wire _1710_;
  wire _1711_;
  wire _1712_;
  wire _1713_;
  wire _1714_;
  wire _1715_;
  wire _1716_;
  wire _1717_;
  wire _1718_;
  wire _1719_;
  wire _1720_;
  wire _1721_;
  wire _1722_;
  wire _1723_;
  wire _1724_;
  wire _1725_;
  wire _1726_;
  wire _1727_;
  wire _1728_;
  wire _1729_;
  wire _1730_;
  wire _1731_;
  wire _1732_;
  wire _1733_;
  wire _1734_;
  wire _1735_;
  wire _1736_;
  wire _1737_;
  wire _1738_;
  wire _1739_;
  wire _1740_;
  wire _1741_;
  wire _1742_;
  wire _1743_;
  wire _1744_;
  wire _1745_;
  wire _1746_;
  wire _1747_;
  wire _1748_;
  wire _1749_;
  wire _1750_;
  wire _1751_;
  wire _1752_;
  wire _1753_;
  wire _1754_;
  wire _1755_;
  wire _1756_;
  wire _1757_;
  wire _1758_;
  wire _1759_;
  wire _1760_;
  wire _1761_;
  wire _1762_;
  wire _1763_;
  wire _1764_;
  wire _1765_;
  wire _1766_;
  wire _1767_;
  wire _1768_;
  wire _1769_;
  wire _1770_;
  wire _1771_;
  wire _1772_;
  wire _1773_;
  wire _1774_;
  wire _1775_;
  wire _1776_;
  wire _1777_;
  wire _1778_;
  wire _1779_;
  wire _1780_;
  wire _1781_;
  wire _1782_;
  wire _1783_;
  wire _1784_;
  wire _1785_;
  wire _1786_;
  wire _1787_;
  wire _1788_;
  wire _1789_;
  wire _1790_;
  wire _1791_;
  wire _1792_;
  wire _1793_;
  wire _1794_;
  wire _1795_;
  wire _1796_;
  wire _1797_;
  wire _1798_;
  wire _1799_;
  wire _1800_;
  wire _1801_;
  wire _1802_;
  wire _1803_;
  wire _1804_;
  wire _1805_;
  wire _1806_;
  wire _1807_;
  wire _1808_;
  wire _1809_;
  wire _1810_;
  wire _1811_;
  wire _1812_;
  wire _1813_;
  wire _1814_;
  wire _1815_;
  wire _1816_;
  wire _1817_;
  wire _1818_;
  wire _1819_;
  wire _1820_;
  wire _1821_;
  wire _1822_;
  wire _1823_;
  wire _1824_;
  wire _1825_;
  wire _1826_;
  wire _1827_;
  wire _1828_;
  wire _1829_;
  wire _1830_;
  wire _1831_;
  wire _1832_;
  wire _1833_;
  wire _1834_;
  wire _1835_;
  wire _1836_;
  wire _1837_;
  wire _1838_;
  wire _1839_;
  wire _1840_;
  wire _1841_;
  wire _1842_;
  wire _1843_;
  wire _1844_;
  wire _1845_;
  wire _1846_;
  wire _1847_;
  wire _1848_;
  wire _1849_;
  wire _1850_;
  wire _1851_;
  wire _1852_;
  wire _1853_;
  wire _1854_;
  wire _1855_;
  wire _1856_;
  wire _1857_;
  wire _1858_;
  wire _1859_;
  wire _1860_;
  wire _1861_;
  wire _1862_;
  wire _1863_;
  wire _1864_;
  wire _1865_;
  wire _1866_;
  wire _1867_;
  wire _1868_;
  wire _1869_;
  wire _1870_;
  wire _1871_;
  wire _1872_;
  wire _1873_;
  wire _1874_;
  wire _1875_;
  wire _1876_;
  wire _1877_;
  wire _1878_;
  wire _1879_;
  wire _1880_;
  wire _1881_;
  wire _1882_;
  wire _1883_;
  wire _1884_;
  wire _1885_;
  wire _1886_;
  wire _1887_;
  wire _1888_;
  wire _1889_;
  wire _1890_;
  wire _1891_;
  wire _1892_;
  wire _1893_;
  wire _1894_;
  wire _1895_;
  wire _1896_;
  wire _1897_;
  wire _1898_;
  wire _1899_;
  wire _1900_;
  wire _1901_;
  wire _1902_;
  wire _1903_;
  wire _1904_;
  wire _1905_;
  wire _1906_;
  wire _1907_;
  wire _1908_;
  wire _1909_;
  wire _1910_;
  wire _1911_;
  wire _1912_;
  wire _1913_;
  wire _1914_;
  wire _1915_;
  wire _1916_;
  wire _1917_;
  wire _1918_;
  wire _1919_;
  wire _1920_;
  wire _1921_;
  wire _1922_;
  wire _1923_;
  wire _1924_;
  wire _1925_;
  wire _1926_;
  wire _1927_;
  wire _1928_;
  wire _1929_;
  wire _1930_;
  wire _1931_;
  wire _1932_;
  wire _1933_;
  wire _1934_;
  wire _1935_;
  wire _1936_;
  wire _1937_;
  wire _1938_;
  wire _1939_;
  wire _1940_;
  wire _1941_;
  wire _1942_;
  wire _1943_;
  wire _1944_;
  wire _1945_;
  wire _1946_;
  wire _1947_;
  wire _1948_;
  wire _1949_;
  wire _1950_;
  wire _1951_;
  wire _1952_;
  wire _1953_;
  wire _1954_;
  wire _1955_;
  wire _1956_;
  wire _1957_;
  wire _1958_;
  wire _1959_;
  wire _1960_;
  wire _1961_;
  wire _1962_;
  wire _1963_;
  wire _1964_;
  wire _1965_;
  wire _1966_;
  wire _1967_;
  wire _1968_;
  wire _1969_;
  wire _1970_;
  wire _1971_;
  wire _1972_;
  wire _1973_;
  wire _1974_;
  wire _1975_;
  wire _1976_;
  wire _1977_;
  wire _1978_;
  wire _1979_;
  wire _1980_;
  wire _1981_;
  wire _1982_;
  wire _1983_;
  wire _1984_;
  wire _1985_;
  wire _1986_;
  wire _1987_;
  wire _1988_;
  wire _1989_;
  wire _1990_;
  wire _1991_;
  wire _1992_;
  wire _1993_;
  wire _1994_;
  wire _1995_;
  wire _1996_;
  wire _1997_;
  wire _1998_;
  wire _1999_;
  wire _2000_;
  wire _2001_;
  wire _2002_;
  wire _2003_;
  wire _2004_;
  wire _2005_;
  wire _2006_;
  wire _2007_;
  wire _2008_;
  wire _2009_;
  wire _2010_;
  wire _2011_;
  wire _2012_;
  wire _2013_;
  wire _2014_;
  wire _2015_;
  wire _2016_;
  wire _2017_;
  wire _2018_;
  wire _2019_;
  wire _2020_;
  wire _2021_;
  wire _2022_;
  wire _2023_;
  wire _2024_;
  wire _2025_;
  wire _2026_;
  wire _2027_;
  wire _2028_;
  wire _2029_;
  wire _2030_;
  wire _2031_;
  wire _2032_;
  wire _2033_;
  wire _2034_;
  wire _2035_;
  wire _2036_;
  wire _2037_;
  wire _2038_;
  wire _2039_;
  wire _2040_;
  wire _2041_;
  wire _2042_;
  wire _2043_;
  wire _2044_;
  wire _2045_;
  wire _2046_;
  wire _2047_;
  wire _2048_;
  wire _2049_;
  wire _2050_;
  wire _2051_;
  wire _2052_;
  wire _2053_;
  wire _2054_;
  wire _2055_;
  wire _2056_;
  wire _2057_;
  wire _2058_;
  wire _2059_;
  wire _2060_;
  wire _2061_;
  wire _2062_;
  wire _2063_;
  wire _2064_;
  wire _2065_;
  wire _2066_;
  wire _2067_;
  wire _2068_;
  wire _2069_;
  wire _2070_;
  wire _2071_;
  wire _2072_;
  wire _2073_;
  wire _2074_;
  wire _2075_;
  wire _2076_;
  wire _2077_;
  wire _2078_;
  wire _2079_;
  wire _2080_;
  wire _2081_;
  wire _2082_;
  wire _2083_;
  wire _2084_;
  wire _2085_;
  wire _2086_;
  wire _2087_;
  wire _2088_;
  wire _2089_;
  wire _2090_;
  wire _2091_;
  wire _2092_;
  wire _2093_;
  wire _2094_;
  wire _2095_;
  wire _2096_;
  wire _2097_;
  wire _2098_;
  wire _2099_;
  wire _2100_;
  wire _2101_;
  wire _2102_;
  wire _2103_;
  wire _2104_;
  wire _2105_;
  wire _2106_;
  wire _2107_;
  wire _2108_;
  wire _2109_;
  wire _2110_;
  wire _2111_;
  wire _2112_;
  wire _2113_;
  wire _2114_;
  wire _2115_;
  wire _2116_;
  wire _2117_;
  wire _2118_;
  wire _2119_;
  wire _2120_;
  wire _2121_;
  wire _2122_;
  wire _2123_;
  wire _2124_;
  wire _2125_;
  wire _2126_;
  wire _2127_;
  wire _2128_;
  wire _2129_;
  wire _2130_;
  wire _2131_;
  wire _2132_;
  wire _2133_;
  wire _2134_;
  wire _2135_;
  wire _2136_;
  wire _2137_;
  wire _2138_;
  wire _2139_;
  wire _2140_;
  wire _2141_;
  wire _2142_;
  wire _2143_;
  wire _2144_;
  wire _2145_;
  wire _2146_;
  wire _2147_;
  wire _2148_;
  wire _2149_;
  wire _2150_;
  wire _2151_;
  wire _2152_;
  wire _2153_;
  wire _2154_;
  wire _2155_;
  wire _2156_;
  wire _2157_;
  wire _2158_;
  wire _2159_;
  wire _2160_;
  wire _2161_;
  wire _2162_;
  wire _2163_;
  wire _2164_;
  wire _2165_;
  wire _2166_;
  wire _2167_;
  wire _2168_;
  wire _2169_;
  wire _2170_;
  wire _2171_;
  wire _2172_;
  wire _2173_;
  wire _2174_;
  wire _2175_;
  wire _2176_;
  wire _2177_;
  wire _2178_;
  wire _2179_;
  wire _2180_;
  wire _2181_;
  wire _2182_;
  wire _2183_;
  wire _2184_;
  wire _2185_;
  wire _2186_;
  wire _2187_;
  wire _2188_;
  wire _2189_;
  wire _2190_;
  wire _2191_;
  wire _2192_;
  wire _2193_;
  wire _2194_;
  wire _2195_;
  wire _2196_;
  wire _2197_;
  wire _2198_;
  wire _2199_;
  wire _2200_;
  wire _2201_;
  wire _2202_;
  wire _2203_;
  wire _2204_;
  wire _2205_;
  wire _2206_;
  wire _2207_;
  wire _2208_;
  wire _2209_;
  wire _2210_;
  wire _2211_;
  wire _2212_;
  wire _2213_;
  wire _2214_;
  wire _2215_;
  wire _2216_;
  wire _2217_;
  wire _2218_;
  wire _2219_;
  wire _2220_;
  wire _2221_;
  wire _2222_;
  wire _2223_;
  wire _2224_;
  wire _2225_;
  wire _2226_;
  wire _2227_;
  wire _2228_;
  wire _2229_;
  wire _2230_;
  wire _2231_;
  wire _2232_;
  wire _2233_;
  wire _2234_;
  wire _2235_;
  wire _2236_;
  wire _2237_;
  wire _2238_;
  wire _2239_;
  wire _2240_;
  wire _2241_;
  wire _2242_;
  wire _2243_;
  wire _2244_;
  wire _2245_;
  wire _2246_;
  wire _2247_;
  wire _2248_;
  wire _2249_;
  wire _2250_;
  wire _2251_;
  wire _2252_;
  wire _2253_;
  wire _2254_;
  wire _2255_;
  wire _2256_;
  wire _2257_;
  wire _2258_;
  wire _2259_;
  wire _2260_;
  wire _2261_;
  wire _2262_;
  wire _2263_;
  wire _2264_;
  wire _2265_;
  wire _2266_;
  wire _2267_;
  wire _2268_;
  wire _2269_;
  wire _2270_;
  wire _2271_;
  wire _2272_;
  wire _2273_;
  wire _2274_;
  wire _2275_;
  wire _2276_;
  wire _2277_;
  wire _2278_;
  wire _2279_;
  wire _2280_;
  wire _2281_;
  wire _2282_;
  wire _2283_;
  wire _2284_;
  wire _2285_;
  wire _2286_;
  wire _2287_;
  wire _2288_;
  wire _2289_;
  wire _2290_;
  wire _2291_;
  wire _2292_;
  wire _2293_;
  wire _2294_;
  wire _2295_;
  wire _2296_;
  wire _2297_;
  wire _2298_;
  wire _2299_;
  wire _2300_;
  wire _2301_;
  wire _2302_;
  wire _2303_;
  wire _2304_;
  wire _2305_;
  wire _2306_;
  wire _2307_;
  wire _2308_;
  wire _2309_;
  wire _2310_;
  wire _2311_;
  wire _2312_;
  wire _2313_;
  wire _2314_;
  wire _2315_;
  wire _2316_;
  wire _2317_;
  wire _2318_;
  wire _2319_;
  wire _2320_;
  wire _2321_;
  wire _2322_;
  wire _2323_;
  wire _2324_;
  wire _2325_;
  wire _2326_;
  wire _2327_;
  wire _2328_;
  wire _2329_;
  wire _2330_;
  wire _2331_;
  wire _2332_;
  wire _2333_;
  wire _2334_;
  wire _2335_;
  wire _2336_;
  wire _2337_;
  wire _2338_;
  wire _2339_;
  wire _2340_;
  wire _2341_;
  wire _2342_;
  wire _2343_;
  wire _2344_;
  wire _2345_;
  wire _2346_;
  wire _2347_;
  wire _2348_;
  wire _2349_;
  wire _2350_;
  wire _2351_;
  wire _2352_;
  wire _2353_;
  wire _2354_;
  wire _2355_;
  wire _2356_;
  wire _2357_;
  wire _2358_;
  wire _2359_;
  wire _2360_;
  wire _2361_;
  wire _2362_;
  wire _2363_;
  wire _2364_;
  wire _2365_;
  wire _2366_;
  wire _2367_;
  wire _2368_;
  wire _2369_;
  wire _2370_;
  wire _2371_;
  wire _2372_;
  wire _2373_;
  wire _2374_;
  wire _2375_;
  wire _2376_;
  wire _2377_;
  wire _2378_;
  wire _2379_;
  wire _2380_;
  wire _2381_;
  wire _2382_;
  wire _2383_;
  wire _2384_;
  wire _2385_;
  wire _2386_;
  wire _2387_;
  wire _2388_;
  wire _2389_;
  wire _2390_;
  wire _2391_;
  wire _2392_;
  wire _2393_;
  wire _2394_;
  wire _2395_;
  wire _2396_;
  wire _2397_;
  wire _2398_;
  wire _2399_;
  wire _2400_;
  wire _2401_;
  wire _2402_;
  wire _2403_;
  wire _2404_;
  wire _2405_;
  wire _2406_;
  wire _2407_;
  wire _2408_;
  wire _2409_;
  wire _2410_;
  wire _2411_;
  wire _2412_;
  wire _2413_;
  wire _2414_;
  wire _2415_;
  wire _2416_;
  wire _2417_;
  wire _2418_;
  wire _2419_;
  wire _2420_;
  wire _2421_;
  wire _2422_;
  wire _2423_;
  wire _2424_;
  wire _2425_;
  wire _2426_;
  wire _2427_;
  wire _2428_;
  wire _2429_;
  wire _2430_;
  wire _2431_;
  wire _2432_;
  wire _2433_;
  wire _2434_;
  wire _2435_;
  wire _2436_;
  wire _2437_;
  wire _2438_;
  wire _2439_;
  wire _2440_;
  wire _2441_;
  wire _2442_;
  wire _2443_;
  wire _2444_;
  wire _2445_;
  wire _2446_;
  wire _2447_;
  wire _2448_;
  wire _2449_;
  wire _2450_;
  wire _2451_;
  wire _2452_;
  wire _2453_;
  wire _2454_;
  wire _2455_;
  wire _2456_;
  wire _2457_;
  wire _2458_;
  wire _2459_;
  wire _2460_;
  wire _2461_;
  wire _2462_;
  wire _2463_;
  wire _2464_;
  wire _2465_;
  wire _2466_;
  wire _2467_;
  wire _2468_;
  wire _2469_;
  wire _2470_;
  wire _2471_;
  wire _2472_;
  wire _2473_;
  wire _2474_;
  wire _2475_;
  wire _2476_;
  wire _2477_;
  wire _2478_;
  wire _2479_;
  wire _2480_;
  wire _2481_;
  wire _2482_;
  wire _2483_;
  wire _2484_;
  wire _2485_;
  wire _2486_;
  wire _2487_;
  wire _2488_;
  wire _2489_;
  wire _2490_;
  wire _2491_;
  wire _2492_;
  wire _2493_;
  wire _2494_;
  wire _2495_;
  wire _2496_;
  wire _2497_;
  wire _2498_;
  wire _2499_;
  wire _2500_;
  wire _2501_;
  wire _2502_;
  wire _2503_;
  wire _2504_;
  wire _2505_;
  wire _2506_;
  wire _2507_;
  wire _2508_;
  wire _2509_;
  wire _2510_;
  wire _2511_;
  wire _2512_;
  wire _2513_;
  wire _2514_;
  wire _2515_;
  wire _2516_;
  wire _2517_;
  wire _2518_;
  wire _2519_;
  wire _2520_;
  wire _2521_;
  wire _2522_;
  wire _2523_;
  wire _2524_;
  wire _2525_;
  wire _2526_;
  wire _2527_;
  wire _2528_;
  wire _2529_;
  wire _2530_;
  wire _2531_;
  wire _2532_;
  wire _2533_;
  wire _2534_;
  wire _2535_;
  wire _2536_;
  wire _2537_;
  wire _2538_;
  wire _2539_;
  wire _2540_;
  wire _2541_;
  wire _2542_;
  wire _2543_;
  wire _2544_;
  wire _2545_;
  wire _2546_;
  wire _2547_;
  wire _2548_;
  wire _2549_;
  wire _2550_;
  wire _2551_;
  wire _2552_;
  wire _2553_;
  wire _2554_;
  wire _2555_;
  wire _2556_;
  wire _2557_;
  wire _2558_;
  wire _2559_;
  wire _2560_;
  wire _2561_;
  wire _2562_;
  wire _2563_;
  wire _2564_;
  wire _2565_;
  wire _2566_;
  wire _2567_;
  wire _2568_;
  wire _2569_;
  wire _2570_;
  wire _2571_;
  wire _2572_;
  wire _2573_;
  wire _2574_;
  wire _2575_;
  wire _2576_;
  wire _2577_;
  wire _2578_;
  wire _2579_;
  wire _2580_;
  wire _2581_;
  wire _2582_;
  wire _2583_;
  wire _2584_;
  wire _2585_;
  wire _2586_;
  wire _2587_;
  wire _2588_;
  wire _2589_;
  wire _2590_;
  wire _2591_;
  wire _2592_;
  wire _2593_;
  wire _2594_;
  wire _2595_;
  wire _2596_;
  wire _2597_;
  wire _2598_;
  wire _2599_;
  wire _2600_;
  wire _2601_;
  wire _2602_;
  wire _2603_;
  wire _2604_;
  wire _2605_;
  wire _2606_;
  wire _2607_;
  wire _2608_;
  wire _2609_;
  wire _2610_;
  wire _2611_;
  wire _2612_;
  wire _2613_;
  wire _2614_;
  wire _2615_;
  wire _2616_;
  wire _2617_;
  wire _2618_;
  wire _2619_;
  wire _2620_;
  wire _2621_;
  wire _2622_;
  wire _2623_;
  wire _2624_;
  wire _2625_;
  wire _2626_;
  wire _2627_;
  wire _2628_;
  wire _2629_;
  wire _2630_;
  wire _2631_;
  wire _2632_;
  wire _2633_;
  wire _2634_;
  wire _2635_;
  wire _2636_;
  wire _2637_;
  wire _2638_;
  wire _2639_;
  wire _2640_;
  wire _2641_;
  wire _2642_;
  wire _2643_;
  wire _2644_;
  wire _2645_;
  wire _2646_;
  wire _2647_;
  wire _2648_;
  wire _2649_;
  wire _2650_;
  wire _2651_;
  wire _2652_;
  wire _2653_;
  wire _2654_;
  wire _2655_;
  wire _2656_;
  wire _2657_;
  wire _2658_;
  wire _2659_;
  wire _2660_;
  wire _2661_;
  wire _2662_;
  wire _2663_;
  wire _2664_;
  wire _2665_;
  wire _2666_;
  wire _2667_;
  wire _2668_;
  wire _2669_;
  wire _2670_;
  wire _2671_;
  wire _2672_;
  wire _2673_;
  wire _2674_;
  wire _2675_;
  wire _2676_;
  wire _2677_;
  wire _2678_;
  wire _2679_;
  wire _2680_;
  wire _2681_;
  wire _2682_;
  wire _2683_;
  wire _2684_;
  wire _2685_;
  wire _2686_;
  wire _2687_;
  wire _2688_;
  wire _2689_;
  wire _2690_;
  wire _2691_;
  wire _2692_;
  wire _2693_;
  wire _2694_;
  wire _2695_;
  wire _2696_;
  wire _2697_;
  wire _2698_;
  wire _2699_;
  wire _2700_;
  wire _2701_;
  wire _2702_;
  wire _2703_;
  wire _2704_;
  wire _2705_;
  wire _2706_;
  wire _2707_;
  wire _2708_;
  wire _2709_;
  wire _2710_;
  wire _2711_;
  wire _2712_;
  wire _2713_;
  wire _2714_;
  wire _2715_;
  wire _2716_;
  wire _2717_;
  wire _2718_;
  wire _2719_;
  wire _2720_;
  wire _2721_;
  wire _2722_;
  wire _2723_;
  wire _2724_;
  wire _2725_;
  wire _2726_;
  wire _2727_;
  wire _2728_;
  wire _2729_;
  wire _2730_;
  wire _2731_;
  wire _2732_;
  wire _2733_;
  wire _2734_;
  wire _2735_;
  wire _2736_;
  wire _2737_;
  wire _2738_;
  wire _2739_;
  wire _2740_;
  wire _2741_;
  wire _2742_;
  wire _2743_;
  wire _2744_;
  wire _2745_;
  wire _2746_;
  wire _2747_;
  wire _2748_;
  wire _2749_;
  wire _2750_;
  wire _2751_;
  wire _2752_;
  wire _2753_;
  wire _2754_;
  wire _2755_;
  wire _2756_;
  wire _2757_;
  wire _2758_;
  wire _2759_;
  wire _2760_;
  wire _2761_;
  wire _2762_;
  wire _2763_;
  wire _2764_;
  wire _2765_;
  wire _2766_;
  wire _2767_;
  wire _2768_;
  wire _2769_;
  wire _2770_;
  wire _2771_;
  wire _2772_;
  wire _2773_;
  wire _2774_;
  wire _2775_;
  wire _2776_;
  wire _2777_;
  wire _2778_;
  wire _2779_;
  wire _2780_;
  wire _2781_;
  wire _2782_;
  wire _2783_;
  wire _2784_;
  wire _2785_;
  wire _2786_;
  wire _2787_;
  wire _2788_;
  wire _2789_;
  wire _2790_;
  wire _2791_;
  wire _2792_;
  wire _2793_;
  wire _2794_;
  wire _2795_;
  wire _2796_;
  wire _2797_;
  wire _2798_;
  wire _2799_;
  wire _2800_;
  wire _2801_;
  wire _2802_;
  wire _2803_;
  wire _2804_;
  wire _2805_;
  wire _2806_;
  wire _2807_;
  wire _2808_;
  wire _2809_;
  wire _2810_;
  wire _2811_;
  wire _2812_;
  wire _2813_;
  wire _2814_;
  wire _2815_;
  wire _2816_;
  wire _2817_;
  wire _2818_;
  wire _2819_;
  wire _2820_;
  wire _2821_;
  wire _2822_;
  wire _2823_;
  wire _2824_;
  wire _2825_;
  wire _2826_;
  wire _2827_;
  wire _2828_;
  wire _2829_;
  wire _2830_;
  wire _2831_;
  wire _2832_;
  wire _2833_;
  wire _2834_;
  wire _2835_;
  wire _2836_;
  wire _2837_;
  wire _2838_;
  wire _2839_;
  wire _2840_;
  wire _2841_;
  wire _2842_;
  wire _2843_;
  wire _2844_;
  wire _2845_;
  wire _2846_;
  wire _2847_;
  wire _2848_;
  wire _2849_;
  wire _2850_;
  wire _2851_;
  wire _2852_;
  wire _2853_;
  wire _2854_;
  wire _2855_;
  wire _2856_;
  wire _2857_;
  wire _2858_;
  wire _2859_;
  wire _2860_;
  wire _2861_;
  wire _2862_;
  wire _2863_;
  wire _2864_;
  wire _2865_;
  wire _2866_;
  wire _2867_;
  wire _2868_;
  wire _2869_;
  wire _2870_;
  wire _2871_;
  wire _2872_;
  wire _2873_;
  wire _2874_;
  wire _2875_;
  wire _2876_;
  wire _2877_;
  wire _2878_;
  wire _2879_;
  wire _2880_;
  wire _2881_;
  wire _2882_;
  wire _2883_;
  wire _2884_;
  wire _2885_;
  wire _2886_;
  wire _2887_;
  wire _2888_;
  wire _2889_;
  wire _2890_;
  wire _2891_;
  wire _2892_;
  wire _2893_;
  wire _2894_;
  wire _2895_;
  wire _2896_;
  wire _2897_;
  wire _2898_;
  wire _2899_;
  wire _2900_;
  wire _2901_;
  wire _2902_;
  wire _2903_;
  wire _2904_;
  wire _2905_;
  wire _2906_;
  wire _2907_;
  wire _2908_;
  wire _2909_;
  wire _2910_;
  wire _2911_;
  wire _2912_;
  wire _2913_;
  wire _2914_;
  wire _2915_;
  wire _2916_;
  wire _2917_;
  wire _2918_;
  wire _2919_;
  wire _2920_;
  wire _2921_;
  wire _2922_;
  wire _2923_;
  wire _2924_;
  wire _2925_;
  wire _2926_;
  wire _2927_;
  wire _2928_;
  wire _2929_;
  wire _2930_;
  wire _2931_;
  wire _2932_;
  wire _2933_;
  wire _2934_;
  wire _2935_;
  wire _2936_;
  wire _2937_;
  wire _2938_;
  wire _2939_;
  wire _2940_;
  wire _2941_;
  wire _2942_;
  wire _2943_;
  wire _2944_;
  wire _2945_;
  wire _2946_;
  wire _2947_;
  wire _2948_;
  wire _2949_;
  wire _2950_;
  wire _2951_;
  wire _2952_;
  wire _2953_;
  wire _2954_;
  wire _2955_;
  wire _2956_;
  wire _2957_;
  wire _2958_;
  wire _2959_;
  wire _2960_;
  wire _2961_;
  wire _2962_;
  wire _2963_;
  wire _2964_;
  wire _2965_;
  wire _2966_;
  wire _2967_;
  wire _2968_;
  wire _2969_;
  wire _2970_;
  wire _2971_;
  wire _2972_;
  wire _2973_;
  wire _2974_;
  wire _2975_;
  wire _2976_;
  wire _2977_;
  wire _2978_;
  wire _2979_;
  wire _2980_;
  wire _2981_;
  wire _2982_;
  wire _2983_;
  wire _2984_;
  wire _2985_;
  wire _2986_;
  wire _2987_;
  wire _2988_;
  wire _2989_;
  wire _2990_;
  wire _2991_;
  wire _2992_;
  wire _2993_;
  wire _2994_;
  wire _2995_;
  wire _2996_;
  wire _2997_;
  wire _2998_;
  wire _2999_;
  wire _3000_;
  wire _3001_;
  wire _3002_;
  wire _3003_;
  wire _3004_;
  wire _3005_;
  wire _3006_;
  wire _3007_;
  wire _3008_;
  wire _3009_;
  wire _3010_;
  wire _3011_;
  wire _3012_;
  wire _3013_;
  wire _3014_;
  wire _3015_;
  wire _3016_;
  wire _3017_;
  wire _3018_;
  wire _3019_;
  wire _3020_;
  wire _3021_;
  wire _3022_;
  wire _3023_;
  wire _3024_;
  wire _3025_;
  wire _3026_;
  wire _3027_;
  wire _3028_;
  wire _3029_;
  wire _3030_;
  wire _3031_;
  wire _3032_;
  wire _3033_;
  wire _3034_;
  wire _3035_;
  wire _3036_;
  wire _3037_;
  wire _3038_;
  wire _3039_;
  wire _3040_;
  wire _3041_;
  wire _3042_;
  wire _3043_;
  wire _3044_;
  wire _3045_;
  wire _3046_;
  wire _3047_;
  wire _3048_;
  wire _3049_;
  wire _3050_;
  wire _3051_;
  wire _3052_;
  wire _3053_;
  wire _3054_;
  wire _3055_;
  wire _3056_;
  wire _3057_;
  wire _3058_;
  wire _3059_;
  wire _3060_;
  wire _3061_;
  wire _3062_;
  wire _3063_;
  wire _3064_;
  wire _3065_;
  wire _3066_;
  wire _3067_;
  wire _3068_;
  wire _3069_;
  wire _3070_;
  wire _3071_;
  wire _3072_;
  wire _3073_;
  wire _3074_;
  wire _3075_;
  wire _3076_;
  wire _3077_;
  wire _3078_;
  wire _3079_;
  wire _3080_;
  wire _3081_;
  wire _3082_;
  wire _3083_;
  wire _3084_;
  wire _3085_;
  wire _3086_;
  wire _3087_;
  wire _3088_;
  wire _3089_;
  wire _3090_;
  wire _3091_;
  wire _3092_;
  wire _3093_;
  wire _3094_;
  wire _3095_;
  wire _3096_;
  wire _3097_;
  wire _3098_;
  wire _3099_;
  wire _3100_;
  wire _3101_;
  wire _3102_;
  wire _3103_;
  wire _3104_;
  wire _3105_;
  wire _3106_;
  wire _3107_;
  wire _3108_;
  wire _3109_;
  wire _3110_;
  wire _3111_;
  wire _3112_;
  wire _3113_;
  wire _3114_;
  wire _3115_;
  wire _3116_;
  wire _3117_;
  wire _3118_;
  wire _3119_;
  wire _3120_;
  wire _3121_;
  wire _3122_;
  wire _3123_;
  wire _3124_;
  wire _3125_;
  wire _3126_;
  wire _3127_;
  wire _3128_;
  wire _3129_;
  wire _3130_;
  wire _3131_;
  wire _3132_;
  wire _3133_;
  wire _3134_;
  wire _3135_;
  wire _3136_;
  wire _3137_;
  wire _3138_;
  wire _3139_;
  wire _3140_;
  wire _3141_;
  wire _3142_;
  wire _3143_;
  wire _3144_;
  wire _3145_;
  wire _3146_;
  wire _3147_;
  wire _3148_;
  wire _3149_;
  wire _3150_;
  wire _3151_;
  wire _3152_;
  wire _3153_;
  wire _3154_;
  wire _3155_;
  wire _3156_;
  wire _3157_;
  wire _3158_;
  wire _3159_;
  wire _3160_;
  wire _3161_;
  wire _3162_;
  wire _3163_;
  wire _3164_;
  wire _3165_;
  wire _3166_;
  wire _3167_;
  wire _3168_;
  wire _3169_;
  wire _3170_;
  wire _3171_;
  wire _3172_;
  wire _3173_;
  wire _3174_;
  wire _3175_;
  wire _3176_;
  wire _3177_;
  wire _3178_;
  wire _3179_;
  wire _3180_;
  wire _3181_;
  wire _3182_;
  wire _3183_;
  wire _3184_;
  wire _3185_;
  wire _3186_;
  wire _3187_;
  wire _3188_;
  wire _3189_;
  wire _3190_;
  wire _3191_;
  wire _3192_;
  wire _3193_;
  wire _3194_;
  wire _3195_;
  wire _3196_;
  wire _3197_;
  wire _3198_;
  wire _3199_;
  wire _3200_;
  wire _3201_;
  wire _3202_;
  wire _3203_;
  wire _3204_;
  wire _3205_;
  wire _3206_;
  wire _3207_;
  wire _3208_;
  wire _3209_;
  wire _3210_;
  wire _3211_;
  wire _3212_;
  wire _3213_;
  wire _3214_;
  wire _3215_;
  wire _3216_;
  wire _3217_;
  wire _3218_;
  wire _3219_;
  wire _3220_;
  wire _3221_;
  wire _3222_;
  wire _3223_;
  wire _3224_;
  wire _3225_;
  wire _3226_;
  wire _3227_;
  wire _3228_;
  wire _3229_;
  wire _3230_;
  wire _3231_;
  wire _3232_;
  wire _3233_;
  wire _3234_;
  wire _3235_;
  wire _3236_;
  wire _3237_;
  wire _3238_;
  wire _3239_;
  wire _3240_;
  wire _3241_;
  wire _3242_;
  wire _3243_;
  wire _3244_;
  wire _3245_;
  wire _3246_;
  wire _3247_;
  wire _3248_;
  wire _3249_;
  wire _3250_;
  wire _3251_;
  wire _3252_;
  wire _3253_;
  wire _3254_;
  wire _3255_;
  wire _3256_;
  wire _3257_;
  wire _3258_;
  wire _3259_;
  wire _3260_;
  wire _3261_;
  wire _3262_;
  wire _3263_;
  wire _3264_;
  wire _3265_;
  wire _3266_;
  wire _3267_;
  wire _3268_;
  wire _3269_;
  wire _3270_;
  wire _3271_;
  wire _3272_;
  wire _3273_;
  wire _3274_;
  wire _3275_;
  wire _3276_;
  wire _3277_;
  wire _3278_;
  wire _3279_;
  wire _3280_;
  wire _3281_;
  wire _3282_;
  wire _3283_;
  wire _3284_;
  wire _3285_;
  wire _3286_;
  wire _3287_;
  wire _3288_;
  wire _3289_;
  wire _3290_;
  wire _3291_;
  wire _3292_;
  wire _3293_;
  wire _3294_;
  wire _3295_;
  wire _3296_;
  wire _3297_;
  wire _3298_;
  wire _3299_;
  wire _3300_;
  wire _3301_;
  wire _3302_;
  wire _3303_;
  wire _3304_;
  wire _3305_;
  wire _3306_;
  wire _3307_;
  wire _3308_;
  wire _3309_;
  wire _3310_;
  wire _3311_;
  wire _3312_;
  wire _3313_;
  wire _3314_;
  wire _3315_;
  wire _3316_;
  wire _3317_;
  wire _3318_;
  wire _3319_;
  wire _3320_;
  wire _3321_;
  wire _3322_;
  wire _3323_;
  wire _3324_;
  wire _3325_;
  wire _3326_;
  wire _3327_;
  wire _3328_;
  wire _3329_;
  wire _3330_;
  wire _3331_;
  wire _3332_;
  wire _3333_;
  wire _3334_;
  wire _3335_;
  wire _3336_;
  wire _3337_;
  wire _3338_;
  wire _3339_;
  wire _3340_;
  wire _3341_;
  wire _3342_;
  wire _3343_;
  wire _3344_;
  wire _3345_;
  wire _3346_;
  wire _3347_;
  wire _3348_;
  wire _3349_;
  wire _3350_;
  wire _3351_;
  wire _3352_;
  wire _3353_;
  wire _3354_;
  wire _3355_;
  wire _3356_;
  wire _3357_;
  wire _3358_;
  wire _3359_;
  wire _3360_;
  wire _3361_;
  wire _3362_;
  wire _3363_;
  wire _3364_;
  wire _3365_;
  wire _3366_;
  wire _3367_;
  wire _3368_;
  wire _3369_;
  wire _3370_;
  wire _3371_;
  wire _3372_;
  wire _3373_;
  wire _3374_;
  wire _3375_;
  wire _3376_;
  wire _3377_;
  wire _3378_;
  wire _3379_;
  wire _3380_;
  wire _3381_;
  wire _3382_;
  wire _3383_;
  wire _3384_;
  wire _3385_;
  wire _3386_;
  wire _3387_;
  wire _3388_;
  wire _3389_;
  wire _3390_;
  wire _3391_;
  wire _3392_;
  wire _3393_;
  wire _3394_;
  wire _3395_;
  wire _3396_;
  wire _3397_;
  wire _3398_;
  wire _3399_;
  wire _3400_;
  wire _3401_;
  wire _3402_;
  wire _3403_;
  wire _3404_;
  wire _3405_;
  wire _3406_;
  wire _3407_;
  wire _3408_;
  wire _3409_;
  wire _3410_;
  wire _3411_;
  wire _3412_;
  wire _3413_;
  wire _3414_;
  wire _3415_;
  wire _3416_;
  wire _3417_;
  wire _3418_;
  wire _3419_;
  wire _3420_;
  wire _3421_;
  wire _3422_;
  wire _3423_;
  wire _3424_;
  wire _3425_;
  wire _3426_;
  wire _3427_;
  wire _3428_;
  wire _3429_;
  wire _3430_;
  wire _3431_;
  wire _3432_;
  wire _3433_;
  wire _3434_;
  wire _3435_;
  wire _3436_;
  wire _3437_;
  wire _3438_;
  wire _3439_;
  wire _3440_;
  wire _3441_;
  wire _3442_;
  wire _3443_;
  wire _3444_;
  wire _3445_;
  wire _3446_;
  wire _3447_;
  wire _3448_;
  wire _3449_;
  wire _3450_;
  wire _3451_;
  wire _3452_;
  wire _3453_;
  wire _3454_;
  wire _3455_;
  wire _3456_;
  wire _3457_;
  wire _3458_;
  wire _3459_;
  wire _3460_;
  wire _3461_;
  wire _3462_;
  wire _3463_;
  wire _3464_;
  wire _3465_;
  wire _3466_;
  wire _3467_;
  wire _3468_;
  wire _3469_;
  wire _3470_;
  wire _3471_;
  wire _3472_;
  wire _3473_;
  wire _3474_;
  wire _3475_;
  wire _3476_;
  wire _3477_;
  wire _3478_;
  wire _3479_;
  wire _3480_;
  wire _3481_;
  wire _3482_;
  wire _3483_;
  wire _3484_;
  wire _3485_;
  wire _3486_;
  wire _3487_;
  wire _3488_;
  wire _3489_;
  wire _3490_;
  wire _3491_;
  wire _3492_;
  wire _3493_;
  wire _3494_;
  wire _3495_;
  wire _3496_;
  wire _3497_;
  wire _3498_;
  wire _3499_;
  wire _3500_;
  wire _3501_;
  wire _3502_;
  wire _3503_;
  wire _3504_;
  wire _3505_;
  wire _3506_;
  wire _3507_;
  wire _3508_;
  wire _3509_;
  wire _3510_;
  wire _3511_;
  wire _3512_;
  wire _3513_;
  wire _3514_;
  wire _3515_;
  wire _3516_;
  wire _3517_;
  wire _3518_;
  wire _3519_;
  wire _3520_;
  wire _3521_;
  wire _3522_;
  wire _3523_;
  wire _3524_;
  wire _3525_;
  wire _3526_;
  wire _3527_;
  wire _3528_;
  wire _3529_;
  wire _3530_;
  wire _3531_;
  wire _3532_;
  wire _3533_;
  wire _3534_;
  wire _3535_;
  wire _3536_;
  wire _3537_;
  wire _3538_;
  wire _3539_;
  wire _3540_;
  wire _3541_;
  wire _3542_;
  wire _3543_;
  wire _3544_;
  wire _3545_;
  wire _3546_;
  wire _3547_;
  wire _3548_;
  wire _3549_;
  wire _3550_;
  wire _3551_;
  wire _3552_;
  wire _3553_;
  wire _3554_;
  wire _3555_;
  wire _3556_;
  wire _3557_;
  wire _3558_;
  wire _3559_;
  wire _3560_;
  wire _3561_;
  wire _3562_;
  wire _3563_;
  wire _3564_;
  wire _3565_;
  wire _3566_;
  wire _3567_;
  wire _3568_;
  wire _3569_;
  wire _3570_;
  wire _3571_;
  wire _3572_;
  wire _3573_;
  wire _3574_;
  wire _3575_;
  wire _3576_;
  wire _3577_;
  wire _3578_;
  wire _3579_;
  wire _3580_;
  wire _3581_;
  wire _3582_;
  wire _3583_;
  wire _3584_;
  wire _3585_;
  wire _3586_;
  wire _3587_;
  wire _3588_;
  wire _3589_;
  wire _3590_;
  wire _3591_;
  wire _3592_;
  wire _3593_;
  wire _3594_;
  wire _3595_;
  wire _3596_;
  wire _3597_;
  wire _3598_;
  wire _3599_;
  wire _3600_;
  wire _3601_;
  wire _3602_;
  wire _3603_;
  wire _3604_;
  wire _3605_;
  wire _3606_;
  wire _3607_;
  wire _3608_;
  wire _3609_;
  wire _3610_;
  wire _3611_;
  wire _3612_;
  wire _3613_;
  wire _3614_;
  wire _3615_;
  wire _3616_;
  wire _3617_;
  wire _3618_;
  wire _3619_;
  wire _3620_;
  wire _3621_;
  wire _3622_;
  wire _3623_;
  wire _3624_;
  wire _3625_;
  wire _3626_;
  wire _3627_;
  wire _3628_;
  wire _3629_;
  wire _3630_;
  wire _3631_;
  wire _3632_;
  wire _3633_;
  wire _3634_;
  wire _3635_;
  wire _3636_;
  wire _3637_;
  wire _3638_;
  wire _3639_;
  wire _3640_;
  wire _3641_;
  wire _3642_;
  wire _3643_;
  wire _3644_;
  wire _3645_;
  wire _3646_;
  wire _3647_;
  wire _3648_;
  wire _3649_;
  wire _3650_;
  wire _3651_;
  wire _3652_;
  wire _3653_;
  wire _3654_;
  wire _3655_;
  wire _3656_;
  wire _3657_;
  wire _3658_;
  wire _3659_;
  wire _3660_;
  wire _3661_;
  wire _3662_;
  wire _3663_;
  wire _3664_;
  wire _3665_;
  wire _3666_;
  wire _3667_;
  wire _3668_;
  wire _3669_;
  wire _3670_;
  wire _3671_;
  wire _3672_;
  wire _3673_;
  wire _3674_;
  wire _3675_;
  wire _3676_;
  wire _3677_;
  wire _3678_;
  wire _3679_;
  wire _3680_;
  wire _3681_;
  wire _3682_;
  wire _3683_;
  wire _3684_;
  wire _3685_;
  wire _3686_;
  wire _3687_;
  wire _3688_;
  wire _3689_;
  wire _3690_;
  wire _3691_;
  wire _3692_;
  wire _3693_;
  wire _3694_;
  wire _3695_;
  wire _3696_;
  wire _3697_;
  wire _3698_;
  wire _3699_;
  wire _3700_;
  wire _3701_;
  wire _3702_;
  wire _3703_;
  wire _3704_;
  wire _3705_;
  wire _3706_;
  wire _3707_;
  wire _3708_;
  wire _3709_;
  wire _3710_;
  wire _3711_;
  wire _3712_;
  wire _3713_;
  wire _3714_;
  wire _3715_;
  wire _3716_;
  wire _3717_;
  wire _3718_;
  wire _3719_;
  wire _3720_;
  wire _3721_;
  wire _3722_;
  wire _3723_;
  wire _3724_;
  wire _3725_;
  wire _3726_;
  wire _3727_;
  wire _3728_;
  wire _3729_;
  wire _3730_;
  wire _3731_;
  wire _3732_;
  wire _3733_;
  wire _3734_;
  wire _3735_;
  wire _3736_;
  wire _3737_;
  wire _3738_;
  wire _3739_;
  wire _3740_;
  wire _3741_;
  wire _3742_;
  wire _3743_;
  wire _3744_;
  wire _3745_;
  wire _3746_;
  wire _3747_;
  wire _3748_;
  wire _3749_;
  wire _3750_;
  wire _3751_;
  wire _3752_;
  wire _3753_;
  wire _3754_;
  wire _3755_;
  wire _3756_;
  wire _3757_;
  wire _3758_;
  wire _3759_;
  wire _3760_;
  wire _3761_;
  wire _3762_;
  wire _3763_;
  wire _3764_;
  wire _3765_;
  wire _3766_;
  wire _3767_;
  wire _3768_;
  wire _3769_;
  wire _3770_;
  wire _3771_;
  wire _3772_;
  wire _3773_;
  wire _3774_;
  wire _3775_;
  wire _3776_;
  wire _3777_;
  wire _3778_;
  wire _3779_;
  wire _3780_;
  wire _3781_;
  wire _3782_;
  wire _3783_;
  wire _3784_;
  wire _3785_;
  wire _3786_;
  wire _3787_;
  wire _3788_;
  wire _3789_;
  wire _3790_;
  wire _3791_;
  wire _3792_;
  wire _3793_;
  wire _3794_;
  wire _3795_;
  wire _3796_;
  wire _3797_;
  wire _3798_;
  wire _3799_;
  wire _3800_;
  wire _3801_;
  wire _3802_;
  wire _3803_;
  wire _3804_;
  wire _3805_;
  wire _3806_;
  wire _3807_;
  wire _3808_;
  wire _3809_;
  wire _3810_;
  wire _3811_;
  wire _3812_;
  wire _3813_;
  wire _3814_;
  wire _3815_;
  wire _3816_;
  wire _3817_;
  wire _3818_;
  wire _3819_;
  wire _3820_;
  wire _3821_;
  wire _3822_;
  wire _3823_;
  wire _3824_;
  wire _3825_;
  wire _3826_;
  wire _3827_;
  wire _3828_;
  wire _3829_;
  wire _3830_;
  wire _3831_;
  wire _3832_;
  wire _3833_;
  wire _3834_;
  wire _3835_;
  wire _3836_;
  wire _3837_;
  wire _3838_;
  wire _3839_;
  wire _3840_;
  wire _3841_;
  wire _3842_;
  wire _3843_;
  wire _3844_;
  wire _3845_;
  wire _3846_;
  wire _3847_;
  wire _3848_;
  wire _3849_;
  wire _3850_;
  wire _3851_;
  wire _3852_;
  wire _3853_;
  wire _3854_;
  wire _3855_;
  wire _3856_;
  wire _3857_;
  wire _3858_;
  wire _3859_;
  wire _3860_;
  wire _3861_;
  wire _3862_;
  wire _3863_;
  wire _3864_;
  wire _3865_;
  wire _3866_;
  wire _3867_;
  wire _3868_;
  wire _3869_;
  wire _3870_;
  wire _3871_;
  wire _3872_;
  wire _3873_;
  wire _3874_;
  wire _3875_;
  wire _3876_;
  wire _3877_;
  wire _3878_;
  wire _3879_;
  wire _3880_;
  wire _3881_;
  wire _3882_;
  wire _3883_;
  wire _3884_;
  wire _3885_;
  wire _3886_;
  wire _3887_;
  wire _3888_;
  wire _3889_;
  wire _3890_;
  wire _3891_;
  wire _3892_;
  wire _3893_;
  wire _3894_;
  wire _3895_;
  wire _3896_;
  wire _3897_;
  wire _3898_;
  wire _3899_;
  wire _3900_;
  wire _3901_;
  wire _3902_;
  wire _3903_;
  wire _3904_;
  wire _3905_;
  wire _3906_;
  wire _3907_;
  wire _3908_;
  wire _3909_;
  wire _3910_;
  wire _3911_;
  wire _3912_;
  wire _3913_;
  wire _3914_;
  wire _3915_;
  wire _3916_;
  wire _3917_;
  wire _3918_;
  wire _3919_;
  wire _3920_;
  wire _3921_;
  wire _3922_;
  wire _3923_;
  wire _3924_;
  wire _3925_;
  wire _3926_;
  wire _3927_;
  wire _3928_;
  wire _3929_;
  wire _3930_;
  wire _3931_;
  wire _3932_;
  wire _3933_;
  wire _3934_;
  wire _3935_;
  wire _3936_;
  wire _3937_;
  wire _3938_;
  wire _3939_;
  wire _3940_;
  wire _3941_;
  wire _3942_;
  wire _3943_;
  wire _3944_;
  wire _3945_;
  wire _3946_;
  wire _3947_;
  wire _3948_;
  wire _3949_;
  wire _3950_;
  wire _3951_;
  wire _3952_;
  wire _3953_;
  wire _3954_;
  wire _3955_;
  wire _3956_;
  wire _3957_;
  wire _3958_;
  wire _3959_;
  wire _3960_;
  wire _3961_;
  wire _3962_;
  wire _3963_;
  wire _3964_;
  wire _3965_;
  wire _3966_;
  wire _3967_;
  wire _3968_;
  wire _3969_;
  wire _3970_;
  wire _3971_;
  wire _3972_;
  wire _3973_;
  wire _3974_;
  wire _3975_;
  wire _3976_;
  wire _3977_;
  wire _3978_;
  wire _3979_;
  wire _3980_;
  wire _3981_;
  wire _3982_;
  wire _3983_;
  wire _3984_;
  wire _3985_;
  wire _3986_;
  wire _3987_;
  wire _3988_;
  wire _3989_;
  wire _3990_;
  wire _3991_;
  wire _3992_;
  wire _3993_;
  wire _3994_;
  wire _3995_;
  wire _3996_;
  wire _3997_;
  wire _3998_;
  wire _3999_;
  wire _4000_;
  wire _4001_;
  wire _4002_;
  wire _4003_;
  wire _4004_;
  wire _4005_;
  wire _4006_;
  wire _4007_;
  wire _4008_;
  wire _4009_;
  wire _4010_;
  wire _4011_;
  wire _4012_;
  wire _4013_;
  wire _4014_;
  wire _4015_;
  wire _4016_;
  wire _4017_;
  wire _4018_;
  wire _4019_;
  wire _4020_;
  wire _4021_;
  wire _4022_;
  wire _4023_;
  wire _4024_;
  wire _4025_;
  wire _4026_;
  wire _4027_;
  wire _4028_;
  wire _4029_;
  wire _4030_;
  wire _4031_;
  wire _4032_;
  wire _4033_;
  wire _4034_;
  wire _4035_;
  wire _4036_;
  wire _4037_;
  wire _4038_;
  wire _4039_;
  wire _4040_;
  wire _4041_;
  wire _4042_;
  wire _4043_;
  wire _4044_;
  wire _4045_;
  wire _4046_;
  wire _4047_;
  wire _4048_;
  wire _4049_;
  wire _4050_;
  wire _4051_;
  wire _4052_;
  wire _4053_;
  wire _4054_;
  wire _4055_;
  wire _4056_;
  wire _4057_;
  wire _4058_;
  wire _4059_;
  wire _4060_;
  wire _4061_;
  wire _4062_;
  wire _4063_;
  wire _4064_;
  wire _4065_;
  wire _4066_;
  wire _4067_;
  wire _4068_;
  wire _4069_;
  wire _4070_;
  wire _4071_;
  wire _4072_;
  wire _4073_;
  wire _4074_;
  wire _4075_;
  wire _4076_;
  wire _4077_;
  wire _4078_;
  wire _4079_;
  wire _4080_;
  wire _4081_;
  wire _4082_;
  wire _4083_;
  wire _4084_;
  wire _4085_;
  wire _4086_;
  wire _4087_;
  wire _4088_;
  wire _4089_;
  wire _4090_;
  wire _4091_;
  wire _4092_;
  wire _4093_;
  wire _4094_;
  wire _4095_;
  wire _4096_;
  wire _4097_;
  wire _4098_;
  wire _4099_;
  wire _4100_;
  wire _4101_;
  wire _4102_;
  wire _4103_;
  wire _4104_;
  wire _4105_;
  wire _4106_;
  wire _4107_;
  wire _4108_;
  wire _4109_;
  wire _4110_;
  wire _4111_;
  wire _4112_;
  wire _4113_;
  wire _4114_;
  wire _4115_;
  wire _4116_;
  wire _4117_;
  wire _4118_;
  wire _4119_;
  wire _4120_;
  wire _4121_;
  wire _4122_;
  wire _4123_;
  wire _4124_;
  wire _4125_;
  wire _4126_;
  wire _4127_;
  wire _4128_;
  wire _4129_;
  wire _4130_;
  wire _4131_;
  wire _4132_;
  wire _4133_;
  wire _4134_;
  wire _4135_;
  wire _4136_;
  wire _4137_;
  wire _4138_;
  wire _4139_;
  wire _4140_;
  wire _4141_;
  wire _4142_;
  wire _4143_;
  wire _4144_;
  wire _4145_;
  wire _4146_;
  wire _4147_;
  wire _4148_;
  wire _4149_;
  wire _4150_;
  wire _4151_;
  wire _4152_;
  wire _4153_;
  wire _4154_;
  wire _4155_;
  wire _4156_;
  wire _4157_;
  wire _4158_;
  wire _4159_;
  wire _4160_;
  wire _4161_;
  wire _4162_;
  wire _4163_;
  wire _4164_;
  wire _4165_;
  wire _4166_;
  wire _4167_;
  wire _4168_;
  wire _4169_;
  wire _4170_;
  wire _4171_;
  wire _4172_;
  wire _4173_;
  wire _4174_;
  wire _4175_;
  wire _4176_;
  wire _4177_;
  wire _4178_;
  wire _4179_;
  wire _4180_;
  wire _4181_;
  wire _4182_;
  wire _4183_;
  wire _4184_;
  wire _4185_;
  wire _4186_;
  wire _4187_;
  wire _4188_;
  wire _4189_;
  wire _4190_;
  wire _4191_;
  wire _4192_;
  wire _4193_;
  wire _4194_;
  wire _4195_;
  wire _4196_;
  wire _4197_;
  wire _4198_;
  wire _4199_;
  wire _4200_;
  wire _4201_;
  wire _4202_;
  wire _4203_;
  wire _4204_;
  wire _4205_;
  wire _4206_;
  wire _4207_;
  wire _4208_;
  wire _4209_;
  wire _4210_;
  wire _4211_;
  wire _4212_;
  wire _4213_;
  wire _4214_;
  wire _4215_;
  wire _4216_;
  wire _4217_;
  wire _4218_;
  wire _4219_;
  wire _4220_;
  wire _4221_;
  wire _4222_;
  wire _4223_;
  wire _4224_;
  wire _4225_;
  wire _4226_;
  wire _4227_;
  wire _4228_;
  wire _4229_;
  wire _4230_;
  wire _4231_;
  wire _4232_;
  wire _4233_;
  wire _4234_;
  wire _4235_;
  wire _4236_;
  wire _4237_;
  wire _4238_;
  wire _4239_;
  wire _4240_;
  wire _4241_;
  wire _4242_;
  wire _4243_;
  wire _4244_;
  wire _4245_;
  wire _4246_;
  wire _4247_;
  wire _4248_;
  wire _4249_;
  wire _4250_;
  wire _4251_;
  wire _4252_;
  wire _4253_;
  wire _4254_;
  wire _4255_;
  wire _4256_;
  wire _4257_;
  wire _4258_;
  wire _4259_;
  wire _4260_;
  wire _4261_;
  wire _4262_;
  wire _4263_;
  wire _4264_;
  wire _4265_;
  wire _4266_;
  wire _4267_;
  wire _4268_;
  wire _4269_;
  wire _4270_;
  wire _4271_;
  wire _4272_;
  wire _4273_;
  wire _4274_;
  wire _4275_;
  wire _4276_;
  wire _4277_;
  wire _4278_;
  wire _4279_;
  wire _4280_;
  wire _4281_;
  wire _4282_;
  wire _4283_;
  wire _4284_;
  wire _4285_;
  wire _4286_;
  wire _4287_;
  wire _4288_;
  wire _4289_;
  wire _4290_;
  wire _4291_;
  wire _4292_;
  wire _4293_;
  wire _4294_;
  wire _4295_;
  wire _4296_;
  wire _4297_;
  wire _4298_;
  wire _4299_;
  wire _4300_;
  wire _4301_;
  wire _4302_;
  wire _4303_;
  wire _4304_;
  wire _4305_;
  wire _4306_;
  wire _4307_;
  wire _4308_;
  wire _4309_;
  wire _4310_;
  wire _4311_;
  wire _4312_;
  wire _4313_;
  wire _4314_;
  wire _4315_;
  wire _4316_;
  wire _4317_;
  wire _4318_;
  wire _4319_;
  wire _4320_;
  wire _4321_;
  wire _4322_;
  wire _4323_;
  wire _4324_;
  wire _4325_;
  wire _4326_;
  wire _4327_;
  wire _4328_;
  wire _4329_;
  wire _4330_;
  wire _4331_;
  wire _4332_;
  wire _4333_;
  wire _4334_;
  wire _4335_;
  wire _4336_;
  wire _4337_;
  wire _4338_;
  wire _4339_;
  wire _4340_;
  wire _4341_;
  wire _4342_;
  wire _4343_;
  wire _4344_;
  wire _4345_;
  wire _4346_;
  wire _4347_;
  wire _4348_;
  wire _4349_;
  wire _4350_;
  wire _4351_;
  wire _4352_;
  wire _4353_;
  wire _4354_;
  wire _4355_;
  wire _4356_;
  wire _4357_;
  wire _4358_;
  wire _4359_;
  wire _4360_;
  wire _4361_;
  wire _4362_;
  wire _4363_;
  wire _4364_;
  wire _4365_;
  wire _4366_;
  wire _4367_;
  wire _4368_;
  wire _4369_;
  wire _4370_;
  wire _4371_;
  wire _4372_;
  wire _4373_;
  wire _4374_;
  wire _4375_;
  wire _4376_;
  wire _4377_;
  wire _4378_;
  wire _4379_;
  wire _4380_;
  wire _4381_;
  wire _4382_;
  wire _4383_;
  wire _4384_;
  wire _4385_;
  wire _4386_;
  wire _4387_;
  wire _4388_;
  wire _4389_;
  wire _4390_;
  wire _4391_;
  wire _4392_;
  wire _4393_;
  wire _4394_;
  wire _4395_;
  wire _4396_;
  wire _4397_;
  wire _4398_;
  wire _4399_;
  wire _4400_;
  wire _4401_;
  wire _4402_;
  wire _4403_;
  wire _4404_;
  wire _4405_;
  wire _4406_;
  wire _4407_;
  wire _4408_;
  wire _4409_;
  wire _4410_;
  wire _4411_;
  wire _4412_;
  wire _4413_;
  wire _4414_;
  wire _4415_;
  wire _4416_;
  wire _4417_;
  wire _4418_;
  wire _4419_;
  wire _4420_;
  wire _4421_;
  wire _4422_;
  wire _4423_;
  wire _4424_;
  wire _4425_;
  wire _4426_;
  wire _4427_;
  wire _4428_;
  wire _4429_;
  wire _4430_;
  wire _4431_;
  wire _4432_;
  wire _4433_;
  wire _4434_;
  wire _4435_;
  wire _4436_;
  wire _4437_;
  wire _4438_;
  wire _4439_;
  wire _4440_;
  wire _4441_;
  wire _4442_;
  wire _4443_;
  wire _4444_;
  wire _4445_;
  wire _4446_;
  wire _4447_;
  wire _4448_;
  wire _4449_;
  wire _4450_;
  wire _4451_;
  wire _4452_;
  wire _4453_;
  wire _4454_;
  wire _4455_;
  wire _4456_;
  wire _4457_;
  wire _4458_;
  wire _4459_;
  wire _4460_;
  wire _4461_;
  wire _4462_;
  wire _4463_;
  wire _4464_;
  wire _4465_;
  wire _4466_;
  wire _4467_;
  wire _4468_;
  wire _4469_;
  wire _4470_;
  wire _4471_;
  wire _4472_;
  wire _4473_;
  wire _4474_;
  wire _4475_;
  wire _4476_;
  wire _4477_;
  wire _4478_;
  wire _4479_;
  wire _4480_;
  wire _4481_;
  wire _4482_;
  wire _4483_;
  wire _4484_;
  wire _4485_;
  wire _4486_;
  wire _4487_;
  wire _4488_;
  wire _4489_;
  wire _4490_;
  wire _4491_;
  wire _4492_;
  wire _4493_;
  wire _4494_;
  wire _4495_;
  wire _4496_;
  wire _4497_;
  wire _4498_;
  wire _4499_;
  wire _4500_;
  wire _4501_;
  wire _4502_;
  wire _4503_;
  wire _4504_;
  wire _4505_;
  wire _4506_;
  wire _4507_;
  wire _4508_;
  wire _4509_;
  wire _4510_;
  wire _4511_;
  wire _4512_;
  wire _4513_;
  wire _4514_;
  wire _4515_;
  wire _4516_;
  wire _4517_;
  wire _4518_;
  wire _4519_;
  wire _4520_;
  wire _4521_;
  wire _4522_;
  wire _4523_;
  wire _4524_;
  wire _4525_;
  wire _4526_;
  wire _4527_;
  wire _4528_;
  wire _4529_;
  wire _4530_;
  wire _4531_;
  wire _4532_;
  wire _4533_;
  wire _4534_;
  wire _4535_;
  wire _4536_;
  wire _4537_;
  wire _4538_;
  wire _4539_;
  wire _4540_;
  wire _4541_;
  wire _4542_;
  wire _4543_;
  wire _4544_;
  wire _4545_;
  wire _4546_;
  wire _4547_;
  wire _4548_;
  wire _4549_;
  wire _4550_;
  wire _4551_;
  wire _4552_;
  wire _4553_;
  wire _4554_;
  wire _4555_;
  wire _4556_;
  wire _4557_;
  wire _4558_;
  wire _4559_;
  wire _4560_;
  wire _4561_;
  wire _4562_;
  wire _4563_;
  wire _4564_;
  wire _4565_;
  wire _4566_;
  wire _4567_;
  wire _4568_;
  wire _4569_;
  wire _4570_;
  wire _4571_;
  wire _4572_;
  wire _4573_;
  wire _4574_;
  wire _4575_;
  wire _4576_;
  wire _4577_;
  wire _4578_;
  wire _4579_;
  wire _4580_;
  wire _4581_;
  wire _4582_;
  wire _4583_;
  wire _4584_;
  wire _4585_;
  wire _4586_;
  wire _4587_;
  wire _4588_;
  wire _4589_;
  wire _4590_;
  wire _4591_;
  wire _4592_;
  wire _4593_;
  wire _4594_;
  wire _4595_;
  wire _4596_;
  wire _4597_;
  wire _4598_;
  wire _4599_;
  wire _4600_;
  wire _4601_;
  wire _4602_;
  wire _4603_;
  wire _4604_;
  wire _4605_;
  wire _4606_;
  wire _4607_;
  wire _4608_;
  wire _4609_;
  wire _4610_;
  wire _4611_;
  wire _4612_;
  wire _4613_;
  wire _4614_;
  wire _4615_;
  wire _4616_;
  wire _4617_;
  wire _4618_;
  wire _4619_;
  wire _4620_;
  wire _4621_;
  wire _4622_;
  wire _4623_;
  wire _4624_;
  wire _4625_;
  wire _4626_;
  wire _4627_;
  wire _4628_;
  wire _4629_;
  wire _4630_;
  wire _4631_;
  wire _4632_;
  wire _4633_;
  wire _4634_;
  wire _4635_;
  wire _4636_;
  wire _4637_;
  wire _4638_;
  wire _4639_;
  wire _4640_;
  wire _4641_;
  wire _4642_;
  wire _4643_;
  wire _4644_;
  wire _4645_;
  wire _4646_;
  wire _4647_;
  wire _4648_;
  wire _4649_;
  wire _4650_;
  wire _4651_;
  wire _4652_;
  wire _4653_;
  wire _4654_;
  wire _4655_;
  wire _4656_;
  wire _4657_;
  wire _4658_;
  wire _4659_;
  wire _4660_;
  wire _4661_;
  wire _4662_;
  wire _4663_;
  wire _4664_;
  wire _4665_;
  wire _4666_;
  wire _4667_;
  wire _4668_;
  wire _4669_;
  wire _4670_;
  wire _4671_;
  wire _4672_;
  wire _4673_;
  wire _4674_;
  wire _4675_;
  wire _4676_;
  wire _4677_;
  wire _4678_;
  wire _4679_;
  wire _4680_;
  wire _4681_;
  wire _4682_;
  wire _4683_;
  wire _4684_;
  wire _4685_;
  wire _4686_;
  wire _4687_;
  wire _4688_;
  wire _4689_;
  wire _4690_;
  wire _4691_;
  wire _4692_;
  wire _4693_;
  wire _4694_;
  wire _4695_;
  wire _4696_;
  wire _4697_;
  wire _4698_;
  wire _4699_;
  wire _4700_;
  wire _4701_;
  wire _4702_;
  wire _4703_;
  wire _4704_;
  wire _4705_;
  wire _4706_;
  wire _4707_;
  wire _4708_;
  wire _4709_;
  wire _4710_;
  wire _4711_;
  wire _4712_;
  wire _4713_;
  wire _4714_;
  wire _4715_;
  wire _4716_;
  wire _4717_;
  wire _4718_;
  wire _4719_;
  wire _4720_;
  wire _4721_;
  wire _4722_;
  wire _4723_;
  wire _4724_;
  wire _4725_;
  wire _4726_;
  wire _4727_;
  wire _4728_;
  wire _4729_;
  wire _4730_;
  wire _4731_;
  wire _4732_;
  wire _4733_;
  wire _4734_;
  wire _4735_;
  wire _4736_;
  wire _4737_;
  wire _4738_;
  wire _4739_;
  wire _4740_;
  wire _4741_;
  wire _4742_;
  wire _4743_;
  wire _4744_;
  wire _4745_;
  wire _4746_;
  wire _4747_;
  wire _4748_;
  wire _4749_;
  wire _4750_;
  wire _4751_;
  wire _4752_;
  wire _4753_;
  wire _4754_;
  wire _4755_;
  wire _4756_;
  wire _4757_;
  wire _4758_;
  wire _4759_;
  wire _4760_;
  wire _4761_;
  wire _4762_;
  wire _4763_;
  wire _4764_;
  wire _4765_;
  wire _4766_;
  wire _4767_;
  wire _4768_;
  wire _4769_;
  wire _4770_;
  wire _4771_;
  wire _4772_;
  wire _4773_;
  wire _4774_;
  wire _4775_;
  wire _4776_;
  wire _4777_;
  wire _4778_;
  wire _4779_;
  wire _4780_;
  wire _4781_;
  wire _4782_;
  wire _4783_;
  wire _4784_;
  wire _4785_;
  wire _4786_;
  wire _4787_;
  wire _4788_;
  wire _4789_;
  wire _4790_;
  wire _4791_;
  wire _4792_;
  wire _4793_;
  wire _4794_;
  wire _4795_;
  wire _4796_;
  wire _4797_;
  wire _4798_;
  wire _4799_;
  wire _4800_;
  wire _4801_;
  wire _4802_;
  wire _4803_;
  wire _4804_;
  wire _4805_;
  wire _4806_;
  wire _4807_;
  wire _4808_;
  wire _4809_;
  wire _4810_;
  wire _4811_;
  wire _4812_;
  wire _4813_;
  wire _4814_;
  wire _4815_;
  wire _4816_;
  wire _4817_;
  wire _4818_;
  wire _4819_;
  wire _4820_;
  wire _4821_;
  wire _4822_;
  wire _4823_;
  wire _4824_;
  wire _4825_;
  wire _4826_;
  wire _4827_;
  wire _4828_;
  wire _4829_;
  wire _4830_;
  wire _4831_;
  wire _4832_;
  wire _4833_;
  wire _4834_;
  wire _4835_;
  wire _4836_;
  wire _4837_;
  wire _4838_;
  wire _4839_;
  wire _4840_;
  wire _4841_;
  wire _4842_;
  wire _4843_;
  wire _4844_;
  wire _4845_;
  wire _4846_;
  wire _4847_;
  wire _4848_;
  wire _4849_;
  wire _4850_;
  wire _4851_;
  wire _4852_;
  wire _4853_;
  wire _4854_;
  wire _4855_;
  wire _4856_;
  wire _4857_;
  wire _4858_;
  wire _4859_;
  wire _4860_;
  wire _4861_;
  wire _4862_;
  wire _4863_;
  wire _4864_;
  wire _4865_;
  wire _4866_;
  wire _4867_;
  wire _4868_;
  wire _4869_;
  wire _4870_;
  wire _4871_;
  wire _4872_;
  wire _4873_;
  wire _4874_;
  wire _4875_;
  wire _4876_;
  wire _4877_;
  wire _4878_;
  wire _4879_;
  wire _4880_;
  wire _4881_;
  wire _4882_;
  wire _4883_;
  wire _4884_;
  wire _4885_;
  wire _4886_;
  wire _4887_;
  wire _4888_;
  wire _4889_;
  wire _4890_;
  wire _4891_;
  wire _4892_;
  wire _4893_;
  wire _4894_;
  wire _4895_;
  wire _4896_;
  wire _4897_;
  wire _4898_;
  wire _4899_;
  wire _4900_;
  wire _4901_;
  wire _4902_;
  wire _4903_;
  wire _4904_;
  wire _4905_;
  wire _4906_;
  wire _4907_;
  wire _4908_;
  wire _4909_;
  wire _4910_;
  wire _4911_;
  wire _4912_;
  wire _4913_;
  wire _4914_;
  wire _4915_;
  wire _4916_;
  wire _4917_;
  wire _4918_;
  wire _4919_;
  wire _4920_;
  wire _4921_;
  wire _4922_;
  wire _4923_;
  wire _4924_;
  wire _4925_;
  wire _4926_;
  wire _4927_;
  wire _4928_;
  wire _4929_;
  wire _4930_;
  wire _4931_;
  wire _4932_;
  wire _4933_;
  wire _4934_;
  wire _4935_;
  wire _4936_;
  wire _4937_;
  wire _4938_;
  wire _4939_;
  wire _4940_;
  wire _4941_;
  wire _4942_;
  wire _4943_;
  wire _4944_;
  wire _4945_;
  wire _4946_;
  wire _4947_;
  wire _4948_;
  wire _4949_;
  wire _4950_;
  wire _4951_;
  wire _4952_;
  wire _4953_;
  wire _4954_;
  wire _4955_;
  wire _4956_;
  wire _4957_;
  wire _4958_;
  wire _4959_;
  wire _4960_;
  wire _4961_;
  wire _4962_;
  wire _4963_;
  wire _4964_;
  wire _4965_;
  wire _4966_;
  wire _4967_;
  wire _4968_;
  wire _4969_;
  wire _4970_;
  wire _4971_;
  wire _4972_;
  wire _4973_;
  wire _4974_;
  wire _4975_;
  wire _4976_;
  wire _4977_;
  wire _4978_;
  wire _4979_;
  wire _4980_;
  wire _4981_;
  wire _4982_;
  wire _4983_;
  wire _4984_;
  wire _4985_;
  wire _4986_;
  wire _4987_;
  wire _4988_;
  wire _4989_;
  wire _4990_;
  wire _4991_;
  wire _4992_;
  wire _4993_;
  wire _4994_;
  wire _4995_;
  wire _4996_;
  wire _4997_;
  wire _4998_;
  wire _4999_;
  wire _5000_;
  wire _5001_;
  wire _5002_;
  wire _5003_;
  wire _5004_;
  wire _5005_;
  wire _5006_;
  wire _5007_;
  wire _5008_;
  wire _5009_;
  wire _5010_;
  wire _5011_;
  wire _5012_;
  wire _5013_;
  wire _5014_;
  wire _5015_;
  wire _5016_;
  wire _5017_;
  wire _5018_;
  wire _5019_;
  wire _5020_;
  wire _5021_;
  wire _5022_;
  wire _5023_;
  wire _5024_;
  wire _5025_;
  wire _5026_;
  wire _5027_;
  wire _5028_;
  wire _5029_;
  wire _5030_;
  wire _5031_;
  wire _5032_;
  wire _5033_;
  wire _5034_;
  wire _5035_;
  wire _5036_;
  wire _5037_;
  wire _5038_;
  wire _5039_;
  wire _5040_;
  wire _5041_;
  wire _5042_;
  wire _5043_;
  wire _5044_;
  wire _5045_;
  wire _5046_;
  wire _5047_;
  wire _5048_;
  wire _5049_;
  wire _5050_;
  wire _5051_;
  wire _5052_;
  wire _5053_;
  wire _5054_;
  wire _5055_;
  wire _5056_;
  wire _5057_;
  wire _5058_;
  wire _5059_;
  wire _5060_;
  wire _5061_;
  wire _5062_;
  wire _5063_;
  wire _5064_;
  wire _5065_;
  wire _5066_;
  wire _5067_;
  wire _5068_;
  wire _5069_;
  wire _5070_;
  wire _5071_;
  wire _5072_;
  wire _5073_;
  wire _5074_;
  wire _5075_;
  wire _5076_;
  wire _5077_;
  wire _5078_;
  wire _5079_;
  wire _5080_;
  wire _5081_;
  wire _5082_;
  wire _5083_;
  wire _5084_;
  wire _5085_;
  wire _5086_;
  wire _5087_;
  wire _5088_;
  wire _5089_;
  wire _5090_;
  wire _5091_;
  wire _5092_;
  wire _5093_;
  wire _5094_;
  wire _5095_;
  wire _5096_;
  wire _5097_;
  wire _5098_;
  wire _5099_;
  wire _5100_;
  wire _5101_;
  wire [1:0] _GEN_170;
  wire [1:0] _GEN_207;
  wire [31:0] _GEN_239;
  wire [5:0] _GEN_34;
  wire [5:0] _GEN_35;
  wire [31:0] _GEN_40;
  wire [31:0] _GEN_41;
  wire _GEN_51;
  wire [31:0] _GEN_586;
  wire [31:0] _GEN_592;
  wire [31:0] _GEN_593;
  wire [31:0] _GEN_594;
  wire [63:0] _GEN_595;
  wire [63:0] _GEN_596;
  wire [63:0] _GEN_597;
  wire [63:0] _GEN_598;
  wire [63:0] _GEN_599;
  wire [63:0] _GEN_600;
  wire [63:0] _GEN_601;
  wire [63:0] _GEN_602;
  wire [63:0] _GEN_603;
  wire [63:0] _GEN_604;
  wire [63:0] _GEN_605;
  wire [63:0] _GEN_606;
  wire [63:0] _GEN_607;
  wire [63:0] _GEN_608;
  wire [63:0] _GEN_609;
  wire [63:0] _GEN_610;
  wire [31:0] _GEN_611;
  wire [1:0] _GEN_73;
  wire _T_14;
  wire _T_15;
  wire [31:0] _T_16;
  wire [31:0] _T_18;
  wire [1:0] _T_20;
  wire [63:0] _T_2000;
  wire [63:0] _T_2003;
  wire [63:0] _T_2005;
  wire [63:0] _T_2008;
  wire [31:0] _T_21;
  wire [31:0] _T_213;
  wire [31:0] _T_22;
  wire [31:0] _T_23;
  wire [31:0] _T_24;
  wire [31:0] _T_27;
  wire [31:0] _T_28;
  wire [7:0] _T_60;
  wire [7:0] _T_62;
  wire [31:0] _T_64;
  wire [7:0] _T_65;
  wire [7:0] _T_67;
  wire [31:0] _T_69;
  wire _any_T_78;
  wire [3:0] _causeIsDebugBreak_T_3;
  wire [3:0] _causeIsDebugBreak_T_4;
  wire [11:0] _debugTVec_T;
  wire [1:0] _decoded_T_10;
  wire [11:0] _decoded_T_14;
  wire [3:0] _decoded_T_16;
  wire [9:0] _decoded_T_18;
  wire [11:0] _decoded_T_2;
  wire [9:0] _decoded_T_20;
  wire [1:0] _decoded_T_22;
  wire [3:0] _decoded_T_4;
  wire [9:0] _decoded_T_6;
  wire [9:0] _decoded_T_8;
  wire [11:0] _decoded_decoded_T;
  wire [10:0] _decoded_decoded_T_10;
  wire [11:0] _decoded_decoded_T_100;
  wire [11:0] _decoded_decoded_T_102;
  wire [11:0] _decoded_decoded_T_104;
  wire [11:0] _decoded_decoded_T_106;
  wire [11:0] _decoded_decoded_T_108;
  wire [11:0] _decoded_decoded_T_110;
  wire [11:0] _decoded_decoded_T_112;
  wire [11:0] _decoded_decoded_T_114;
  wire [11:0] _decoded_decoded_T_116;
  wire [11:0] _decoded_decoded_T_118;
  wire [11:0] _decoded_decoded_T_12;
  wire [11:0] _decoded_decoded_T_120;
  wire [11:0] _decoded_decoded_T_122;
  wire [11:0] _decoded_decoded_T_124;
  wire [11:0] _decoded_decoded_T_126;
  wire [11:0] _decoded_decoded_T_128;
  wire [10:0] _decoded_decoded_T_130;
  wire [5:0] _decoded_decoded_T_132;
  wire [10:0] _decoded_decoded_T_134;
  wire [11:0] _decoded_decoded_T_136;
  wire [11:0] _decoded_decoded_T_138;
  wire [11:0] _decoded_decoded_T_14;
  wire [11:0] _decoded_decoded_T_140;
  wire [11:0] _decoded_decoded_T_142;
  wire [11:0] _decoded_decoded_T_144;
  wire [11:0] _decoded_decoded_T_146;
  wire [11:0] _decoded_decoded_T_148;
  wire [11:0] _decoded_decoded_T_150;
  wire [11:0] _decoded_decoded_T_152;
  wire [11:0] _decoded_decoded_T_154;
  wire [11:0] _decoded_decoded_T_156;
  wire [11:0] _decoded_decoded_T_158;
  wire [11:0] _decoded_decoded_T_16;
  wire [11:0] _decoded_decoded_T_160;
  wire [11:0] _decoded_decoded_T_162;
  wire [11:0] _decoded_decoded_T_164;
  wire [11:0] _decoded_decoded_T_166;
  wire [11:0] _decoded_decoded_T_168;
  wire [11:0] _decoded_decoded_T_170;
  wire [11:0] _decoded_decoded_T_172;
  wire [11:0] _decoded_decoded_T_174;
  wire [11:0] _decoded_decoded_T_176;
  wire [11:0] _decoded_decoded_T_178;
  wire [11:0] _decoded_decoded_T_18;
  wire [11:0] _decoded_decoded_T_180;
  wire [11:0] _decoded_decoded_T_182;
  wire [11:0] _decoded_decoded_T_184;
  wire [11:0] _decoded_decoded_T_186;
  wire [11:0] _decoded_decoded_T_188;
  wire [11:0] _decoded_decoded_T_190;
  wire [11:0] _decoded_decoded_T_192;
  wire [11:0] _decoded_decoded_T_194;
  wire [10:0] _decoded_decoded_T_196;
  wire [11:0] _decoded_decoded_T_198;
  wire [11:0] _decoded_decoded_T_2;
  wire [11:0] _decoded_decoded_T_20;
  wire [11:0] _decoded_decoded_T_200;
  wire [11:0] _decoded_decoded_T_202;
  wire [11:0] _decoded_decoded_T_204;
  wire [11:0] _decoded_decoded_T_206;
  wire [11:0] _decoded_decoded_T_208;
  wire [11:0] _decoded_decoded_T_210;
  wire [11:0] _decoded_decoded_T_212;
  wire [11:0] _decoded_decoded_T_214;
  wire [11:0] _decoded_decoded_T_216;
  wire [11:0] _decoded_decoded_T_218;
  wire [11:0] _decoded_decoded_T_22;
  wire [11:0] _decoded_decoded_T_220;
  wire [11:0] _decoded_decoded_T_222;
  wire [11:0] _decoded_decoded_T_224;
  wire [11:0] _decoded_decoded_T_226;
  wire [11:0] _decoded_decoded_T_228;
  wire [11:0] _decoded_decoded_T_230;
  wire [11:0] _decoded_decoded_T_232;
  wire [11:0] _decoded_decoded_T_234;
  wire [11:0] _decoded_decoded_T_236;
  wire [11:0] _decoded_decoded_T_238;
  wire [11:0] _decoded_decoded_T_24;
  wire [11:0] _decoded_decoded_T_240;
  wire [11:0] _decoded_decoded_T_242;
  wire [11:0] _decoded_decoded_T_244;
  wire [11:0] _decoded_decoded_T_246;
  wire [11:0] _decoded_decoded_T_248;
  wire [11:0] _decoded_decoded_T_250;
  wire [11:0] _decoded_decoded_T_252;
  wire [11:0] _decoded_decoded_T_254;
  wire [11:0] _decoded_decoded_T_256;
  wire [10:0] _decoded_decoded_T_258;
  wire [11:0] _decoded_decoded_T_26;
  wire [11:0] _decoded_decoded_T_260;
  wire _decoded_decoded_T_261;
  wire [11:0] _decoded_decoded_T_262;
  wire _decoded_decoded_T_263;
  wire [9:0] _decoded_decoded_T_264;
  wire [11:0] _decoded_decoded_T_28;
  wire [11:0] _decoded_decoded_T_30;
  wire [11:0] _decoded_decoded_T_32;
  wire [11:0] _decoded_decoded_T_34;
  wire [11:0] _decoded_decoded_T_36;
  wire [11:0] _decoded_decoded_T_38;
  wire [11:0] _decoded_decoded_T_4;
  wire [11:0] _decoded_decoded_T_40;
  wire [11:0] _decoded_decoded_T_42;
  wire [11:0] _decoded_decoded_T_44;
  wire [11:0] _decoded_decoded_T_46;
  wire [11:0] _decoded_decoded_T_48;
  wire [11:0] _decoded_decoded_T_50;
  wire [11:0] _decoded_decoded_T_52;
  wire [11:0] _decoded_decoded_T_54;
  wire [11:0] _decoded_decoded_T_56;
  wire [11:0] _decoded_decoded_T_58;
  wire [11:0] _decoded_decoded_T_6;
  wire [11:0] _decoded_decoded_T_60;
  wire [11:0] _decoded_decoded_T_62;
  wire [11:0] _decoded_decoded_T_64;
  wire [11:0] _decoded_decoded_T_66;
  wire [11:0] _decoded_decoded_T_68;
  wire [11:0] _decoded_decoded_T_70;
  wire [11:0] _decoded_decoded_T_72;
  wire [11:0] _decoded_decoded_T_74;
  wire [9:0] _decoded_decoded_T_76;
  wire [11:0] _decoded_decoded_T_78;
  wire [10:0] _decoded_decoded_T_8;
  wire [11:0] _decoded_decoded_T_80;
  wire [11:0] _decoded_decoded_T_82;
  wire [11:0] _decoded_decoded_T_84;
  wire [11:0] _decoded_decoded_T_86;
  wire [11:0] _decoded_decoded_T_88;
  wire [11:0] _decoded_decoded_T_90;
  wire [11:0] _decoded_decoded_T_92;
  wire [11:0] _decoded_decoded_T_94;
  wire [11:0] _decoded_decoded_T_96;
  wire [11:0] _decoded_decoded_T_98;
  wire _decoded_decoded_orMatrixOutputs_T;
  wire _decoded_decoded_orMatrixOutputs_T_2;
  wire [31:0] _epc_T_1;
  wire [7:0] _io_decode_0_read_illegal_T_12;
  wire _io_decode_0_read_illegal_T_15;
  wire _io_decode_0_read_illegal_T_17;
  wire _io_decode_0_read_illegal_T_21;
  wire [31:0] _io_rw_rdata_T_1;
  wire [31:0] _io_rw_rdata_T_10;
  wire [31:0] _io_rw_rdata_T_107;
  wire [31:0] _io_rw_rdata_T_108;
  wire [31:0] _io_rw_rdata_T_109;
  wire [31:0] _io_rw_rdata_T_110;
  wire [29:0] _io_rw_rdata_T_113;
  wire [29:0] _io_rw_rdata_T_114;
  wire [29:0] _io_rw_rdata_T_115;
  wire [29:0] _io_rw_rdata_T_116;
  wire [29:0] _io_rw_rdata_T_117;
  wire [29:0] _io_rw_rdata_T_118;
  wire [29:0] _io_rw_rdata_T_119;
  wire [29:0] _io_rw_rdata_T_120;
  wire [31:0] _io_rw_rdata_T_129;
  wire _io_rw_rdata_T_13;
  wire [31:0] _io_rw_rdata_T_130;
  wire [31:0] _io_rw_rdata_T_132;
  wire [31:0] _io_rw_rdata_T_14;
  wire [31:0] _io_rw_rdata_T_148;
  wire [31:0] _io_rw_rdata_T_149;
  wire [31:0] _io_rw_rdata_T_15;
  wire [2:0] _io_rw_rdata_T_17;
  wire [63:0] _io_rw_rdata_T_240;
  wire [63:0] _io_rw_rdata_T_241;
  wire [63:0] _io_rw_rdata_T_242;
  wire [63:0] _io_rw_rdata_T_245;
  wire [63:0] _io_rw_rdata_T_246;
  wire [63:0] _io_rw_rdata_T_247;
  wire [63:0] _io_rw_rdata_T_248;
  wire [63:0] _io_rw_rdata_T_249;
  wire [63:0] _io_rw_rdata_T_250;
  wire [63:0] _io_rw_rdata_T_251;
  wire [63:0] _io_rw_rdata_T_252;
  wire [63:0] _io_rw_rdata_T_261;
  wire [63:0] _io_rw_rdata_T_262;
  wire [63:0] _io_rw_rdata_T_264;
  wire [31:0] _io_rw_rdata_T_4;
  wire [31:0] _io_rw_rdata_T_5;
  wire [31:0] _io_rw_rdata_T_6;
  wire [15:0] _io_rw_rdata_T_7;
  wire [31:0] _io_rw_rdata_T_8;
  wire [57:0] _large_r_T_1;
  wire [57:0] _large_r_T_3;
  wire [31:0] _m_interrupts_T_3;
  wire [31:0] _m_interrupts_T_5;
  wire [31:0] _newBPC_T_2;
  wire [31:0] _newBPC_T_3;
  wire [104:0] _new_mstatus_WIRE;
  wire [31:0] _notDebugTVec_T_1;
  wire [30:0] _pmp_mask_T_12;
  wire [30:0] _pmp_mask_T_13;
  wire [32:0] _pmp_mask_T_14;
  wire [30:0] _pmp_mask_T_17;
  wire [30:0] _pmp_mask_T_18;
  wire [32:0] _pmp_mask_T_19;
  wire [30:0] _pmp_mask_T_2;
  wire [30:0] _pmp_mask_T_22;
  wire [30:0] _pmp_mask_T_23;
  wire [32:0] _pmp_mask_T_24;
  wire [30:0] _pmp_mask_T_27;
  wire [30:0] _pmp_mask_T_28;
  wire [32:0] _pmp_mask_T_29;
  wire [30:0] _pmp_mask_T_3;
  wire [30:0] _pmp_mask_T_32;
  wire [30:0] _pmp_mask_T_33;
  wire [32:0] _pmp_mask_T_34;
  wire [30:0] _pmp_mask_T_37;
  wire [30:0] _pmp_mask_T_38;
  wire [32:0] _pmp_mask_T_39;
  wire [32:0] _pmp_mask_T_4;
  wire [30:0] _pmp_mask_T_7;
  wire [30:0] _pmp_mask_T_8;
  wire [32:0] _pmp_mask_T_9;
  wire [15:0] _read_mip_T;
  wire [104:0] _read_mstatus_T;
  wire [6:0] _read_mtvec_T_1;
  wire [31:0] _read_mtvec_T_3;
  wire [31:0] _read_mtvec_T_4;
  wire [31:0] _reg_custom_0_T;
  wire [31:0] _reg_custom_0_T_2;
  wire [31:0] _reg_custom_0_T_3;
  wire [2:0] _reg_dcsr_cause_T_2;
  wire [31:0] _reg_mcause_T;
  wire [31:0] _reg_mcountinhibit_T_1;
  wire [31:0] _reg_mepc_T_1;
  wire [31:0] _reg_mepc_T_2;
  wire [31:0] _reg_mie_T;
  wire [31:0] _reg_misa_T;
  wire _reg_misa_T_1;
  wire [3:0] _reg_misa_T_2;
  wire [31:0] _reg_misa_T_3;
  wire [31:0] _reg_misa_T_4;
  wire [31:0] _reg_misa_T_5;
  wire [31:0] _reg_misa_T_7;
  wire [31:0] _reg_misa_T_8;
  wire [3:0] _which_T_100;
  wire [3:0] _which_T_101;
  wire [3:0] _which_T_102;
  wire [3:0] _which_T_103;
  wire [3:0] _which_T_104;
  wire [3:0] _which_T_105;
  wire [3:0] _which_T_106;
  wire [3:0] _which_T_107;
  wire [3:0] _which_T_108;
  wire [3:0] _which_T_109;
  wire [3:0] _which_T_111;
  wire [3:0] _which_T_112;
  wire [3:0] _which_T_113;
  wire [3:0] _which_T_114;
  wire [3:0] _which_T_115;
  wire [3:0] _which_T_116;
  wire [3:0] _which_T_117;
  wire [3:0] _which_T_118;
  wire [3:0] _which_T_119;
  wire [3:0] _which_T_120;
  wire [3:0] _which_T_121;
  wire [3:0] _which_T_122;
  wire [3:0] _which_T_123;
  wire [3:0] _which_T_124;
  wire [3:0] _which_T_95;
  wire [3:0] _which_T_96;
  wire [3:0] _which_T_97;
  wire [3:0] _which_T_98;
  wire [3:0] _which_T_99;
  wire [12:0] addr;
  wire [11:0] addr_1;
  input clock;
  wire clock;
  wire [14:0] d_interrupts;
  wire [11:0] debugTVec;
  wire decoded_130;
  wire decoded_132;
  wire decoded_andMatrixInput_0_1;
  wire decoded_andMatrixInput_0_10;
  wire decoded_andMatrixInput_0_11;
  wire decoded_andMatrixInput_0_2;
  wire decoded_andMatrixInput_0_4;
  wire decoded_andMatrixInput_0_5;
  wire decoded_andMatrixInput_0_7;
  wire decoded_andMatrixInput_0_8;
  wire decoded_andMatrixInput_7_2;
  wire decoded_andMatrixInput_7_6;
  wire decoded_decoded_andMatrixInput_0_1;
  wire decoded_decoded_andMatrixInput_0_5;
  wire decoded_decoded_andMatrixInput_10_58;
  wire decoded_decoded_andMatrixInput_10_65;
  wire decoded_decoded_andMatrixInput_2_2;
  wire decoded_decoded_andMatrixInput_3_10;
  wire decoded_decoded_andMatrixInput_4_18;
  wire decoded_decoded_andMatrixInput_4_4;
  wire decoded_decoded_andMatrixInput_6_34;
  wire decoded_decoded_andMatrixInput_7_39;
  wire decoded_decoded_andMatrixInput_8;
  wire decoded_decoded_andMatrixInput_9;
  wire [132:0] decoded_decoded_invMatrixOutputs;
  wire [32:0] decoded_decoded_invMatrixOutputs_lo_lo;
  wire [7:0] decoded_decoded_invMatrixOutputs_lo_lo_lo_lo;
  wire [5:0] decoded_decoded_lo;
  wire [4:0] decoded_decoded_lo_129;
  wire [5:0] decoded_decoded_lo_130;
  wire [5:0] decoded_decoded_lo_34;
  wire [5:0] decoded_decoded_lo_39;
  wire [4:0] decoded_decoded_lo_4;
  wire [5:0] decoded_decoded_lo_59;
  wire [4:0] decoded_decoded_lo_65;
  wire [4:0] decoded_decoded_lo_67;
  wire [5:0] decoded_decoded_lo_68;
  wire [4:0] decoded_decoded_lo_98;
  wire [5:0] decoded_decoded_lo_99;
  wire [132:0] decoded_decoded_orMatrixOutputs;
  wire [32:0] decoded_decoded_orMatrixOutputs_lo_lo;
  wire [7:0] decoded_decoded_orMatrixOutputs_lo_lo_lo_lo;
  wire [11:0] decoded_decoded_plaInput;
  wire [31:0] decoded_invInputs;
  wire [8:0] decoded_invMatrixOutputs;
  wire [8:0] decoded_invMatrixOutputs_1;
  wire [8:0] decoded_orMatrixOutputs;
  wire [8:0] decoded_orMatrixOutputs_1;
  wire [31:0] decoded_plaInput;
  wire [31:0] epc;
  wire exception;
  wire f;
  output [31:0] io_bp_0_address;
  wire [31:0] io_bp_0_address;
  output io_bp_0_control_action;
  wire io_bp_0_control_action;
  output io_bp_0_control_r;
  wire io_bp_0_control_r;
  output [1:0] io_bp_0_control_tmatch;
  wire [1:0] io_bp_0_control_tmatch;
  output io_bp_0_control_w;
  wire io_bp_0_control_w;
  output io_bp_0_control_x;
  wire io_bp_0_control_x;
  input [31:0] io_cause;
  wire [31:0] io_cause;
  output io_csr_stall;
  wire io_csr_stall;
  output [31:0] io_customCSRs_0_value;
  wire [31:0] io_customCSRs_0_value;
  output io_decode_0_fp_csr;
  wire io_decode_0_fp_csr;
  output io_decode_0_fp_illegal;
  wire io_decode_0_fp_illegal;
  input [31:0] io_decode_0_inst;
  wire [31:0] io_decode_0_inst;
  output io_decode_0_read_illegal;
  wire io_decode_0_read_illegal;
  wire io_decode_0_read_illegal_andMatrixInput_0;
  wire io_decode_0_read_illegal_andMatrixInput_1;
  wire io_decode_0_read_illegal_andMatrixInput_3;
  wire io_decode_0_read_illegal_andMatrixInput_4;
  wire io_decode_0_read_illegal_andMatrixInput_5;
  wire io_decode_0_read_illegal_andMatrixInput_6;
  output io_decode_0_rocc_illegal;
  wire io_decode_0_rocc_illegal;
  output io_decode_0_system_illegal;
  wire io_decode_0_system_illegal;
  output io_decode_0_write_flush;
  wire io_decode_0_write_flush;
  wire [11:0] io_decode_0_write_flush_addr_m;
  output io_decode_0_write_illegal;
  wire io_decode_0_write_illegal;
  output io_eret;
  wire io_eret;
  output [31:0] io_evec;
  wire [31:0] io_evec;
  input io_exception;
  wire io_exception;
  input io_gva;
  wire io_gva;
  input io_hartid;
  wire io_hartid;
  output io_inhibit_cycle;
  wire io_inhibit_cycle;
  input [31:0] io_inst_0;
  wire [31:0] io_inst_0;
  output io_interrupt;
  wire io_interrupt;
  output [31:0] io_interrupt_cause;
  wire [31:0] io_interrupt_cause;
  input io_interrupts_debug;
  wire io_interrupts_debug;
  input io_interrupts_meip;
  wire io_interrupts_meip;
  input io_interrupts_msip;
  wire io_interrupts_msip;
  input io_interrupts_mtip;
  wire io_interrupts_mtip;
  input [31:0] io_pc;
  wire [31:0] io_pc;
  output [29:0] io_pmp_0_addr;
  wire [29:0] io_pmp_0_addr;
  output [1:0] io_pmp_0_cfg_a;
  wire [1:0] io_pmp_0_cfg_a;
  output io_pmp_0_cfg_l;
  wire io_pmp_0_cfg_l;
  output io_pmp_0_cfg_r;
  wire io_pmp_0_cfg_r;
  output io_pmp_0_cfg_w;
  wire io_pmp_0_cfg_w;
  output io_pmp_0_cfg_x;
  wire io_pmp_0_cfg_x;
  output [31:0] io_pmp_0_mask;
  wire [31:0] io_pmp_0_mask;
  output [29:0] io_pmp_1_addr;
  wire [29:0] io_pmp_1_addr;
  output [1:0] io_pmp_1_cfg_a;
  wire [1:0] io_pmp_1_cfg_a;
  output io_pmp_1_cfg_l;
  wire io_pmp_1_cfg_l;
  output io_pmp_1_cfg_r;
  wire io_pmp_1_cfg_r;
  output io_pmp_1_cfg_w;
  wire io_pmp_1_cfg_w;
  output io_pmp_1_cfg_x;
  wire io_pmp_1_cfg_x;
  output [31:0] io_pmp_1_mask;
  wire [31:0] io_pmp_1_mask;
  output [29:0] io_pmp_2_addr;
  wire [29:0] io_pmp_2_addr;
  output [1:0] io_pmp_2_cfg_a;
  wire [1:0] io_pmp_2_cfg_a;
  output io_pmp_2_cfg_l;
  wire io_pmp_2_cfg_l;
  output io_pmp_2_cfg_r;
  wire io_pmp_2_cfg_r;
  output io_pmp_2_cfg_w;
  wire io_pmp_2_cfg_w;
  output io_pmp_2_cfg_x;
  wire io_pmp_2_cfg_x;
  output [31:0] io_pmp_2_mask;
  wire [31:0] io_pmp_2_mask;
  output [29:0] io_pmp_3_addr;
  wire [29:0] io_pmp_3_addr;
  output [1:0] io_pmp_3_cfg_a;
  wire [1:0] io_pmp_3_cfg_a;
  output io_pmp_3_cfg_l;
  wire io_pmp_3_cfg_l;
  output io_pmp_3_cfg_r;
  wire io_pmp_3_cfg_r;
  output io_pmp_3_cfg_w;
  wire io_pmp_3_cfg_w;
  output io_pmp_3_cfg_x;
  wire io_pmp_3_cfg_x;
  output [31:0] io_pmp_3_mask;
  wire [31:0] io_pmp_3_mask;
  output [29:0] io_pmp_4_addr;
  wire [29:0] io_pmp_4_addr;
  output [1:0] io_pmp_4_cfg_a;
  wire [1:0] io_pmp_4_cfg_a;
  output io_pmp_4_cfg_l;
  wire io_pmp_4_cfg_l;
  output io_pmp_4_cfg_r;
  wire io_pmp_4_cfg_r;
  output io_pmp_4_cfg_w;
  wire io_pmp_4_cfg_w;
  output io_pmp_4_cfg_x;
  wire io_pmp_4_cfg_x;
  output [31:0] io_pmp_4_mask;
  wire [31:0] io_pmp_4_mask;
  output [29:0] io_pmp_5_addr;
  wire [29:0] io_pmp_5_addr;
  output [1:0] io_pmp_5_cfg_a;
  wire [1:0] io_pmp_5_cfg_a;
  output io_pmp_5_cfg_l;
  wire io_pmp_5_cfg_l;
  output io_pmp_5_cfg_r;
  wire io_pmp_5_cfg_r;
  output io_pmp_5_cfg_w;
  wire io_pmp_5_cfg_w;
  output io_pmp_5_cfg_x;
  wire io_pmp_5_cfg_x;
  output [31:0] io_pmp_5_mask;
  wire [31:0] io_pmp_5_mask;
  output [29:0] io_pmp_6_addr;
  wire [29:0] io_pmp_6_addr;
  output [1:0] io_pmp_6_cfg_a;
  wire [1:0] io_pmp_6_cfg_a;
  output io_pmp_6_cfg_l;
  wire io_pmp_6_cfg_l;
  output io_pmp_6_cfg_r;
  wire io_pmp_6_cfg_r;
  output io_pmp_6_cfg_w;
  wire io_pmp_6_cfg_w;
  output io_pmp_6_cfg_x;
  wire io_pmp_6_cfg_x;
  output [31:0] io_pmp_6_mask;
  wire [31:0] io_pmp_6_mask;
  output [29:0] io_pmp_7_addr;
  wire [29:0] io_pmp_7_addr;
  output [1:0] io_pmp_7_cfg_a;
  wire [1:0] io_pmp_7_cfg_a;
  output io_pmp_7_cfg_l;
  wire io_pmp_7_cfg_l;
  output io_pmp_7_cfg_r;
  wire io_pmp_7_cfg_r;
  output io_pmp_7_cfg_w;
  wire io_pmp_7_cfg_w;
  output io_pmp_7_cfg_x;
  wire io_pmp_7_cfg_x;
  output [31:0] io_pmp_7_mask;
  wire [31:0] io_pmp_7_mask;
  input io_retire;
  wire io_retire;
  input [11:0] io_rw_addr;
  wire [11:0] io_rw_addr;
  input [2:0] io_rw_cmd;
  wire [2:0] io_rw_cmd;
  output [31:0] io_rw_rdata;
  wire [31:0] io_rw_rdata;
  input [31:0] io_rw_wdata;
  wire [31:0] io_rw_wdata;
  output io_singleStep;
  wire io_singleStep;
  output io_status_cease;
  wire io_status_cease;
  wire io_status_cease_r;
  output io_status_debug;
  wire io_status_debug;
  output [1:0] io_status_dprv;
  wire [1:0] io_status_dprv;
  output io_status_dv;
  wire io_status_dv;
  output [1:0] io_status_fs;
  wire [1:0] io_status_fs;
  output io_status_gva;
  wire io_status_gva;
  output io_status_hie;
  wire io_status_hie;
  output [31:0] io_status_isa;
  wire [31:0] io_status_isa;
  output io_status_mbe;
  wire io_status_mbe;
  output io_status_mie;
  wire io_status_mie;
  output io_status_mpie;
  wire io_status_mpie;
  output [1:0] io_status_mpp;
  wire [1:0] io_status_mpp;
  output io_status_mprv;
  wire io_status_mprv;
  output io_status_mpv;
  wire io_status_mpv;
  output io_status_mxr;
  wire io_status_mxr;
  output [1:0] io_status_prv;
  wire [1:0] io_status_prv;
  output io_status_sbe;
  wire io_status_sbe;
  output io_status_sd;
  wire io_status_sd;
  output io_status_sd_rv32;
  wire io_status_sd_rv32;
  output io_status_sie;
  wire io_status_sie;
  output io_status_spie;
  wire io_status_spie;
  output io_status_spp;
  wire io_status_spp;
  output io_status_sum;
  wire io_status_sum;
  output [1:0] io_status_sxl;
  wire [1:0] io_status_sxl;
  output io_status_tsr;
  wire io_status_tsr;
  output io_status_tvm;
  wire io_status_tvm;
  output io_status_tw;
  wire io_status_tw;
  output io_status_ube;
  wire io_status_ube;
  output io_status_uie;
  wire io_status_uie;
  output io_status_upie;
  wire io_status_upie;
  output [1:0] io_status_uxl;
  wire [1:0] io_status_uxl;
  output io_status_v;
  wire io_status_v;
  output [1:0] io_status_vs;
  wire [1:0] io_status_vs;
  output io_status_wfi;
  wire io_status_wfi;
  output [1:0] io_status_xs;
  wire [1:0] io_status_xs;
  output [7:0] io_status_zero1;
  wire [7:0] io_status_zero1;
  output [22:0] io_status_zero2;
  wire [22:0] io_status_zero2;
  output [31:0] io_time;
  wire [31:0] io_time;
  output io_trace_0_exception;
  wire io_trace_0_exception;
  output [31:0] io_trace_0_iaddr;
  wire [31:0] io_trace_0_iaddr;
  output [31:0] io_trace_0_insn;
  wire [31:0] io_trace_0_insn;
  output io_trace_0_valid;
  wire io_trace_0_valid;
  input [31:0] io_tval;
  wire [31:0] io_tval;
  input io_ungated_clock;
  wire io_ungated_clock;
  wire [57:0] large_;
  wire [57:0] large_1;
  wire [15:0] lo_11;
  wire [15:0] lo_16;
  wire [6:0] lo_4;
  wire [31:0] m_interrupts;
  wire [1:0] newCfg_1_a;
  wire newCfg_1_l;
  wire newCfg_1_r;
  wire newCfg_1_w;
  wire newCfg_1_x;
  wire [1:0] newCfg_2_a;
  wire newCfg_2_l;
  wire newCfg_2_r;
  wire newCfg_2_w;
  wire newCfg_2_x;
  wire [1:0] newCfg_3_a;
  wire newCfg_3_l;
  wire newCfg_3_r;
  wire newCfg_3_w;
  wire newCfg_3_x;
  wire [1:0] newCfg_a;
  wire newCfg_l;
  wire newCfg_r;
  wire newCfg_w;
  wire newCfg_x;
  wire new_dcsr_ebreakm;
  wire new_mstatus_mie;
  wire new_mstatus_mpie;
  wire [31:0] notDebugTVec;
  wire [6:0] notDebugTVec_interruptOffset;
  wire [31:0] notDebugTVec_interruptVec;
  wire [31:0] pending_interrupts;
  wire [30:0] pmp_mask_base;
  wire [30:0] pmp_mask_base_1;
  wire [30:0] pmp_mask_base_2;
  wire [30:0] pmp_mask_base_3;
  wire [30:0] pmp_mask_base_4;
  wire [30:0] pmp_mask_base_5;
  wire [30:0] pmp_mask_base_6;
  wire [30:0] pmp_mask_base_7;
  wire [15:0] read_mip;
  wire [31:0] read_mstatus;
  wire [82:0] read_mstatus_hi;
  wire [64:0] read_mstatus_hi_hi;
  wire [21:0] read_mstatus_lo;
  wire [8:0] read_mstatus_lo_lo;
  wire [31:0] read_mtvec;
  wire [31:0] reg_bp_0_address;
  wire reg_bp_0_control_action;
  wire reg_bp_0_control_dmode;
  wire reg_bp_0_control_r;
  wire [1:0] reg_bp_0_control_tmatch;
  wire reg_bp_0_control_w;
  wire reg_bp_0_control_x;
  wire [31:0] reg_custom_0;
  wire [2:0] reg_dcsr_cause;
  wire reg_dcsr_ebreakm;
  wire reg_dcsr_step;
  wire reg_debug;
  wire [31:0] reg_dpc;
  wire [31:0] reg_dscratch0;
  wire [31:0] reg_mcause;
  wire [2:0] reg_mcountinhibit;
  wire [31:0] reg_mepc;
  wire [31:0] reg_mie;
  wire [31:0] reg_misa;
  wire [31:0] reg_mscratch;
  wire reg_mstatus_gva;
  wire reg_mstatus_mie;
  wire reg_mstatus_mpie;
  wire reg_mstatus_spp;
  wire [31:0] reg_mtval;
  wire [31:0] reg_mtvec;
  wire [29:0] reg_pmp_0_addr;
  wire [1:0] reg_pmp_0_cfg_a;
  wire reg_pmp_0_cfg_l;
  wire reg_pmp_0_cfg_r;
  wire reg_pmp_0_cfg_w;
  wire reg_pmp_0_cfg_x;
  wire [29:0] reg_pmp_1_addr;
  wire [1:0] reg_pmp_1_cfg_a;
  wire reg_pmp_1_cfg_l;
  wire reg_pmp_1_cfg_r;
  wire reg_pmp_1_cfg_w;
  wire reg_pmp_1_cfg_x;
  wire [29:0] reg_pmp_2_addr;
  wire [1:0] reg_pmp_2_cfg_a;
  wire reg_pmp_2_cfg_l;
  wire reg_pmp_2_cfg_r;
  wire reg_pmp_2_cfg_w;
  wire reg_pmp_2_cfg_x;
  wire [29:0] reg_pmp_3_addr;
  wire [1:0] reg_pmp_3_cfg_a;
  wire reg_pmp_3_cfg_l;
  wire reg_pmp_3_cfg_r;
  wire reg_pmp_3_cfg_w;
  wire reg_pmp_3_cfg_x;
  wire [29:0] reg_pmp_4_addr;
  wire [1:0] reg_pmp_4_cfg_a;
  wire reg_pmp_4_cfg_l;
  wire reg_pmp_4_cfg_r;
  wire reg_pmp_4_cfg_w;
  wire reg_pmp_4_cfg_x;
  wire [29:0] reg_pmp_5_addr;
  wire [1:0] reg_pmp_5_cfg_a;
  wire reg_pmp_5_cfg_l;
  wire reg_pmp_5_cfg_r;
  wire reg_pmp_5_cfg_w;
  wire reg_pmp_5_cfg_x;
  wire [29:0] reg_pmp_6_addr;
  wire [1:0] reg_pmp_6_cfg_a;
  wire reg_pmp_6_cfg_l;
  wire reg_pmp_6_cfg_r;
  wire reg_pmp_6_cfg_w;
  wire reg_pmp_6_cfg_x;
  wire [29:0] reg_pmp_7_addr;
  wire [1:0] reg_pmp_7_cfg_a;
  wire reg_pmp_7_cfg_l;
  wire reg_pmp_7_cfg_r;
  wire reg_pmp_7_cfg_w;
  wire reg_pmp_7_cfg_x;
  wire reg_singleStepped;
  wire reg_wfi;
  input reset;
  wire reset;
  wire [5:0] small_;
  wire [5:0] small_1;
  wire [31:0] tvec;
  wire [63:0] value;
  wire [63:0] value_1;
  wire [31:0] wdata;
  wire [3:0] whichInterrupt;
  wire x79;
  wire x86;
  MUX2_X1 _5102_ (
    .A(_2195_),
    .B(reg_pmp_1_addr[27]),
    .S(_3031_),
    .Z(_0392_)
  );
  MUX2_X1 _5103_ (
    .A(_2241_),
    .B(reg_pmp_1_addr[28]),
    .S(_3031_),
    .Z(_0393_)
  );
  MUX2_X1 _5104_ (
    .A(_2285_),
    .B(reg_pmp_1_addr[29]),
    .S(_3031_),
    .Z(_0394_)
  );
  AND2_X1 _5105_ (
    .A1(reg_pmp_7_cfg_l),
    .A2(reg_pmp_7_cfg_a[0]),
    .ZN(_3032_)
  );
  AND2_X1 _5106_ (
    .A1(_0004_),
    .A2(_3032_),
    .ZN(_3033_)
  );
  OR2_X1 _5107_ (
    .A1(reg_pmp_6_cfg_l),
    .A2(_3033_),
    .ZN(_3034_)
  );
  OR2_X1 _5108_ (
    .A1(_0737_),
    .A2(_3034_),
    .ZN(_3035_)
  );
  OR2_X1 _5109_ (
    .A1(_0815_),
    .A2(_3035_),
    .ZN(_3036_)
  );
  MUX2_X1 _5110_ (
    .A(_1241_),
    .B(reg_pmp_6_addr[0]),
    .S(_3036_),
    .Z(_0395_)
  );
  MUX2_X1 _5111_ (
    .A(_1290_),
    .B(reg_pmp_6_addr[1]),
    .S(_3036_),
    .Z(_0396_)
  );
  MUX2_X1 _5112_ (
    .A(_1346_),
    .B(reg_pmp_6_addr[2]),
    .S(_3036_),
    .Z(_0397_)
  );
  MUX2_X1 _5113_ (
    .A(_1409_),
    .B(reg_pmp_6_addr[3]),
    .S(_3036_),
    .Z(_0398_)
  );
  MUX2_X1 _5114_ (
    .A(_1456_),
    .B(reg_pmp_6_addr[4]),
    .S(_3036_),
    .Z(_0399_)
  );
  MUX2_X1 _5115_ (
    .A(_1499_),
    .B(reg_pmp_6_addr[5]),
    .S(_3036_),
    .Z(_0400_)
  );
  MUX2_X1 _5116_ (
    .A(_1545_),
    .B(reg_pmp_6_addr[6]),
    .S(_3036_),
    .Z(_0401_)
  );
  MUX2_X1 _5117_ (
    .A(_1601_),
    .B(reg_pmp_6_addr[7]),
    .S(_3036_),
    .Z(_0402_)
  );
  MUX2_X1 _5118_ (
    .A(_1129_),
    .B(reg_pmp_6_addr[8]),
    .S(_3036_),
    .Z(_0403_)
  );
  MUX2_X1 _5119_ (
    .A(_1175_),
    .B(reg_pmp_6_addr[9]),
    .S(_3036_),
    .Z(_0404_)
  );
  MUX2_X1 _5120_ (
    .A(_1647_),
    .B(reg_pmp_6_addr[10]),
    .S(_3036_),
    .Z(_0405_)
  );
  MUX2_X1 _5121_ (
    .A(_1698_),
    .B(reg_pmp_6_addr[11]),
    .S(_3036_),
    .Z(_0406_)
  );
  MUX2_X1 _5122_ (
    .A(_1748_),
    .B(reg_pmp_6_addr[12]),
    .S(_3036_),
    .Z(_0407_)
  );
  MUX2_X1 _5123_ (
    .A(_1790_),
    .B(reg_pmp_6_addr[13]),
    .S(_3036_),
    .Z(_0408_)
  );
  MUX2_X1 _5124_ (
    .A(_1832_),
    .B(reg_pmp_6_addr[14]),
    .S(_3036_),
    .Z(_0409_)
  );
  MUX2_X1 _5125_ (
    .A(_1880_),
    .B(reg_pmp_6_addr[15]),
    .S(_3036_),
    .Z(_0410_)
  );
  MUX2_X1 _5126_ (
    .A(_0862_),
    .B(reg_pmp_6_addr[16]),
    .S(_3036_),
    .Z(_0411_)
  );
  MUX2_X1 _5127_ (
    .A(_1926_),
    .B(reg_pmp_6_addr[17]),
    .S(_3036_),
    .Z(_0412_)
  );
  MUX2_X1 _5128_ (
    .A(_0908_),
    .B(reg_pmp_6_addr[18]),
    .S(_3036_),
    .Z(_0413_)
  );
  MUX2_X1 _5129_ (
    .A(_0967_),
    .B(reg_pmp_6_addr[19]),
    .S(_3036_),
    .Z(_0414_)
  );
  MUX2_X1 _5130_ (
    .A(_1017_),
    .B(reg_pmp_6_addr[20]),
    .S(_3036_),
    .Z(_0415_)
  );
  MUX2_X1 _5131_ (
    .A(_1968_),
    .B(reg_pmp_6_addr[21]),
    .S(_3036_),
    .Z(_0416_)
  );
  MUX2_X1 _5132_ (
    .A(_2010_),
    .B(reg_pmp_6_addr[22]),
    .S(_3036_),
    .Z(_0417_)
  );
  MUX2_X1 _5133_ (
    .A(_1071_),
    .B(reg_pmp_6_addr[23]),
    .S(_3036_),
    .Z(_0418_)
  );
  MUX2_X1 _5134_ (
    .A(_2056_),
    .B(reg_pmp_6_addr[24]),
    .S(_3036_),
    .Z(_0419_)
  );
  MUX2_X1 _5135_ (
    .A(_2102_),
    .B(reg_pmp_6_addr[25]),
    .S(_3036_),
    .Z(_0420_)
  );
  MUX2_X1 _5136_ (
    .A(_2148_),
    .B(reg_pmp_6_addr[26]),
    .S(_3036_),
    .Z(_0421_)
  );
  MUX2_X1 _5137_ (
    .A(_2195_),
    .B(reg_pmp_6_addr[27]),
    .S(_3036_),
    .Z(_0422_)
  );
  MUX2_X1 _5138_ (
    .A(_2241_),
    .B(reg_pmp_6_addr[28]),
    .S(_3036_),
    .Z(_0423_)
  );
  MUX2_X1 _5139_ (
    .A(_2285_),
    .B(reg_pmp_6_addr[29]),
    .S(_3036_),
    .Z(_0424_)
  );
  AND2_X1 _5140_ (
    .A1(_0736_),
    .A2(_1394_),
    .ZN(_3037_)
  );
  INV_X1 _5141_ (
    .A(_3037_),
    .ZN(_3038_)
  );
  AND2_X1 _5142_ (
    .A1(_1409_),
    .A2(_3037_),
    .ZN(_3039_)
  );
  AND2_X1 _5143_ (
    .A1(reg_custom_0[3]),
    .A2(_3038_),
    .ZN(_3040_)
  );
  OR2_X1 _5144_ (
    .A1(reset),
    .A2(_3040_),
    .ZN(_3041_)
  );
  OR2_X1 _5145_ (
    .A1(_3039_),
    .A2(_3041_),
    .ZN(_0425_)
  );
  AND2_X1 _5146_ (
    .A1(io_pc[1]),
    .A2(_1347_),
    .ZN(_3042_)
  );
  AND2_X1 _5147_ (
    .A1(_0736_),
    .A2(_1057_),
    .ZN(_3043_)
  );
  INV_X1 _5148_ (
    .A(_3043_),
    .ZN(_3044_)
  );
  OR2_X1 _5149_ (
    .A1(_3042_),
    .A2(_3044_),
    .ZN(_3045_)
  );
  MUX2_X1 _5150_ (
    .A(_1241_),
    .B(reg_misa[0]),
    .S(_3045_),
    .Z(_3046_)
  );
  OR2_X1 _5151_ (
    .A1(reset),
    .A2(_3046_),
    .ZN(_0426_)
  );
  MUX2_X1 _5152_ (
    .A(_1346_),
    .B(reg_misa[2]),
    .S(_3045_),
    .Z(_3047_)
  );
  OR2_X1 _5153_ (
    .A1(reset),
    .A2(_3047_),
    .ZN(_0427_)
  );
  MUX2_X1 _5154_ (
    .A(_1748_),
    .B(reg_misa[12]),
    .S(_3045_),
    .Z(_3048_)
  );
  OR2_X1 _5155_ (
    .A1(reset),
    .A2(_3048_),
    .ZN(_0428_)
  );
  AND2_X1 _5156_ (
    .A1(large_[16]),
    .A2(large_[15]),
    .ZN(_3049_)
  );
  AND2_X1 _5157_ (
    .A1(large_[17]),
    .A2(large_[14]),
    .ZN(_3050_)
  );
  AND2_X1 _5158_ (
    .A1(_3049_),
    .A2(_3050_),
    .ZN(_3051_)
  );
  AND2_X1 _5159_ (
    .A1(large_[19]),
    .A2(large_[18]),
    .ZN(_3052_)
  );
  AND2_X1 _5160_ (
    .A1(_3051_),
    .A2(_3052_),
    .ZN(_3053_)
  );
  AND2_X1 _5161_ (
    .A1(large_[11]),
    .A2(large_[10]),
    .ZN(_3054_)
  );
  AND2_X1 _5162_ (
    .A1(small_[4]),
    .A2(small_[3]),
    .ZN(_3055_)
  );
  AND2_X1 _5163_ (
    .A1(small_[5]),
    .A2(_T_14),
    .ZN(_3056_)
  );
  AND2_X1 _5164_ (
    .A1(_3055_),
    .A2(_3056_),
    .ZN(_3057_)
  );
  AND2_X1 _5165_ (
    .A1(small_[0]),
    .A2(io_retire),
    .ZN(_3058_)
  );
  AND2_X1 _5166_ (
    .A1(small_[2]),
    .A2(small_[1]),
    .ZN(_3059_)
  );
  AND2_X1 _5167_ (
    .A1(_3058_),
    .A2(_3059_),
    .ZN(_3060_)
  );
  AND2_X1 _5168_ (
    .A1(_3057_),
    .A2(_3060_),
    .ZN(_3061_)
  );
  AND2_X1 _5169_ (
    .A1(large_[1]),
    .A2(large_[0]),
    .ZN(_3062_)
  );
  AND2_X1 _5170_ (
    .A1(_3061_),
    .A2(_3062_),
    .ZN(_3063_)
  );
  INV_X1 _5171_ (
    .A(_3063_),
    .ZN(_3064_)
  );
  AND2_X1 _5172_ (
    .A1(large_[5]),
    .A2(large_[4]),
    .ZN(_3065_)
  );
  AND2_X1 _5173_ (
    .A1(large_[6]),
    .A2(large_[2]),
    .ZN(_3066_)
  );
  AND2_X1 _5174_ (
    .A1(_3065_),
    .A2(_3066_),
    .ZN(_3067_)
  );
  AND2_X1 _5175_ (
    .A1(large_[3]),
    .A2(_3067_),
    .ZN(_3068_)
  );
  AND2_X1 _5176_ (
    .A1(_3063_),
    .A2(_3068_),
    .ZN(_3069_)
  );
  AND2_X1 _5177_ (
    .A1(large_[7]),
    .A2(_3069_),
    .ZN(_3070_)
  );
  AND2_X1 _5178_ (
    .A1(large_[8]),
    .A2(_3070_),
    .ZN(_3071_)
  );
  AND2_X1 _5179_ (
    .A1(large_[9]),
    .A2(_3071_),
    .ZN(_3072_)
  );
  AND2_X1 _5180_ (
    .A1(_3054_),
    .A2(_3072_),
    .ZN(_3073_)
  );
  INV_X1 _5181_ (
    .A(_3073_),
    .ZN(_3074_)
  );
  AND2_X1 _5182_ (
    .A1(large_[12]),
    .A2(_3073_),
    .ZN(_3075_)
  );
  INV_X1 _5183_ (
    .A(_3075_),
    .ZN(_3076_)
  );
  AND2_X1 _5184_ (
    .A1(large_[13]),
    .A2(_3075_),
    .ZN(_3077_)
  );
  OR2_X1 _5185_ (
    .A1(_0625_),
    .A2(_3076_),
    .ZN(_3078_)
  );
  AND2_X1 _5186_ (
    .A1(_3053_),
    .A2(_3077_),
    .ZN(_3079_)
  );
  INV_X1 _5187_ (
    .A(_3079_),
    .ZN(_3080_)
  );
  AND2_X1 _5188_ (
    .A1(large_[20]),
    .A2(_3079_),
    .ZN(_3081_)
  );
  INV_X1 _5189_ (
    .A(_3081_),
    .ZN(_3082_)
  );
  AND2_X1 _5190_ (
    .A1(large_[21]),
    .A2(_3081_),
    .ZN(_3083_)
  );
  AND2_X1 _5191_ (
    .A1(large_[22]),
    .A2(_3083_),
    .ZN(_3084_)
  );
  INV_X1 _5192_ (
    .A(_3084_),
    .ZN(_3085_)
  );
  AND2_X1 _5193_ (
    .A1(large_[23]),
    .A2(_3084_),
    .ZN(_3086_)
  );
  INV_X1 _5194_ (
    .A(_3086_),
    .ZN(_3087_)
  );
  AND2_X1 _5195_ (
    .A1(large_[24]),
    .A2(_3086_),
    .ZN(_3088_)
  );
  INV_X1 _5196_ (
    .A(_3088_),
    .ZN(_3089_)
  );
  AND2_X1 _5197_ (
    .A1(large_[25]),
    .A2(_3088_),
    .ZN(_3090_)
  );
  INV_X1 _5198_ (
    .A(_3090_),
    .ZN(_3091_)
  );
  AND2_X1 _5199_ (
    .A1(large_[21]),
    .A2(large_[20]),
    .ZN(_3092_)
  );
  AND2_X1 _5200_ (
    .A1(_3079_),
    .A2(_3092_),
    .ZN(_3093_)
  );
  INV_X1 _5201_ (
    .A(_3093_),
    .ZN(_3094_)
  );
  AND2_X1 _5202_ (
    .A1(large_[23]),
    .A2(large_[22]),
    .ZN(_3095_)
  );
  AND2_X1 _5203_ (
    .A1(large_[25]),
    .A2(large_[24]),
    .ZN(_3096_)
  );
  AND2_X1 _5204_ (
    .A1(_3095_),
    .A2(_3096_),
    .ZN(_3097_)
  );
  AND2_X1 _5205_ (
    .A1(_3093_),
    .A2(_3097_),
    .ZN(_3098_)
  );
  AND2_X1 _5206_ (
    .A1(large_[3]),
    .A2(large_[2]),
    .ZN(_3099_)
  );
  AND2_X1 _5207_ (
    .A1(_3062_),
    .A2(_3099_),
    .ZN(_3100_)
  );
  AND2_X1 _5208_ (
    .A1(large_[6]),
    .A2(_3065_),
    .ZN(_3101_)
  );
  AND2_X1 _5209_ (
    .A1(_3100_),
    .A2(_3101_),
    .ZN(_3102_)
  );
  AND2_X1 _5210_ (
    .A1(_3061_),
    .A2(_3102_),
    .ZN(_3103_)
  );
  AND2_X1 _5211_ (
    .A1(large_[9]),
    .A2(large_[7]),
    .ZN(_3104_)
  );
  AND2_X1 _5212_ (
    .A1(large_[8]),
    .A2(_3104_),
    .ZN(_3105_)
  );
  AND2_X1 _5213_ (
    .A1(_3103_),
    .A2(_3105_),
    .ZN(_3106_)
  );
  AND2_X1 _5214_ (
    .A1(large_[12]),
    .A2(_3054_),
    .ZN(_3107_)
  );
  AND2_X1 _5215_ (
    .A1(_3106_),
    .A2(_3107_),
    .ZN(_3108_)
  );
  AND2_X1 _5216_ (
    .A1(large_[13]),
    .A2(_3108_),
    .ZN(_3109_)
  );
  AND2_X1 _5217_ (
    .A1(_3053_),
    .A2(_3109_),
    .ZN(_3110_)
  );
  OR2_X1 _5218_ (
    .A1(large_[26]),
    .A2(_3098_),
    .ZN(_3111_)
  );
  AND2_X1 _5219_ (
    .A1(large_[26]),
    .A2(_3090_),
    .ZN(_3112_)
  );
  INV_X1 _5220_ (
    .A(_3112_),
    .ZN(_3113_)
  );
  AND2_X1 _5221_ (
    .A1(_0736_),
    .A2(_0827_),
    .ZN(_3114_)
  );
  OR2_X1 _5222_ (
    .A1(_0737_),
    .A2(_0828_),
    .ZN(_3115_)
  );
  AND2_X1 _5223_ (
    .A1(_0736_),
    .A2(_0828_),
    .ZN(_3116_)
  );
  AND2_X1 _5224_ (
    .A1(_0858_),
    .A2(_3116_),
    .ZN(_3117_)
  );
  OR2_X1 _5225_ (
    .A1(_0737_),
    .A2(_3117_),
    .ZN(_3118_)
  );
  AND2_X1 _5226_ (
    .A1(_3113_),
    .A2(_3118_),
    .ZN(_3119_)
  );
  AND2_X1 _5227_ (
    .A1(_0736_),
    .A2(_0857_),
    .ZN(_3120_)
  );
  INV_X1 _5228_ (
    .A(_3120_),
    .ZN(_3121_)
  );
  AND2_X1 _5229_ (
    .A1(_3115_),
    .A2(_3121_),
    .ZN(_3122_)
  );
  OR2_X1 _5230_ (
    .A1(_3114_),
    .A2(_3120_),
    .ZN(_3123_)
  );
  AND2_X1 _5231_ (
    .A1(large_[26]),
    .A2(_3098_),
    .ZN(_3124_)
  );
  AND2_X1 _5232_ (
    .A1(_3111_),
    .A2(_3119_),
    .ZN(_3125_)
  );
  AND2_X1 _5233_ (
    .A1(_1241_),
    .A2(_3114_),
    .ZN(_3126_)
  );
  AND2_X1 _5234_ (
    .A1(large_[26]),
    .A2(_3120_),
    .ZN(_3127_)
  );
  OR2_X1 _5235_ (
    .A1(_3125_),
    .A2(_3126_),
    .ZN(_3128_)
  );
  OR2_X1 _5236_ (
    .A1(_3127_),
    .A2(_3128_),
    .ZN(_3129_)
  );
  AND2_X1 _5237_ (
    .A1(_0654_),
    .A2(_3129_),
    .ZN(_0429_)
  );
  XOR2_X1 _5238_ (
    .A(large_[27]),
    .B(_3124_),
    .Z(_3130_)
  );
  AND2_X1 _5239_ (
    .A1(_3122_),
    .A2(_3130_),
    .ZN(_3131_)
  );
  AND2_X1 _5240_ (
    .A1(_1290_),
    .A2(_3114_),
    .ZN(_3132_)
  );
  AND2_X1 _5241_ (
    .A1(large_[27]),
    .A2(_3120_),
    .ZN(_3133_)
  );
  OR2_X1 _5242_ (
    .A1(_3131_),
    .A2(_3133_),
    .ZN(_3134_)
  );
  OR2_X1 _5243_ (
    .A1(_3132_),
    .A2(_3134_),
    .ZN(_3135_)
  );
  AND2_X1 _5244_ (
    .A1(_0654_),
    .A2(_3135_),
    .ZN(_0430_)
  );
  AND2_X1 _5245_ (
    .A1(large_[27]),
    .A2(large_[26]),
    .ZN(_3136_)
  );
  AND2_X1 _5246_ (
    .A1(_3092_),
    .A2(_3136_),
    .ZN(_3137_)
  );
  AND2_X1 _5247_ (
    .A1(_3097_),
    .A2(_3137_),
    .ZN(_3138_)
  );
  AND2_X1 _5248_ (
    .A1(_3110_),
    .A2(_3138_),
    .ZN(_3139_)
  );
  INV_X1 _5249_ (
    .A(_3139_),
    .ZN(_3140_)
  );
  AND2_X1 _5250_ (
    .A1(large_[28]),
    .A2(_3139_),
    .ZN(_3141_)
  );
  OR2_X1 _5251_ (
    .A1(_0635_),
    .A2(_3140_),
    .ZN(_3142_)
  );
  OR2_X1 _5252_ (
    .A1(large_[28]),
    .A2(_3139_),
    .ZN(_3143_)
  );
  AND2_X1 _5253_ (
    .A1(_3122_),
    .A2(_3143_),
    .ZN(_3144_)
  );
  AND2_X1 _5254_ (
    .A1(_3142_),
    .A2(_3144_),
    .ZN(_3145_)
  );
  AND2_X1 _5255_ (
    .A1(_1346_),
    .A2(_3114_),
    .ZN(_3146_)
  );
  AND2_X1 _5256_ (
    .A1(large_[28]),
    .A2(_3120_),
    .ZN(_3147_)
  );
  OR2_X1 _5257_ (
    .A1(_3145_),
    .A2(_3146_),
    .ZN(_3148_)
  );
  OR2_X1 _5258_ (
    .A1(_3147_),
    .A2(_3148_),
    .ZN(_3149_)
  );
  AND2_X1 _5259_ (
    .A1(_0654_),
    .A2(_3149_),
    .ZN(_0431_)
  );
  AND2_X1 _5260_ (
    .A1(large_[29]),
    .A2(_3141_),
    .ZN(_3150_)
  );
  INV_X1 _5261_ (
    .A(_3150_),
    .ZN(_3151_)
  );
  OR2_X1 _5262_ (
    .A1(large_[29]),
    .A2(_3141_),
    .ZN(_3152_)
  );
  AND2_X1 _5263_ (
    .A1(_3118_),
    .A2(_3152_),
    .ZN(_3153_)
  );
  AND2_X1 _5264_ (
    .A1(large_[29]),
    .A2(large_[28]),
    .ZN(_3154_)
  );
  AND2_X1 _5265_ (
    .A1(_3139_),
    .A2(_3154_),
    .ZN(_3155_)
  );
  AND2_X1 _5266_ (
    .A1(_3151_),
    .A2(_3153_),
    .ZN(_3156_)
  );
  AND2_X1 _5267_ (
    .A1(_1409_),
    .A2(_3114_),
    .ZN(_3157_)
  );
  AND2_X1 _5268_ (
    .A1(large_[29]),
    .A2(_3120_),
    .ZN(_3158_)
  );
  OR2_X1 _5269_ (
    .A1(_3156_),
    .A2(_3158_),
    .ZN(_3159_)
  );
  OR2_X1 _5270_ (
    .A1(_3157_),
    .A2(_3159_),
    .ZN(_3160_)
  );
  AND2_X1 _5271_ (
    .A1(_0654_),
    .A2(_3160_),
    .ZN(_0432_)
  );
  AND2_X1 _5272_ (
    .A1(large_[30]),
    .A2(_3155_),
    .ZN(_3161_)
  );
  XOR2_X1 _5273_ (
    .A(large_[30]),
    .B(_3150_),
    .Z(_3162_)
  );
  AND2_X1 _5274_ (
    .A1(_3122_),
    .A2(_3162_),
    .ZN(_3163_)
  );
  AND2_X1 _5275_ (
    .A1(_1456_),
    .A2(_3114_),
    .ZN(_3164_)
  );
  AND2_X1 _5276_ (
    .A1(large_[30]),
    .A2(_3120_),
    .ZN(_3165_)
  );
  OR2_X1 _5277_ (
    .A1(_3163_),
    .A2(_3164_),
    .ZN(_3166_)
  );
  OR2_X1 _5278_ (
    .A1(_3165_),
    .A2(_3166_),
    .ZN(_3167_)
  );
  AND2_X1 _5279_ (
    .A1(_0654_),
    .A2(_3167_),
    .ZN(_0433_)
  );
  OR2_X1 _5280_ (
    .A1(large_[31]),
    .A2(_3161_),
    .ZN(_3168_)
  );
  AND2_X1 _5281_ (
    .A1(large_[31]),
    .A2(_3161_),
    .ZN(_3169_)
  );
  INV_X1 _5282_ (
    .A(_3169_),
    .ZN(_3170_)
  );
  AND2_X1 _5283_ (
    .A1(_3122_),
    .A2(_3170_),
    .ZN(_3171_)
  );
  AND2_X1 _5284_ (
    .A1(_3168_),
    .A2(_3171_),
    .ZN(_3172_)
  );
  AND2_X1 _5285_ (
    .A1(_1499_),
    .A2(_3114_),
    .ZN(_3173_)
  );
  AND2_X1 _5286_ (
    .A1(large_[31]),
    .A2(_3120_),
    .ZN(_3174_)
  );
  OR2_X1 _5287_ (
    .A1(_3172_),
    .A2(_3174_),
    .ZN(_3175_)
  );
  OR2_X1 _5288_ (
    .A1(_3173_),
    .A2(_3175_),
    .ZN(_3176_)
  );
  AND2_X1 _5289_ (
    .A1(_0654_),
    .A2(_3176_),
    .ZN(_0434_)
  );
  AND2_X1 _5290_ (
    .A1(large_[31]),
    .A2(_3154_),
    .ZN(_3177_)
  );
  AND2_X1 _5291_ (
    .A1(large_[30]),
    .A2(_3177_),
    .ZN(_3178_)
  );
  AND2_X1 _5292_ (
    .A1(_3139_),
    .A2(_3178_),
    .ZN(_3179_)
  );
  AND2_X1 _5293_ (
    .A1(large_[32]),
    .A2(_3169_),
    .ZN(_3180_)
  );
  AND2_X1 _5294_ (
    .A1(large_[32]),
    .A2(_3179_),
    .ZN(_3181_)
  );
  XOR2_X1 _5295_ (
    .A(large_[32]),
    .B(_3179_),
    .Z(_3182_)
  );
  AND2_X1 _5296_ (
    .A1(_3122_),
    .A2(_3182_),
    .ZN(_3183_)
  );
  AND2_X1 _5297_ (
    .A1(_1545_),
    .A2(_3114_),
    .ZN(_3184_)
  );
  AND2_X1 _5298_ (
    .A1(large_[32]),
    .A2(_3120_),
    .ZN(_3185_)
  );
  OR2_X1 _5299_ (
    .A1(_3183_),
    .A2(_3184_),
    .ZN(_3186_)
  );
  OR2_X1 _5300_ (
    .A1(_3185_),
    .A2(_3186_),
    .ZN(_3187_)
  );
  AND2_X1 _5301_ (
    .A1(_0654_),
    .A2(_3187_),
    .ZN(_0435_)
  );
  OR2_X1 _5302_ (
    .A1(large_[33]),
    .A2(_3181_),
    .ZN(_3188_)
  );
  AND2_X1 _5303_ (
    .A1(large_[33]),
    .A2(_3180_),
    .ZN(_3189_)
  );
  INV_X1 _5304_ (
    .A(_3189_),
    .ZN(_3190_)
  );
  AND2_X1 _5305_ (
    .A1(_3122_),
    .A2(_3188_),
    .ZN(_3191_)
  );
  AND2_X1 _5306_ (
    .A1(_3190_),
    .A2(_3191_),
    .ZN(_3192_)
  );
  AND2_X1 _5307_ (
    .A1(_1601_),
    .A2(_3114_),
    .ZN(_3193_)
  );
  AND2_X1 _5308_ (
    .A1(large_[33]),
    .A2(_3120_),
    .ZN(_3194_)
  );
  OR2_X1 _5309_ (
    .A1(_3192_),
    .A2(_3194_),
    .ZN(_3195_)
  );
  OR2_X1 _5310_ (
    .A1(_3193_),
    .A2(_3195_),
    .ZN(_3196_)
  );
  AND2_X1 _5311_ (
    .A1(_0654_),
    .A2(_3196_),
    .ZN(_0436_)
  );
  OR2_X1 _5312_ (
    .A1(large_[34]),
    .A2(_3189_),
    .ZN(_3197_)
  );
  AND2_X1 _5313_ (
    .A1(large_[34]),
    .A2(_3189_),
    .ZN(_3198_)
  );
  INV_X1 _5314_ (
    .A(_3198_),
    .ZN(_3199_)
  );
  AND2_X1 _5315_ (
    .A1(_3122_),
    .A2(_3199_),
    .ZN(_3200_)
  );
  AND2_X1 _5316_ (
    .A1(large_[34]),
    .A2(large_[33]),
    .ZN(_3201_)
  );
  AND2_X1 _5317_ (
    .A1(_3197_),
    .A2(_3200_),
    .ZN(_3202_)
  );
  AND2_X1 _5318_ (
    .A1(_1129_),
    .A2(_3114_),
    .ZN(_3203_)
  );
  AND2_X1 _5319_ (
    .A1(large_[34]),
    .A2(_3120_),
    .ZN(_3204_)
  );
  OR2_X1 _5320_ (
    .A1(_3202_),
    .A2(_3204_),
    .ZN(_3205_)
  );
  OR2_X1 _5321_ (
    .A1(_3203_),
    .A2(_3205_),
    .ZN(_3206_)
  );
  AND2_X1 _5322_ (
    .A1(_0654_),
    .A2(_3206_),
    .ZN(_0437_)
  );
  OR2_X1 _5323_ (
    .A1(large_[35]),
    .A2(_3198_),
    .ZN(_3207_)
  );
  AND2_X1 _5324_ (
    .A1(large_[35]),
    .A2(_3198_),
    .ZN(_3208_)
  );
  AND2_X1 _5325_ (
    .A1(large_[35]),
    .A2(_3201_),
    .ZN(_3209_)
  );
  AND2_X1 _5326_ (
    .A1(_3181_),
    .A2(_3209_),
    .ZN(_3210_)
  );
  INV_X1 _5327_ (
    .A(_3210_),
    .ZN(_3211_)
  );
  AND2_X1 _5328_ (
    .A1(_3122_),
    .A2(_3211_),
    .ZN(_3212_)
  );
  AND2_X1 _5329_ (
    .A1(_3207_),
    .A2(_3212_),
    .ZN(_3213_)
  );
  AND2_X1 _5330_ (
    .A1(_1175_),
    .A2(_3114_),
    .ZN(_3214_)
  );
  AND2_X1 _5331_ (
    .A1(large_[35]),
    .A2(_3120_),
    .ZN(_3215_)
  );
  OR2_X1 _5332_ (
    .A1(_3214_),
    .A2(_3215_),
    .ZN(_3216_)
  );
  OR2_X1 _5333_ (
    .A1(_3213_),
    .A2(_3216_),
    .ZN(_3217_)
  );
  AND2_X1 _5334_ (
    .A1(_0654_),
    .A2(_3217_),
    .ZN(_0438_)
  );
  AND2_X1 _5335_ (
    .A1(large_[36]),
    .A2(_3208_),
    .ZN(_3218_)
  );
  AND2_X1 _5336_ (
    .A1(large_[36]),
    .A2(_3210_),
    .ZN(_3219_)
  );
  XOR2_X1 _5337_ (
    .A(large_[36]),
    .B(_3210_),
    .Z(_3220_)
  );
  AND2_X1 _5338_ (
    .A1(_3122_),
    .A2(_3220_),
    .ZN(_3221_)
  );
  AND2_X1 _5339_ (
    .A1(_1647_),
    .A2(_3114_),
    .ZN(_3222_)
  );
  AND2_X1 _5340_ (
    .A1(large_[36]),
    .A2(_3120_),
    .ZN(_3223_)
  );
  OR2_X1 _5341_ (
    .A1(_3221_),
    .A2(_3222_),
    .ZN(_3224_)
  );
  OR2_X1 _5342_ (
    .A1(_3223_),
    .A2(_3224_),
    .ZN(_3225_)
  );
  AND2_X1 _5343_ (
    .A1(_0654_),
    .A2(_3225_),
    .ZN(_0439_)
  );
  AND2_X1 _5344_ (
    .A1(large_[37]),
    .A2(large_[36]),
    .ZN(_3226_)
  );
  AND2_X1 _5345_ (
    .A1(large_[37]),
    .A2(_3218_),
    .ZN(_3227_)
  );
  XOR2_X1 _5346_ (
    .A(large_[37]),
    .B(_3219_),
    .Z(_3228_)
  );
  AND2_X1 _5347_ (
    .A1(_3122_),
    .A2(_3228_),
    .ZN(_3229_)
  );
  AND2_X1 _5348_ (
    .A1(_1698_),
    .A2(_3114_),
    .ZN(_3230_)
  );
  AND2_X1 _5349_ (
    .A1(large_[37]),
    .A2(_3120_),
    .ZN(_3231_)
  );
  OR2_X1 _5350_ (
    .A1(_3229_),
    .A2(_3230_),
    .ZN(_3232_)
  );
  OR2_X1 _5351_ (
    .A1(_3231_),
    .A2(_3232_),
    .ZN(_3233_)
  );
  AND2_X1 _5352_ (
    .A1(_0654_),
    .A2(_3233_),
    .ZN(_0440_)
  );
  OR2_X1 _5353_ (
    .A1(large_[38]),
    .A2(_3227_),
    .ZN(_3234_)
  );
  AND2_X1 _5354_ (
    .A1(large_[38]),
    .A2(_3227_),
    .ZN(_3235_)
  );
  INV_X1 _5355_ (
    .A(_3235_),
    .ZN(_3236_)
  );
  AND2_X1 _5356_ (
    .A1(_3122_),
    .A2(_3236_),
    .ZN(_3237_)
  );
  AND2_X1 _5357_ (
    .A1(large_[38]),
    .A2(_3226_),
    .ZN(_3238_)
  );
  AND2_X1 _5358_ (
    .A1(_3234_),
    .A2(_3237_),
    .ZN(_3239_)
  );
  AND2_X1 _5359_ (
    .A1(_1748_),
    .A2(_3114_),
    .ZN(_3240_)
  );
  AND2_X1 _5360_ (
    .A1(large_[38]),
    .A2(_3120_),
    .ZN(_3241_)
  );
  OR2_X1 _5361_ (
    .A1(_3239_),
    .A2(_3240_),
    .ZN(_3242_)
  );
  OR2_X1 _5362_ (
    .A1(_3241_),
    .A2(_3242_),
    .ZN(_3243_)
  );
  AND2_X1 _5363_ (
    .A1(_0654_),
    .A2(_3243_),
    .ZN(_0441_)
  );
  OR2_X1 _5364_ (
    .A1(large_[39]),
    .A2(_3235_),
    .ZN(_3244_)
  );
  AND2_X1 _5365_ (
    .A1(_3122_),
    .A2(_3244_),
    .ZN(_3245_)
  );
  AND2_X1 _5366_ (
    .A1(large_[39]),
    .A2(_3235_),
    .ZN(_3246_)
  );
  INV_X1 _5367_ (
    .A(_3246_),
    .ZN(_3247_)
  );
  AND2_X1 _5368_ (
    .A1(_3245_),
    .A2(_3247_),
    .ZN(_3248_)
  );
  AND2_X1 _5369_ (
    .A1(_1790_),
    .A2(_3114_),
    .ZN(_3249_)
  );
  AND2_X1 _5370_ (
    .A1(large_[39]),
    .A2(_3120_),
    .ZN(_3250_)
  );
  OR2_X1 _5371_ (
    .A1(_3248_),
    .A2(_3249_),
    .ZN(_3251_)
  );
  OR2_X1 _5372_ (
    .A1(_3250_),
    .A2(_3251_),
    .ZN(_3252_)
  );
  AND2_X1 _5373_ (
    .A1(_0654_),
    .A2(_3252_),
    .ZN(_0442_)
  );
  AND2_X1 _5374_ (
    .A1(large_[39]),
    .A2(large_[32]),
    .ZN(_3253_)
  );
  AND2_X1 _5375_ (
    .A1(large_[30]),
    .A2(_3253_),
    .ZN(_3254_)
  );
  AND2_X1 _5376_ (
    .A1(_3177_),
    .A2(_3254_),
    .ZN(_3255_)
  );
  AND2_X1 _5377_ (
    .A1(_3209_),
    .A2(_3238_),
    .ZN(_3256_)
  );
  AND2_X1 _5378_ (
    .A1(_3255_),
    .A2(_3256_),
    .ZN(_3257_)
  );
  AND2_X1 _5379_ (
    .A1(_3138_),
    .A2(_3257_),
    .ZN(_3258_)
  );
  AND2_X1 _5380_ (
    .A1(_3079_),
    .A2(_3258_),
    .ZN(_3259_)
  );
  AND2_X1 _5381_ (
    .A1(_3209_),
    .A2(_3253_),
    .ZN(_3260_)
  );
  AND2_X1 _5382_ (
    .A1(_3178_),
    .A2(_3260_),
    .ZN(_3261_)
  );
  AND2_X1 _5383_ (
    .A1(_3138_),
    .A2(_3238_),
    .ZN(_3262_)
  );
  AND2_X1 _5384_ (
    .A1(_3261_),
    .A2(_3262_),
    .ZN(_3263_)
  );
  AND2_X1 _5385_ (
    .A1(_3110_),
    .A2(_3263_),
    .ZN(_3264_)
  );
  AND2_X1 _5386_ (
    .A1(large_[40]),
    .A2(_3264_),
    .ZN(_3265_)
  );
  XOR2_X1 _5387_ (
    .A(large_[40]),
    .B(_3264_),
    .Z(_3266_)
  );
  AND2_X1 _5388_ (
    .A1(_3122_),
    .A2(_3266_),
    .ZN(_3267_)
  );
  AND2_X1 _5389_ (
    .A1(_1832_),
    .A2(_3114_),
    .ZN(_3268_)
  );
  AND2_X1 _5390_ (
    .A1(large_[40]),
    .A2(_3120_),
    .ZN(_3269_)
  );
  OR2_X1 _5391_ (
    .A1(_3267_),
    .A2(_3268_),
    .ZN(_3270_)
  );
  OR2_X1 _5392_ (
    .A1(_3269_),
    .A2(_3270_),
    .ZN(_3271_)
  );
  AND2_X1 _5393_ (
    .A1(_0654_),
    .A2(_3271_),
    .ZN(_0443_)
  );
  AND2_X1 _5394_ (
    .A1(large_[41]),
    .A2(large_[40]),
    .ZN(_3272_)
  );
  AND2_X1 _5395_ (
    .A1(large_[41]),
    .A2(_3265_),
    .ZN(_3273_)
  );
  XOR2_X1 _5396_ (
    .A(large_[41]),
    .B(_3265_),
    .Z(_3274_)
  );
  AND2_X1 _5397_ (
    .A1(_3122_),
    .A2(_3274_),
    .ZN(_3275_)
  );
  AND2_X1 _5398_ (
    .A1(_1880_),
    .A2(_3114_),
    .ZN(_3276_)
  );
  AND2_X1 _5399_ (
    .A1(large_[41]),
    .A2(_3120_),
    .ZN(_3277_)
  );
  OR2_X1 _5400_ (
    .A1(_3276_),
    .A2(_3277_),
    .ZN(_3278_)
  );
  OR2_X1 _5401_ (
    .A1(_3275_),
    .A2(_3278_),
    .ZN(_3279_)
  );
  AND2_X1 _5402_ (
    .A1(_0654_),
    .A2(_3279_),
    .ZN(_0444_)
  );
  AND2_X1 _5403_ (
    .A1(large_[42]),
    .A2(_3273_),
    .ZN(_3280_)
  );
  XOR2_X1 _5404_ (
    .A(large_[42]),
    .B(_3273_),
    .Z(_3281_)
  );
  AND2_X1 _5405_ (
    .A1(_3122_),
    .A2(_3281_),
    .ZN(_3282_)
  );
  AND2_X1 _5406_ (
    .A1(_0862_),
    .A2(_3114_),
    .ZN(_3283_)
  );
  AND2_X1 _5407_ (
    .A1(large_[42]),
    .A2(_3120_),
    .ZN(_3284_)
  );
  OR2_X1 _5408_ (
    .A1(_3282_),
    .A2(_3283_),
    .ZN(_3285_)
  );
  OR2_X1 _5409_ (
    .A1(_3284_),
    .A2(_3285_),
    .ZN(_3286_)
  );
  AND2_X1 _5410_ (
    .A1(_0654_),
    .A2(_3286_),
    .ZN(_0445_)
  );
  OR2_X1 _5411_ (
    .A1(large_[43]),
    .A2(_3280_),
    .ZN(_3287_)
  );
  AND2_X1 _5412_ (
    .A1(large_[43]),
    .A2(large_[42]),
    .ZN(_3288_)
  );
  AND2_X1 _5413_ (
    .A1(_3272_),
    .A2(_3288_),
    .ZN(_3289_)
  );
  AND2_X1 _5414_ (
    .A1(_3259_),
    .A2(_3289_),
    .ZN(_3290_)
  );
  AND2_X1 _5415_ (
    .A1(large_[43]),
    .A2(_3280_),
    .ZN(_3291_)
  );
  INV_X1 _5416_ (
    .A(_3291_),
    .ZN(_3292_)
  );
  AND2_X1 _5417_ (
    .A1(_3122_),
    .A2(_3292_),
    .ZN(_3293_)
  );
  AND2_X1 _5418_ (
    .A1(_3287_),
    .A2(_3293_),
    .ZN(_3294_)
  );
  AND2_X1 _5419_ (
    .A1(_1926_),
    .A2(_3114_),
    .ZN(_3295_)
  );
  AND2_X1 _5420_ (
    .A1(large_[43]),
    .A2(_3120_),
    .ZN(_3296_)
  );
  OR2_X1 _5421_ (
    .A1(_3295_),
    .A2(_3296_),
    .ZN(_3297_)
  );
  OR2_X1 _5422_ (
    .A1(_3294_),
    .A2(_3297_),
    .ZN(_3298_)
  );
  AND2_X1 _5423_ (
    .A1(_0654_),
    .A2(_3298_),
    .ZN(_0446_)
  );
  AND2_X1 _5424_ (
    .A1(_3264_),
    .A2(_3289_),
    .ZN(_3299_)
  );
  AND2_X1 _5425_ (
    .A1(large_[44]),
    .A2(_3290_),
    .ZN(_3300_)
  );
  INV_X1 _5426_ (
    .A(_3300_),
    .ZN(_3301_)
  );
  AND2_X1 _5427_ (
    .A1(large_[44]),
    .A2(_3299_),
    .ZN(_3302_)
  );
  XOR2_X1 _5428_ (
    .A(large_[44]),
    .B(_3299_),
    .Z(_3303_)
  );
  AND2_X1 _5429_ (
    .A1(_3122_),
    .A2(_3303_),
    .ZN(_3304_)
  );
  AND2_X1 _5430_ (
    .A1(_0908_),
    .A2(_3114_),
    .ZN(_3305_)
  );
  AND2_X1 _5431_ (
    .A1(large_[44]),
    .A2(_3120_),
    .ZN(_3306_)
  );
  OR2_X1 _5432_ (
    .A1(_3304_),
    .A2(_3305_),
    .ZN(_3307_)
  );
  OR2_X1 _5433_ (
    .A1(_3306_),
    .A2(_3307_),
    .ZN(_3308_)
  );
  AND2_X1 _5434_ (
    .A1(_0654_),
    .A2(_3308_),
    .ZN(_0447_)
  );
  OR2_X1 _5435_ (
    .A1(large_[45]),
    .A2(_3302_),
    .ZN(_3309_)
  );
  AND2_X1 _5436_ (
    .A1(_3122_),
    .A2(_3309_),
    .ZN(_3310_)
  );
  AND2_X1 _5437_ (
    .A1(large_[45]),
    .A2(_3300_),
    .ZN(_3311_)
  );
  INV_X1 _5438_ (
    .A(_3311_),
    .ZN(_3312_)
  );
  AND2_X1 _5439_ (
    .A1(_3310_),
    .A2(_3312_),
    .ZN(_3313_)
  );
  AND2_X1 _5440_ (
    .A1(_0967_),
    .A2(_3114_),
    .ZN(_3314_)
  );
  AND2_X1 _5441_ (
    .A1(large_[45]),
    .A2(_3120_),
    .ZN(_3315_)
  );
  OR2_X1 _5442_ (
    .A1(_3313_),
    .A2(_3315_),
    .ZN(_3316_)
  );
  OR2_X1 _5443_ (
    .A1(_3314_),
    .A2(_3316_),
    .ZN(_3317_)
  );
  AND2_X1 _5444_ (
    .A1(_0654_),
    .A2(_3317_),
    .ZN(_0448_)
  );
  OR2_X1 _5445_ (
    .A1(large_[46]),
    .A2(_3311_),
    .ZN(_3318_)
  );
  AND2_X1 _5446_ (
    .A1(large_[46]),
    .A2(large_[45]),
    .ZN(_3319_)
  );
  INV_X1 _5447_ (
    .A(_3319_),
    .ZN(_3320_)
  );
  OR2_X1 _5448_ (
    .A1(_3301_),
    .A2(_3320_),
    .ZN(_3321_)
  );
  AND2_X1 _5449_ (
    .A1(_3122_),
    .A2(_3321_),
    .ZN(_3322_)
  );
  AND2_X1 _5450_ (
    .A1(_3302_),
    .A2(_3319_),
    .ZN(_3323_)
  );
  AND2_X1 _5451_ (
    .A1(_3318_),
    .A2(_3322_),
    .ZN(_3324_)
  );
  AND2_X1 _5452_ (
    .A1(_1017_),
    .A2(_3114_),
    .ZN(_3325_)
  );
  AND2_X1 _5453_ (
    .A1(large_[46]),
    .A2(_3120_),
    .ZN(_3326_)
  );
  OR2_X1 _5454_ (
    .A1(_3324_),
    .A2(_3326_),
    .ZN(_3327_)
  );
  OR2_X1 _5455_ (
    .A1(_3325_),
    .A2(_3327_),
    .ZN(_3328_)
  );
  AND2_X1 _5456_ (
    .A1(_0654_),
    .A2(_3328_),
    .ZN(_0449_)
  );
  OR2_X1 _5457_ (
    .A1(large_[47]),
    .A2(_3323_),
    .ZN(_3329_)
  );
  AND2_X1 _5458_ (
    .A1(_3122_),
    .A2(_3329_),
    .ZN(_3330_)
  );
  OR2_X1 _5459_ (
    .A1(_0634_),
    .A2(_3321_),
    .ZN(_3331_)
  );
  AND2_X1 _5460_ (
    .A1(large_[47]),
    .A2(_3323_),
    .ZN(_3332_)
  );
  AND2_X1 _5461_ (
    .A1(_3330_),
    .A2(_3331_),
    .ZN(_3333_)
  );
  AND2_X1 _5462_ (
    .A1(_1968_),
    .A2(_3114_),
    .ZN(_3334_)
  );
  AND2_X1 _5463_ (
    .A1(large_[47]),
    .A2(_3120_),
    .ZN(_3335_)
  );
  OR2_X1 _5464_ (
    .A1(_3333_),
    .A2(_3335_),
    .ZN(_3336_)
  );
  OR2_X1 _5465_ (
    .A1(_3334_),
    .A2(_3336_),
    .ZN(_3337_)
  );
  AND2_X1 _5466_ (
    .A1(_0654_),
    .A2(_3337_),
    .ZN(_0450_)
  );
  AND2_X1 _5467_ (
    .A1(large_[48]),
    .A2(_3332_),
    .ZN(_3338_)
  );
  XOR2_X1 _5468_ (
    .A(large_[48]),
    .B(_3332_),
    .Z(_3339_)
  );
  AND2_X1 _5469_ (
    .A1(_3122_),
    .A2(_3339_),
    .ZN(_3340_)
  );
  AND2_X1 _5470_ (
    .A1(_2010_),
    .A2(_3114_),
    .ZN(_3341_)
  );
  AND2_X1 _5471_ (
    .A1(large_[48]),
    .A2(_3120_),
    .ZN(_3342_)
  );
  OR2_X1 _5472_ (
    .A1(_3341_),
    .A2(_3342_),
    .ZN(_3343_)
  );
  OR2_X1 _5473_ (
    .A1(_3340_),
    .A2(_3343_),
    .ZN(_3344_)
  );
  AND2_X1 _5474_ (
    .A1(_0654_),
    .A2(_3344_),
    .ZN(_0451_)
  );
  AND2_X1 _5475_ (
    .A1(large_[49]),
    .A2(_3338_),
    .ZN(_3345_)
  );
  XOR2_X1 _5476_ (
    .A(large_[49]),
    .B(_3338_),
    .Z(_3346_)
  );
  AND2_X1 _5477_ (
    .A1(_3122_),
    .A2(_3346_),
    .ZN(_3347_)
  );
  AND2_X1 _5478_ (
    .A1(_1071_),
    .A2(_3114_),
    .ZN(_3348_)
  );
  AND2_X1 _5479_ (
    .A1(large_[49]),
    .A2(_3120_),
    .ZN(_3349_)
  );
  OR2_X1 _5480_ (
    .A1(_3348_),
    .A2(_3349_),
    .ZN(_3350_)
  );
  OR2_X1 _5481_ (
    .A1(_3347_),
    .A2(_3350_),
    .ZN(_3351_)
  );
  AND2_X1 _5482_ (
    .A1(_0654_),
    .A2(_3351_),
    .ZN(_0452_)
  );
  AND2_X1 _5483_ (
    .A1(large_[50]),
    .A2(_3345_),
    .ZN(_3352_)
  );
  XOR2_X1 _5484_ (
    .A(_0633_),
    .B(_3345_),
    .Z(_3353_)
  );
  OR2_X1 _5485_ (
    .A1(_3123_),
    .A2(_3353_),
    .ZN(_3354_)
  );
  INV_X1 _5486_ (
    .A(_3354_),
    .ZN(_3355_)
  );
  AND2_X1 _5487_ (
    .A1(_2056_),
    .A2(_3114_),
    .ZN(_3356_)
  );
  AND2_X1 _5488_ (
    .A1(large_[50]),
    .A2(_3120_),
    .ZN(_3357_)
  );
  OR2_X1 _5489_ (
    .A1(_3355_),
    .A2(_3356_),
    .ZN(_3358_)
  );
  OR2_X1 _5490_ (
    .A1(_3357_),
    .A2(_3358_),
    .ZN(_3359_)
  );
  AND2_X1 _5491_ (
    .A1(_0654_),
    .A2(_3359_),
    .ZN(_0453_)
  );
  OR2_X1 _5492_ (
    .A1(large_[51]),
    .A2(_3352_),
    .ZN(_3360_)
  );
  AND2_X1 _5493_ (
    .A1(large_[51]),
    .A2(_3352_),
    .ZN(_3361_)
  );
  INV_X1 _5494_ (
    .A(_3361_),
    .ZN(_3362_)
  );
  AND2_X1 _5495_ (
    .A1(_3122_),
    .A2(_3362_),
    .ZN(_3363_)
  );
  AND2_X1 _5496_ (
    .A1(_3360_),
    .A2(_3363_),
    .ZN(_3364_)
  );
  AND2_X1 _5497_ (
    .A1(_2102_),
    .A2(_3114_),
    .ZN(_3365_)
  );
  AND2_X1 _5498_ (
    .A1(large_[51]),
    .A2(_3120_),
    .ZN(_3366_)
  );
  OR2_X1 _5499_ (
    .A1(_3364_),
    .A2(_3365_),
    .ZN(_3367_)
  );
  OR2_X1 _5500_ (
    .A1(_3366_),
    .A2(_3367_),
    .ZN(_3368_)
  );
  AND2_X1 _5501_ (
    .A1(_0654_),
    .A2(_3368_),
    .ZN(_0454_)
  );
  AND2_X1 _5502_ (
    .A1(large_[52]),
    .A2(_3361_),
    .ZN(_3369_)
  );
  XOR2_X1 _5503_ (
    .A(large_[52]),
    .B(_3361_),
    .Z(_3370_)
  );
  AND2_X1 _5504_ (
    .A1(_3122_),
    .A2(_3370_),
    .ZN(_3371_)
  );
  AND2_X1 _5505_ (
    .A1(_2148_),
    .A2(_3114_),
    .ZN(_3372_)
  );
  AND2_X1 _5506_ (
    .A1(large_[52]),
    .A2(_3120_),
    .ZN(_3373_)
  );
  OR2_X1 _5507_ (
    .A1(_3371_),
    .A2(_3372_),
    .ZN(_3374_)
  );
  OR2_X1 _5508_ (
    .A1(_3373_),
    .A2(_3374_),
    .ZN(_3375_)
  );
  AND2_X1 _5509_ (
    .A1(_0654_),
    .A2(_3375_),
    .ZN(_0455_)
  );
  AND2_X1 _5510_ (
    .A1(large_[53]),
    .A2(_3369_),
    .ZN(_3376_)
  );
  XOR2_X1 _5511_ (
    .A(large_[53]),
    .B(_3369_),
    .Z(_3377_)
  );
  AND2_X1 _5512_ (
    .A1(_3122_),
    .A2(_3377_),
    .ZN(_3378_)
  );
  AND2_X1 _5513_ (
    .A1(_2195_),
    .A2(_3114_),
    .ZN(_3379_)
  );
  AND2_X1 _5514_ (
    .A1(large_[53]),
    .A2(_3120_),
    .ZN(_3380_)
  );
  OR2_X1 _5515_ (
    .A1(_3378_),
    .A2(_3379_),
    .ZN(_3381_)
  );
  OR2_X1 _5516_ (
    .A1(_3380_),
    .A2(_3381_),
    .ZN(_3382_)
  );
  AND2_X1 _5517_ (
    .A1(_0654_),
    .A2(_3382_),
    .ZN(_0456_)
  );
  OR2_X1 _5518_ (
    .A1(large_[54]),
    .A2(_3376_),
    .ZN(_3383_)
  );
  AND2_X1 _5519_ (
    .A1(large_[54]),
    .A2(_3376_),
    .ZN(_3384_)
  );
  INV_X1 _5520_ (
    .A(_3384_),
    .ZN(_3385_)
  );
  AND2_X1 _5521_ (
    .A1(_3122_),
    .A2(_3385_),
    .ZN(_3386_)
  );
  AND2_X1 _5522_ (
    .A1(_3383_),
    .A2(_3386_),
    .ZN(_3387_)
  );
  AND2_X1 _5523_ (
    .A1(_2241_),
    .A2(_3114_),
    .ZN(_3388_)
  );
  AND2_X1 _5524_ (
    .A1(large_[54]),
    .A2(_3120_),
    .ZN(_3389_)
  );
  OR2_X1 _5525_ (
    .A1(_3387_),
    .A2(_3388_),
    .ZN(_3390_)
  );
  OR2_X1 _5526_ (
    .A1(_3389_),
    .A2(_3390_),
    .ZN(_3391_)
  );
  AND2_X1 _5527_ (
    .A1(_0654_),
    .A2(_3391_),
    .ZN(_0457_)
  );
  OR2_X1 _5528_ (
    .A1(large_[55]),
    .A2(_3384_),
    .ZN(_3392_)
  );
  AND2_X1 _5529_ (
    .A1(large_[55]),
    .A2(_3384_),
    .ZN(_3393_)
  );
  INV_X1 _5530_ (
    .A(_3393_),
    .ZN(_3394_)
  );
  AND2_X1 _5531_ (
    .A1(_3122_),
    .A2(_3394_),
    .ZN(_3395_)
  );
  AND2_X1 _5532_ (
    .A1(_3392_),
    .A2(_3395_),
    .ZN(_3396_)
  );
  AND2_X1 _5533_ (
    .A1(_2285_),
    .A2(_3114_),
    .ZN(_3397_)
  );
  AND2_X1 _5534_ (
    .A1(large_[55]),
    .A2(_3120_),
    .ZN(_3398_)
  );
  OR2_X1 _5535_ (
    .A1(_3396_),
    .A2(_3397_),
    .ZN(_3399_)
  );
  OR2_X1 _5536_ (
    .A1(_3398_),
    .A2(_3399_),
    .ZN(_3400_)
  );
  AND2_X1 _5537_ (
    .A1(_0654_),
    .A2(_3400_),
    .ZN(_0458_)
  );
  OR2_X1 _5538_ (
    .A1(large_[56]),
    .A2(_3393_),
    .ZN(_3401_)
  );
  AND2_X1 _5539_ (
    .A1(large_[56]),
    .A2(_3393_),
    .ZN(_3402_)
  );
  INV_X1 _5540_ (
    .A(_3402_),
    .ZN(_3403_)
  );
  AND2_X1 _5541_ (
    .A1(_3122_),
    .A2(_3403_),
    .ZN(_3404_)
  );
  AND2_X1 _5542_ (
    .A1(_3401_),
    .A2(_3404_),
    .ZN(_3405_)
  );
  AND2_X1 _5543_ (
    .A1(_2435_),
    .A2(_3114_),
    .ZN(_3406_)
  );
  AND2_X1 _5544_ (
    .A1(large_[56]),
    .A2(_3120_),
    .ZN(_3407_)
  );
  OR2_X1 _5545_ (
    .A1(_3405_),
    .A2(_3406_),
    .ZN(_3408_)
  );
  OR2_X1 _5546_ (
    .A1(_3407_),
    .A2(_3408_),
    .ZN(_3409_)
  );
  AND2_X1 _5547_ (
    .A1(_0654_),
    .A2(_3409_),
    .ZN(_0459_)
  );
  XOR2_X1 _5548_ (
    .A(large_[57]),
    .B(_3402_),
    .Z(_3410_)
  );
  AND2_X1 _5549_ (
    .A1(_3122_),
    .A2(_3410_),
    .ZN(_3411_)
  );
  AND2_X1 _5550_ (
    .A1(_2365_),
    .A2(_3114_),
    .ZN(_3412_)
  );
  AND2_X1 _5551_ (
    .A1(large_[57]),
    .A2(_3120_),
    .ZN(_3413_)
  );
  OR2_X1 _5552_ (
    .A1(_3412_),
    .A2(_3413_),
    .ZN(_3414_)
  );
  OR2_X1 _5553_ (
    .A1(_3411_),
    .A2(_3414_),
    .ZN(_3415_)
  );
  AND2_X1 _5554_ (
    .A1(_0654_),
    .A2(_3415_),
    .ZN(_0460_)
  );
  AND2_X1 _5555_ (
    .A1(_0652_),
    .A2(io_retire),
    .ZN(_3416_)
  );
  AND2_X1 _5556_ (
    .A1(_0652_),
    .A2(_3058_),
    .ZN(_3417_)
  );
  XOR2_X1 _5557_ (
    .A(small_[0]),
    .B(_3416_),
    .Z(_3418_)
  );
  AND2_X1 _5558_ (
    .A1(_3117_),
    .A2(_3418_),
    .ZN(_3419_)
  );
  AND2_X1 _5559_ (
    .A1(small_[0]),
    .A2(_3114_),
    .ZN(_3420_)
  );
  AND2_X1 _5560_ (
    .A1(_0737_),
    .A2(_3418_),
    .ZN(_3421_)
  );
  OR2_X1 _5561_ (
    .A1(_3420_),
    .A2(_3421_),
    .ZN(_3422_)
  );
  OR2_X1 _5562_ (
    .A1(_3419_),
    .A2(_3422_),
    .ZN(_3423_)
  );
  AND2_X1 _5563_ (
    .A1(_1241_),
    .A2(_3120_),
    .ZN(_3424_)
  );
  OR2_X1 _5564_ (
    .A1(_3423_),
    .A2(_3424_),
    .ZN(_3425_)
  );
  AND2_X1 _5565_ (
    .A1(_0654_),
    .A2(_3425_),
    .ZN(_0461_)
  );
  OR2_X1 _5566_ (
    .A1(small_[1]),
    .A2(_3417_),
    .ZN(_3426_)
  );
  AND2_X1 _5567_ (
    .A1(small_[1]),
    .A2(_3114_),
    .ZN(_3427_)
  );
  AND2_X1 _5568_ (
    .A1(small_[1]),
    .A2(_3417_),
    .ZN(_3428_)
  );
  INV_X1 _5569_ (
    .A(_3428_),
    .ZN(_3429_)
  );
  AND2_X1 _5570_ (
    .A1(_3118_),
    .A2(_3429_),
    .ZN(_3430_)
  );
  OR2_X1 _5571_ (
    .A1(_3427_),
    .A2(_3430_),
    .ZN(_3431_)
  );
  AND2_X1 _5572_ (
    .A1(_3426_),
    .A2(_3431_),
    .ZN(_3432_)
  );
  AND2_X1 _5573_ (
    .A1(_1290_),
    .A2(_3120_),
    .ZN(_3433_)
  );
  OR2_X1 _5574_ (
    .A1(_3432_),
    .A2(_3433_),
    .ZN(_3434_)
  );
  AND2_X1 _5575_ (
    .A1(_0654_),
    .A2(_3434_),
    .ZN(_0462_)
  );
  AND2_X1 _5576_ (
    .A1(small_[2]),
    .A2(_3114_),
    .ZN(_3435_)
  );
  AND2_X1 _5577_ (
    .A1(_0652_),
    .A2(_3060_),
    .ZN(_3436_)
  );
  XOR2_X1 _5578_ (
    .A(small_[2]),
    .B(_3428_),
    .Z(_3437_)
  );
  AND2_X1 _5579_ (
    .A1(_3118_),
    .A2(_3437_),
    .ZN(_3438_)
  );
  OR2_X1 _5580_ (
    .A1(_3435_),
    .A2(_3438_),
    .ZN(_3439_)
  );
  AND2_X1 _5581_ (
    .A1(_1346_),
    .A2(_3120_),
    .ZN(_3440_)
  );
  OR2_X1 _5582_ (
    .A1(_3439_),
    .A2(_3440_),
    .ZN(_3441_)
  );
  AND2_X1 _5583_ (
    .A1(_0654_),
    .A2(_3441_),
    .ZN(_0463_)
  );
  OR2_X1 _5584_ (
    .A1(small_[3]),
    .A2(_3436_),
    .ZN(_3442_)
  );
  AND2_X1 _5585_ (
    .A1(small_[3]),
    .A2(_3114_),
    .ZN(_3443_)
  );
  AND2_X1 _5586_ (
    .A1(small_[3]),
    .A2(_3436_),
    .ZN(_3444_)
  );
  INV_X1 _5587_ (
    .A(_3444_),
    .ZN(_3445_)
  );
  AND2_X1 _5588_ (
    .A1(_3122_),
    .A2(_3445_),
    .ZN(_3446_)
  );
  OR2_X1 _5589_ (
    .A1(_3443_),
    .A2(_3446_),
    .ZN(_3447_)
  );
  AND2_X1 _5590_ (
    .A1(_3442_),
    .A2(_3447_),
    .ZN(_3448_)
  );
  AND2_X1 _5591_ (
    .A1(_1409_),
    .A2(_3120_),
    .ZN(_3449_)
  );
  OR2_X1 _5592_ (
    .A1(_3448_),
    .A2(_3449_),
    .ZN(_3450_)
  );
  AND2_X1 _5593_ (
    .A1(_0654_),
    .A2(_3450_),
    .ZN(_0464_)
  );
  OR2_X1 _5594_ (
    .A1(small_[4]),
    .A2(_3444_),
    .ZN(_3451_)
  );
  AND2_X1 _5595_ (
    .A1(small_[4]),
    .A2(_3114_),
    .ZN(_3452_)
  );
  AND2_X1 _5596_ (
    .A1(_3055_),
    .A2(_3436_),
    .ZN(_3453_)
  );
  INV_X1 _5597_ (
    .A(_3453_),
    .ZN(_3454_)
  );
  AND2_X1 _5598_ (
    .A1(_3118_),
    .A2(_3454_),
    .ZN(_3455_)
  );
  OR2_X1 _5599_ (
    .A1(_3452_),
    .A2(_3455_),
    .ZN(_3456_)
  );
  AND2_X1 _5600_ (
    .A1(_3451_),
    .A2(_3456_),
    .ZN(_3457_)
  );
  AND2_X1 _5601_ (
    .A1(_1456_),
    .A2(_3120_),
    .ZN(_3458_)
  );
  OR2_X1 _5602_ (
    .A1(_3457_),
    .A2(_3458_),
    .ZN(_3459_)
  );
  AND2_X1 _5603_ (
    .A1(_0654_),
    .A2(_3459_),
    .ZN(_0465_)
  );
  AND2_X1 _5604_ (
    .A1(small_[5]),
    .A2(_3114_),
    .ZN(_3460_)
  );
  XOR2_X1 _5605_ (
    .A(small_[5]),
    .B(_3453_),
    .Z(_3461_)
  );
  AND2_X1 _5606_ (
    .A1(_3122_),
    .A2(_3461_),
    .ZN(_3462_)
  );
  OR2_X1 _5607_ (
    .A1(_3460_),
    .A2(_3462_),
    .ZN(_3463_)
  );
  AND2_X1 _5608_ (
    .A1(_1499_),
    .A2(_3120_),
    .ZN(_3464_)
  );
  OR2_X1 _5609_ (
    .A1(_3463_),
    .A2(_3464_),
    .ZN(_3465_)
  );
  AND2_X1 _5610_ (
    .A1(_0654_),
    .A2(_3465_),
    .ZN(_0466_)
  );
  AND2_X1 _5611_ (
    .A1(_0736_),
    .A2(_0780_),
    .ZN(_3466_)
  );
  OR2_X1 _5612_ (
    .A1(_0737_),
    .A2(_0781_),
    .ZN(_3467_)
  );
  OR2_X1 _5613_ (
    .A1(_1241_),
    .A2(_3467_),
    .ZN(_3468_)
  );
  OR2_X1 _5614_ (
    .A1(reg_mtvec[0]),
    .A2(_3466_),
    .ZN(_3469_)
  );
  AND2_X1 _5615_ (
    .A1(_0654_),
    .A2(_3469_),
    .ZN(_3470_)
  );
  AND2_X1 _5616_ (
    .A1(_3468_),
    .A2(_3470_),
    .ZN(_0467_)
  );
  OR2_X1 _5617_ (
    .A1(_1346_),
    .A2(_3467_),
    .ZN(_3471_)
  );
  OR2_X1 _5618_ (
    .A1(reg_mtvec[2]),
    .A2(_3466_),
    .ZN(_3472_)
  );
  AND2_X1 _5619_ (
    .A1(_0654_),
    .A2(_3472_),
    .ZN(_3473_)
  );
  AND2_X1 _5620_ (
    .A1(_3471_),
    .A2(_3473_),
    .ZN(_0468_)
  );
  OR2_X1 _5621_ (
    .A1(_1409_),
    .A2(_3467_),
    .ZN(_3474_)
  );
  OR2_X1 _5622_ (
    .A1(reg_mtvec[3]),
    .A2(_3466_),
    .ZN(_3475_)
  );
  AND2_X1 _5623_ (
    .A1(_0654_),
    .A2(_3475_),
    .ZN(_3476_)
  );
  AND2_X1 _5624_ (
    .A1(_3474_),
    .A2(_3476_),
    .ZN(_0469_)
  );
  OR2_X1 _5625_ (
    .A1(_1456_),
    .A2(_3467_),
    .ZN(_3477_)
  );
  OR2_X1 _5626_ (
    .A1(reg_mtvec[4]),
    .A2(_3466_),
    .ZN(_3478_)
  );
  AND2_X1 _5627_ (
    .A1(_0654_),
    .A2(_3478_),
    .ZN(_3479_)
  );
  AND2_X1 _5628_ (
    .A1(_3477_),
    .A2(_3479_),
    .ZN(_0470_)
  );
  OR2_X1 _5629_ (
    .A1(_1499_),
    .A2(_3467_),
    .ZN(_3480_)
  );
  OR2_X1 _5630_ (
    .A1(reg_mtvec[5]),
    .A2(_3466_),
    .ZN(_3481_)
  );
  AND2_X1 _5631_ (
    .A1(_0654_),
    .A2(_3481_),
    .ZN(_3482_)
  );
  AND2_X1 _5632_ (
    .A1(_3480_),
    .A2(_3482_),
    .ZN(_0471_)
  );
  OR2_X1 _5633_ (
    .A1(_1545_),
    .A2(_3467_),
    .ZN(_3483_)
  );
  OR2_X1 _5634_ (
    .A1(reg_mtvec[6]),
    .A2(_3466_),
    .ZN(_3484_)
  );
  AND2_X1 _5635_ (
    .A1(_0654_),
    .A2(_3484_),
    .ZN(_3485_)
  );
  AND2_X1 _5636_ (
    .A1(_3483_),
    .A2(_3485_),
    .ZN(_0472_)
  );
  OR2_X1 _5637_ (
    .A1(_1601_),
    .A2(_3467_),
    .ZN(_3486_)
  );
  OR2_X1 _5638_ (
    .A1(reg_mtvec[7]),
    .A2(_3466_),
    .ZN(_3487_)
  );
  AND2_X1 _5639_ (
    .A1(_0654_),
    .A2(_3487_),
    .ZN(_3488_)
  );
  AND2_X1 _5640_ (
    .A1(_3486_),
    .A2(_3488_),
    .ZN(_0473_)
  );
  OR2_X1 _5641_ (
    .A1(_1129_),
    .A2(_3467_),
    .ZN(_3489_)
  );
  OR2_X1 _5642_ (
    .A1(reg_mtvec[8]),
    .A2(_3466_),
    .ZN(_3490_)
  );
  AND2_X1 _5643_ (
    .A1(_0654_),
    .A2(_3490_),
    .ZN(_3491_)
  );
  AND2_X1 _5644_ (
    .A1(_3489_),
    .A2(_3491_),
    .ZN(_0474_)
  );
  OR2_X1 _5645_ (
    .A1(_1175_),
    .A2(_3467_),
    .ZN(_3492_)
  );
  OR2_X1 _5646_ (
    .A1(reg_mtvec[9]),
    .A2(_3466_),
    .ZN(_3493_)
  );
  AND2_X1 _5647_ (
    .A1(_0654_),
    .A2(_3493_),
    .ZN(_3494_)
  );
  AND2_X1 _5648_ (
    .A1(_3492_),
    .A2(_3494_),
    .ZN(_0475_)
  );
  OR2_X1 _5649_ (
    .A1(_1647_),
    .A2(_3467_),
    .ZN(_3495_)
  );
  OR2_X1 _5650_ (
    .A1(reg_mtvec[10]),
    .A2(_3466_),
    .ZN(_3496_)
  );
  AND2_X1 _5651_ (
    .A1(_0654_),
    .A2(_3496_),
    .ZN(_3497_)
  );
  AND2_X1 _5652_ (
    .A1(_3495_),
    .A2(_3497_),
    .ZN(_0476_)
  );
  OR2_X1 _5653_ (
    .A1(_1698_),
    .A2(_3467_),
    .ZN(_3498_)
  );
  OR2_X1 _5654_ (
    .A1(reg_mtvec[11]),
    .A2(_3466_),
    .ZN(_3499_)
  );
  AND2_X1 _5655_ (
    .A1(_0654_),
    .A2(_3499_),
    .ZN(_3500_)
  );
  AND2_X1 _5656_ (
    .A1(_3498_),
    .A2(_3500_),
    .ZN(_0477_)
  );
  OR2_X1 _5657_ (
    .A1(_1748_),
    .A2(_3467_),
    .ZN(_3501_)
  );
  OR2_X1 _5658_ (
    .A1(reg_mtvec[12]),
    .A2(_3466_),
    .ZN(_3502_)
  );
  AND2_X1 _5659_ (
    .A1(_0654_),
    .A2(_3502_),
    .ZN(_3503_)
  );
  AND2_X1 _5660_ (
    .A1(_3501_),
    .A2(_3503_),
    .ZN(_0478_)
  );
  OR2_X1 _5661_ (
    .A1(_1790_),
    .A2(_3467_),
    .ZN(_3504_)
  );
  OR2_X1 _5662_ (
    .A1(reg_mtvec[13]),
    .A2(_3466_),
    .ZN(_3505_)
  );
  AND2_X1 _5663_ (
    .A1(_0654_),
    .A2(_3505_),
    .ZN(_3506_)
  );
  AND2_X1 _5664_ (
    .A1(_3504_),
    .A2(_3506_),
    .ZN(_0479_)
  );
  OR2_X1 _5665_ (
    .A1(_1832_),
    .A2(_3467_),
    .ZN(_3507_)
  );
  OR2_X1 _5666_ (
    .A1(reg_mtvec[14]),
    .A2(_3466_),
    .ZN(_3508_)
  );
  AND2_X1 _5667_ (
    .A1(_0654_),
    .A2(_3508_),
    .ZN(_3509_)
  );
  AND2_X1 _5668_ (
    .A1(_3507_),
    .A2(_3509_),
    .ZN(_0480_)
  );
  OR2_X1 _5669_ (
    .A1(_1880_),
    .A2(_3467_),
    .ZN(_3510_)
  );
  OR2_X1 _5670_ (
    .A1(reg_mtvec[15]),
    .A2(_3466_),
    .ZN(_3511_)
  );
  AND2_X1 _5671_ (
    .A1(_0654_),
    .A2(_3511_),
    .ZN(_3512_)
  );
  AND2_X1 _5672_ (
    .A1(_3510_),
    .A2(_3512_),
    .ZN(_0481_)
  );
  OR2_X1 _5673_ (
    .A1(_0862_),
    .A2(_3467_),
    .ZN(_3513_)
  );
  OR2_X1 _5674_ (
    .A1(reg_mtvec[16]),
    .A2(_3466_),
    .ZN(_3514_)
  );
  AND2_X1 _5675_ (
    .A1(_0654_),
    .A2(_3514_),
    .ZN(_3515_)
  );
  AND2_X1 _5676_ (
    .A1(_3513_),
    .A2(_3515_),
    .ZN(_0482_)
  );
  OR2_X1 _5677_ (
    .A1(_1926_),
    .A2(_3467_),
    .ZN(_3516_)
  );
  OR2_X1 _5678_ (
    .A1(reg_mtvec[17]),
    .A2(_3466_),
    .ZN(_3517_)
  );
  AND2_X1 _5679_ (
    .A1(_0654_),
    .A2(_3517_),
    .ZN(_3518_)
  );
  AND2_X1 _5680_ (
    .A1(_3516_),
    .A2(_3518_),
    .ZN(_0483_)
  );
  OR2_X1 _5681_ (
    .A1(_0908_),
    .A2(_3467_),
    .ZN(_3519_)
  );
  OR2_X1 _5682_ (
    .A1(reg_mtvec[18]),
    .A2(_3466_),
    .ZN(_3520_)
  );
  AND2_X1 _5683_ (
    .A1(_0654_),
    .A2(_3520_),
    .ZN(_3521_)
  );
  AND2_X1 _5684_ (
    .A1(_3519_),
    .A2(_3521_),
    .ZN(_0484_)
  );
  OR2_X1 _5685_ (
    .A1(_0967_),
    .A2(_3467_),
    .ZN(_3522_)
  );
  OR2_X1 _5686_ (
    .A1(reg_mtvec[19]),
    .A2(_3466_),
    .ZN(_3523_)
  );
  AND2_X1 _5687_ (
    .A1(_0654_),
    .A2(_3523_),
    .ZN(_3524_)
  );
  AND2_X1 _5688_ (
    .A1(_3522_),
    .A2(_3524_),
    .ZN(_0485_)
  );
  OR2_X1 _5689_ (
    .A1(_1017_),
    .A2(_3467_),
    .ZN(_3525_)
  );
  OR2_X1 _5690_ (
    .A1(reg_mtvec[20]),
    .A2(_3466_),
    .ZN(_3526_)
  );
  AND2_X1 _5691_ (
    .A1(_0654_),
    .A2(_3526_),
    .ZN(_3527_)
  );
  AND2_X1 _5692_ (
    .A1(_3525_),
    .A2(_3527_),
    .ZN(_0486_)
  );
  OR2_X1 _5693_ (
    .A1(_1968_),
    .A2(_3467_),
    .ZN(_3528_)
  );
  OR2_X1 _5694_ (
    .A1(reg_mtvec[21]),
    .A2(_3466_),
    .ZN(_3529_)
  );
  AND2_X1 _5695_ (
    .A1(_0654_),
    .A2(_3529_),
    .ZN(_3530_)
  );
  AND2_X1 _5696_ (
    .A1(_3528_),
    .A2(_3530_),
    .ZN(_0487_)
  );
  OR2_X1 _5697_ (
    .A1(_2010_),
    .A2(_3467_),
    .ZN(_3531_)
  );
  OR2_X1 _5698_ (
    .A1(reg_mtvec[22]),
    .A2(_3466_),
    .ZN(_3532_)
  );
  AND2_X1 _5699_ (
    .A1(_0654_),
    .A2(_3532_),
    .ZN(_3533_)
  );
  AND2_X1 _5700_ (
    .A1(_3531_),
    .A2(_3533_),
    .ZN(_0488_)
  );
  OR2_X1 _5701_ (
    .A1(_1071_),
    .A2(_3467_),
    .ZN(_3534_)
  );
  OR2_X1 _5702_ (
    .A1(reg_mtvec[23]),
    .A2(_3466_),
    .ZN(_3535_)
  );
  AND2_X1 _5703_ (
    .A1(_0654_),
    .A2(_3535_),
    .ZN(_3536_)
  );
  AND2_X1 _5704_ (
    .A1(_3534_),
    .A2(_3536_),
    .ZN(_0489_)
  );
  OR2_X1 _5705_ (
    .A1(_2056_),
    .A2(_3467_),
    .ZN(_3537_)
  );
  OR2_X1 _5706_ (
    .A1(reg_mtvec[24]),
    .A2(_3466_),
    .ZN(_3538_)
  );
  AND2_X1 _5707_ (
    .A1(_0654_),
    .A2(_3538_),
    .ZN(_3539_)
  );
  AND2_X1 _5708_ (
    .A1(_3537_),
    .A2(_3539_),
    .ZN(_0490_)
  );
  OR2_X1 _5709_ (
    .A1(_2102_),
    .A2(_3467_),
    .ZN(_3540_)
  );
  OR2_X1 _5710_ (
    .A1(reg_mtvec[25]),
    .A2(_3466_),
    .ZN(_3541_)
  );
  AND2_X1 _5711_ (
    .A1(_0654_),
    .A2(_3541_),
    .ZN(_3542_)
  );
  AND2_X1 _5712_ (
    .A1(_3540_),
    .A2(_3542_),
    .ZN(_0491_)
  );
  OR2_X1 _5713_ (
    .A1(_2148_),
    .A2(_3467_),
    .ZN(_3543_)
  );
  OR2_X1 _5714_ (
    .A1(reg_mtvec[26]),
    .A2(_3466_),
    .ZN(_3544_)
  );
  AND2_X1 _5715_ (
    .A1(_0654_),
    .A2(_3544_),
    .ZN(_3545_)
  );
  AND2_X1 _5716_ (
    .A1(_3543_),
    .A2(_3545_),
    .ZN(_0492_)
  );
  OR2_X1 _5717_ (
    .A1(_2195_),
    .A2(_3467_),
    .ZN(_3546_)
  );
  OR2_X1 _5718_ (
    .A1(reg_mtvec[27]),
    .A2(_3466_),
    .ZN(_3547_)
  );
  AND2_X1 _5719_ (
    .A1(_0654_),
    .A2(_3547_),
    .ZN(_3548_)
  );
  AND2_X1 _5720_ (
    .A1(_3546_),
    .A2(_3548_),
    .ZN(_0493_)
  );
  OR2_X1 _5721_ (
    .A1(_2241_),
    .A2(_3467_),
    .ZN(_3549_)
  );
  OR2_X1 _5722_ (
    .A1(reg_mtvec[28]),
    .A2(_3466_),
    .ZN(_3550_)
  );
  AND2_X1 _5723_ (
    .A1(_0654_),
    .A2(_3550_),
    .ZN(_3551_)
  );
  AND2_X1 _5724_ (
    .A1(_3549_),
    .A2(_3551_),
    .ZN(_0494_)
  );
  OR2_X1 _5725_ (
    .A1(_2285_),
    .A2(_3467_),
    .ZN(_3552_)
  );
  OR2_X1 _5726_ (
    .A1(reg_mtvec[29]),
    .A2(_3466_),
    .ZN(_3553_)
  );
  AND2_X1 _5727_ (
    .A1(_0654_),
    .A2(_3553_),
    .ZN(_3554_)
  );
  AND2_X1 _5728_ (
    .A1(_3552_),
    .A2(_3554_),
    .ZN(_0495_)
  );
  OR2_X1 _5729_ (
    .A1(_2435_),
    .A2(_3467_),
    .ZN(_3555_)
  );
  OR2_X1 _5730_ (
    .A1(reg_mtvec[30]),
    .A2(_3466_),
    .ZN(_3556_)
  );
  AND2_X1 _5731_ (
    .A1(_0654_),
    .A2(_3556_),
    .ZN(_3557_)
  );
  AND2_X1 _5732_ (
    .A1(_3555_),
    .A2(_3557_),
    .ZN(_0496_)
  );
  OR2_X1 _5733_ (
    .A1(_2365_),
    .A2(_3467_),
    .ZN(_3558_)
  );
  OR2_X1 _5734_ (
    .A1(reg_mtvec[31]),
    .A2(_3466_),
    .ZN(_3559_)
  );
  AND2_X1 _5735_ (
    .A1(_0654_),
    .A2(_3559_),
    .ZN(_3560_)
  );
  AND2_X1 _5736_ (
    .A1(_3558_),
    .A2(_3560_),
    .ZN(_0497_)
  );
  AND2_X1 _5737_ (
    .A1(_0736_),
    .A2(_0834_),
    .ZN(_3561_)
  );
  OR2_X1 _5738_ (
    .A1(_0737_),
    .A2(_0835_),
    .ZN(_3562_)
  );
  MUX2_X1 _5739_ (
    .A(_2490_),
    .B(reg_mcause[0]),
    .S(_2507_),
    .Z(_3563_)
  );
  MUX2_X1 _5740_ (
    .A(_1241_),
    .B(_3563_),
    .S(_3562_),
    .Z(_3564_)
  );
  AND2_X1 _5741_ (
    .A1(_0654_),
    .A2(_3564_),
    .ZN(_0498_)
  );
  OR2_X1 _5742_ (
    .A1(io_cause[1]),
    .A2(_2468_),
    .ZN(_3565_)
  );
  MUX2_X1 _5743_ (
    .A(_3565_),
    .B(reg_mcause[1]),
    .S(_2507_),
    .Z(_3566_)
  );
  OR2_X1 _5744_ (
    .A1(_3561_),
    .A2(_3566_),
    .ZN(_3567_)
  );
  OR2_X1 _5745_ (
    .A1(_1290_),
    .A2(_3562_),
    .ZN(_3568_)
  );
  AND2_X1 _5746_ (
    .A1(_0654_),
    .A2(_3568_),
    .ZN(_3569_)
  );
  AND2_X1 _5747_ (
    .A1(_3567_),
    .A2(_3569_),
    .ZN(_0499_)
  );
  MUX2_X1 _5748_ (
    .A(_2492_),
    .B(reg_mcause[2]),
    .S(_2507_),
    .Z(_3570_)
  );
  OR2_X1 _5749_ (
    .A1(_3561_),
    .A2(_3570_),
    .ZN(_3571_)
  );
  OR2_X1 _5750_ (
    .A1(_1346_),
    .A2(_3562_),
    .ZN(_3572_)
  );
  AND2_X1 _5751_ (
    .A1(_0654_),
    .A2(_3572_),
    .ZN(_3573_)
  );
  AND2_X1 _5752_ (
    .A1(_3571_),
    .A2(_3573_),
    .ZN(_0500_)
  );
  MUX2_X1 _5753_ (
    .A(_2497_),
    .B(reg_mcause[3]),
    .S(_2507_),
    .Z(_3574_)
  );
  OR2_X1 _5754_ (
    .A1(_3561_),
    .A2(_3574_),
    .ZN(_3575_)
  );
  OR2_X1 _5755_ (
    .A1(_1409_),
    .A2(_3562_),
    .ZN(_3576_)
  );
  AND2_X1 _5756_ (
    .A1(_0654_),
    .A2(_3576_),
    .ZN(_3577_)
  );
  AND2_X1 _5757_ (
    .A1(_3575_),
    .A2(_3577_),
    .ZN(_0501_)
  );
  AND2_X1 _5758_ (
    .A1(_0654_),
    .A2(_3562_),
    .ZN(_3578_)
  );
  AND2_X1 _5759_ (
    .A1(io_cause[4]),
    .A2(_2467_),
    .ZN(_3579_)
  );
  MUX2_X1 _5760_ (
    .A(_3579_),
    .B(reg_mcause[4]),
    .S(_2507_),
    .Z(_3580_)
  );
  AND2_X1 _5761_ (
    .A1(_3578_),
    .A2(_3580_),
    .ZN(_0502_)
  );
  MUX2_X1 _5762_ (
    .A(_2483_),
    .B(reg_mcause[5]),
    .S(_2507_),
    .Z(_3581_)
  );
  AND2_X1 _5763_ (
    .A1(_3578_),
    .A2(_3581_),
    .ZN(_0503_)
  );
  MUX2_X1 _5764_ (
    .A(_2486_),
    .B(reg_mcause[6]),
    .S(_2507_),
    .Z(_3582_)
  );
  AND2_X1 _5765_ (
    .A1(_3578_),
    .A2(_3582_),
    .ZN(_0504_)
  );
  MUX2_X1 _5766_ (
    .A(_2485_),
    .B(reg_mcause[7]),
    .S(_2507_),
    .Z(_3583_)
  );
  AND2_X1 _5767_ (
    .A1(_3578_),
    .A2(_3583_),
    .ZN(_0505_)
  );
  AND2_X1 _5768_ (
    .A1(io_cause[8]),
    .A2(_2467_),
    .ZN(_3584_)
  );
  MUX2_X1 _5769_ (
    .A(_3584_),
    .B(reg_mcause[8]),
    .S(_2507_),
    .Z(_3585_)
  );
  AND2_X1 _5770_ (
    .A1(_3578_),
    .A2(_3585_),
    .ZN(_0506_)
  );
  AND2_X1 _5771_ (
    .A1(io_cause[9]),
    .A2(_2467_),
    .ZN(_3586_)
  );
  MUX2_X1 _5772_ (
    .A(_3586_),
    .B(reg_mcause[9]),
    .S(_2507_),
    .Z(_3587_)
  );
  AND2_X1 _5773_ (
    .A1(_3578_),
    .A2(_3587_),
    .ZN(_0507_)
  );
  AND2_X1 _5774_ (
    .A1(io_cause[10]),
    .A2(_2467_),
    .ZN(_3588_)
  );
  MUX2_X1 _5775_ (
    .A(_3588_),
    .B(reg_mcause[10]),
    .S(_2507_),
    .Z(_3589_)
  );
  AND2_X1 _5776_ (
    .A1(_3578_),
    .A2(_3589_),
    .ZN(_0508_)
  );
  AND2_X1 _5777_ (
    .A1(io_cause[11]),
    .A2(_2467_),
    .ZN(_3590_)
  );
  MUX2_X1 _5778_ (
    .A(_3590_),
    .B(reg_mcause[11]),
    .S(_2507_),
    .Z(_3591_)
  );
  AND2_X1 _5779_ (
    .A1(_3578_),
    .A2(_3591_),
    .ZN(_0509_)
  );
  AND2_X1 _5780_ (
    .A1(io_cause[12]),
    .A2(_2467_),
    .ZN(_3592_)
  );
  MUX2_X1 _5781_ (
    .A(_3592_),
    .B(reg_mcause[12]),
    .S(_2507_),
    .Z(_3593_)
  );
  AND2_X1 _5782_ (
    .A1(_3578_),
    .A2(_3593_),
    .ZN(_0510_)
  );
  AND2_X1 _5783_ (
    .A1(io_cause[13]),
    .A2(_2467_),
    .ZN(_3594_)
  );
  MUX2_X1 _5784_ (
    .A(_3594_),
    .B(reg_mcause[13]),
    .S(_2507_),
    .Z(_3595_)
  );
  AND2_X1 _5785_ (
    .A1(_3578_),
    .A2(_3595_),
    .ZN(_0511_)
  );
  AND2_X1 _5786_ (
    .A1(io_cause[14]),
    .A2(_2467_),
    .ZN(_3596_)
  );
  MUX2_X1 _5787_ (
    .A(_3596_),
    .B(reg_mcause[14]),
    .S(_2507_),
    .Z(_3597_)
  );
  AND2_X1 _5788_ (
    .A1(_3578_),
    .A2(_3597_),
    .ZN(_0512_)
  );
  AND2_X1 _5789_ (
    .A1(io_cause[15]),
    .A2(_2467_),
    .ZN(_3598_)
  );
  MUX2_X1 _5790_ (
    .A(_3598_),
    .B(reg_mcause[15]),
    .S(_2507_),
    .Z(_3599_)
  );
  AND2_X1 _5791_ (
    .A1(_3578_),
    .A2(_3599_),
    .ZN(_0513_)
  );
  AND2_X1 _5792_ (
    .A1(io_cause[16]),
    .A2(_2467_),
    .ZN(_3600_)
  );
  MUX2_X1 _5793_ (
    .A(_3600_),
    .B(reg_mcause[16]),
    .S(_2507_),
    .Z(_3601_)
  );
  AND2_X1 _5794_ (
    .A1(_3578_),
    .A2(_3601_),
    .ZN(_0514_)
  );
  AND2_X1 _5795_ (
    .A1(io_cause[17]),
    .A2(_2467_),
    .ZN(_3602_)
  );
  MUX2_X1 _5796_ (
    .A(_3602_),
    .B(reg_mcause[17]),
    .S(_2507_),
    .Z(_3603_)
  );
  AND2_X1 _5797_ (
    .A1(_3578_),
    .A2(_3603_),
    .ZN(_0515_)
  );
  AND2_X1 _5798_ (
    .A1(io_cause[18]),
    .A2(_2467_),
    .ZN(_3604_)
  );
  MUX2_X1 _5799_ (
    .A(_3604_),
    .B(reg_mcause[18]),
    .S(_2507_),
    .Z(_3605_)
  );
  AND2_X1 _5800_ (
    .A1(_3578_),
    .A2(_3605_),
    .ZN(_0516_)
  );
  AND2_X1 _5801_ (
    .A1(io_cause[19]),
    .A2(_2467_),
    .ZN(_3606_)
  );
  MUX2_X1 _5802_ (
    .A(_3606_),
    .B(reg_mcause[19]),
    .S(_2507_),
    .Z(_3607_)
  );
  AND2_X1 _5803_ (
    .A1(_3578_),
    .A2(_3607_),
    .ZN(_0517_)
  );
  AND2_X1 _5804_ (
    .A1(io_cause[20]),
    .A2(_2467_),
    .ZN(_3608_)
  );
  MUX2_X1 _5805_ (
    .A(_3608_),
    .B(reg_mcause[20]),
    .S(_2507_),
    .Z(_3609_)
  );
  AND2_X1 _5806_ (
    .A1(_3578_),
    .A2(_3609_),
    .ZN(_0518_)
  );
  AND2_X1 _5807_ (
    .A1(io_cause[21]),
    .A2(_2467_),
    .ZN(_3610_)
  );
  MUX2_X1 _5808_ (
    .A(_3610_),
    .B(reg_mcause[21]),
    .S(_2507_),
    .Z(_3611_)
  );
  AND2_X1 _5809_ (
    .A1(_3578_),
    .A2(_3611_),
    .ZN(_0519_)
  );
  AND2_X1 _5810_ (
    .A1(io_cause[22]),
    .A2(_2467_),
    .ZN(_3612_)
  );
  MUX2_X1 _5811_ (
    .A(_3612_),
    .B(reg_mcause[22]),
    .S(_2507_),
    .Z(_3613_)
  );
  AND2_X1 _5812_ (
    .A1(_3578_),
    .A2(_3613_),
    .ZN(_0520_)
  );
  AND2_X1 _5813_ (
    .A1(io_cause[23]),
    .A2(_2467_),
    .ZN(_3614_)
  );
  MUX2_X1 _5814_ (
    .A(_3614_),
    .B(reg_mcause[23]),
    .S(_2507_),
    .Z(_3615_)
  );
  AND2_X1 _5815_ (
    .A1(_3578_),
    .A2(_3615_),
    .ZN(_0521_)
  );
  AND2_X1 _5816_ (
    .A1(io_cause[24]),
    .A2(_2467_),
    .ZN(_3616_)
  );
  MUX2_X1 _5817_ (
    .A(_3616_),
    .B(reg_mcause[24]),
    .S(_2507_),
    .Z(_3617_)
  );
  AND2_X1 _5818_ (
    .A1(_3578_),
    .A2(_3617_),
    .ZN(_0522_)
  );
  AND2_X1 _5819_ (
    .A1(io_cause[25]),
    .A2(_2467_),
    .ZN(_3618_)
  );
  MUX2_X1 _5820_ (
    .A(_3618_),
    .B(reg_mcause[25]),
    .S(_2507_),
    .Z(_3619_)
  );
  AND2_X1 _5821_ (
    .A1(_3578_),
    .A2(_3619_),
    .ZN(_0523_)
  );
  AND2_X1 _5822_ (
    .A1(io_cause[26]),
    .A2(_2467_),
    .ZN(_3620_)
  );
  MUX2_X1 _5823_ (
    .A(_3620_),
    .B(reg_mcause[26]),
    .S(_2507_),
    .Z(_3621_)
  );
  AND2_X1 _5824_ (
    .A1(_3578_),
    .A2(_3621_),
    .ZN(_0524_)
  );
  AND2_X1 _5825_ (
    .A1(io_cause[27]),
    .A2(_2467_),
    .ZN(_3622_)
  );
  MUX2_X1 _5826_ (
    .A(_3622_),
    .B(reg_mcause[27]),
    .S(_2507_),
    .Z(_3623_)
  );
  AND2_X1 _5827_ (
    .A1(_3578_),
    .A2(_3623_),
    .ZN(_0525_)
  );
  AND2_X1 _5828_ (
    .A1(io_cause[28]),
    .A2(_2467_),
    .ZN(_3624_)
  );
  MUX2_X1 _5829_ (
    .A(_3624_),
    .B(reg_mcause[28]),
    .S(_2507_),
    .Z(_3625_)
  );
  AND2_X1 _5830_ (
    .A1(_3578_),
    .A2(_3625_),
    .ZN(_0526_)
  );
  AND2_X1 _5831_ (
    .A1(io_cause[29]),
    .A2(_2467_),
    .ZN(_3626_)
  );
  MUX2_X1 _5832_ (
    .A(_3626_),
    .B(reg_mcause[29]),
    .S(_2507_),
    .Z(_3627_)
  );
  AND2_X1 _5833_ (
    .A1(_3578_),
    .A2(_3627_),
    .ZN(_0527_)
  );
  AND2_X1 _5834_ (
    .A1(io_cause[30]),
    .A2(_2467_),
    .ZN(_3628_)
  );
  MUX2_X1 _5835_ (
    .A(_3628_),
    .B(reg_mcause[30]),
    .S(_2507_),
    .Z(_3629_)
  );
  AND2_X1 _5836_ (
    .A1(_3578_),
    .A2(_3629_),
    .ZN(_0528_)
  );
  MUX2_X1 _5837_ (
    .A(_2539_),
    .B(reg_mcause[31]),
    .S(_2507_),
    .Z(_3630_)
  );
  OR2_X1 _5838_ (
    .A1(_3561_),
    .A2(_3630_),
    .ZN(_3631_)
  );
  OR2_X1 _5839_ (
    .A1(_2365_),
    .A2(_3562_),
    .ZN(_3632_)
  );
  AND2_X1 _5840_ (
    .A1(_0654_),
    .A2(_3632_),
    .ZN(_3633_)
  );
  AND2_X1 _5841_ (
    .A1(_3631_),
    .A2(_3633_),
    .ZN(_0529_)
  );
  OR2_X1 _5842_ (
    .A1(_0737_),
    .A2(_1353_),
    .ZN(_3634_)
  );
  MUX2_X1 _5843_ (
    .A(_1409_),
    .B(reg_mie[3]),
    .S(_3634_),
    .Z(_0530_)
  );
  MUX2_X1 _5844_ (
    .A(_1601_),
    .B(reg_mie[7]),
    .S(_3634_),
    .Z(_0531_)
  );
  MUX2_X1 _5845_ (
    .A(_1698_),
    .B(reg_mie[11]),
    .S(_3634_),
    .Z(_0532_)
  );
  AND2_X1 _5846_ (
    .A1(_0003_),
    .A2(_0733_),
    .ZN(_3635_)
  );
  INV_X1 _5847_ (
    .A(_3635_),
    .ZN(_3636_)
  );
  AND2_X1 _5848_ (
    .A1(_0736_),
    .A2(_3635_),
    .ZN(_3637_)
  );
  OR2_X1 _5849_ (
    .A1(_0737_),
    .A2(_3636_),
    .ZN(_3638_)
  );
  MUX2_X1 _5850_ (
    .A(reg_pmp_7_cfg_r),
    .B(_2056_),
    .S(_3637_),
    .Z(_0533_)
  );
  MUX2_X1 _5851_ (
    .A(reg_pmp_7_cfg_w),
    .B(_2322_),
    .S(_3637_),
    .Z(_0534_)
  );
  MUX2_X1 _5852_ (
    .A(reg_pmp_7_cfg_x),
    .B(_2148_),
    .S(_3637_),
    .Z(_0535_)
  );
  AND2_X1 _5853_ (
    .A1(_0736_),
    .A2(_0849_),
    .ZN(_3639_)
  );
  INV_X1 _5854_ (
    .A(_3639_),
    .ZN(_3640_)
  );
  OR2_X1 _5855_ (
    .A1(reg_pmp_7_cfg_l),
    .A2(_3640_),
    .ZN(_3641_)
  );
  MUX2_X1 _5856_ (
    .A(_1241_),
    .B(reg_pmp_7_addr[0]),
    .S(_3641_),
    .Z(_0536_)
  );
  MUX2_X1 _5857_ (
    .A(_1290_),
    .B(reg_pmp_7_addr[1]),
    .S(_3641_),
    .Z(_0537_)
  );
  MUX2_X1 _5858_ (
    .A(_1346_),
    .B(reg_pmp_7_addr[2]),
    .S(_3641_),
    .Z(_0538_)
  );
  MUX2_X1 _5859_ (
    .A(_1409_),
    .B(reg_pmp_7_addr[3]),
    .S(_3641_),
    .Z(_0539_)
  );
  MUX2_X1 _5860_ (
    .A(_1456_),
    .B(reg_pmp_7_addr[4]),
    .S(_3641_),
    .Z(_0540_)
  );
  MUX2_X1 _5861_ (
    .A(_1499_),
    .B(reg_pmp_7_addr[5]),
    .S(_3641_),
    .Z(_0541_)
  );
  MUX2_X1 _5862_ (
    .A(_1545_),
    .B(reg_pmp_7_addr[6]),
    .S(_3641_),
    .Z(_0542_)
  );
  MUX2_X1 _5863_ (
    .A(_1601_),
    .B(reg_pmp_7_addr[7]),
    .S(_3641_),
    .Z(_0543_)
  );
  MUX2_X1 _5864_ (
    .A(_1129_),
    .B(reg_pmp_7_addr[8]),
    .S(_3641_),
    .Z(_0544_)
  );
  MUX2_X1 _5865_ (
    .A(_1175_),
    .B(reg_pmp_7_addr[9]),
    .S(_3641_),
    .Z(_0545_)
  );
  MUX2_X1 _5866_ (
    .A(_1647_),
    .B(reg_pmp_7_addr[10]),
    .S(_3641_),
    .Z(_0546_)
  );
  MUX2_X1 _5867_ (
    .A(_1698_),
    .B(reg_pmp_7_addr[11]),
    .S(_3641_),
    .Z(_0547_)
  );
  MUX2_X1 _5868_ (
    .A(_1748_),
    .B(reg_pmp_7_addr[12]),
    .S(_3641_),
    .Z(_0548_)
  );
  MUX2_X1 _5869_ (
    .A(_1790_),
    .B(reg_pmp_7_addr[13]),
    .S(_3641_),
    .Z(_0549_)
  );
  MUX2_X1 _5870_ (
    .A(_1832_),
    .B(reg_pmp_7_addr[14]),
    .S(_3641_),
    .Z(_0550_)
  );
  MUX2_X1 _5871_ (
    .A(_1880_),
    .B(reg_pmp_7_addr[15]),
    .S(_3641_),
    .Z(_0551_)
  );
  MUX2_X1 _5872_ (
    .A(_0862_),
    .B(reg_pmp_7_addr[16]),
    .S(_3641_),
    .Z(_0552_)
  );
  MUX2_X1 _5873_ (
    .A(_1926_),
    .B(reg_pmp_7_addr[17]),
    .S(_3641_),
    .Z(_0553_)
  );
  MUX2_X1 _5874_ (
    .A(_0908_),
    .B(reg_pmp_7_addr[18]),
    .S(_3641_),
    .Z(_0554_)
  );
  MUX2_X1 _5875_ (
    .A(_0967_),
    .B(reg_pmp_7_addr[19]),
    .S(_3641_),
    .Z(_0555_)
  );
  MUX2_X1 _5876_ (
    .A(_1017_),
    .B(reg_pmp_7_addr[20]),
    .S(_3641_),
    .Z(_0556_)
  );
  MUX2_X1 _5877_ (
    .A(_1968_),
    .B(reg_pmp_7_addr[21]),
    .S(_3641_),
    .Z(_0557_)
  );
  MUX2_X1 _5878_ (
    .A(_2010_),
    .B(reg_pmp_7_addr[22]),
    .S(_3641_),
    .Z(_0558_)
  );
  MUX2_X1 _5879_ (
    .A(_1071_),
    .B(reg_pmp_7_addr[23]),
    .S(_3641_),
    .Z(_0559_)
  );
  MUX2_X1 _5880_ (
    .A(_2056_),
    .B(reg_pmp_7_addr[24]),
    .S(_3641_),
    .Z(_0560_)
  );
  MUX2_X1 _5881_ (
    .A(_2102_),
    .B(reg_pmp_7_addr[25]),
    .S(_3641_),
    .Z(_0561_)
  );
  MUX2_X1 _5882_ (
    .A(_2148_),
    .B(reg_pmp_7_addr[26]),
    .S(_3641_),
    .Z(_0562_)
  );
  MUX2_X1 _5883_ (
    .A(_2195_),
    .B(reg_pmp_7_addr[27]),
    .S(_3641_),
    .Z(_0563_)
  );
  MUX2_X1 _5884_ (
    .A(_2241_),
    .B(reg_pmp_7_addr[28]),
    .S(_3641_),
    .Z(_0564_)
  );
  MUX2_X1 _5885_ (
    .A(_2285_),
    .B(reg_pmp_7_addr[29]),
    .S(_3641_),
    .Z(_0565_)
  );
  OR2_X1 _5886_ (
    .A1(reg_pmp_7_cfg_a[0]),
    .A2(_3637_),
    .ZN(_3642_)
  );
  AND2_X1 _5887_ (
    .A1(_0654_),
    .A2(_3642_),
    .ZN(_3643_)
  );
  OR2_X1 _5888_ (
    .A1(_2195_),
    .A2(_3638_),
    .ZN(_3644_)
  );
  AND2_X1 _5889_ (
    .A1(_3643_),
    .A2(_3644_),
    .ZN(_0566_)
  );
  OR2_X1 _5890_ (
    .A1(reg_pmp_7_cfg_a[1]),
    .A2(_3637_),
    .ZN(_3645_)
  );
  AND2_X1 _5891_ (
    .A1(_0654_),
    .A2(_3645_),
    .ZN(_3646_)
  );
  OR2_X1 _5892_ (
    .A1(_2241_),
    .A2(_3638_),
    .ZN(_3647_)
  );
  AND2_X1 _5893_ (
    .A1(_3646_),
    .A2(_3647_),
    .ZN(_0567_)
  );
  OR2_X1 _5894_ (
    .A1(reg_pmp_7_cfg_l),
    .A2(_3637_),
    .ZN(_3648_)
  );
  AND2_X1 _5895_ (
    .A1(_0654_),
    .A2(_3648_),
    .ZN(_3649_)
  );
  OR2_X1 _5896_ (
    .A1(_2365_),
    .A2(_3638_),
    .ZN(_3650_)
  );
  AND2_X1 _5897_ (
    .A1(_3649_),
    .A2(_3650_),
    .ZN(_0568_)
  );
  AND2_X1 _5898_ (
    .A1(large_1[0]),
    .A2(_2660_),
    .ZN(_3651_)
  );
  MUX2_X1 _5899_ (
    .A(_large_r_T_3[0]),
    .B(large_1[0]),
    .S(_2627_),
    .Z(_3652_)
  );
  AND2_X1 _5900_ (
    .A1(_2669_),
    .A2(_3652_),
    .ZN(_3653_)
  );
  OR2_X1 _5901_ (
    .A1(_3651_),
    .A2(_3653_),
    .ZN(_3654_)
  );
  AND2_X1 _5902_ (
    .A1(_1545_),
    .A2(_2662_),
    .ZN(_3655_)
  );
  OR2_X1 _5903_ (
    .A1(_3654_),
    .A2(_3655_),
    .ZN(_3656_)
  );
  AND2_X1 _5904_ (
    .A1(_0654_),
    .A2(_3656_),
    .ZN(_0569_)
  );
  OR2_X1 _5905_ (
    .A1(large_1[1]),
    .A2(_2616_),
    .ZN(_3657_)
  );
  AND2_X1 _5906_ (
    .A1(large_1[1]),
    .A2(_2660_),
    .ZN(_3658_)
  );
  AND2_X1 _5907_ (
    .A1(_2669_),
    .A2(_3657_),
    .ZN(_3659_)
  );
  INV_X1 _5908_ (
    .A(_3659_),
    .ZN(_3660_)
  );
  OR2_X1 _5909_ (
    .A1(_2629_),
    .A2(_3660_),
    .ZN(_3661_)
  );
  INV_X1 _5910_ (
    .A(_3661_),
    .ZN(_3662_)
  );
  OR2_X1 _5911_ (
    .A1(_3658_),
    .A2(_3662_),
    .ZN(_3663_)
  );
  AND2_X1 _5912_ (
    .A1(_1601_),
    .A2(_2662_),
    .ZN(_3664_)
  );
  OR2_X1 _5913_ (
    .A1(_3663_),
    .A2(_3664_),
    .ZN(_3665_)
  );
  AND2_X1 _5914_ (
    .A1(_0654_),
    .A2(_3665_),
    .ZN(_0570_)
  );
  AND2_X1 _5915_ (
    .A1(_1129_),
    .A2(_2662_),
    .ZN(_3666_)
  );
  OR2_X1 _5916_ (
    .A1(large_1[2]),
    .A2(_2617_),
    .ZN(_3667_)
  );
  AND2_X1 _5917_ (
    .A1(large_1[2]),
    .A2(_2660_),
    .ZN(_3668_)
  );
  AND2_X1 _5918_ (
    .A1(large_1[2]),
    .A2(_2617_),
    .ZN(_3669_)
  );
  INV_X1 _5919_ (
    .A(_3669_),
    .ZN(_3670_)
  );
  AND2_X1 _5920_ (
    .A1(_2666_),
    .A2(_3670_),
    .ZN(_3671_)
  );
  OR2_X1 _5921_ (
    .A1(_3668_),
    .A2(_3671_),
    .ZN(_3672_)
  );
  AND2_X1 _5922_ (
    .A1(_3667_),
    .A2(_3672_),
    .ZN(_3673_)
  );
  OR2_X1 _5923_ (
    .A1(_3666_),
    .A2(_3673_),
    .ZN(_3674_)
  );
  AND2_X1 _5924_ (
    .A1(_0654_),
    .A2(_3674_),
    .ZN(_0571_)
  );
  AND2_X1 _5925_ (
    .A1(_1175_),
    .A2(_2662_),
    .ZN(_3675_)
  );
  OR2_X1 _5926_ (
    .A1(large_1[3]),
    .A2(_3669_),
    .ZN(_3676_)
  );
  AND2_X1 _5927_ (
    .A1(large_1[3]),
    .A2(_2660_),
    .ZN(_3677_)
  );
  AND2_X1 _5928_ (
    .A1(large_1[3]),
    .A2(_3669_),
    .ZN(_3678_)
  );
  INV_X1 _5929_ (
    .A(_3678_),
    .ZN(_3679_)
  );
  AND2_X1 _5930_ (
    .A1(_2666_),
    .A2(_3679_),
    .ZN(_3680_)
  );
  OR2_X1 _5931_ (
    .A1(_3677_),
    .A2(_3680_),
    .ZN(_3681_)
  );
  AND2_X1 _5932_ (
    .A1(_3676_),
    .A2(_3681_),
    .ZN(_3682_)
  );
  OR2_X1 _5933_ (
    .A1(_3675_),
    .A2(_3682_),
    .ZN(_3683_)
  );
  AND2_X1 _5934_ (
    .A1(_0654_),
    .A2(_3683_),
    .ZN(_0572_)
  );
  OR2_X1 _5935_ (
    .A1(large_1[4]),
    .A2(_3678_),
    .ZN(_3684_)
  );
  AND2_X1 _5936_ (
    .A1(_2598_),
    .A2(_3669_),
    .ZN(_3685_)
  );
  INV_X1 _5937_ (
    .A(_3685_),
    .ZN(_3686_)
  );
  AND2_X1 _5938_ (
    .A1(_2666_),
    .A2(_3686_),
    .ZN(_3687_)
  );
  AND2_X1 _5939_ (
    .A1(_3684_),
    .A2(_3687_),
    .ZN(_3688_)
  );
  AND2_X1 _5940_ (
    .A1(large_1[4]),
    .A2(_2660_),
    .ZN(_3689_)
  );
  OR2_X1 _5941_ (
    .A1(_3688_),
    .A2(_3689_),
    .ZN(_3690_)
  );
  AND2_X1 _5942_ (
    .A1(_1647_),
    .A2(_2662_),
    .ZN(_3691_)
  );
  OR2_X1 _5943_ (
    .A1(_3690_),
    .A2(_3691_),
    .ZN(_3692_)
  );
  AND2_X1 _5944_ (
    .A1(_0654_),
    .A2(_3692_),
    .ZN(_0573_)
  );
  AND2_X1 _5945_ (
    .A1(_1698_),
    .A2(_2662_),
    .ZN(_3693_)
  );
  OR2_X1 _5946_ (
    .A1(large_1[5]),
    .A2(_3685_),
    .ZN(_3694_)
  );
  AND2_X1 _5947_ (
    .A1(large_1[5]),
    .A2(_2660_),
    .ZN(_3695_)
  );
  AND2_X1 _5948_ (
    .A1(large_1[5]),
    .A2(_3685_),
    .ZN(_3696_)
  );
  INV_X1 _5949_ (
    .A(_3696_),
    .ZN(_3697_)
  );
  AND2_X1 _5950_ (
    .A1(_2666_),
    .A2(_3697_),
    .ZN(_3698_)
  );
  OR2_X1 _5951_ (
    .A1(_3695_),
    .A2(_3698_),
    .ZN(_3699_)
  );
  AND2_X1 _5952_ (
    .A1(_3694_),
    .A2(_3699_),
    .ZN(_3700_)
  );
  OR2_X1 _5953_ (
    .A1(_3693_),
    .A2(_3700_),
    .ZN(_3701_)
  );
  AND2_X1 _5954_ (
    .A1(_0654_),
    .A2(_3701_),
    .ZN(_0574_)
  );
  OR2_X1 _5955_ (
    .A1(large_1[6]),
    .A2(_3696_),
    .ZN(_3702_)
  );
  AND2_X1 _5956_ (
    .A1(large_1[6]),
    .A2(_2660_),
    .ZN(_3703_)
  );
  OR2_X1 _5957_ (
    .A1(_2630_),
    .A2(_2670_),
    .ZN(_3704_)
  );
  INV_X1 _5958_ (
    .A(_3704_),
    .ZN(_3705_)
  );
  AND2_X1 _5959_ (
    .A1(_3702_),
    .A2(_3705_),
    .ZN(_3706_)
  );
  OR2_X1 _5960_ (
    .A1(_3703_),
    .A2(_3706_),
    .ZN(_3707_)
  );
  AND2_X1 _5961_ (
    .A1(_1748_),
    .A2(_2662_),
    .ZN(_3708_)
  );
  OR2_X1 _5962_ (
    .A1(_3707_),
    .A2(_3708_),
    .ZN(_3709_)
  );
  AND2_X1 _5963_ (
    .A1(_0654_),
    .A2(_3709_),
    .ZN(_0575_)
  );
  OR2_X1 _5964_ (
    .A1(large_1[7]),
    .A2(_2618_),
    .ZN(_3710_)
  );
  AND2_X1 _5965_ (
    .A1(_2669_),
    .A2(_3710_),
    .ZN(_3711_)
  );
  AND2_X1 _5966_ (
    .A1(large_1[7]),
    .A2(_2618_),
    .ZN(_3712_)
  );
  INV_X1 _5967_ (
    .A(_3712_),
    .ZN(_3713_)
  );
  AND2_X1 _5968_ (
    .A1(_3711_),
    .A2(_3713_),
    .ZN(_3714_)
  );
  AND2_X1 _5969_ (
    .A1(large_1[7]),
    .A2(_2660_),
    .ZN(_3715_)
  );
  AND2_X1 _5970_ (
    .A1(_1790_),
    .A2(_2667_),
    .ZN(_3716_)
  );
  OR2_X1 _5971_ (
    .A1(_3715_),
    .A2(_3716_),
    .ZN(_3717_)
  );
  OR2_X1 _5972_ (
    .A1(_3714_),
    .A2(_3717_),
    .ZN(_3718_)
  );
  AND2_X1 _5973_ (
    .A1(_0654_),
    .A2(_3718_),
    .ZN(_0576_)
  );
  OR2_X1 _5974_ (
    .A1(large_1[8]),
    .A2(_3712_),
    .ZN(_3719_)
  );
  AND2_X1 _5975_ (
    .A1(large_1[8]),
    .A2(_2660_),
    .ZN(_3720_)
  );
  AND2_X1 _5976_ (
    .A1(large_1[8]),
    .A2(_3712_),
    .ZN(_3721_)
  );
  INV_X1 _5977_ (
    .A(_3721_),
    .ZN(_3722_)
  );
  AND2_X1 _5978_ (
    .A1(_2666_),
    .A2(_3722_),
    .ZN(_3723_)
  );
  OR2_X1 _5979_ (
    .A1(_3720_),
    .A2(_3723_),
    .ZN(_3724_)
  );
  AND2_X1 _5980_ (
    .A1(_3719_),
    .A2(_3724_),
    .ZN(_3725_)
  );
  AND2_X1 _5981_ (
    .A1(_1832_),
    .A2(_2662_),
    .ZN(_3726_)
  );
  OR2_X1 _5982_ (
    .A1(_3725_),
    .A2(_3726_),
    .ZN(_3727_)
  );
  AND2_X1 _5983_ (
    .A1(_0654_),
    .A2(_3727_),
    .ZN(_0577_)
  );
  OR2_X1 _5984_ (
    .A1(large_1[9]),
    .A2(_3721_),
    .ZN(_3728_)
  );
  OR2_X1 _5985_ (
    .A1(_2645_),
    .A2(_2670_),
    .ZN(_3729_)
  );
  INV_X1 _5986_ (
    .A(_3729_),
    .ZN(_3730_)
  );
  AND2_X1 _5987_ (
    .A1(_3728_),
    .A2(_3730_),
    .ZN(_3731_)
  );
  AND2_X1 _5988_ (
    .A1(large_1[9]),
    .A2(_2660_),
    .ZN(_3732_)
  );
  AND2_X1 _5989_ (
    .A1(_1880_),
    .A2(_2662_),
    .ZN(_3733_)
  );
  OR2_X1 _5990_ (
    .A1(_3732_),
    .A2(_3733_),
    .ZN(_3734_)
  );
  OR2_X1 _5991_ (
    .A1(_3731_),
    .A2(_3734_),
    .ZN(_3735_)
  );
  AND2_X1 _5992_ (
    .A1(_0654_),
    .A2(_3735_),
    .ZN(_0578_)
  );
  OR2_X1 _5993_ (
    .A1(large_1[10]),
    .A2(_2619_),
    .ZN(_3736_)
  );
  AND2_X1 _5994_ (
    .A1(large_1[10]),
    .A2(_2660_),
    .ZN(_3737_)
  );
  AND2_X1 _5995_ (
    .A1(_2669_),
    .A2(_3736_),
    .ZN(_3738_)
  );
  AND2_X1 _5996_ (
    .A1(_2648_),
    .A2(_3738_),
    .ZN(_3739_)
  );
  AND2_X1 _5997_ (
    .A1(_0862_),
    .A2(_2667_),
    .ZN(_3740_)
  );
  OR2_X1 _5998_ (
    .A1(_3739_),
    .A2(_3740_),
    .ZN(_3741_)
  );
  OR2_X1 _5999_ (
    .A1(_3737_),
    .A2(_3741_),
    .ZN(_3742_)
  );
  AND2_X1 _6000_ (
    .A1(_0654_),
    .A2(_3742_),
    .ZN(_0579_)
  );
  OR2_X1 _6001_ (
    .A1(large_1[11]),
    .A2(_2620_),
    .ZN(_3743_)
  );
  OR2_X1 _6002_ (
    .A1(_2649_),
    .A2(_2670_),
    .ZN(_3744_)
  );
  INV_X1 _6003_ (
    .A(_3744_),
    .ZN(_3745_)
  );
  AND2_X1 _6004_ (
    .A1(_3743_),
    .A2(_3745_),
    .ZN(_3746_)
  );
  AND2_X1 _6005_ (
    .A1(large_1[11]),
    .A2(_2660_),
    .ZN(_3747_)
  );
  AND2_X1 _6006_ (
    .A1(_1926_),
    .A2(_2662_),
    .ZN(_3748_)
  );
  OR2_X1 _6007_ (
    .A1(_3747_),
    .A2(_3748_),
    .ZN(_3749_)
  );
  OR2_X1 _6008_ (
    .A1(_3746_),
    .A2(_3749_),
    .ZN(_3750_)
  );
  AND2_X1 _6009_ (
    .A1(_0654_),
    .A2(_3750_),
    .ZN(_0580_)
  );
  OR2_X1 _6010_ (
    .A1(large_1[12]),
    .A2(_2621_),
    .ZN(_3751_)
  );
  AND2_X1 _6011_ (
    .A1(_2669_),
    .A2(_3751_),
    .ZN(_3752_)
  );
  AND2_X1 _6012_ (
    .A1(large_1[12]),
    .A2(_2633_),
    .ZN(_3753_)
  );
  INV_X1 _6013_ (
    .A(_3753_),
    .ZN(_3754_)
  );
  AND2_X1 _6014_ (
    .A1(_3752_),
    .A2(_3754_),
    .ZN(_3755_)
  );
  AND2_X1 _6015_ (
    .A1(large_1[12]),
    .A2(_2660_),
    .ZN(_3756_)
  );
  AND2_X1 _6016_ (
    .A1(_0908_),
    .A2(_2667_),
    .ZN(_3757_)
  );
  OR2_X1 _6017_ (
    .A1(_3756_),
    .A2(_3757_),
    .ZN(_3758_)
  );
  OR2_X1 _6018_ (
    .A1(_3755_),
    .A2(_3758_),
    .ZN(_3759_)
  );
  AND2_X1 _6019_ (
    .A1(_0654_),
    .A2(_3759_),
    .ZN(_0581_)
  );
  OR2_X1 _6020_ (
    .A1(large_1[13]),
    .A2(_3753_),
    .ZN(_3760_)
  );
  AND2_X1 _6021_ (
    .A1(large_1[13]),
    .A2(_3753_),
    .ZN(_3761_)
  );
  INV_X1 _6022_ (
    .A(_3761_),
    .ZN(_3762_)
  );
  AND2_X1 _6023_ (
    .A1(_2669_),
    .A2(_3762_),
    .ZN(_3763_)
  );
  AND2_X1 _6024_ (
    .A1(_3760_),
    .A2(_3763_),
    .ZN(_3764_)
  );
  AND2_X1 _6025_ (
    .A1(large_1[13]),
    .A2(_2660_),
    .ZN(_3765_)
  );
  AND2_X1 _6026_ (
    .A1(_0967_),
    .A2(_2667_),
    .ZN(_3766_)
  );
  OR2_X1 _6027_ (
    .A1(_3765_),
    .A2(_3766_),
    .ZN(_3767_)
  );
  OR2_X1 _6028_ (
    .A1(_3764_),
    .A2(_3767_),
    .ZN(_3768_)
  );
  AND2_X1 _6029_ (
    .A1(_0654_),
    .A2(_3768_),
    .ZN(_0582_)
  );
  OR2_X1 _6030_ (
    .A1(large_1[14]),
    .A2(_3761_),
    .ZN(_3769_)
  );
  OR2_X1 _6031_ (
    .A1(_2651_),
    .A2(_2670_),
    .ZN(_3770_)
  );
  INV_X1 _6032_ (
    .A(_3770_),
    .ZN(_3771_)
  );
  AND2_X1 _6033_ (
    .A1(_3769_),
    .A2(_3771_),
    .ZN(_3772_)
  );
  AND2_X1 _6034_ (
    .A1(large_1[14]),
    .A2(_2660_),
    .ZN(_3773_)
  );
  AND2_X1 _6035_ (
    .A1(_1017_),
    .A2(_2662_),
    .ZN(_3774_)
  );
  OR2_X1 _6036_ (
    .A1(_3773_),
    .A2(_3774_),
    .ZN(_3775_)
  );
  OR2_X1 _6037_ (
    .A1(_3772_),
    .A2(_3775_),
    .ZN(_3776_)
  );
  AND2_X1 _6038_ (
    .A1(_0654_),
    .A2(_3776_),
    .ZN(_0583_)
  );
  OR2_X1 _6039_ (
    .A1(large_1[15]),
    .A2(_2622_),
    .ZN(_3777_)
  );
  AND2_X1 _6040_ (
    .A1(large_1[15]),
    .A2(_2634_),
    .ZN(_3778_)
  );
  OR2_X1 _6041_ (
    .A1(_2670_),
    .A2(_3778_),
    .ZN(_3779_)
  );
  INV_X1 _6042_ (
    .A(_3779_),
    .ZN(_3780_)
  );
  AND2_X1 _6043_ (
    .A1(_3777_),
    .A2(_3780_),
    .ZN(_3781_)
  );
  AND2_X1 _6044_ (
    .A1(large_1[15]),
    .A2(_2660_),
    .ZN(_3782_)
  );
  AND2_X1 _6045_ (
    .A1(_1968_),
    .A2(_2667_),
    .ZN(_3783_)
  );
  OR2_X1 _6046_ (
    .A1(_3782_),
    .A2(_3783_),
    .ZN(_3784_)
  );
  OR2_X1 _6047_ (
    .A1(_3781_),
    .A2(_3784_),
    .ZN(_3785_)
  );
  AND2_X1 _6048_ (
    .A1(_0654_),
    .A2(_3785_),
    .ZN(_0584_)
  );
  OR2_X1 _6049_ (
    .A1(large_1[16]),
    .A2(_3778_),
    .ZN(_3786_)
  );
  AND2_X1 _6050_ (
    .A1(large_1[16]),
    .A2(_3778_),
    .ZN(_3787_)
  );
  INV_X1 _6051_ (
    .A(_3787_),
    .ZN(_3788_)
  );
  AND2_X1 _6052_ (
    .A1(_2669_),
    .A2(_3788_),
    .ZN(_3789_)
  );
  AND2_X1 _6053_ (
    .A1(_3786_),
    .A2(_3789_),
    .ZN(_3790_)
  );
  AND2_X1 _6054_ (
    .A1(large_1[16]),
    .A2(_2660_),
    .ZN(_3791_)
  );
  AND2_X1 _6055_ (
    .A1(_2010_),
    .A2(_2662_),
    .ZN(_3792_)
  );
  OR2_X1 _6056_ (
    .A1(_3791_),
    .A2(_3792_),
    .ZN(_3793_)
  );
  OR2_X1 _6057_ (
    .A1(_3790_),
    .A2(_3793_),
    .ZN(_3794_)
  );
  AND2_X1 _6058_ (
    .A1(_0654_),
    .A2(_3794_),
    .ZN(_0585_)
  );
  OR2_X1 _6059_ (
    .A1(large_1[17]),
    .A2(_3787_),
    .ZN(_3795_)
  );
  AND2_X1 _6060_ (
    .A1(large_1[17]),
    .A2(_3787_),
    .ZN(_3796_)
  );
  INV_X1 _6061_ (
    .A(_3796_),
    .ZN(_3797_)
  );
  AND2_X1 _6062_ (
    .A1(_2669_),
    .A2(_3797_),
    .ZN(_3798_)
  );
  AND2_X1 _6063_ (
    .A1(_3795_),
    .A2(_3798_),
    .ZN(_3799_)
  );
  AND2_X1 _6064_ (
    .A1(large_1[17]),
    .A2(_2660_),
    .ZN(_3800_)
  );
  AND2_X1 _6065_ (
    .A1(_1071_),
    .A2(_2662_),
    .ZN(_3801_)
  );
  OR2_X1 _6066_ (
    .A1(_3800_),
    .A2(_3801_),
    .ZN(_3802_)
  );
  OR2_X1 _6067_ (
    .A1(_3799_),
    .A2(_3802_),
    .ZN(_3803_)
  );
  AND2_X1 _6068_ (
    .A1(_0654_),
    .A2(_3803_),
    .ZN(_0586_)
  );
  OR2_X1 _6069_ (
    .A1(large_1[18]),
    .A2(_3796_),
    .ZN(_3804_)
  );
  AND2_X1 _6070_ (
    .A1(_2669_),
    .A2(_3804_),
    .ZN(_3805_)
  );
  AND2_X1 _6071_ (
    .A1(large_1[18]),
    .A2(_3796_),
    .ZN(_3806_)
  );
  INV_X1 _6072_ (
    .A(_3806_),
    .ZN(_3807_)
  );
  AND2_X1 _6073_ (
    .A1(_3805_),
    .A2(_3807_),
    .ZN(_3808_)
  );
  AND2_X1 _6074_ (
    .A1(large_1[18]),
    .A2(_2660_),
    .ZN(_3809_)
  );
  AND2_X1 _6075_ (
    .A1(_2056_),
    .A2(_2662_),
    .ZN(_3810_)
  );
  OR2_X1 _6076_ (
    .A1(_3809_),
    .A2(_3810_),
    .ZN(_3811_)
  );
  OR2_X1 _6077_ (
    .A1(_3808_),
    .A2(_3811_),
    .ZN(_3812_)
  );
  AND2_X1 _6078_ (
    .A1(_0654_),
    .A2(_3812_),
    .ZN(_0587_)
  );
  OR2_X1 _6079_ (
    .A1(large_1[19]),
    .A2(_3806_),
    .ZN(_3813_)
  );
  AND2_X1 _6080_ (
    .A1(large_1[19]),
    .A2(_3806_),
    .ZN(_3814_)
  );
  INV_X1 _6081_ (
    .A(_3814_),
    .ZN(_3815_)
  );
  AND2_X1 _6082_ (
    .A1(_2669_),
    .A2(_3815_),
    .ZN(_3816_)
  );
  AND2_X1 _6083_ (
    .A1(_3813_),
    .A2(_3816_),
    .ZN(_3817_)
  );
  AND2_X1 _6084_ (
    .A1(large_1[19]),
    .A2(_2660_),
    .ZN(_3818_)
  );
  AND2_X1 _6085_ (
    .A1(_2102_),
    .A2(_2667_),
    .ZN(_3819_)
  );
  OR2_X1 _6086_ (
    .A1(_3818_),
    .A2(_3819_),
    .ZN(_3820_)
  );
  OR2_X1 _6087_ (
    .A1(_3817_),
    .A2(_3820_),
    .ZN(_3821_)
  );
  AND2_X1 _6088_ (
    .A1(_0654_),
    .A2(_3821_),
    .ZN(_0588_)
  );
  OR2_X1 _6089_ (
    .A1(large_1[20]),
    .A2(_3814_),
    .ZN(_3822_)
  );
  AND2_X1 _6090_ (
    .A1(large_1[20]),
    .A2(_3814_),
    .ZN(_3823_)
  );
  OR2_X1 _6091_ (
    .A1(_0628_),
    .A2(_3815_),
    .ZN(_3824_)
  );
  AND2_X1 _6092_ (
    .A1(_2669_),
    .A2(_3824_),
    .ZN(_3825_)
  );
  AND2_X1 _6093_ (
    .A1(_3822_),
    .A2(_3825_),
    .ZN(_3826_)
  );
  AND2_X1 _6094_ (
    .A1(large_1[20]),
    .A2(_2660_),
    .ZN(_3827_)
  );
  AND2_X1 _6095_ (
    .A1(_2148_),
    .A2(_2662_),
    .ZN(_3828_)
  );
  OR2_X1 _6096_ (
    .A1(_3827_),
    .A2(_3828_),
    .ZN(_3829_)
  );
  OR2_X1 _6097_ (
    .A1(_3826_),
    .A2(_3829_),
    .ZN(_3830_)
  );
  AND2_X1 _6098_ (
    .A1(_0654_),
    .A2(_3830_),
    .ZN(_0589_)
  );
  OR2_X1 _6099_ (
    .A1(large_1[21]),
    .A2(_3823_),
    .ZN(_3831_)
  );
  AND2_X1 _6100_ (
    .A1(_2669_),
    .A2(_3831_),
    .ZN(_3832_)
  );
  AND2_X1 _6101_ (
    .A1(large_1[21]),
    .A2(_3823_),
    .ZN(_3833_)
  );
  INV_X1 _6102_ (
    .A(_3833_),
    .ZN(_3834_)
  );
  AND2_X1 _6103_ (
    .A1(_3832_),
    .A2(_3834_),
    .ZN(_3835_)
  );
  AND2_X1 _6104_ (
    .A1(large_1[21]),
    .A2(_2660_),
    .ZN(_3836_)
  );
  AND2_X1 _6105_ (
    .A1(_2195_),
    .A2(_2667_),
    .ZN(_3837_)
  );
  OR2_X1 _6106_ (
    .A1(_3836_),
    .A2(_3837_),
    .ZN(_3838_)
  );
  OR2_X1 _6107_ (
    .A1(_3835_),
    .A2(_3838_),
    .ZN(_3839_)
  );
  AND2_X1 _6108_ (
    .A1(_0654_),
    .A2(_3839_),
    .ZN(_0590_)
  );
  OR2_X1 _6109_ (
    .A1(large_1[22]),
    .A2(_3833_),
    .ZN(_3840_)
  );
  INV_X1 _6110_ (
    .A(_3840_),
    .ZN(_3841_)
  );
  AND2_X1 _6111_ (
    .A1(large_1[22]),
    .A2(_3833_),
    .ZN(_3842_)
  );
  OR2_X1 _6112_ (
    .A1(_0627_),
    .A2(_3834_),
    .ZN(_3843_)
  );
  OR2_X1 _6113_ (
    .A1(_2670_),
    .A2(_3842_),
    .ZN(_3844_)
  );
  OR2_X1 _6114_ (
    .A1(_3841_),
    .A2(_3844_),
    .ZN(_3845_)
  );
  AND2_X1 _6115_ (
    .A1(large_1[22]),
    .A2(_2660_),
    .ZN(_3846_)
  );
  AND2_X1 _6116_ (
    .A1(_2241_),
    .A2(_2662_),
    .ZN(_3847_)
  );
  OR2_X1 _6117_ (
    .A1(_3846_),
    .A2(_3847_),
    .ZN(_3848_)
  );
  INV_X1 _6118_ (
    .A(_3848_),
    .ZN(_3849_)
  );
  AND2_X1 _6119_ (
    .A1(_3845_),
    .A2(_3849_),
    .ZN(_3850_)
  );
  OR2_X1 _6120_ (
    .A1(reset),
    .A2(_3850_),
    .ZN(_3851_)
  );
  INV_X1 _6121_ (
    .A(_3851_),
    .ZN(_0591_)
  );
  OR2_X1 _6122_ (
    .A1(large_1[23]),
    .A2(_3842_),
    .ZN(_3852_)
  );
  OR2_X1 _6123_ (
    .A1(_0626_),
    .A2(_3843_),
    .ZN(_3853_)
  );
  AND2_X1 _6124_ (
    .A1(_2669_),
    .A2(_3852_),
    .ZN(_3854_)
  );
  AND2_X1 _6125_ (
    .A1(_3853_),
    .A2(_3854_),
    .ZN(_3855_)
  );
  AND2_X1 _6126_ (
    .A1(large_1[23]),
    .A2(_2660_),
    .ZN(_3856_)
  );
  AND2_X1 _6127_ (
    .A1(_2285_),
    .A2(_2662_),
    .ZN(_3857_)
  );
  OR2_X1 _6128_ (
    .A1(_3856_),
    .A2(_3857_),
    .ZN(_3858_)
  );
  OR2_X1 _6129_ (
    .A1(_3855_),
    .A2(_3858_),
    .ZN(_3859_)
  );
  AND2_X1 _6130_ (
    .A1(_0654_),
    .A2(_3859_),
    .ZN(_0592_)
  );
  OR2_X1 _6131_ (
    .A1(large_1[24]),
    .A2(_2653_),
    .ZN(_3860_)
  );
  AND2_X1 _6132_ (
    .A1(_2669_),
    .A2(_3860_),
    .ZN(_3861_)
  );
  AND2_X1 _6133_ (
    .A1(_2656_),
    .A2(_3861_),
    .ZN(_3862_)
  );
  AND2_X1 _6134_ (
    .A1(large_1[24]),
    .A2(_2660_),
    .ZN(_3863_)
  );
  AND2_X1 _6135_ (
    .A1(_2435_),
    .A2(_2662_),
    .ZN(_3864_)
  );
  OR2_X1 _6136_ (
    .A1(_3863_),
    .A2(_3864_),
    .ZN(_3865_)
  );
  OR2_X1 _6137_ (
    .A1(_3862_),
    .A2(_3865_),
    .ZN(_3866_)
  );
  AND2_X1 _6138_ (
    .A1(_0654_),
    .A2(_3866_),
    .ZN(_0593_)
  );
  OR2_X1 _6139_ (
    .A1(large_1[25]),
    .A2(_2655_),
    .ZN(_3867_)
  );
  AND2_X1 _6140_ (
    .A1(_2669_),
    .A2(_3867_),
    .ZN(_3868_)
  );
  AND2_X1 _6141_ (
    .A1(_2658_),
    .A2(_3868_),
    .ZN(_3869_)
  );
  AND2_X1 _6142_ (
    .A1(large_1[25]),
    .A2(_2660_),
    .ZN(_3870_)
  );
  AND2_X1 _6143_ (
    .A1(_2365_),
    .A2(_2667_),
    .ZN(_3871_)
  );
  OR2_X1 _6144_ (
    .A1(_3870_),
    .A2(_3871_),
    .ZN(_3872_)
  );
  OR2_X1 _6145_ (
    .A1(_3869_),
    .A2(_3872_),
    .ZN(_3873_)
  );
  AND2_X1 _6146_ (
    .A1(_0654_),
    .A2(_3873_),
    .ZN(_0594_)
  );
  AND2_X1 _6147_ (
    .A1(large_[0]),
    .A2(_3114_),
    .ZN(_3874_)
  );
  MUX2_X1 _6148_ (
    .A(large_[0]),
    .B(_large_r_T_1[0]),
    .S(_3061_),
    .Z(_3875_)
  );
  AND2_X1 _6149_ (
    .A1(_3122_),
    .A2(_3875_),
    .ZN(_3876_)
  );
  OR2_X1 _6150_ (
    .A1(_3874_),
    .A2(_3876_),
    .ZN(_3877_)
  );
  AND2_X1 _6151_ (
    .A1(_1545_),
    .A2(_3120_),
    .ZN(_3878_)
  );
  OR2_X1 _6152_ (
    .A1(_3877_),
    .A2(_3878_),
    .ZN(_3879_)
  );
  AND2_X1 _6153_ (
    .A1(_0654_),
    .A2(_3879_),
    .ZN(_0595_)
  );
  AND2_X1 _6154_ (
    .A1(large_[0]),
    .A2(_3061_),
    .ZN(_3880_)
  );
  OR2_X1 _6155_ (
    .A1(large_[1]),
    .A2(_3880_),
    .ZN(_3881_)
  );
  AND2_X1 _6156_ (
    .A1(large_[1]),
    .A2(_3114_),
    .ZN(_3882_)
  );
  AND2_X1 _6157_ (
    .A1(_3064_),
    .A2(_3118_),
    .ZN(_3883_)
  );
  OR2_X1 _6158_ (
    .A1(_3882_),
    .A2(_3883_),
    .ZN(_3884_)
  );
  AND2_X1 _6159_ (
    .A1(_3881_),
    .A2(_3884_),
    .ZN(_3885_)
  );
  AND2_X1 _6160_ (
    .A1(_1601_),
    .A2(_3120_),
    .ZN(_3886_)
  );
  OR2_X1 _6161_ (
    .A1(_3885_),
    .A2(_3886_),
    .ZN(_3887_)
  );
  AND2_X1 _6162_ (
    .A1(_0654_),
    .A2(_3887_),
    .ZN(_0596_)
  );
  AND2_X1 _6163_ (
    .A1(large_[2]),
    .A2(_3063_),
    .ZN(_3888_)
  );
  XOR2_X1 _6164_ (
    .A(large_[2]),
    .B(_3063_),
    .Z(_3889_)
  );
  AND2_X1 _6165_ (
    .A1(_3117_),
    .A2(_3889_),
    .ZN(_3890_)
  );
  AND2_X1 _6166_ (
    .A1(large_[2]),
    .A2(_3114_),
    .ZN(_3891_)
  );
  AND2_X1 _6167_ (
    .A1(_0737_),
    .A2(_3889_),
    .ZN(_3892_)
  );
  OR2_X1 _6168_ (
    .A1(_3891_),
    .A2(_3892_),
    .ZN(_3893_)
  );
  OR2_X1 _6169_ (
    .A1(_3890_),
    .A2(_3893_),
    .ZN(_3894_)
  );
  AND2_X1 _6170_ (
    .A1(_1129_),
    .A2(_3120_),
    .ZN(_3895_)
  );
  OR2_X1 _6171_ (
    .A1(_3894_),
    .A2(_3895_),
    .ZN(_3896_)
  );
  AND2_X1 _6172_ (
    .A1(_0654_),
    .A2(_3896_),
    .ZN(_0597_)
  );
  AND2_X1 _6173_ (
    .A1(large_[3]),
    .A2(_3114_),
    .ZN(_3897_)
  );
  AND2_X1 _6174_ (
    .A1(large_[3]),
    .A2(_3888_),
    .ZN(_3898_)
  );
  AND2_X1 _6175_ (
    .A1(_1175_),
    .A2(_3120_),
    .ZN(_3899_)
  );
  XOR2_X1 _6176_ (
    .A(large_[3]),
    .B(_3888_),
    .Z(_3900_)
  );
  AND2_X1 _6177_ (
    .A1(_3122_),
    .A2(_3900_),
    .ZN(_3901_)
  );
  OR2_X1 _6178_ (
    .A1(_3899_),
    .A2(_3901_),
    .ZN(_3902_)
  );
  OR2_X1 _6179_ (
    .A1(_3897_),
    .A2(_3902_),
    .ZN(_3903_)
  );
  AND2_X1 _6180_ (
    .A1(_0654_),
    .A2(_3903_),
    .ZN(_0598_)
  );
  AND2_X1 _6181_ (
    .A1(large_[4]),
    .A2(_3114_),
    .ZN(_3904_)
  );
  AND2_X1 _6182_ (
    .A1(large_[4]),
    .A2(_3898_),
    .ZN(_3905_)
  );
  XOR2_X1 _6183_ (
    .A(large_[4]),
    .B(_3898_),
    .Z(_3906_)
  );
  AND2_X1 _6184_ (
    .A1(_3122_),
    .A2(_3906_),
    .ZN(_3907_)
  );
  OR2_X1 _6185_ (
    .A1(_3904_),
    .A2(_3907_),
    .ZN(_3908_)
  );
  AND2_X1 _6186_ (
    .A1(_1647_),
    .A2(_3120_),
    .ZN(_3909_)
  );
  OR2_X1 _6187_ (
    .A1(_3908_),
    .A2(_3909_),
    .ZN(_3910_)
  );
  AND2_X1 _6188_ (
    .A1(_0654_),
    .A2(_3910_),
    .ZN(_0599_)
  );
  AND2_X1 _6189_ (
    .A1(large_[5]),
    .A2(_3114_),
    .ZN(_3911_)
  );
  AND2_X1 _6190_ (
    .A1(_3065_),
    .A2(_3898_),
    .ZN(_3912_)
  );
  XOR2_X1 _6191_ (
    .A(large_[5]),
    .B(_3905_),
    .Z(_3913_)
  );
  AND2_X1 _6192_ (
    .A1(_1698_),
    .A2(_3120_),
    .ZN(_3914_)
  );
  OR2_X1 _6193_ (
    .A1(_3913_),
    .A2(_3914_),
    .ZN(_3915_)
  );
  AND2_X1 _6194_ (
    .A1(_1698_),
    .A2(_3115_),
    .ZN(_3916_)
  );
  OR2_X1 _6195_ (
    .A1(_3122_),
    .A2(_3916_),
    .ZN(_3917_)
  );
  AND2_X1 _6196_ (
    .A1(_3915_),
    .A2(_3917_),
    .ZN(_3918_)
  );
  OR2_X1 _6197_ (
    .A1(_3911_),
    .A2(_3918_),
    .ZN(_3919_)
  );
  AND2_X1 _6198_ (
    .A1(_0654_),
    .A2(_3919_),
    .ZN(_0600_)
  );
  AND2_X1 _6199_ (
    .A1(large_[6]),
    .A2(_3114_),
    .ZN(_3920_)
  );
  XOR2_X1 _6200_ (
    .A(large_[6]),
    .B(_3912_),
    .Z(_3921_)
  );
  AND2_X1 _6201_ (
    .A1(_1748_),
    .A2(_3120_),
    .ZN(_3922_)
  );
  OR2_X1 _6202_ (
    .A1(_3921_),
    .A2(_3922_),
    .ZN(_3923_)
  );
  AND2_X1 _6203_ (
    .A1(_1748_),
    .A2(_3115_),
    .ZN(_3924_)
  );
  OR2_X1 _6204_ (
    .A1(_3122_),
    .A2(_3924_),
    .ZN(_3925_)
  );
  AND2_X1 _6205_ (
    .A1(_3923_),
    .A2(_3925_),
    .ZN(_3926_)
  );
  OR2_X1 _6206_ (
    .A1(_3920_),
    .A2(_3926_),
    .ZN(_3927_)
  );
  AND2_X1 _6207_ (
    .A1(_0654_),
    .A2(_3927_),
    .ZN(_0601_)
  );
  AND2_X1 _6208_ (
    .A1(large_[7]),
    .A2(_3103_),
    .ZN(_3928_)
  );
  XOR2_X1 _6209_ (
    .A(large_[7]),
    .B(_3103_),
    .Z(_3929_)
  );
  OR2_X1 _6210_ (
    .A1(_0857_),
    .A2(_3929_),
    .ZN(_3930_)
  );
  AND2_X1 _6211_ (
    .A1(_3116_),
    .A2(_3930_),
    .ZN(_3931_)
  );
  OR2_X1 _6212_ (
    .A1(_0858_),
    .A2(_1790_),
    .ZN(_3932_)
  );
  AND2_X1 _6213_ (
    .A1(_3931_),
    .A2(_3932_),
    .ZN(_3933_)
  );
  AND2_X1 _6214_ (
    .A1(_0737_),
    .A2(_3929_),
    .ZN(_3934_)
  );
  AND2_X1 _6215_ (
    .A1(large_[7]),
    .A2(_3114_),
    .ZN(_3935_)
  );
  OR2_X1 _6216_ (
    .A1(_3934_),
    .A2(_3935_),
    .ZN(_3936_)
  );
  OR2_X1 _6217_ (
    .A1(_3933_),
    .A2(_3936_),
    .ZN(_3937_)
  );
  AND2_X1 _6218_ (
    .A1(_0654_),
    .A2(_3937_),
    .ZN(_0602_)
  );
  AND2_X1 _6219_ (
    .A1(large_[8]),
    .A2(_3114_),
    .ZN(_3938_)
  );
  AND2_X1 _6220_ (
    .A1(large_[8]),
    .A2(_3928_),
    .ZN(_3939_)
  );
  XOR2_X1 _6221_ (
    .A(large_[8]),
    .B(_3928_),
    .Z(_3940_)
  );
  AND2_X1 _6222_ (
    .A1(_1832_),
    .A2(_3120_),
    .ZN(_3941_)
  );
  OR2_X1 _6223_ (
    .A1(_3940_),
    .A2(_3941_),
    .ZN(_3942_)
  );
  AND2_X1 _6224_ (
    .A1(_1832_),
    .A2(_3115_),
    .ZN(_3943_)
  );
  OR2_X1 _6225_ (
    .A1(_3122_),
    .A2(_3943_),
    .ZN(_3944_)
  );
  AND2_X1 _6226_ (
    .A1(_3942_),
    .A2(_3944_),
    .ZN(_3945_)
  );
  OR2_X1 _6227_ (
    .A1(_3938_),
    .A2(_3945_),
    .ZN(_3946_)
  );
  AND2_X1 _6228_ (
    .A1(_0654_),
    .A2(_3946_),
    .ZN(_0603_)
  );
  AND2_X1 _6229_ (
    .A1(large_[9]),
    .A2(_3114_),
    .ZN(_3947_)
  );
  XOR2_X1 _6230_ (
    .A(large_[9]),
    .B(_3939_),
    .Z(_3948_)
  );
  AND2_X1 _6231_ (
    .A1(_3122_),
    .A2(_3948_),
    .ZN(_3949_)
  );
  OR2_X1 _6232_ (
    .A1(_3947_),
    .A2(_3949_),
    .ZN(_3950_)
  );
  AND2_X1 _6233_ (
    .A1(_1880_),
    .A2(_3120_),
    .ZN(_3951_)
  );
  OR2_X1 _6234_ (
    .A1(_3950_),
    .A2(_3951_),
    .ZN(_3952_)
  );
  AND2_X1 _6235_ (
    .A1(_0654_),
    .A2(_3952_),
    .ZN(_0604_)
  );
  OR2_X1 _6236_ (
    .A1(large_[10]),
    .A2(_3106_),
    .ZN(_3953_)
  );
  AND2_X1 _6237_ (
    .A1(large_[10]),
    .A2(_3072_),
    .ZN(_3954_)
  );
  INV_X1 _6238_ (
    .A(_3954_),
    .ZN(_3955_)
  );
  AND2_X1 _6239_ (
    .A1(_3118_),
    .A2(_3955_),
    .ZN(_3956_)
  );
  AND2_X1 _6240_ (
    .A1(_3953_),
    .A2(_3956_),
    .ZN(_3957_)
  );
  AND2_X1 _6241_ (
    .A1(large_[10]),
    .A2(_3114_),
    .ZN(_3958_)
  );
  OR2_X1 _6242_ (
    .A1(_3957_),
    .A2(_3958_),
    .ZN(_3959_)
  );
  AND2_X1 _6243_ (
    .A1(_0862_),
    .A2(_3120_),
    .ZN(_3960_)
  );
  OR2_X1 _6244_ (
    .A1(_3959_),
    .A2(_3960_),
    .ZN(_3961_)
  );
  AND2_X1 _6245_ (
    .A1(_0654_),
    .A2(_3961_),
    .ZN(_0605_)
  );
  AND2_X1 _6246_ (
    .A1(_3074_),
    .A2(_3118_),
    .ZN(_3962_)
  );
  OR2_X1 _6247_ (
    .A1(_3114_),
    .A2(_3962_),
    .ZN(_3963_)
  );
  AND2_X1 _6248_ (
    .A1(_3954_),
    .A2(_3962_),
    .ZN(_3964_)
  );
  OR2_X1 _6249_ (
    .A1(large_[11]),
    .A2(_3964_),
    .ZN(_3965_)
  );
  AND2_X1 _6250_ (
    .A1(_3963_),
    .A2(_3965_),
    .ZN(_3966_)
  );
  AND2_X1 _6251_ (
    .A1(_1926_),
    .A2(_3120_),
    .ZN(_3967_)
  );
  OR2_X1 _6252_ (
    .A1(_3966_),
    .A2(_3967_),
    .ZN(_3968_)
  );
  AND2_X1 _6253_ (
    .A1(_0654_),
    .A2(_3968_),
    .ZN(_0606_)
  );
  AND2_X1 _6254_ (
    .A1(_3073_),
    .A2(_3118_),
    .ZN(_3969_)
  );
  MUX2_X1 _6255_ (
    .A(_3969_),
    .B(_3963_),
    .S(large_[12]),
    .Z(_3970_)
  );
  AND2_X1 _6256_ (
    .A1(_0908_),
    .A2(_3120_),
    .ZN(_3971_)
  );
  OR2_X1 _6257_ (
    .A1(_3970_),
    .A2(_3971_),
    .ZN(_3972_)
  );
  AND2_X1 _6258_ (
    .A1(_0654_),
    .A2(_3972_),
    .ZN(_0607_)
  );
  AND2_X1 _6259_ (
    .A1(large_[13]),
    .A2(_3114_),
    .ZN(_3973_)
  );
  XOR2_X1 _6260_ (
    .A(large_[13]),
    .B(_3108_),
    .Z(_3974_)
  );
  AND2_X1 _6261_ (
    .A1(_3122_),
    .A2(_3974_),
    .ZN(_3975_)
  );
  OR2_X1 _6262_ (
    .A1(_3973_),
    .A2(_3975_),
    .ZN(_3976_)
  );
  AND2_X1 _6263_ (
    .A1(_0967_),
    .A2(_3120_),
    .ZN(_3977_)
  );
  OR2_X1 _6264_ (
    .A1(_3976_),
    .A2(_3977_),
    .ZN(_3978_)
  );
  AND2_X1 _6265_ (
    .A1(_0654_),
    .A2(_3978_),
    .ZN(_0608_)
  );
  OR2_X1 _6266_ (
    .A1(large_[14]),
    .A2(_3109_),
    .ZN(_3979_)
  );
  AND2_X1 _6267_ (
    .A1(large_[14]),
    .A2(_3114_),
    .ZN(_3980_)
  );
  AND2_X1 _6268_ (
    .A1(large_[14]),
    .A2(_3077_),
    .ZN(_3981_)
  );
  OR2_X1 _6269_ (
    .A1(_0624_),
    .A2(_3078_),
    .ZN(_3982_)
  );
  AND2_X1 _6270_ (
    .A1(_3122_),
    .A2(_3982_),
    .ZN(_3983_)
  );
  AND2_X1 _6271_ (
    .A1(_3979_),
    .A2(_3983_),
    .ZN(_3984_)
  );
  OR2_X1 _6272_ (
    .A1(_3980_),
    .A2(_3984_),
    .ZN(_3985_)
  );
  AND2_X1 _6273_ (
    .A1(_1017_),
    .A2(_3120_),
    .ZN(_3986_)
  );
  OR2_X1 _6274_ (
    .A1(_3985_),
    .A2(_3986_),
    .ZN(_3987_)
  );
  AND2_X1 _6275_ (
    .A1(_0654_),
    .A2(_3987_),
    .ZN(_0609_)
  );
  OR2_X1 _6276_ (
    .A1(large_[15]),
    .A2(_3981_),
    .ZN(_3988_)
  );
  AND2_X1 _6277_ (
    .A1(large_[15]),
    .A2(_3114_),
    .ZN(_3989_)
  );
  AND2_X1 _6278_ (
    .A1(large_[15]),
    .A2(_3981_),
    .ZN(_3990_)
  );
  OR2_X1 _6279_ (
    .A1(_0623_),
    .A2(_3982_),
    .ZN(_3991_)
  );
  AND2_X1 _6280_ (
    .A1(_3122_),
    .A2(_3988_),
    .ZN(_3992_)
  );
  AND2_X1 _6281_ (
    .A1(_3991_),
    .A2(_3992_),
    .ZN(_3993_)
  );
  OR2_X1 _6282_ (
    .A1(_3989_),
    .A2(_3993_),
    .ZN(_3994_)
  );
  AND2_X1 _6283_ (
    .A1(_1968_),
    .A2(_3120_),
    .ZN(_3995_)
  );
  OR2_X1 _6284_ (
    .A1(_3994_),
    .A2(_3995_),
    .ZN(_3996_)
  );
  AND2_X1 _6285_ (
    .A1(_0654_),
    .A2(_3996_),
    .ZN(_0610_)
  );
  OR2_X1 _6286_ (
    .A1(large_[16]),
    .A2(_3990_),
    .ZN(_3997_)
  );
  AND2_X1 _6287_ (
    .A1(large_[16]),
    .A2(_3990_),
    .ZN(_3998_)
  );
  OR2_X1 _6288_ (
    .A1(_0622_),
    .A2(_3991_),
    .ZN(_3999_)
  );
  AND2_X1 _6289_ (
    .A1(_3122_),
    .A2(_3999_),
    .ZN(_4000_)
  );
  AND2_X1 _6290_ (
    .A1(_3997_),
    .A2(_4000_),
    .ZN(_4001_)
  );
  AND2_X1 _6291_ (
    .A1(large_[16]),
    .A2(_3114_),
    .ZN(_4002_)
  );
  AND2_X1 _6292_ (
    .A1(_2010_),
    .A2(_3120_),
    .ZN(_4003_)
  );
  OR2_X1 _6293_ (
    .A1(_4001_),
    .A2(_4002_),
    .ZN(_4004_)
  );
  OR2_X1 _6294_ (
    .A1(_4003_),
    .A2(_4004_),
    .ZN(_4005_)
  );
  AND2_X1 _6295_ (
    .A1(_0654_),
    .A2(_4005_),
    .ZN(_0611_)
  );
  OR2_X1 _6296_ (
    .A1(large_[17]),
    .A2(_3998_),
    .ZN(_4006_)
  );
  AND2_X1 _6297_ (
    .A1(large_[17]),
    .A2(_3998_),
    .ZN(_4007_)
  );
  INV_X1 _6298_ (
    .A(_4007_),
    .ZN(_4008_)
  );
  AND2_X1 _6299_ (
    .A1(_3122_),
    .A2(_4006_),
    .ZN(_4009_)
  );
  AND2_X1 _6300_ (
    .A1(_4008_),
    .A2(_4009_),
    .ZN(_4010_)
  );
  AND2_X1 _6301_ (
    .A1(large_[17]),
    .A2(_3114_),
    .ZN(_4011_)
  );
  AND2_X1 _6302_ (
    .A1(_1071_),
    .A2(_3120_),
    .ZN(_4012_)
  );
  OR2_X1 _6303_ (
    .A1(_4011_),
    .A2(_4012_),
    .ZN(_4013_)
  );
  OR2_X1 _6304_ (
    .A1(_4010_),
    .A2(_4013_),
    .ZN(_4014_)
  );
  AND2_X1 _6305_ (
    .A1(_0654_),
    .A2(_4014_),
    .ZN(_0612_)
  );
  OR2_X1 _6306_ (
    .A1(large_[18]),
    .A2(_4007_),
    .ZN(_4015_)
  );
  AND2_X1 _6307_ (
    .A1(large_[18]),
    .A2(_4007_),
    .ZN(_4016_)
  );
  INV_X1 _6308_ (
    .A(_4016_),
    .ZN(_4017_)
  );
  AND2_X1 _6309_ (
    .A1(_3122_),
    .A2(_4017_),
    .ZN(_4018_)
  );
  AND2_X1 _6310_ (
    .A1(_4015_),
    .A2(_4018_),
    .ZN(_4019_)
  );
  AND2_X1 _6311_ (
    .A1(large_[18]),
    .A2(_3114_),
    .ZN(_4020_)
  );
  AND2_X1 _6312_ (
    .A1(_2056_),
    .A2(_3120_),
    .ZN(_4021_)
  );
  OR2_X1 _6313_ (
    .A1(_4019_),
    .A2(_4020_),
    .ZN(_4022_)
  );
  OR2_X1 _6314_ (
    .A1(_4021_),
    .A2(_4022_),
    .ZN(_4023_)
  );
  AND2_X1 _6315_ (
    .A1(_0654_),
    .A2(_4023_),
    .ZN(_0613_)
  );
  OR2_X1 _6316_ (
    .A1(large_[19]),
    .A2(_4016_),
    .ZN(_4024_)
  );
  AND2_X1 _6317_ (
    .A1(_3080_),
    .A2(_3118_),
    .ZN(_4025_)
  );
  AND2_X1 _6318_ (
    .A1(_4024_),
    .A2(_4025_),
    .ZN(_4026_)
  );
  AND2_X1 _6319_ (
    .A1(large_[19]),
    .A2(_3114_),
    .ZN(_4027_)
  );
  AND2_X1 _6320_ (
    .A1(_2102_),
    .A2(_3120_),
    .ZN(_4028_)
  );
  OR2_X1 _6321_ (
    .A1(_4027_),
    .A2(_4028_),
    .ZN(_4029_)
  );
  OR2_X1 _6322_ (
    .A1(_4026_),
    .A2(_4029_),
    .ZN(_4030_)
  );
  AND2_X1 _6323_ (
    .A1(_0654_),
    .A2(_4030_),
    .ZN(_0614_)
  );
  OR2_X1 _6324_ (
    .A1(large_[20]),
    .A2(_3110_),
    .ZN(_4031_)
  );
  AND2_X1 _6325_ (
    .A1(_3082_),
    .A2(_3118_),
    .ZN(_4032_)
  );
  AND2_X1 _6326_ (
    .A1(_4031_),
    .A2(_4032_),
    .ZN(_4033_)
  );
  AND2_X1 _6327_ (
    .A1(large_[20]),
    .A2(_3114_),
    .ZN(_4034_)
  );
  AND2_X1 _6328_ (
    .A1(_2148_),
    .A2(_3120_),
    .ZN(_4035_)
  );
  OR2_X1 _6329_ (
    .A1(_4034_),
    .A2(_4035_),
    .ZN(_4036_)
  );
  OR2_X1 _6330_ (
    .A1(_4033_),
    .A2(_4036_),
    .ZN(_4037_)
  );
  AND2_X1 _6331_ (
    .A1(_0654_),
    .A2(_4037_),
    .ZN(_0615_)
  );
  OR2_X1 _6332_ (
    .A1(large_[21]),
    .A2(_3081_),
    .ZN(_4038_)
  );
  AND2_X1 _6333_ (
    .A1(_3122_),
    .A2(_4038_),
    .ZN(_4039_)
  );
  AND2_X1 _6334_ (
    .A1(_3094_),
    .A2(_4039_),
    .ZN(_4040_)
  );
  AND2_X1 _6335_ (
    .A1(large_[21]),
    .A2(_3114_),
    .ZN(_4041_)
  );
  AND2_X1 _6336_ (
    .A1(_2195_),
    .A2(_3120_),
    .ZN(_4042_)
  );
  OR2_X1 _6337_ (
    .A1(_4041_),
    .A2(_4042_),
    .ZN(_4043_)
  );
  OR2_X1 _6338_ (
    .A1(_4040_),
    .A2(_4043_),
    .ZN(_4044_)
  );
  AND2_X1 _6339_ (
    .A1(_0654_),
    .A2(_4044_),
    .ZN(_0616_)
  );
  OR2_X1 _6340_ (
    .A1(large_[22]),
    .A2(_3093_),
    .ZN(_4045_)
  );
  AND2_X1 _6341_ (
    .A1(_3085_),
    .A2(_3118_),
    .ZN(_4046_)
  );
  AND2_X1 _6342_ (
    .A1(_4045_),
    .A2(_4046_),
    .ZN(_4047_)
  );
  AND2_X1 _6343_ (
    .A1(large_[22]),
    .A2(_3114_),
    .ZN(_4048_)
  );
  AND2_X1 _6344_ (
    .A1(_2241_),
    .A2(_3120_),
    .ZN(_4049_)
  );
  OR2_X1 _6345_ (
    .A1(_4048_),
    .A2(_4049_),
    .ZN(_4050_)
  );
  OR2_X1 _6346_ (
    .A1(_4047_),
    .A2(_4050_),
    .ZN(_4051_)
  );
  AND2_X1 _6347_ (
    .A1(_0654_),
    .A2(_4051_),
    .ZN(_0617_)
  );
  OR2_X1 _6348_ (
    .A1(large_[23]),
    .A2(_3084_),
    .ZN(_4052_)
  );
  AND2_X1 _6349_ (
    .A1(_3087_),
    .A2(_3118_),
    .ZN(_4053_)
  );
  AND2_X1 _6350_ (
    .A1(_4052_),
    .A2(_4053_),
    .ZN(_4054_)
  );
  AND2_X1 _6351_ (
    .A1(large_[23]),
    .A2(_3114_),
    .ZN(_4055_)
  );
  AND2_X1 _6352_ (
    .A1(_2285_),
    .A2(_3120_),
    .ZN(_4056_)
  );
  OR2_X1 _6353_ (
    .A1(_4055_),
    .A2(_4056_),
    .ZN(_4057_)
  );
  OR2_X1 _6354_ (
    .A1(_4054_),
    .A2(_4057_),
    .ZN(_4058_)
  );
  AND2_X1 _6355_ (
    .A1(_0654_),
    .A2(_4058_),
    .ZN(_0618_)
  );
  OR2_X1 _6356_ (
    .A1(large_[24]),
    .A2(_3086_),
    .ZN(_4059_)
  );
  AND2_X1 _6357_ (
    .A1(_3089_),
    .A2(_3118_),
    .ZN(_4060_)
  );
  AND2_X1 _6358_ (
    .A1(_4059_),
    .A2(_4060_),
    .ZN(_4061_)
  );
  AND2_X1 _6359_ (
    .A1(large_[24]),
    .A2(_3114_),
    .ZN(_4062_)
  );
  AND2_X1 _6360_ (
    .A1(_2435_),
    .A2(_3120_),
    .ZN(_4063_)
  );
  OR2_X1 _6361_ (
    .A1(_4061_),
    .A2(_4063_),
    .ZN(_4064_)
  );
  OR2_X1 _6362_ (
    .A1(_4062_),
    .A2(_4064_),
    .ZN(_4065_)
  );
  AND2_X1 _6363_ (
    .A1(_0654_),
    .A2(_4065_),
    .ZN(_0619_)
  );
  OR2_X1 _6364_ (
    .A1(large_[25]),
    .A2(_3088_),
    .ZN(_4066_)
  );
  AND2_X1 _6365_ (
    .A1(_3091_),
    .A2(_3118_),
    .ZN(_4067_)
  );
  AND2_X1 _6366_ (
    .A1(_4066_),
    .A2(_4067_),
    .ZN(_4068_)
  );
  AND2_X1 _6367_ (
    .A1(large_[25]),
    .A2(_3114_),
    .ZN(_4069_)
  );
  AND2_X1 _6368_ (
    .A1(_2365_),
    .A2(_3120_),
    .ZN(_4070_)
  );
  OR2_X1 _6369_ (
    .A1(_4068_),
    .A2(_4070_),
    .ZN(_4071_)
  );
  OR2_X1 _6370_ (
    .A1(_4069_),
    .A2(_4071_),
    .ZN(_4072_)
  );
  AND2_X1 _6371_ (
    .A1(_0654_),
    .A2(_4072_),
    .ZN(_0620_)
  );
  MUX2_X1 _6372_ (
    .A(reg_pmp_6_cfg_w),
    .B(_2327_),
    .S(_0740_),
    .Z(_0621_)
  );
  AND2_X1 _6373_ (
    .A1(io_decode_0_inst[31]),
    .A2(io_decode_0_inst[30]),
    .ZN(io_decode_0_write_illegal)
  );
  OR2_X1 _6374_ (
    .A1(_0737_),
    .A2(_0751_),
    .ZN(_4073_)
  );
  OR2_X1 _6375_ (
    .A1(reg_debug),
    .A2(_2469_),
    .ZN(_4074_)
  );
  OR2_X1 _6376_ (
    .A1(_2505_),
    .A2(_4074_),
    .ZN(_4075_)
  );
  MUX2_X1 _6377_ (
    .A(io_pc[1]),
    .B(reg_dpc[1]),
    .S(_4075_),
    .Z(_4076_)
  );
  MUX2_X1 _6378_ (
    .A(_1290_),
    .B(_4076_),
    .S(_4073_),
    .Z(_0000_[1])
  );
  MUX2_X1 _6379_ (
    .A(io_pc[2]),
    .B(reg_dpc[2]),
    .S(_4075_),
    .Z(_4077_)
  );
  MUX2_X1 _6380_ (
    .A(_1346_),
    .B(_4077_),
    .S(_4073_),
    .Z(_0000_[2])
  );
  MUX2_X1 _6381_ (
    .A(io_pc[3]),
    .B(reg_dpc[3]),
    .S(_4075_),
    .Z(_4078_)
  );
  MUX2_X1 _6382_ (
    .A(_1409_),
    .B(_4078_),
    .S(_4073_),
    .Z(_0000_[3])
  );
  MUX2_X1 _6383_ (
    .A(io_pc[4]),
    .B(reg_dpc[4]),
    .S(_4075_),
    .Z(_4079_)
  );
  MUX2_X1 _6384_ (
    .A(_1456_),
    .B(_4079_),
    .S(_4073_),
    .Z(_0000_[4])
  );
  MUX2_X1 _6385_ (
    .A(io_pc[5]),
    .B(reg_dpc[5]),
    .S(_4075_),
    .Z(_4080_)
  );
  MUX2_X1 _6386_ (
    .A(_1499_),
    .B(_4080_),
    .S(_4073_),
    .Z(_0000_[5])
  );
  MUX2_X1 _6387_ (
    .A(io_pc[6]),
    .B(reg_dpc[6]),
    .S(_4075_),
    .Z(_4081_)
  );
  MUX2_X1 _6388_ (
    .A(_1545_),
    .B(_4081_),
    .S(_4073_),
    .Z(_0000_[6])
  );
  MUX2_X1 _6389_ (
    .A(io_pc[7]),
    .B(reg_dpc[7]),
    .S(_4075_),
    .Z(_4082_)
  );
  MUX2_X1 _6390_ (
    .A(_1601_),
    .B(_4082_),
    .S(_4073_),
    .Z(_0000_[7])
  );
  MUX2_X1 _6391_ (
    .A(io_pc[8]),
    .B(reg_dpc[8]),
    .S(_4075_),
    .Z(_4083_)
  );
  MUX2_X1 _6392_ (
    .A(_1129_),
    .B(_4083_),
    .S(_4073_),
    .Z(_0000_[8])
  );
  MUX2_X1 _6393_ (
    .A(io_pc[9]),
    .B(reg_dpc[9]),
    .S(_4075_),
    .Z(_4084_)
  );
  MUX2_X1 _6394_ (
    .A(_1175_),
    .B(_4084_),
    .S(_4073_),
    .Z(_0000_[9])
  );
  MUX2_X1 _6395_ (
    .A(io_pc[10]),
    .B(reg_dpc[10]),
    .S(_4075_),
    .Z(_4085_)
  );
  MUX2_X1 _6396_ (
    .A(_1647_),
    .B(_4085_),
    .S(_4073_),
    .Z(_0000_[10])
  );
  MUX2_X1 _6397_ (
    .A(io_pc[11]),
    .B(reg_dpc[11]),
    .S(_4075_),
    .Z(_4086_)
  );
  MUX2_X1 _6398_ (
    .A(_1698_),
    .B(_4086_),
    .S(_4073_),
    .Z(_0000_[11])
  );
  MUX2_X1 _6399_ (
    .A(io_pc[12]),
    .B(reg_dpc[12]),
    .S(_4075_),
    .Z(_4087_)
  );
  MUX2_X1 _6400_ (
    .A(_1748_),
    .B(_4087_),
    .S(_4073_),
    .Z(_0000_[12])
  );
  MUX2_X1 _6401_ (
    .A(io_pc[13]),
    .B(reg_dpc[13]),
    .S(_4075_),
    .Z(_4088_)
  );
  MUX2_X1 _6402_ (
    .A(_1790_),
    .B(_4088_),
    .S(_4073_),
    .Z(_0000_[13])
  );
  MUX2_X1 _6403_ (
    .A(io_pc[14]),
    .B(reg_dpc[14]),
    .S(_4075_),
    .Z(_4089_)
  );
  MUX2_X1 _6404_ (
    .A(_1832_),
    .B(_4089_),
    .S(_4073_),
    .Z(_0000_[14])
  );
  MUX2_X1 _6405_ (
    .A(io_pc[15]),
    .B(reg_dpc[15]),
    .S(_4075_),
    .Z(_4090_)
  );
  MUX2_X1 _6406_ (
    .A(_1880_),
    .B(_4090_),
    .S(_4073_),
    .Z(_0000_[15])
  );
  MUX2_X1 _6407_ (
    .A(io_pc[16]),
    .B(reg_dpc[16]),
    .S(_4075_),
    .Z(_4091_)
  );
  MUX2_X1 _6408_ (
    .A(_0862_),
    .B(_4091_),
    .S(_4073_),
    .Z(_0000_[16])
  );
  MUX2_X1 _6409_ (
    .A(io_pc[17]),
    .B(reg_dpc[17]),
    .S(_4075_),
    .Z(_4092_)
  );
  MUX2_X1 _6410_ (
    .A(_1926_),
    .B(_4092_),
    .S(_4073_),
    .Z(_0000_[17])
  );
  MUX2_X1 _6411_ (
    .A(io_pc[18]),
    .B(reg_dpc[18]),
    .S(_4075_),
    .Z(_4093_)
  );
  MUX2_X1 _6412_ (
    .A(_0908_),
    .B(_4093_),
    .S(_4073_),
    .Z(_0000_[18])
  );
  MUX2_X1 _6413_ (
    .A(io_pc[19]),
    .B(reg_dpc[19]),
    .S(_4075_),
    .Z(_4094_)
  );
  MUX2_X1 _6414_ (
    .A(_0967_),
    .B(_4094_),
    .S(_4073_),
    .Z(_0000_[19])
  );
  MUX2_X1 _6415_ (
    .A(io_pc[20]),
    .B(reg_dpc[20]),
    .S(_4075_),
    .Z(_4095_)
  );
  MUX2_X1 _6416_ (
    .A(_1017_),
    .B(_4095_),
    .S(_4073_),
    .Z(_0000_[20])
  );
  MUX2_X1 _6417_ (
    .A(io_pc[21]),
    .B(reg_dpc[21]),
    .S(_4075_),
    .Z(_4096_)
  );
  MUX2_X1 _6418_ (
    .A(_1968_),
    .B(_4096_),
    .S(_4073_),
    .Z(_0000_[21])
  );
  MUX2_X1 _6419_ (
    .A(io_pc[22]),
    .B(reg_dpc[22]),
    .S(_4075_),
    .Z(_4097_)
  );
  MUX2_X1 _6420_ (
    .A(_2010_),
    .B(_4097_),
    .S(_4073_),
    .Z(_0000_[22])
  );
  MUX2_X1 _6421_ (
    .A(io_pc[23]),
    .B(reg_dpc[23]),
    .S(_4075_),
    .Z(_4098_)
  );
  MUX2_X1 _6422_ (
    .A(_1071_),
    .B(_4098_),
    .S(_4073_),
    .Z(_0000_[23])
  );
  MUX2_X1 _6423_ (
    .A(io_pc[24]),
    .B(reg_dpc[24]),
    .S(_4075_),
    .Z(_4099_)
  );
  MUX2_X1 _6424_ (
    .A(_2056_),
    .B(_4099_),
    .S(_4073_),
    .Z(_0000_[24])
  );
  MUX2_X1 _6425_ (
    .A(io_pc[25]),
    .B(reg_dpc[25]),
    .S(_4075_),
    .Z(_4100_)
  );
  MUX2_X1 _6426_ (
    .A(_2102_),
    .B(_4100_),
    .S(_4073_),
    .Z(_0000_[25])
  );
  MUX2_X1 _6427_ (
    .A(io_pc[26]),
    .B(reg_dpc[26]),
    .S(_4075_),
    .Z(_4101_)
  );
  MUX2_X1 _6428_ (
    .A(_2148_),
    .B(_4101_),
    .S(_4073_),
    .Z(_0000_[26])
  );
  MUX2_X1 _6429_ (
    .A(io_pc[27]),
    .B(reg_dpc[27]),
    .S(_4075_),
    .Z(_4102_)
  );
  MUX2_X1 _6430_ (
    .A(_2195_),
    .B(_4102_),
    .S(_4073_),
    .Z(_0000_[27])
  );
  MUX2_X1 _6431_ (
    .A(io_pc[28]),
    .B(reg_dpc[28]),
    .S(_4075_),
    .Z(_4103_)
  );
  MUX2_X1 _6432_ (
    .A(_2241_),
    .B(_4103_),
    .S(_4073_),
    .Z(_0000_[28])
  );
  MUX2_X1 _6433_ (
    .A(io_pc[29]),
    .B(reg_dpc[29]),
    .S(_4075_),
    .Z(_4104_)
  );
  MUX2_X1 _6434_ (
    .A(_2285_),
    .B(_4104_),
    .S(_4073_),
    .Z(_0000_[29])
  );
  MUX2_X1 _6435_ (
    .A(io_pc[30]),
    .B(reg_dpc[30]),
    .S(_4075_),
    .Z(_4105_)
  );
  MUX2_X1 _6436_ (
    .A(_2435_),
    .B(_4105_),
    .S(_4073_),
    .Z(_0000_[30])
  );
  MUX2_X1 _6437_ (
    .A(io_pc[31]),
    .B(reg_dpc[31]),
    .S(_4075_),
    .Z(_4106_)
  );
  MUX2_X1 _6438_ (
    .A(_2365_),
    .B(_4106_),
    .S(_4073_),
    .Z(_0000_[31])
  );
  OR2_X1 _6439_ (
    .A1(_0737_),
    .A2(_0784_),
    .ZN(_4107_)
  );
  MUX2_X1 _6440_ (
    .A(io_pc[1]),
    .B(reg_mepc[1]),
    .S(_2507_),
    .Z(_4108_)
  );
  MUX2_X1 _6441_ (
    .A(_1290_),
    .B(_4108_),
    .S(_4107_),
    .Z(_0001_[1])
  );
  MUX2_X1 _6442_ (
    .A(io_pc[2]),
    .B(reg_mepc[2]),
    .S(_2507_),
    .Z(_4109_)
  );
  MUX2_X1 _6443_ (
    .A(_1346_),
    .B(_4109_),
    .S(_4107_),
    .Z(_0001_[2])
  );
  MUX2_X1 _6444_ (
    .A(io_pc[3]),
    .B(reg_mepc[3]),
    .S(_2507_),
    .Z(_4110_)
  );
  MUX2_X1 _6445_ (
    .A(_1409_),
    .B(_4110_),
    .S(_4107_),
    .Z(_0001_[3])
  );
  MUX2_X1 _6446_ (
    .A(io_pc[4]),
    .B(reg_mepc[4]),
    .S(_2507_),
    .Z(_4111_)
  );
  MUX2_X1 _6447_ (
    .A(_1456_),
    .B(_4111_),
    .S(_4107_),
    .Z(_0001_[4])
  );
  MUX2_X1 _6448_ (
    .A(io_pc[5]),
    .B(reg_mepc[5]),
    .S(_2507_),
    .Z(_4112_)
  );
  MUX2_X1 _6449_ (
    .A(_1499_),
    .B(_4112_),
    .S(_4107_),
    .Z(_0001_[5])
  );
  MUX2_X1 _6450_ (
    .A(io_pc[6]),
    .B(reg_mepc[6]),
    .S(_2507_),
    .Z(_4113_)
  );
  MUX2_X1 _6451_ (
    .A(_1545_),
    .B(_4113_),
    .S(_4107_),
    .Z(_0001_[6])
  );
  MUX2_X1 _6452_ (
    .A(io_pc[7]),
    .B(reg_mepc[7]),
    .S(_2507_),
    .Z(_4114_)
  );
  MUX2_X1 _6453_ (
    .A(_1601_),
    .B(_4114_),
    .S(_4107_),
    .Z(_0001_[7])
  );
  MUX2_X1 _6454_ (
    .A(io_pc[8]),
    .B(reg_mepc[8]),
    .S(_2507_),
    .Z(_4115_)
  );
  MUX2_X1 _6455_ (
    .A(_1129_),
    .B(_4115_),
    .S(_4107_),
    .Z(_0001_[8])
  );
  MUX2_X1 _6456_ (
    .A(io_pc[9]),
    .B(reg_mepc[9]),
    .S(_2507_),
    .Z(_4116_)
  );
  MUX2_X1 _6457_ (
    .A(_1175_),
    .B(_4116_),
    .S(_4107_),
    .Z(_0001_[9])
  );
  MUX2_X1 _6458_ (
    .A(io_pc[10]),
    .B(reg_mepc[10]),
    .S(_2507_),
    .Z(_4117_)
  );
  MUX2_X1 _6459_ (
    .A(_1647_),
    .B(_4117_),
    .S(_4107_),
    .Z(_0001_[10])
  );
  MUX2_X1 _6460_ (
    .A(io_pc[11]),
    .B(reg_mepc[11]),
    .S(_2507_),
    .Z(_4118_)
  );
  MUX2_X1 _6461_ (
    .A(_1698_),
    .B(_4118_),
    .S(_4107_),
    .Z(_0001_[11])
  );
  MUX2_X1 _6462_ (
    .A(io_pc[12]),
    .B(reg_mepc[12]),
    .S(_2507_),
    .Z(_4119_)
  );
  MUX2_X1 _6463_ (
    .A(_1748_),
    .B(_4119_),
    .S(_4107_),
    .Z(_0001_[12])
  );
  MUX2_X1 _6464_ (
    .A(io_pc[13]),
    .B(reg_mepc[13]),
    .S(_2507_),
    .Z(_4120_)
  );
  MUX2_X1 _6465_ (
    .A(_1790_),
    .B(_4120_),
    .S(_4107_),
    .Z(_0001_[13])
  );
  MUX2_X1 _6466_ (
    .A(io_pc[14]),
    .B(reg_mepc[14]),
    .S(_2507_),
    .Z(_4121_)
  );
  MUX2_X1 _6467_ (
    .A(_1832_),
    .B(_4121_),
    .S(_4107_),
    .Z(_0001_[14])
  );
  MUX2_X1 _6468_ (
    .A(io_pc[15]),
    .B(reg_mepc[15]),
    .S(_2507_),
    .Z(_4122_)
  );
  MUX2_X1 _6469_ (
    .A(_1880_),
    .B(_4122_),
    .S(_4107_),
    .Z(_0001_[15])
  );
  MUX2_X1 _6470_ (
    .A(io_pc[16]),
    .B(reg_mepc[16]),
    .S(_2507_),
    .Z(_4123_)
  );
  MUX2_X1 _6471_ (
    .A(_0862_),
    .B(_4123_),
    .S(_4107_),
    .Z(_0001_[16])
  );
  MUX2_X1 _6472_ (
    .A(io_pc[17]),
    .B(reg_mepc[17]),
    .S(_2507_),
    .Z(_4124_)
  );
  MUX2_X1 _6473_ (
    .A(_1926_),
    .B(_4124_),
    .S(_4107_),
    .Z(_0001_[17])
  );
  MUX2_X1 _6474_ (
    .A(io_pc[18]),
    .B(reg_mepc[18]),
    .S(_2507_),
    .Z(_4125_)
  );
  MUX2_X1 _6475_ (
    .A(_0908_),
    .B(_4125_),
    .S(_4107_),
    .Z(_0001_[18])
  );
  MUX2_X1 _6476_ (
    .A(io_pc[19]),
    .B(reg_mepc[19]),
    .S(_2507_),
    .Z(_4126_)
  );
  MUX2_X1 _6477_ (
    .A(_0967_),
    .B(_4126_),
    .S(_4107_),
    .Z(_0001_[19])
  );
  MUX2_X1 _6478_ (
    .A(io_pc[20]),
    .B(reg_mepc[20]),
    .S(_2507_),
    .Z(_4127_)
  );
  MUX2_X1 _6479_ (
    .A(_1017_),
    .B(_4127_),
    .S(_4107_),
    .Z(_0001_[20])
  );
  MUX2_X1 _6480_ (
    .A(io_pc[21]),
    .B(reg_mepc[21]),
    .S(_2507_),
    .Z(_4128_)
  );
  MUX2_X1 _6481_ (
    .A(_1968_),
    .B(_4128_),
    .S(_4107_),
    .Z(_0001_[21])
  );
  MUX2_X1 _6482_ (
    .A(io_pc[22]),
    .B(reg_mepc[22]),
    .S(_2507_),
    .Z(_4129_)
  );
  MUX2_X1 _6483_ (
    .A(_2010_),
    .B(_4129_),
    .S(_4107_),
    .Z(_0001_[22])
  );
  MUX2_X1 _6484_ (
    .A(io_pc[23]),
    .B(reg_mepc[23]),
    .S(_2507_),
    .Z(_4130_)
  );
  MUX2_X1 _6485_ (
    .A(_1071_),
    .B(_4130_),
    .S(_4107_),
    .Z(_0001_[23])
  );
  MUX2_X1 _6486_ (
    .A(io_pc[24]),
    .B(reg_mepc[24]),
    .S(_2507_),
    .Z(_4131_)
  );
  MUX2_X1 _6487_ (
    .A(_2056_),
    .B(_4131_),
    .S(_4107_),
    .Z(_0001_[24])
  );
  MUX2_X1 _6488_ (
    .A(io_pc[25]),
    .B(reg_mepc[25]),
    .S(_2507_),
    .Z(_4132_)
  );
  MUX2_X1 _6489_ (
    .A(_2102_),
    .B(_4132_),
    .S(_4107_),
    .Z(_0001_[25])
  );
  MUX2_X1 _6490_ (
    .A(io_pc[26]),
    .B(reg_mepc[26]),
    .S(_2507_),
    .Z(_4133_)
  );
  MUX2_X1 _6491_ (
    .A(_2148_),
    .B(_4133_),
    .S(_4107_),
    .Z(_0001_[26])
  );
  MUX2_X1 _6492_ (
    .A(io_pc[27]),
    .B(reg_mepc[27]),
    .S(_2507_),
    .Z(_4134_)
  );
  MUX2_X1 _6493_ (
    .A(_2195_),
    .B(_4134_),
    .S(_4107_),
    .Z(_0001_[27])
  );
  MUX2_X1 _6494_ (
    .A(io_pc[28]),
    .B(reg_mepc[28]),
    .S(_2507_),
    .Z(_4135_)
  );
  MUX2_X1 _6495_ (
    .A(_2241_),
    .B(_4135_),
    .S(_4107_),
    .Z(_0001_[28])
  );
  MUX2_X1 _6496_ (
    .A(io_pc[29]),
    .B(reg_mepc[29]),
    .S(_2507_),
    .Z(_4136_)
  );
  MUX2_X1 _6497_ (
    .A(_2285_),
    .B(_4136_),
    .S(_4107_),
    .Z(_0001_[29])
  );
  MUX2_X1 _6498_ (
    .A(io_pc[30]),
    .B(reg_mepc[30]),
    .S(_2507_),
    .Z(_4137_)
  );
  MUX2_X1 _6499_ (
    .A(_2435_),
    .B(_4137_),
    .S(_4107_),
    .Z(_0001_[30])
  );
  MUX2_X1 _6500_ (
    .A(io_pc[31]),
    .B(reg_mepc[31]),
    .S(_2507_),
    .Z(_4138_)
  );
  MUX2_X1 _6501_ (
    .A(_2365_),
    .B(_4138_),
    .S(_4107_),
    .Z(_0001_[31])
  );
  OR2_X1 _6502_ (
    .A1(_0737_),
    .A2(_0765_),
    .ZN(_4139_)
  );
  MUX2_X1 _6503_ (
    .A(io_tval[0]),
    .B(reg_mtval[0]),
    .S(_2507_),
    .Z(_4140_)
  );
  MUX2_X1 _6504_ (
    .A(_1241_),
    .B(_4140_),
    .S(_4139_),
    .Z(_0002_[0])
  );
  MUX2_X1 _6505_ (
    .A(io_tval[1]),
    .B(reg_mtval[1]),
    .S(_2507_),
    .Z(_4141_)
  );
  MUX2_X1 _6506_ (
    .A(_1290_),
    .B(_4141_),
    .S(_4139_),
    .Z(_0002_[1])
  );
  MUX2_X1 _6507_ (
    .A(io_tval[2]),
    .B(reg_mtval[2]),
    .S(_2507_),
    .Z(_4142_)
  );
  MUX2_X1 _6508_ (
    .A(_1346_),
    .B(_4142_),
    .S(_4139_),
    .Z(_0002_[2])
  );
  MUX2_X1 _6509_ (
    .A(io_tval[3]),
    .B(reg_mtval[3]),
    .S(_2507_),
    .Z(_4143_)
  );
  MUX2_X1 _6510_ (
    .A(_1409_),
    .B(_4143_),
    .S(_4139_),
    .Z(_0002_[3])
  );
  MUX2_X1 _6511_ (
    .A(io_tval[4]),
    .B(reg_mtval[4]),
    .S(_2507_),
    .Z(_4144_)
  );
  MUX2_X1 _6512_ (
    .A(_1456_),
    .B(_4144_),
    .S(_4139_),
    .Z(_0002_[4])
  );
  MUX2_X1 _6513_ (
    .A(io_tval[5]),
    .B(reg_mtval[5]),
    .S(_2507_),
    .Z(_4145_)
  );
  MUX2_X1 _6514_ (
    .A(_1499_),
    .B(_4145_),
    .S(_4139_),
    .Z(_0002_[5])
  );
  MUX2_X1 _6515_ (
    .A(io_tval[6]),
    .B(reg_mtval[6]),
    .S(_2507_),
    .Z(_4146_)
  );
  MUX2_X1 _6516_ (
    .A(_1545_),
    .B(_4146_),
    .S(_4139_),
    .Z(_0002_[6])
  );
  MUX2_X1 _6517_ (
    .A(io_tval[7]),
    .B(reg_mtval[7]),
    .S(_2507_),
    .Z(_4147_)
  );
  MUX2_X1 _6518_ (
    .A(_1601_),
    .B(_4147_),
    .S(_4139_),
    .Z(_0002_[7])
  );
  MUX2_X1 _6519_ (
    .A(io_tval[8]),
    .B(reg_mtval[8]),
    .S(_2507_),
    .Z(_4148_)
  );
  MUX2_X1 _6520_ (
    .A(_1129_),
    .B(_4148_),
    .S(_4139_),
    .Z(_0002_[8])
  );
  MUX2_X1 _6521_ (
    .A(io_tval[9]),
    .B(reg_mtval[9]),
    .S(_2507_),
    .Z(_4149_)
  );
  MUX2_X1 _6522_ (
    .A(_1175_),
    .B(_4149_),
    .S(_4139_),
    .Z(_0002_[9])
  );
  MUX2_X1 _6523_ (
    .A(io_tval[10]),
    .B(reg_mtval[10]),
    .S(_2507_),
    .Z(_4150_)
  );
  MUX2_X1 _6524_ (
    .A(_1647_),
    .B(_4150_),
    .S(_4139_),
    .Z(_0002_[10])
  );
  MUX2_X1 _6525_ (
    .A(io_tval[11]),
    .B(reg_mtval[11]),
    .S(_2507_),
    .Z(_4151_)
  );
  MUX2_X1 _6526_ (
    .A(_1698_),
    .B(_4151_),
    .S(_4139_),
    .Z(_0002_[11])
  );
  MUX2_X1 _6527_ (
    .A(io_tval[12]),
    .B(reg_mtval[12]),
    .S(_2507_),
    .Z(_4152_)
  );
  MUX2_X1 _6528_ (
    .A(_1748_),
    .B(_4152_),
    .S(_4139_),
    .Z(_0002_[12])
  );
  MUX2_X1 _6529_ (
    .A(io_tval[13]),
    .B(reg_mtval[13]),
    .S(_2507_),
    .Z(_4153_)
  );
  MUX2_X1 _6530_ (
    .A(_1790_),
    .B(_4153_),
    .S(_4139_),
    .Z(_0002_[13])
  );
  MUX2_X1 _6531_ (
    .A(io_tval[14]),
    .B(reg_mtval[14]),
    .S(_2507_),
    .Z(_4154_)
  );
  MUX2_X1 _6532_ (
    .A(_1832_),
    .B(_4154_),
    .S(_4139_),
    .Z(_0002_[14])
  );
  MUX2_X1 _6533_ (
    .A(io_tval[15]),
    .B(reg_mtval[15]),
    .S(_2507_),
    .Z(_4155_)
  );
  MUX2_X1 _6534_ (
    .A(_1880_),
    .B(_4155_),
    .S(_4139_),
    .Z(_0002_[15])
  );
  MUX2_X1 _6535_ (
    .A(io_tval[16]),
    .B(reg_mtval[16]),
    .S(_2507_),
    .Z(_4156_)
  );
  MUX2_X1 _6536_ (
    .A(_0862_),
    .B(_4156_),
    .S(_4139_),
    .Z(_0002_[16])
  );
  MUX2_X1 _6537_ (
    .A(io_tval[17]),
    .B(reg_mtval[17]),
    .S(_2507_),
    .Z(_4157_)
  );
  MUX2_X1 _6538_ (
    .A(_1926_),
    .B(_4157_),
    .S(_4139_),
    .Z(_0002_[17])
  );
  MUX2_X1 _6539_ (
    .A(io_tval[18]),
    .B(reg_mtval[18]),
    .S(_2507_),
    .Z(_4158_)
  );
  MUX2_X1 _6540_ (
    .A(_0908_),
    .B(_4158_),
    .S(_4139_),
    .Z(_0002_[18])
  );
  MUX2_X1 _6541_ (
    .A(io_tval[19]),
    .B(reg_mtval[19]),
    .S(_2507_),
    .Z(_4159_)
  );
  MUX2_X1 _6542_ (
    .A(_0967_),
    .B(_4159_),
    .S(_4139_),
    .Z(_0002_[19])
  );
  MUX2_X1 _6543_ (
    .A(io_tval[20]),
    .B(reg_mtval[20]),
    .S(_2507_),
    .Z(_4160_)
  );
  MUX2_X1 _6544_ (
    .A(_1017_),
    .B(_4160_),
    .S(_4139_),
    .Z(_0002_[20])
  );
  MUX2_X1 _6545_ (
    .A(io_tval[21]),
    .B(reg_mtval[21]),
    .S(_2507_),
    .Z(_4161_)
  );
  MUX2_X1 _6546_ (
    .A(_1968_),
    .B(_4161_),
    .S(_4139_),
    .Z(_0002_[21])
  );
  MUX2_X1 _6547_ (
    .A(io_tval[22]),
    .B(reg_mtval[22]),
    .S(_2507_),
    .Z(_4162_)
  );
  MUX2_X1 _6548_ (
    .A(_2010_),
    .B(_4162_),
    .S(_4139_),
    .Z(_0002_[22])
  );
  MUX2_X1 _6549_ (
    .A(io_tval[23]),
    .B(reg_mtval[23]),
    .S(_2507_),
    .Z(_4163_)
  );
  MUX2_X1 _6550_ (
    .A(_1071_),
    .B(_4163_),
    .S(_4139_),
    .Z(_0002_[23])
  );
  MUX2_X1 _6551_ (
    .A(io_tval[24]),
    .B(reg_mtval[24]),
    .S(_2507_),
    .Z(_4164_)
  );
  MUX2_X1 _6552_ (
    .A(_2056_),
    .B(_4164_),
    .S(_4139_),
    .Z(_0002_[24])
  );
  MUX2_X1 _6553_ (
    .A(io_tval[25]),
    .B(reg_mtval[25]),
    .S(_2507_),
    .Z(_4165_)
  );
  MUX2_X1 _6554_ (
    .A(_2102_),
    .B(_4165_),
    .S(_4139_),
    .Z(_0002_[25])
  );
  MUX2_X1 _6555_ (
    .A(io_tval[26]),
    .B(reg_mtval[26]),
    .S(_2507_),
    .Z(_4166_)
  );
  MUX2_X1 _6556_ (
    .A(_2148_),
    .B(_4166_),
    .S(_4139_),
    .Z(_0002_[26])
  );
  MUX2_X1 _6557_ (
    .A(io_tval[27]),
    .B(reg_mtval[27]),
    .S(_2507_),
    .Z(_4167_)
  );
  MUX2_X1 _6558_ (
    .A(_2195_),
    .B(_4167_),
    .S(_4139_),
    .Z(_0002_[27])
  );
  MUX2_X1 _6559_ (
    .A(io_tval[28]),
    .B(reg_mtval[28]),
    .S(_2507_),
    .Z(_4168_)
  );
  MUX2_X1 _6560_ (
    .A(_2241_),
    .B(_4168_),
    .S(_4139_),
    .Z(_0002_[28])
  );
  MUX2_X1 _6561_ (
    .A(io_tval[29]),
    .B(reg_mtval[29]),
    .S(_2507_),
    .Z(_4169_)
  );
  MUX2_X1 _6562_ (
    .A(_2285_),
    .B(_4169_),
    .S(_4139_),
    .Z(_0002_[29])
  );
  MUX2_X1 _6563_ (
    .A(io_tval[30]),
    .B(reg_mtval[30]),
    .S(_2507_),
    .Z(_4170_)
  );
  MUX2_X1 _6564_ (
    .A(_2435_),
    .B(_4170_),
    .S(_4139_),
    .Z(_0002_[30])
  );
  MUX2_X1 _6565_ (
    .A(io_tval[31]),
    .B(reg_mtval[31]),
    .S(_2507_),
    .Z(_4171_)
  );
  MUX2_X1 _6566_ (
    .A(_2365_),
    .B(_4171_),
    .S(_4139_),
    .Z(_0002_[31])
  );
  AND2_X1 _6567_ (
    .A1(reg_mstatus_mie),
    .A2(_0677_),
    .ZN(_4172_)
  );
  OR2_X1 _6568_ (
    .A1(_0676_),
    .A2(io_interrupts_debug),
    .ZN(_4173_)
  );
  AND2_X1 _6569_ (
    .A1(_2575_),
    .A2(_4172_),
    .ZN(io_interrupt_cause[0])
  );
  OR2_X1 _6570_ (
    .A1(io_interrupts_debug),
    .A2(io_interrupt_cause[0]),
    .ZN(io_interrupt_cause[1])
  );
  OR2_X1 _6571_ (
    .A1(_2574_),
    .A2(_4173_),
    .ZN(io_interrupt_cause[2])
  );
  AND2_X1 _6572_ (
    .A1(reg_mstatus_mie),
    .A2(_2572_),
    .ZN(_4174_)
  );
  OR2_X1 _6573_ (
    .A1(io_interrupts_debug),
    .A2(_4174_),
    .ZN(io_interrupt_cause[3])
  );
  AND2_X1 _6574_ (
    .A1(_1260_),
    .A2(_2519_),
    .ZN(_4175_)
  );
  AND2_X1 _6575_ (
    .A1(_1252_),
    .A2(_2515_),
    .ZN(_4176_)
  );
  OR2_X1 _6576_ (
    .A1(_4175_),
    .A2(_4176_),
    .ZN(io_evec[1])
  );
  AND2_X1 _6577_ (
    .A1(_2505_),
    .A2(_2511_),
    .ZN(_4177_)
  );
  AND2_X1 _6578_ (
    .A1(reg_mtvec[0]),
    .A2(_2539_),
    .ZN(_4178_)
  );
  AND2_X1 _6579_ (
    .A1(_2489_),
    .A2(_4178_),
    .ZN(_4179_)
  );
  MUX2_X1 _6580_ (
    .A(_1308_),
    .B(io_cause[0]),
    .S(_4179_),
    .Z(_4180_)
  );
  AND2_X1 _6581_ (
    .A1(_4177_),
    .A2(_4180_),
    .ZN(_4181_)
  );
  AND2_X1 _6582_ (
    .A1(reg_mepc[2]),
    .A2(_2519_),
    .ZN(_4182_)
  );
  AND2_X1 _6583_ (
    .A1(reg_dpc[2]),
    .A2(_2515_),
    .ZN(_4183_)
  );
  OR2_X1 _6584_ (
    .A1(_4182_),
    .A2(_4183_),
    .ZN(_4184_)
  );
  OR2_X1 _6585_ (
    .A1(_4181_),
    .A2(_4184_),
    .ZN(io_evec[2])
  );
  AND2_X1 _6586_ (
    .A1(reg_debug),
    .A2(_2465_),
    .ZN(_4185_)
  );
  MUX2_X1 _6587_ (
    .A(_1397_),
    .B(io_cause[1]),
    .S(_4179_),
    .Z(_4186_)
  );
  AND2_X1 _6588_ (
    .A1(_2505_),
    .A2(_4186_),
    .ZN(_4187_)
  );
  OR2_X1 _6589_ (
    .A1(_4185_),
    .A2(_4187_),
    .ZN(_4188_)
  );
  AND2_X1 _6590_ (
    .A1(_2511_),
    .A2(_4188_),
    .ZN(_4189_)
  );
  AND2_X1 _6591_ (
    .A1(reg_dpc[3]),
    .A2(_2515_),
    .ZN(_4190_)
  );
  AND2_X1 _6592_ (
    .A1(reg_mepc[3]),
    .A2(_2519_),
    .ZN(_4191_)
  );
  OR2_X1 _6593_ (
    .A1(_4190_),
    .A2(_4191_),
    .ZN(_4192_)
  );
  OR2_X1 _6594_ (
    .A1(_4189_),
    .A2(_4192_),
    .ZN(io_evec[3])
  );
  MUX2_X1 _6595_ (
    .A(_1418_),
    .B(io_cause[2]),
    .S(_4179_),
    .Z(_4193_)
  );
  AND2_X1 _6596_ (
    .A1(_4177_),
    .A2(_4193_),
    .ZN(_4194_)
  );
  AND2_X1 _6597_ (
    .A1(reg_mepc[4]),
    .A2(_2519_),
    .ZN(_4195_)
  );
  AND2_X1 _6598_ (
    .A1(reg_dpc[4]),
    .A2(_2515_),
    .ZN(_4196_)
  );
  OR2_X1 _6599_ (
    .A1(_4195_),
    .A2(_4196_),
    .ZN(_4197_)
  );
  OR2_X1 _6600_ (
    .A1(_4194_),
    .A2(_4197_),
    .ZN(io_evec[4])
  );
  MUX2_X1 _6601_ (
    .A(_1465_),
    .B(_2497_),
    .S(_4179_),
    .Z(_4198_)
  );
  AND2_X1 _6602_ (
    .A1(_4177_),
    .A2(_4198_),
    .ZN(_4199_)
  );
  AND2_X1 _6603_ (
    .A1(reg_mepc[5]),
    .A2(_2519_),
    .ZN(_4200_)
  );
  AND2_X1 _6604_ (
    .A1(reg_dpc[5]),
    .A2(_2515_),
    .ZN(_4201_)
  );
  OR2_X1 _6605_ (
    .A1(_4200_),
    .A2(_4201_),
    .ZN(_4202_)
  );
  OR2_X1 _6606_ (
    .A1(_4199_),
    .A2(_4202_),
    .ZN(io_evec[5])
  );
  MUX2_X1 _6607_ (
    .A(_1517_),
    .B(io_cause[4]),
    .S(_4179_),
    .Z(_4203_)
  );
  AND2_X1 _6608_ (
    .A1(_4177_),
    .A2(_4203_),
    .ZN(_4204_)
  );
  AND2_X1 _6609_ (
    .A1(reg_mepc[6]),
    .A2(_2519_),
    .ZN(_4205_)
  );
  AND2_X1 _6610_ (
    .A1(reg_dpc[6]),
    .A2(_2515_),
    .ZN(_4206_)
  );
  OR2_X1 _6611_ (
    .A1(_4205_),
    .A2(_4206_),
    .ZN(_4207_)
  );
  OR2_X1 _6612_ (
    .A1(_4204_),
    .A2(_4207_),
    .ZN(io_evec[6])
  );
  AND2_X1 _6613_ (
    .A1(reg_mtvec[7]),
    .A2(_4177_),
    .ZN(_4208_)
  );
  AND2_X1 _6614_ (
    .A1(reg_mepc[7]),
    .A2(_2519_),
    .ZN(_4209_)
  );
  AND2_X1 _6615_ (
    .A1(reg_dpc[7]),
    .A2(_2515_),
    .ZN(_4210_)
  );
  OR2_X1 _6616_ (
    .A1(_4209_),
    .A2(_4210_),
    .ZN(_4211_)
  );
  OR2_X1 _6617_ (
    .A1(_4208_),
    .A2(_4211_),
    .ZN(io_evec[7])
  );
  AND2_X1 _6618_ (
    .A1(reg_mtvec[8]),
    .A2(_4177_),
    .ZN(_4212_)
  );
  AND2_X1 _6619_ (
    .A1(reg_mepc[8]),
    .A2(_2519_),
    .ZN(_4213_)
  );
  AND2_X1 _6620_ (
    .A1(reg_dpc[8]),
    .A2(_2515_),
    .ZN(_4214_)
  );
  OR2_X1 _6621_ (
    .A1(_4213_),
    .A2(_4214_),
    .ZN(_4215_)
  );
  OR2_X1 _6622_ (
    .A1(_4212_),
    .A2(_4215_),
    .ZN(io_evec[8])
  );
  AND2_X1 _6623_ (
    .A1(reg_mtvec[9]),
    .A2(_4177_),
    .ZN(_4216_)
  );
  AND2_X1 _6624_ (
    .A1(reg_dpc[9]),
    .A2(_2515_),
    .ZN(_4217_)
  );
  AND2_X1 _6625_ (
    .A1(reg_mepc[9]),
    .A2(_2519_),
    .ZN(_4218_)
  );
  OR2_X1 _6626_ (
    .A1(_4217_),
    .A2(_4218_),
    .ZN(_4219_)
  );
  OR2_X1 _6627_ (
    .A1(_4216_),
    .A2(_4219_),
    .ZN(io_evec[9])
  );
  AND2_X1 _6628_ (
    .A1(reg_mtvec[10]),
    .A2(_4177_),
    .ZN(_4220_)
  );
  AND2_X1 _6629_ (
    .A1(reg_mepc[10]),
    .A2(_2519_),
    .ZN(_4221_)
  );
  AND2_X1 _6630_ (
    .A1(reg_dpc[10]),
    .A2(_2515_),
    .ZN(_4222_)
  );
  OR2_X1 _6631_ (
    .A1(_4221_),
    .A2(_4222_),
    .ZN(_4223_)
  );
  OR2_X1 _6632_ (
    .A1(_4220_),
    .A2(_4223_),
    .ZN(io_evec[10])
  );
  OR2_X1 _6633_ (
    .A1(reg_mtvec[11]),
    .A2(_2506_),
    .ZN(_4224_)
  );
  AND2_X1 _6634_ (
    .A1(_2511_),
    .A2(_4224_),
    .ZN(_4225_)
  );
  AND2_X1 _6635_ (
    .A1(reg_mepc[11]),
    .A2(_2519_),
    .ZN(_4226_)
  );
  AND2_X1 _6636_ (
    .A1(reg_dpc[11]),
    .A2(_2515_),
    .ZN(_4227_)
  );
  OR2_X1 _6637_ (
    .A1(_4226_),
    .A2(_4227_),
    .ZN(_4228_)
  );
  OR2_X1 _6638_ (
    .A1(_4225_),
    .A2(_4228_),
    .ZN(io_evec[11])
  );
  AND2_X1 _6639_ (
    .A1(reg_mtvec[12]),
    .A2(_4177_),
    .ZN(_4229_)
  );
  AND2_X1 _6640_ (
    .A1(reg_mepc[12]),
    .A2(_2519_),
    .ZN(_4230_)
  );
  AND2_X1 _6641_ (
    .A1(reg_dpc[12]),
    .A2(_2515_),
    .ZN(_4231_)
  );
  OR2_X1 _6642_ (
    .A1(_4230_),
    .A2(_4231_),
    .ZN(_4232_)
  );
  OR2_X1 _6643_ (
    .A1(_4229_),
    .A2(_4232_),
    .ZN(io_evec[12])
  );
  AND2_X1 _6644_ (
    .A1(reg_mtvec[13]),
    .A2(_4177_),
    .ZN(_4233_)
  );
  AND2_X1 _6645_ (
    .A1(reg_mepc[13]),
    .A2(_2519_),
    .ZN(_4234_)
  );
  AND2_X1 _6646_ (
    .A1(reg_dpc[13]),
    .A2(_2515_),
    .ZN(_4235_)
  );
  OR2_X1 _6647_ (
    .A1(_4234_),
    .A2(_4235_),
    .ZN(_4236_)
  );
  OR2_X1 _6648_ (
    .A1(_4233_),
    .A2(_4236_),
    .ZN(io_evec[13])
  );
  AND2_X1 _6649_ (
    .A1(reg_mtvec[14]),
    .A2(_4177_),
    .ZN(_4237_)
  );
  AND2_X1 _6650_ (
    .A1(reg_mepc[14]),
    .A2(_2519_),
    .ZN(_4238_)
  );
  AND2_X1 _6651_ (
    .A1(reg_dpc[14]),
    .A2(_2515_),
    .ZN(_4239_)
  );
  OR2_X1 _6652_ (
    .A1(_4238_),
    .A2(_4239_),
    .ZN(_4240_)
  );
  OR2_X1 _6653_ (
    .A1(_4237_),
    .A2(_4240_),
    .ZN(io_evec[14])
  );
  AND2_X1 _6654_ (
    .A1(reg_mtvec[15]),
    .A2(_4177_),
    .ZN(_4241_)
  );
  AND2_X1 _6655_ (
    .A1(reg_mepc[15]),
    .A2(_2519_),
    .ZN(_4242_)
  );
  AND2_X1 _6656_ (
    .A1(reg_dpc[15]),
    .A2(_2515_),
    .ZN(_4243_)
  );
  OR2_X1 _6657_ (
    .A1(_4242_),
    .A2(_4243_),
    .ZN(_4244_)
  );
  OR2_X1 _6658_ (
    .A1(_4241_),
    .A2(_4244_),
    .ZN(io_evec[15])
  );
  AND2_X1 _6659_ (
    .A1(reg_mtvec[16]),
    .A2(_4177_),
    .ZN(_4245_)
  );
  AND2_X1 _6660_ (
    .A1(reg_mepc[16]),
    .A2(_2519_),
    .ZN(_4246_)
  );
  AND2_X1 _6661_ (
    .A1(reg_dpc[16]),
    .A2(_2515_),
    .ZN(_4247_)
  );
  OR2_X1 _6662_ (
    .A1(_4246_),
    .A2(_4247_),
    .ZN(_4248_)
  );
  OR2_X1 _6663_ (
    .A1(_4245_),
    .A2(_4248_),
    .ZN(io_evec[16])
  );
  AND2_X1 _6664_ (
    .A1(reg_mtvec[17]),
    .A2(_4177_),
    .ZN(_4249_)
  );
  AND2_X1 _6665_ (
    .A1(reg_mepc[17]),
    .A2(_2519_),
    .ZN(_4250_)
  );
  AND2_X1 _6666_ (
    .A1(reg_dpc[17]),
    .A2(_2515_),
    .ZN(_4251_)
  );
  OR2_X1 _6667_ (
    .A1(_4250_),
    .A2(_4251_),
    .ZN(_4252_)
  );
  OR2_X1 _6668_ (
    .A1(_4249_),
    .A2(_4252_),
    .ZN(io_evec[17])
  );
  AND2_X1 _6669_ (
    .A1(reg_mtvec[18]),
    .A2(_4177_),
    .ZN(_4253_)
  );
  AND2_X1 _6670_ (
    .A1(reg_mepc[18]),
    .A2(_2519_),
    .ZN(_4254_)
  );
  AND2_X1 _6671_ (
    .A1(reg_dpc[18]),
    .A2(_2515_),
    .ZN(_4255_)
  );
  OR2_X1 _6672_ (
    .A1(_4254_),
    .A2(_4255_),
    .ZN(_4256_)
  );
  OR2_X1 _6673_ (
    .A1(_4253_),
    .A2(_4256_),
    .ZN(io_evec[18])
  );
  AND2_X1 _6674_ (
    .A1(reg_mtvec[19]),
    .A2(_4177_),
    .ZN(_4257_)
  );
  AND2_X1 _6675_ (
    .A1(reg_dpc[19]),
    .A2(_2515_),
    .ZN(_4258_)
  );
  AND2_X1 _6676_ (
    .A1(reg_mepc[19]),
    .A2(_2519_),
    .ZN(_4259_)
  );
  OR2_X1 _6677_ (
    .A1(_4258_),
    .A2(_4259_),
    .ZN(_4260_)
  );
  OR2_X1 _6678_ (
    .A1(_4257_),
    .A2(_4260_),
    .ZN(io_evec[19])
  );
  AND2_X1 _6679_ (
    .A1(reg_mtvec[20]),
    .A2(_4177_),
    .ZN(_4261_)
  );
  AND2_X1 _6680_ (
    .A1(reg_dpc[20]),
    .A2(_2515_),
    .ZN(_4262_)
  );
  AND2_X1 _6681_ (
    .A1(reg_mepc[20]),
    .A2(_2519_),
    .ZN(_4263_)
  );
  OR2_X1 _6682_ (
    .A1(_4262_),
    .A2(_4263_),
    .ZN(_4264_)
  );
  OR2_X1 _6683_ (
    .A1(_4261_),
    .A2(_4264_),
    .ZN(io_evec[20])
  );
  AND2_X1 _6684_ (
    .A1(reg_mtvec[21]),
    .A2(_4177_),
    .ZN(_4265_)
  );
  AND2_X1 _6685_ (
    .A1(reg_mepc[21]),
    .A2(_2519_),
    .ZN(_4266_)
  );
  AND2_X1 _6686_ (
    .A1(reg_dpc[21]),
    .A2(_2515_),
    .ZN(_4267_)
  );
  OR2_X1 _6687_ (
    .A1(_4266_),
    .A2(_4267_),
    .ZN(_4268_)
  );
  OR2_X1 _6688_ (
    .A1(_4265_),
    .A2(_4268_),
    .ZN(io_evec[21])
  );
  AND2_X1 _6689_ (
    .A1(reg_mtvec[22]),
    .A2(_4177_),
    .ZN(_4269_)
  );
  AND2_X1 _6690_ (
    .A1(reg_mepc[22]),
    .A2(_2519_),
    .ZN(_4270_)
  );
  AND2_X1 _6691_ (
    .A1(reg_dpc[22]),
    .A2(_2515_),
    .ZN(_4271_)
  );
  OR2_X1 _6692_ (
    .A1(_4270_),
    .A2(_4271_),
    .ZN(_4272_)
  );
  OR2_X1 _6693_ (
    .A1(_4269_),
    .A2(_4272_),
    .ZN(io_evec[22])
  );
  AND2_X1 _6694_ (
    .A1(reg_mtvec[23]),
    .A2(_4177_),
    .ZN(_4273_)
  );
  AND2_X1 _6695_ (
    .A1(reg_dpc[23]),
    .A2(_2515_),
    .ZN(_4274_)
  );
  AND2_X1 _6696_ (
    .A1(reg_mepc[23]),
    .A2(_2519_),
    .ZN(_4275_)
  );
  OR2_X1 _6697_ (
    .A1(_4274_),
    .A2(_4275_),
    .ZN(_4276_)
  );
  OR2_X1 _6698_ (
    .A1(_4273_),
    .A2(_4276_),
    .ZN(io_evec[23])
  );
  AND2_X1 _6699_ (
    .A1(reg_mtvec[24]),
    .A2(_4177_),
    .ZN(_4277_)
  );
  AND2_X1 _6700_ (
    .A1(reg_dpc[24]),
    .A2(_2515_),
    .ZN(_4278_)
  );
  AND2_X1 _6701_ (
    .A1(reg_mepc[24]),
    .A2(_2519_),
    .ZN(_4279_)
  );
  OR2_X1 _6702_ (
    .A1(_4278_),
    .A2(_4279_),
    .ZN(_4280_)
  );
  OR2_X1 _6703_ (
    .A1(_4277_),
    .A2(_4280_),
    .ZN(io_evec[24])
  );
  AND2_X1 _6704_ (
    .A1(reg_mtvec[25]),
    .A2(_4177_),
    .ZN(_4281_)
  );
  AND2_X1 _6705_ (
    .A1(reg_dpc[25]),
    .A2(_2515_),
    .ZN(_4282_)
  );
  AND2_X1 _6706_ (
    .A1(reg_mepc[25]),
    .A2(_2519_),
    .ZN(_4283_)
  );
  OR2_X1 _6707_ (
    .A1(_4282_),
    .A2(_4283_),
    .ZN(_4284_)
  );
  OR2_X1 _6708_ (
    .A1(_4281_),
    .A2(_4284_),
    .ZN(io_evec[25])
  );
  AND2_X1 _6709_ (
    .A1(reg_mtvec[26]),
    .A2(_4177_),
    .ZN(_4285_)
  );
  AND2_X1 _6710_ (
    .A1(reg_mepc[26]),
    .A2(_2519_),
    .ZN(_4286_)
  );
  AND2_X1 _6711_ (
    .A1(reg_dpc[26]),
    .A2(_2515_),
    .ZN(_4287_)
  );
  OR2_X1 _6712_ (
    .A1(_4286_),
    .A2(_4287_),
    .ZN(_4288_)
  );
  OR2_X1 _6713_ (
    .A1(_4285_),
    .A2(_4288_),
    .ZN(io_evec[26])
  );
  AND2_X1 _6714_ (
    .A1(reg_mtvec[27]),
    .A2(_4177_),
    .ZN(_4289_)
  );
  AND2_X1 _6715_ (
    .A1(reg_mepc[27]),
    .A2(_2519_),
    .ZN(_4290_)
  );
  AND2_X1 _6716_ (
    .A1(reg_dpc[27]),
    .A2(_2515_),
    .ZN(_4291_)
  );
  OR2_X1 _6717_ (
    .A1(_4290_),
    .A2(_4291_),
    .ZN(_4292_)
  );
  OR2_X1 _6718_ (
    .A1(_4289_),
    .A2(_4292_),
    .ZN(io_evec[27])
  );
  AND2_X1 _6719_ (
    .A1(reg_mtvec[28]),
    .A2(_4177_),
    .ZN(_4293_)
  );
  AND2_X1 _6720_ (
    .A1(reg_dpc[28]),
    .A2(_2515_),
    .ZN(_4294_)
  );
  AND2_X1 _6721_ (
    .A1(reg_mepc[28]),
    .A2(_2519_),
    .ZN(_4295_)
  );
  OR2_X1 _6722_ (
    .A1(_4294_),
    .A2(_4295_),
    .ZN(_4296_)
  );
  OR2_X1 _6723_ (
    .A1(_4293_),
    .A2(_4296_),
    .ZN(io_evec[28])
  );
  AND2_X1 _6724_ (
    .A1(reg_mtvec[29]),
    .A2(_4177_),
    .ZN(_4297_)
  );
  AND2_X1 _6725_ (
    .A1(reg_mepc[29]),
    .A2(_2519_),
    .ZN(_4298_)
  );
  AND2_X1 _6726_ (
    .A1(reg_dpc[29]),
    .A2(_2515_),
    .ZN(_4299_)
  );
  OR2_X1 _6727_ (
    .A1(_4298_),
    .A2(_4299_),
    .ZN(_4300_)
  );
  OR2_X1 _6728_ (
    .A1(_4297_),
    .A2(_4300_),
    .ZN(io_evec[29])
  );
  AND2_X1 _6729_ (
    .A1(reg_mtvec[30]),
    .A2(_4177_),
    .ZN(_4301_)
  );
  AND2_X1 _6730_ (
    .A1(reg_mepc[30]),
    .A2(_2519_),
    .ZN(_4302_)
  );
  AND2_X1 _6731_ (
    .A1(reg_dpc[30]),
    .A2(_2515_),
    .ZN(_4303_)
  );
  OR2_X1 _6732_ (
    .A1(_4302_),
    .A2(_4303_),
    .ZN(_4304_)
  );
  OR2_X1 _6733_ (
    .A1(_4301_),
    .A2(_4304_),
    .ZN(io_evec[30])
  );
  AND2_X1 _6734_ (
    .A1(reg_mtvec[31]),
    .A2(_4177_),
    .ZN(_4305_)
  );
  AND2_X1 _6735_ (
    .A1(reg_mepc[31]),
    .A2(_2519_),
    .ZN(_4306_)
  );
  AND2_X1 _6736_ (
    .A1(reg_dpc[31]),
    .A2(_2515_),
    .ZN(_4307_)
  );
  OR2_X1 _6737_ (
    .A1(_4306_),
    .A2(_4307_),
    .ZN(_4308_)
  );
  OR2_X1 _6738_ (
    .A1(_4305_),
    .A2(_4308_),
    .ZN(io_evec[31])
  );
  OR2_X1 _6739_ (
    .A1(io_decode_0_inst[25]),
    .A2(io_decode_0_inst[24]),
    .ZN(_4309_)
  );
  OR2_X1 _6740_ (
    .A1(_0659_),
    .A2(_4309_),
    .ZN(_4310_)
  );
  OR2_X1 _6741_ (
    .A1(io_decode_0_inst[27]),
    .A2(_4310_),
    .ZN(_4311_)
  );
  OR2_X1 _6742_ (
    .A1(io_decode_0_inst[22]),
    .A2(io_decode_0_inst[23]),
    .ZN(_4312_)
  );
  INV_X1 _6743_ (
    .A(_4312_),
    .ZN(_4313_)
  );
  OR2_X1 _6744_ (
    .A1(io_decode_0_inst[31]),
    .A2(io_decode_0_inst[30]),
    .ZN(_4314_)
  );
  OR2_X1 _6745_ (
    .A1(_4312_),
    .A2(_4314_),
    .ZN(_4315_)
  );
  OR2_X1 _6746_ (
    .A1(_0661_),
    .A2(_4312_),
    .ZN(_4316_)
  );
  OR2_X1 _6747_ (
    .A1(io_decode_0_inst[26]),
    .A2(io_decode_0_inst[27]),
    .ZN(_4317_)
  );
  OR2_X1 _6748_ (
    .A1(_4311_),
    .A2(_4315_),
    .ZN(io_decode_0_write_flush)
  );
  AND2_X1 _6749_ (
    .A1(reg_pmp_0_cfg_a[0]),
    .A2(reg_pmp_0_addr[0]),
    .ZN(io_pmp_0_mask[3])
  );
  AND2_X1 _6750_ (
    .A1(reg_pmp_0_addr[1]),
    .A2(io_pmp_0_mask[3]),
    .ZN(io_pmp_0_mask[4])
  );
  AND2_X1 _6751_ (
    .A1(reg_pmp_0_addr[2]),
    .A2(io_pmp_0_mask[4]),
    .ZN(io_pmp_0_mask[5])
  );
  AND2_X1 _6752_ (
    .A1(reg_pmp_0_addr[3]),
    .A2(io_pmp_0_mask[5]),
    .ZN(io_pmp_0_mask[6])
  );
  AND2_X1 _6753_ (
    .A1(reg_pmp_0_addr[4]),
    .A2(io_pmp_0_mask[6]),
    .ZN(io_pmp_0_mask[7])
  );
  AND2_X1 _6754_ (
    .A1(reg_pmp_0_addr[5]),
    .A2(io_pmp_0_mask[7]),
    .ZN(io_pmp_0_mask[8])
  );
  AND2_X1 _6755_ (
    .A1(reg_pmp_0_addr[6]),
    .A2(io_pmp_0_mask[8]),
    .ZN(io_pmp_0_mask[9])
  );
  AND2_X1 _6756_ (
    .A1(reg_pmp_0_addr[7]),
    .A2(io_pmp_0_mask[9]),
    .ZN(io_pmp_0_mask[10])
  );
  AND2_X1 _6757_ (
    .A1(reg_pmp_0_addr[8]),
    .A2(io_pmp_0_mask[10]),
    .ZN(io_pmp_0_mask[11])
  );
  AND2_X1 _6758_ (
    .A1(reg_pmp_0_addr[9]),
    .A2(io_pmp_0_mask[11]),
    .ZN(io_pmp_0_mask[12])
  );
  AND2_X1 _6759_ (
    .A1(reg_pmp_0_addr[10]),
    .A2(io_pmp_0_mask[12]),
    .ZN(io_pmp_0_mask[13])
  );
  AND2_X1 _6760_ (
    .A1(reg_pmp_0_addr[11]),
    .A2(io_pmp_0_mask[13]),
    .ZN(io_pmp_0_mask[14])
  );
  AND2_X1 _6761_ (
    .A1(reg_pmp_0_addr[12]),
    .A2(io_pmp_0_mask[14]),
    .ZN(io_pmp_0_mask[15])
  );
  AND2_X1 _6762_ (
    .A1(reg_pmp_0_addr[13]),
    .A2(io_pmp_0_mask[15]),
    .ZN(io_pmp_0_mask[16])
  );
  AND2_X1 _6763_ (
    .A1(reg_pmp_0_addr[14]),
    .A2(io_pmp_0_mask[16]),
    .ZN(io_pmp_0_mask[17])
  );
  AND2_X1 _6764_ (
    .A1(reg_pmp_0_addr[15]),
    .A2(io_pmp_0_mask[17]),
    .ZN(io_pmp_0_mask[18])
  );
  AND2_X1 _6765_ (
    .A1(reg_pmp_0_addr[16]),
    .A2(io_pmp_0_mask[18]),
    .ZN(io_pmp_0_mask[19])
  );
  AND2_X1 _6766_ (
    .A1(reg_pmp_0_addr[17]),
    .A2(io_pmp_0_mask[19]),
    .ZN(io_pmp_0_mask[20])
  );
  AND2_X1 _6767_ (
    .A1(reg_pmp_0_addr[18]),
    .A2(io_pmp_0_mask[20]),
    .ZN(io_pmp_0_mask[21])
  );
  AND2_X1 _6768_ (
    .A1(reg_pmp_0_addr[19]),
    .A2(io_pmp_0_mask[21]),
    .ZN(io_pmp_0_mask[22])
  );
  AND2_X1 _6769_ (
    .A1(reg_pmp_0_addr[20]),
    .A2(io_pmp_0_mask[22]),
    .ZN(io_pmp_0_mask[23])
  );
  AND2_X1 _6770_ (
    .A1(reg_pmp_0_addr[21]),
    .A2(io_pmp_0_mask[23]),
    .ZN(io_pmp_0_mask[24])
  );
  AND2_X1 _6771_ (
    .A1(reg_pmp_0_addr[22]),
    .A2(io_pmp_0_mask[24]),
    .ZN(io_pmp_0_mask[25])
  );
  AND2_X1 _6772_ (
    .A1(reg_pmp_0_addr[23]),
    .A2(io_pmp_0_mask[25]),
    .ZN(io_pmp_0_mask[26])
  );
  AND2_X1 _6773_ (
    .A1(reg_pmp_0_addr[24]),
    .A2(io_pmp_0_mask[26]),
    .ZN(io_pmp_0_mask[27])
  );
  AND2_X1 _6774_ (
    .A1(reg_pmp_0_addr[25]),
    .A2(io_pmp_0_mask[27]),
    .ZN(io_pmp_0_mask[28])
  );
  AND2_X1 _6775_ (
    .A1(reg_pmp_0_addr[26]),
    .A2(io_pmp_0_mask[28]),
    .ZN(io_pmp_0_mask[29])
  );
  AND2_X1 _6776_ (
    .A1(reg_pmp_0_addr[27]),
    .A2(io_pmp_0_mask[29]),
    .ZN(io_pmp_0_mask[30])
  );
  AND2_X1 _6777_ (
    .A1(reg_pmp_0_addr[28]),
    .A2(io_pmp_0_mask[30]),
    .ZN(io_pmp_0_mask[31])
  );
  AND2_X1 _6778_ (
    .A1(reg_pmp_1_cfg_a[0]),
    .A2(reg_pmp_1_addr[0]),
    .ZN(io_pmp_1_mask[3])
  );
  AND2_X1 _6779_ (
    .A1(reg_pmp_1_addr[1]),
    .A2(io_pmp_1_mask[3]),
    .ZN(io_pmp_1_mask[4])
  );
  AND2_X1 _6780_ (
    .A1(reg_pmp_1_addr[2]),
    .A2(io_pmp_1_mask[4]),
    .ZN(io_pmp_1_mask[5])
  );
  AND2_X1 _6781_ (
    .A1(reg_pmp_1_addr[3]),
    .A2(io_pmp_1_mask[5]),
    .ZN(io_pmp_1_mask[6])
  );
  AND2_X1 _6782_ (
    .A1(reg_pmp_1_addr[4]),
    .A2(io_pmp_1_mask[6]),
    .ZN(io_pmp_1_mask[7])
  );
  AND2_X1 _6783_ (
    .A1(reg_pmp_1_addr[5]),
    .A2(io_pmp_1_mask[7]),
    .ZN(io_pmp_1_mask[8])
  );
  AND2_X1 _6784_ (
    .A1(reg_pmp_1_addr[6]),
    .A2(io_pmp_1_mask[8]),
    .ZN(io_pmp_1_mask[9])
  );
  AND2_X1 _6785_ (
    .A1(reg_pmp_1_addr[7]),
    .A2(io_pmp_1_mask[9]),
    .ZN(io_pmp_1_mask[10])
  );
  AND2_X1 _6786_ (
    .A1(reg_pmp_1_addr[8]),
    .A2(io_pmp_1_mask[10]),
    .ZN(io_pmp_1_mask[11])
  );
  AND2_X1 _6787_ (
    .A1(reg_pmp_1_addr[9]),
    .A2(io_pmp_1_mask[11]),
    .ZN(io_pmp_1_mask[12])
  );
  AND2_X1 _6788_ (
    .A1(reg_pmp_1_addr[10]),
    .A2(io_pmp_1_mask[12]),
    .ZN(io_pmp_1_mask[13])
  );
  AND2_X1 _6789_ (
    .A1(reg_pmp_1_addr[11]),
    .A2(io_pmp_1_mask[13]),
    .ZN(io_pmp_1_mask[14])
  );
  AND2_X1 _6790_ (
    .A1(reg_pmp_1_addr[12]),
    .A2(io_pmp_1_mask[14]),
    .ZN(io_pmp_1_mask[15])
  );
  AND2_X1 _6791_ (
    .A1(reg_pmp_1_addr[13]),
    .A2(io_pmp_1_mask[15]),
    .ZN(io_pmp_1_mask[16])
  );
  AND2_X1 _6792_ (
    .A1(reg_pmp_1_addr[14]),
    .A2(io_pmp_1_mask[16]),
    .ZN(io_pmp_1_mask[17])
  );
  AND2_X1 _6793_ (
    .A1(reg_pmp_1_addr[15]),
    .A2(io_pmp_1_mask[17]),
    .ZN(io_pmp_1_mask[18])
  );
  AND2_X1 _6794_ (
    .A1(reg_pmp_1_addr[16]),
    .A2(io_pmp_1_mask[18]),
    .ZN(io_pmp_1_mask[19])
  );
  AND2_X1 _6795_ (
    .A1(reg_pmp_1_addr[17]),
    .A2(io_pmp_1_mask[19]),
    .ZN(io_pmp_1_mask[20])
  );
  AND2_X1 _6796_ (
    .A1(reg_pmp_1_addr[18]),
    .A2(io_pmp_1_mask[20]),
    .ZN(io_pmp_1_mask[21])
  );
  AND2_X1 _6797_ (
    .A1(reg_pmp_1_addr[19]),
    .A2(io_pmp_1_mask[21]),
    .ZN(io_pmp_1_mask[22])
  );
  AND2_X1 _6798_ (
    .A1(reg_pmp_1_addr[20]),
    .A2(io_pmp_1_mask[22]),
    .ZN(io_pmp_1_mask[23])
  );
  AND2_X1 _6799_ (
    .A1(reg_pmp_1_addr[21]),
    .A2(io_pmp_1_mask[23]),
    .ZN(io_pmp_1_mask[24])
  );
  AND2_X1 _6800_ (
    .A1(reg_pmp_1_addr[22]),
    .A2(io_pmp_1_mask[24]),
    .ZN(io_pmp_1_mask[25])
  );
  AND2_X1 _6801_ (
    .A1(reg_pmp_1_addr[23]),
    .A2(io_pmp_1_mask[25]),
    .ZN(io_pmp_1_mask[26])
  );
  AND2_X1 _6802_ (
    .A1(reg_pmp_1_addr[24]),
    .A2(io_pmp_1_mask[26]),
    .ZN(io_pmp_1_mask[27])
  );
  AND2_X1 _6803_ (
    .A1(reg_pmp_1_addr[25]),
    .A2(io_pmp_1_mask[27]),
    .ZN(io_pmp_1_mask[28])
  );
  AND2_X1 _6804_ (
    .A1(reg_pmp_1_addr[26]),
    .A2(io_pmp_1_mask[28]),
    .ZN(io_pmp_1_mask[29])
  );
  AND2_X1 _6805_ (
    .A1(reg_pmp_1_addr[27]),
    .A2(io_pmp_1_mask[29]),
    .ZN(io_pmp_1_mask[30])
  );
  AND2_X1 _6806_ (
    .A1(reg_pmp_1_addr[28]),
    .A2(io_pmp_1_mask[30]),
    .ZN(io_pmp_1_mask[31])
  );
  AND2_X1 _6807_ (
    .A1(reg_pmp_2_cfg_a[0]),
    .A2(reg_pmp_2_addr[0]),
    .ZN(io_pmp_2_mask[3])
  );
  AND2_X1 _6808_ (
    .A1(reg_pmp_2_addr[1]),
    .A2(io_pmp_2_mask[3]),
    .ZN(io_pmp_2_mask[4])
  );
  AND2_X1 _6809_ (
    .A1(reg_pmp_2_addr[2]),
    .A2(io_pmp_2_mask[4]),
    .ZN(io_pmp_2_mask[5])
  );
  AND2_X1 _6810_ (
    .A1(reg_pmp_2_addr[3]),
    .A2(io_pmp_2_mask[5]),
    .ZN(io_pmp_2_mask[6])
  );
  AND2_X1 _6811_ (
    .A1(reg_pmp_2_addr[4]),
    .A2(io_pmp_2_mask[6]),
    .ZN(io_pmp_2_mask[7])
  );
  AND2_X1 _6812_ (
    .A1(reg_pmp_2_addr[5]),
    .A2(io_pmp_2_mask[7]),
    .ZN(io_pmp_2_mask[8])
  );
  AND2_X1 _6813_ (
    .A1(reg_pmp_2_addr[6]),
    .A2(io_pmp_2_mask[8]),
    .ZN(io_pmp_2_mask[9])
  );
  AND2_X1 _6814_ (
    .A1(reg_pmp_2_addr[7]),
    .A2(io_pmp_2_mask[9]),
    .ZN(io_pmp_2_mask[10])
  );
  AND2_X1 _6815_ (
    .A1(reg_pmp_2_addr[8]),
    .A2(io_pmp_2_mask[10]),
    .ZN(io_pmp_2_mask[11])
  );
  AND2_X1 _6816_ (
    .A1(reg_pmp_2_addr[9]),
    .A2(io_pmp_2_mask[11]),
    .ZN(io_pmp_2_mask[12])
  );
  AND2_X1 _6817_ (
    .A1(reg_pmp_2_addr[10]),
    .A2(io_pmp_2_mask[12]),
    .ZN(io_pmp_2_mask[13])
  );
  AND2_X1 _6818_ (
    .A1(reg_pmp_2_addr[11]),
    .A2(io_pmp_2_mask[13]),
    .ZN(io_pmp_2_mask[14])
  );
  AND2_X1 _6819_ (
    .A1(reg_pmp_2_addr[12]),
    .A2(io_pmp_2_mask[14]),
    .ZN(io_pmp_2_mask[15])
  );
  AND2_X1 _6820_ (
    .A1(reg_pmp_2_addr[13]),
    .A2(io_pmp_2_mask[15]),
    .ZN(io_pmp_2_mask[16])
  );
  AND2_X1 _6821_ (
    .A1(reg_pmp_2_addr[14]),
    .A2(io_pmp_2_mask[16]),
    .ZN(io_pmp_2_mask[17])
  );
  AND2_X1 _6822_ (
    .A1(reg_pmp_2_addr[15]),
    .A2(io_pmp_2_mask[17]),
    .ZN(io_pmp_2_mask[18])
  );
  AND2_X1 _6823_ (
    .A1(reg_pmp_2_addr[16]),
    .A2(io_pmp_2_mask[18]),
    .ZN(io_pmp_2_mask[19])
  );
  AND2_X1 _6824_ (
    .A1(reg_pmp_2_addr[17]),
    .A2(io_pmp_2_mask[19]),
    .ZN(io_pmp_2_mask[20])
  );
  AND2_X1 _6825_ (
    .A1(reg_pmp_2_addr[18]),
    .A2(io_pmp_2_mask[20]),
    .ZN(io_pmp_2_mask[21])
  );
  AND2_X1 _6826_ (
    .A1(reg_pmp_2_addr[19]),
    .A2(io_pmp_2_mask[21]),
    .ZN(io_pmp_2_mask[22])
  );
  AND2_X1 _6827_ (
    .A1(reg_pmp_2_addr[20]),
    .A2(io_pmp_2_mask[22]),
    .ZN(io_pmp_2_mask[23])
  );
  AND2_X1 _6828_ (
    .A1(reg_pmp_2_addr[21]),
    .A2(io_pmp_2_mask[23]),
    .ZN(io_pmp_2_mask[24])
  );
  AND2_X1 _6829_ (
    .A1(reg_pmp_2_addr[22]),
    .A2(io_pmp_2_mask[24]),
    .ZN(io_pmp_2_mask[25])
  );
  AND2_X1 _6830_ (
    .A1(reg_pmp_2_addr[23]),
    .A2(io_pmp_2_mask[25]),
    .ZN(io_pmp_2_mask[26])
  );
  AND2_X1 _6831_ (
    .A1(reg_pmp_2_addr[24]),
    .A2(io_pmp_2_mask[26]),
    .ZN(io_pmp_2_mask[27])
  );
  AND2_X1 _6832_ (
    .A1(reg_pmp_2_addr[25]),
    .A2(io_pmp_2_mask[27]),
    .ZN(io_pmp_2_mask[28])
  );
  AND2_X1 _6833_ (
    .A1(reg_pmp_2_addr[26]),
    .A2(io_pmp_2_mask[28]),
    .ZN(io_pmp_2_mask[29])
  );
  AND2_X1 _6834_ (
    .A1(reg_pmp_2_addr[27]),
    .A2(io_pmp_2_mask[29]),
    .ZN(io_pmp_2_mask[30])
  );
  AND2_X1 _6835_ (
    .A1(reg_pmp_2_addr[28]),
    .A2(io_pmp_2_mask[30]),
    .ZN(io_pmp_2_mask[31])
  );
  AND2_X1 _6836_ (
    .A1(reg_pmp_3_cfg_a[0]),
    .A2(reg_pmp_3_addr[0]),
    .ZN(io_pmp_3_mask[3])
  );
  AND2_X1 _6837_ (
    .A1(reg_pmp_3_addr[1]),
    .A2(io_pmp_3_mask[3]),
    .ZN(io_pmp_3_mask[4])
  );
  AND2_X1 _6838_ (
    .A1(reg_pmp_3_addr[2]),
    .A2(io_pmp_3_mask[4]),
    .ZN(io_pmp_3_mask[5])
  );
  AND2_X1 _6839_ (
    .A1(reg_pmp_3_addr[3]),
    .A2(io_pmp_3_mask[5]),
    .ZN(io_pmp_3_mask[6])
  );
  AND2_X1 _6840_ (
    .A1(reg_pmp_3_addr[4]),
    .A2(io_pmp_3_mask[6]),
    .ZN(io_pmp_3_mask[7])
  );
  AND2_X1 _6841_ (
    .A1(reg_pmp_3_addr[5]),
    .A2(io_pmp_3_mask[7]),
    .ZN(io_pmp_3_mask[8])
  );
  AND2_X1 _6842_ (
    .A1(reg_pmp_3_addr[6]),
    .A2(io_pmp_3_mask[8]),
    .ZN(io_pmp_3_mask[9])
  );
  AND2_X1 _6843_ (
    .A1(reg_pmp_3_addr[7]),
    .A2(io_pmp_3_mask[9]),
    .ZN(io_pmp_3_mask[10])
  );
  AND2_X1 _6844_ (
    .A1(reg_pmp_3_addr[8]),
    .A2(io_pmp_3_mask[10]),
    .ZN(io_pmp_3_mask[11])
  );
  AND2_X1 _6845_ (
    .A1(reg_pmp_3_addr[9]),
    .A2(io_pmp_3_mask[11]),
    .ZN(io_pmp_3_mask[12])
  );
  AND2_X1 _6846_ (
    .A1(reg_pmp_3_addr[10]),
    .A2(io_pmp_3_mask[12]),
    .ZN(io_pmp_3_mask[13])
  );
  AND2_X1 _6847_ (
    .A1(reg_pmp_3_addr[11]),
    .A2(io_pmp_3_mask[13]),
    .ZN(io_pmp_3_mask[14])
  );
  AND2_X1 _6848_ (
    .A1(reg_pmp_3_addr[12]),
    .A2(io_pmp_3_mask[14]),
    .ZN(io_pmp_3_mask[15])
  );
  AND2_X1 _6849_ (
    .A1(reg_pmp_3_addr[13]),
    .A2(io_pmp_3_mask[15]),
    .ZN(io_pmp_3_mask[16])
  );
  AND2_X1 _6850_ (
    .A1(reg_pmp_3_addr[14]),
    .A2(io_pmp_3_mask[16]),
    .ZN(io_pmp_3_mask[17])
  );
  AND2_X1 _6851_ (
    .A1(reg_pmp_3_addr[15]),
    .A2(io_pmp_3_mask[17]),
    .ZN(io_pmp_3_mask[18])
  );
  AND2_X1 _6852_ (
    .A1(reg_pmp_3_addr[16]),
    .A2(io_pmp_3_mask[18]),
    .ZN(io_pmp_3_mask[19])
  );
  AND2_X1 _6853_ (
    .A1(reg_pmp_3_addr[17]),
    .A2(io_pmp_3_mask[19]),
    .ZN(io_pmp_3_mask[20])
  );
  AND2_X1 _6854_ (
    .A1(reg_pmp_3_addr[18]),
    .A2(io_pmp_3_mask[20]),
    .ZN(io_pmp_3_mask[21])
  );
  AND2_X1 _6855_ (
    .A1(reg_pmp_3_addr[19]),
    .A2(io_pmp_3_mask[21]),
    .ZN(io_pmp_3_mask[22])
  );
  AND2_X1 _6856_ (
    .A1(reg_pmp_3_addr[20]),
    .A2(io_pmp_3_mask[22]),
    .ZN(io_pmp_3_mask[23])
  );
  AND2_X1 _6857_ (
    .A1(reg_pmp_3_addr[21]),
    .A2(io_pmp_3_mask[23]),
    .ZN(io_pmp_3_mask[24])
  );
  AND2_X1 _6858_ (
    .A1(reg_pmp_3_addr[22]),
    .A2(io_pmp_3_mask[24]),
    .ZN(io_pmp_3_mask[25])
  );
  AND2_X1 _6859_ (
    .A1(reg_pmp_3_addr[23]),
    .A2(io_pmp_3_mask[25]),
    .ZN(io_pmp_3_mask[26])
  );
  AND2_X1 _6860_ (
    .A1(reg_pmp_3_addr[24]),
    .A2(io_pmp_3_mask[26]),
    .ZN(io_pmp_3_mask[27])
  );
  AND2_X1 _6861_ (
    .A1(reg_pmp_3_addr[25]),
    .A2(io_pmp_3_mask[27]),
    .ZN(io_pmp_3_mask[28])
  );
  AND2_X1 _6862_ (
    .A1(reg_pmp_3_addr[26]),
    .A2(io_pmp_3_mask[28]),
    .ZN(io_pmp_3_mask[29])
  );
  AND2_X1 _6863_ (
    .A1(reg_pmp_3_addr[27]),
    .A2(io_pmp_3_mask[29]),
    .ZN(io_pmp_3_mask[30])
  );
  AND2_X1 _6864_ (
    .A1(reg_pmp_3_addr[28]),
    .A2(io_pmp_3_mask[30]),
    .ZN(io_pmp_3_mask[31])
  );
  AND2_X1 _6865_ (
    .A1(reg_pmp_4_cfg_a[0]),
    .A2(reg_pmp_4_addr[0]),
    .ZN(io_pmp_4_mask[3])
  );
  AND2_X1 _6866_ (
    .A1(reg_pmp_4_addr[1]),
    .A2(io_pmp_4_mask[3]),
    .ZN(io_pmp_4_mask[4])
  );
  AND2_X1 _6867_ (
    .A1(reg_pmp_4_addr[2]),
    .A2(io_pmp_4_mask[4]),
    .ZN(io_pmp_4_mask[5])
  );
  AND2_X1 _6868_ (
    .A1(reg_pmp_4_addr[3]),
    .A2(io_pmp_4_mask[5]),
    .ZN(io_pmp_4_mask[6])
  );
  AND2_X1 _6869_ (
    .A1(reg_pmp_4_addr[4]),
    .A2(io_pmp_4_mask[6]),
    .ZN(io_pmp_4_mask[7])
  );
  AND2_X1 _6870_ (
    .A1(reg_pmp_4_addr[5]),
    .A2(io_pmp_4_mask[7]),
    .ZN(io_pmp_4_mask[8])
  );
  AND2_X1 _6871_ (
    .A1(reg_pmp_4_addr[6]),
    .A2(io_pmp_4_mask[8]),
    .ZN(io_pmp_4_mask[9])
  );
  AND2_X1 _6872_ (
    .A1(reg_pmp_4_addr[7]),
    .A2(io_pmp_4_mask[9]),
    .ZN(io_pmp_4_mask[10])
  );
  AND2_X1 _6873_ (
    .A1(reg_pmp_4_addr[8]),
    .A2(io_pmp_4_mask[10]),
    .ZN(io_pmp_4_mask[11])
  );
  AND2_X1 _6874_ (
    .A1(reg_pmp_4_addr[9]),
    .A2(io_pmp_4_mask[11]),
    .ZN(io_pmp_4_mask[12])
  );
  AND2_X1 _6875_ (
    .A1(reg_pmp_4_addr[10]),
    .A2(io_pmp_4_mask[12]),
    .ZN(io_pmp_4_mask[13])
  );
  AND2_X1 _6876_ (
    .A1(reg_pmp_4_addr[11]),
    .A2(io_pmp_4_mask[13]),
    .ZN(io_pmp_4_mask[14])
  );
  AND2_X1 _6877_ (
    .A1(reg_pmp_4_addr[12]),
    .A2(io_pmp_4_mask[14]),
    .ZN(io_pmp_4_mask[15])
  );
  AND2_X1 _6878_ (
    .A1(reg_pmp_4_addr[13]),
    .A2(io_pmp_4_mask[15]),
    .ZN(io_pmp_4_mask[16])
  );
  AND2_X1 _6879_ (
    .A1(reg_pmp_4_addr[14]),
    .A2(io_pmp_4_mask[16]),
    .ZN(io_pmp_4_mask[17])
  );
  AND2_X1 _6880_ (
    .A1(reg_pmp_4_addr[15]),
    .A2(io_pmp_4_mask[17]),
    .ZN(io_pmp_4_mask[18])
  );
  AND2_X1 _6881_ (
    .A1(reg_pmp_4_addr[16]),
    .A2(io_pmp_4_mask[18]),
    .ZN(io_pmp_4_mask[19])
  );
  AND2_X1 _6882_ (
    .A1(reg_pmp_4_addr[17]),
    .A2(io_pmp_4_mask[19]),
    .ZN(io_pmp_4_mask[20])
  );
  AND2_X1 _6883_ (
    .A1(reg_pmp_4_addr[18]),
    .A2(io_pmp_4_mask[20]),
    .ZN(io_pmp_4_mask[21])
  );
  AND2_X1 _6884_ (
    .A1(reg_pmp_4_addr[19]),
    .A2(io_pmp_4_mask[21]),
    .ZN(io_pmp_4_mask[22])
  );
  AND2_X1 _6885_ (
    .A1(reg_pmp_4_addr[20]),
    .A2(io_pmp_4_mask[22]),
    .ZN(io_pmp_4_mask[23])
  );
  AND2_X1 _6886_ (
    .A1(reg_pmp_4_addr[21]),
    .A2(io_pmp_4_mask[23]),
    .ZN(io_pmp_4_mask[24])
  );
  AND2_X1 _6887_ (
    .A1(reg_pmp_4_addr[22]),
    .A2(io_pmp_4_mask[24]),
    .ZN(io_pmp_4_mask[25])
  );
  AND2_X1 _6888_ (
    .A1(reg_pmp_4_addr[23]),
    .A2(io_pmp_4_mask[25]),
    .ZN(io_pmp_4_mask[26])
  );
  AND2_X1 _6889_ (
    .A1(reg_pmp_4_addr[24]),
    .A2(io_pmp_4_mask[26]),
    .ZN(io_pmp_4_mask[27])
  );
  AND2_X1 _6890_ (
    .A1(reg_pmp_4_addr[25]),
    .A2(io_pmp_4_mask[27]),
    .ZN(io_pmp_4_mask[28])
  );
  AND2_X1 _6891_ (
    .A1(reg_pmp_4_addr[26]),
    .A2(io_pmp_4_mask[28]),
    .ZN(io_pmp_4_mask[29])
  );
  AND2_X1 _6892_ (
    .A1(reg_pmp_4_addr[27]),
    .A2(io_pmp_4_mask[29]),
    .ZN(io_pmp_4_mask[30])
  );
  AND2_X1 _6893_ (
    .A1(reg_pmp_4_addr[28]),
    .A2(io_pmp_4_mask[30]),
    .ZN(io_pmp_4_mask[31])
  );
  AND2_X1 _6894_ (
    .A1(reg_pmp_5_cfg_a[0]),
    .A2(reg_pmp_5_addr[0]),
    .ZN(io_pmp_5_mask[3])
  );
  AND2_X1 _6895_ (
    .A1(reg_pmp_5_addr[1]),
    .A2(io_pmp_5_mask[3]),
    .ZN(io_pmp_5_mask[4])
  );
  AND2_X1 _6896_ (
    .A1(reg_pmp_5_addr[2]),
    .A2(io_pmp_5_mask[4]),
    .ZN(io_pmp_5_mask[5])
  );
  AND2_X1 _6897_ (
    .A1(reg_pmp_5_addr[3]),
    .A2(io_pmp_5_mask[5]),
    .ZN(io_pmp_5_mask[6])
  );
  AND2_X1 _6898_ (
    .A1(reg_pmp_5_addr[4]),
    .A2(io_pmp_5_mask[6]),
    .ZN(io_pmp_5_mask[7])
  );
  AND2_X1 _6899_ (
    .A1(reg_pmp_5_addr[5]),
    .A2(io_pmp_5_mask[7]),
    .ZN(io_pmp_5_mask[8])
  );
  AND2_X1 _6900_ (
    .A1(reg_pmp_5_addr[6]),
    .A2(io_pmp_5_mask[8]),
    .ZN(io_pmp_5_mask[9])
  );
  AND2_X1 _6901_ (
    .A1(reg_pmp_5_addr[7]),
    .A2(io_pmp_5_mask[9]),
    .ZN(io_pmp_5_mask[10])
  );
  AND2_X1 _6902_ (
    .A1(reg_pmp_5_addr[8]),
    .A2(io_pmp_5_mask[10]),
    .ZN(io_pmp_5_mask[11])
  );
  AND2_X1 _6903_ (
    .A1(reg_pmp_5_addr[9]),
    .A2(io_pmp_5_mask[11]),
    .ZN(io_pmp_5_mask[12])
  );
  AND2_X1 _6904_ (
    .A1(reg_pmp_5_addr[10]),
    .A2(io_pmp_5_mask[12]),
    .ZN(io_pmp_5_mask[13])
  );
  AND2_X1 _6905_ (
    .A1(reg_pmp_5_addr[11]),
    .A2(io_pmp_5_mask[13]),
    .ZN(io_pmp_5_mask[14])
  );
  AND2_X1 _6906_ (
    .A1(reg_pmp_5_addr[12]),
    .A2(io_pmp_5_mask[14]),
    .ZN(io_pmp_5_mask[15])
  );
  AND2_X1 _6907_ (
    .A1(reg_pmp_5_addr[13]),
    .A2(io_pmp_5_mask[15]),
    .ZN(io_pmp_5_mask[16])
  );
  AND2_X1 _6908_ (
    .A1(reg_pmp_5_addr[14]),
    .A2(io_pmp_5_mask[16]),
    .ZN(io_pmp_5_mask[17])
  );
  AND2_X1 _6909_ (
    .A1(reg_pmp_5_addr[15]),
    .A2(io_pmp_5_mask[17]),
    .ZN(io_pmp_5_mask[18])
  );
  AND2_X1 _6910_ (
    .A1(reg_pmp_5_addr[16]),
    .A2(io_pmp_5_mask[18]),
    .ZN(io_pmp_5_mask[19])
  );
  AND2_X1 _6911_ (
    .A1(reg_pmp_5_addr[17]),
    .A2(io_pmp_5_mask[19]),
    .ZN(io_pmp_5_mask[20])
  );
  AND2_X1 _6912_ (
    .A1(reg_pmp_5_addr[18]),
    .A2(io_pmp_5_mask[20]),
    .ZN(io_pmp_5_mask[21])
  );
  AND2_X1 _6913_ (
    .A1(reg_pmp_5_addr[19]),
    .A2(io_pmp_5_mask[21]),
    .ZN(io_pmp_5_mask[22])
  );
  AND2_X1 _6914_ (
    .A1(reg_pmp_5_addr[20]),
    .A2(io_pmp_5_mask[22]),
    .ZN(io_pmp_5_mask[23])
  );
  AND2_X1 _6915_ (
    .A1(reg_pmp_5_addr[21]),
    .A2(io_pmp_5_mask[23]),
    .ZN(io_pmp_5_mask[24])
  );
  AND2_X1 _6916_ (
    .A1(reg_pmp_5_addr[22]),
    .A2(io_pmp_5_mask[24]),
    .ZN(io_pmp_5_mask[25])
  );
  AND2_X1 _6917_ (
    .A1(reg_pmp_5_addr[23]),
    .A2(io_pmp_5_mask[25]),
    .ZN(io_pmp_5_mask[26])
  );
  AND2_X1 _6918_ (
    .A1(reg_pmp_5_addr[24]),
    .A2(io_pmp_5_mask[26]),
    .ZN(io_pmp_5_mask[27])
  );
  AND2_X1 _6919_ (
    .A1(reg_pmp_5_addr[25]),
    .A2(io_pmp_5_mask[27]),
    .ZN(io_pmp_5_mask[28])
  );
  AND2_X1 _6920_ (
    .A1(reg_pmp_5_addr[26]),
    .A2(io_pmp_5_mask[28]),
    .ZN(io_pmp_5_mask[29])
  );
  AND2_X1 _6921_ (
    .A1(reg_pmp_5_addr[27]),
    .A2(io_pmp_5_mask[29]),
    .ZN(io_pmp_5_mask[30])
  );
  AND2_X1 _6922_ (
    .A1(reg_pmp_5_addr[28]),
    .A2(io_pmp_5_mask[30]),
    .ZN(io_pmp_5_mask[31])
  );
  AND2_X1 _6923_ (
    .A1(reg_pmp_6_cfg_a[0]),
    .A2(reg_pmp_6_addr[0]),
    .ZN(io_pmp_6_mask[3])
  );
  AND2_X1 _6924_ (
    .A1(reg_pmp_6_addr[1]),
    .A2(io_pmp_6_mask[3]),
    .ZN(io_pmp_6_mask[4])
  );
  AND2_X1 _6925_ (
    .A1(reg_pmp_6_addr[2]),
    .A2(io_pmp_6_mask[4]),
    .ZN(io_pmp_6_mask[5])
  );
  AND2_X1 _6926_ (
    .A1(reg_pmp_6_addr[3]),
    .A2(io_pmp_6_mask[5]),
    .ZN(io_pmp_6_mask[6])
  );
  AND2_X1 _6927_ (
    .A1(reg_pmp_6_addr[4]),
    .A2(io_pmp_6_mask[6]),
    .ZN(io_pmp_6_mask[7])
  );
  AND2_X1 _6928_ (
    .A1(reg_pmp_6_addr[5]),
    .A2(io_pmp_6_mask[7]),
    .ZN(io_pmp_6_mask[8])
  );
  AND2_X1 _6929_ (
    .A1(reg_pmp_6_addr[6]),
    .A2(io_pmp_6_mask[8]),
    .ZN(io_pmp_6_mask[9])
  );
  AND2_X1 _6930_ (
    .A1(reg_pmp_6_addr[7]),
    .A2(io_pmp_6_mask[9]),
    .ZN(io_pmp_6_mask[10])
  );
  AND2_X1 _6931_ (
    .A1(reg_pmp_6_addr[8]),
    .A2(io_pmp_6_mask[10]),
    .ZN(io_pmp_6_mask[11])
  );
  AND2_X1 _6932_ (
    .A1(reg_pmp_6_addr[9]),
    .A2(io_pmp_6_mask[11]),
    .ZN(io_pmp_6_mask[12])
  );
  AND2_X1 _6933_ (
    .A1(reg_pmp_6_addr[10]),
    .A2(io_pmp_6_mask[12]),
    .ZN(io_pmp_6_mask[13])
  );
  AND2_X1 _6934_ (
    .A1(reg_pmp_6_addr[11]),
    .A2(io_pmp_6_mask[13]),
    .ZN(io_pmp_6_mask[14])
  );
  AND2_X1 _6935_ (
    .A1(reg_pmp_6_addr[12]),
    .A2(io_pmp_6_mask[14]),
    .ZN(io_pmp_6_mask[15])
  );
  AND2_X1 _6936_ (
    .A1(reg_pmp_6_addr[13]),
    .A2(io_pmp_6_mask[15]),
    .ZN(io_pmp_6_mask[16])
  );
  AND2_X1 _6937_ (
    .A1(reg_pmp_6_addr[14]),
    .A2(io_pmp_6_mask[16]),
    .ZN(io_pmp_6_mask[17])
  );
  AND2_X1 _6938_ (
    .A1(reg_pmp_6_addr[15]),
    .A2(io_pmp_6_mask[17]),
    .ZN(io_pmp_6_mask[18])
  );
  AND2_X1 _6939_ (
    .A1(reg_pmp_6_addr[16]),
    .A2(io_pmp_6_mask[18]),
    .ZN(io_pmp_6_mask[19])
  );
  AND2_X1 _6940_ (
    .A1(reg_pmp_6_addr[17]),
    .A2(io_pmp_6_mask[19]),
    .ZN(io_pmp_6_mask[20])
  );
  AND2_X1 _6941_ (
    .A1(reg_pmp_6_addr[18]),
    .A2(io_pmp_6_mask[20]),
    .ZN(io_pmp_6_mask[21])
  );
  AND2_X1 _6942_ (
    .A1(reg_pmp_6_addr[19]),
    .A2(io_pmp_6_mask[21]),
    .ZN(io_pmp_6_mask[22])
  );
  AND2_X1 _6943_ (
    .A1(reg_pmp_6_addr[20]),
    .A2(io_pmp_6_mask[22]),
    .ZN(io_pmp_6_mask[23])
  );
  AND2_X1 _6944_ (
    .A1(reg_pmp_6_addr[21]),
    .A2(io_pmp_6_mask[23]),
    .ZN(io_pmp_6_mask[24])
  );
  AND2_X1 _6945_ (
    .A1(reg_pmp_6_addr[22]),
    .A2(io_pmp_6_mask[24]),
    .ZN(io_pmp_6_mask[25])
  );
  AND2_X1 _6946_ (
    .A1(reg_pmp_6_addr[23]),
    .A2(io_pmp_6_mask[25]),
    .ZN(io_pmp_6_mask[26])
  );
  AND2_X1 _6947_ (
    .A1(reg_pmp_6_addr[24]),
    .A2(io_pmp_6_mask[26]),
    .ZN(io_pmp_6_mask[27])
  );
  AND2_X1 _6948_ (
    .A1(reg_pmp_6_addr[25]),
    .A2(io_pmp_6_mask[27]),
    .ZN(io_pmp_6_mask[28])
  );
  AND2_X1 _6949_ (
    .A1(reg_pmp_6_addr[26]),
    .A2(io_pmp_6_mask[28]),
    .ZN(io_pmp_6_mask[29])
  );
  AND2_X1 _6950_ (
    .A1(reg_pmp_6_addr[27]),
    .A2(io_pmp_6_mask[29]),
    .ZN(io_pmp_6_mask[30])
  );
  AND2_X1 _6951_ (
    .A1(reg_pmp_6_addr[28]),
    .A2(io_pmp_6_mask[30]),
    .ZN(io_pmp_6_mask[31])
  );
  AND2_X1 _6952_ (
    .A1(reg_pmp_7_cfg_a[0]),
    .A2(reg_pmp_7_addr[0]),
    .ZN(io_pmp_7_mask[3])
  );
  AND2_X1 _6953_ (
    .A1(reg_pmp_7_addr[1]),
    .A2(io_pmp_7_mask[3]),
    .ZN(io_pmp_7_mask[4])
  );
  AND2_X1 _6954_ (
    .A1(reg_pmp_7_addr[2]),
    .A2(io_pmp_7_mask[4]),
    .ZN(io_pmp_7_mask[5])
  );
  AND2_X1 _6955_ (
    .A1(reg_pmp_7_addr[3]),
    .A2(io_pmp_7_mask[5]),
    .ZN(io_pmp_7_mask[6])
  );
  AND2_X1 _6956_ (
    .A1(reg_pmp_7_addr[4]),
    .A2(io_pmp_7_mask[6]),
    .ZN(io_pmp_7_mask[7])
  );
  AND2_X1 _6957_ (
    .A1(reg_pmp_7_addr[5]),
    .A2(io_pmp_7_mask[7]),
    .ZN(io_pmp_7_mask[8])
  );
  AND2_X1 _6958_ (
    .A1(reg_pmp_7_addr[6]),
    .A2(io_pmp_7_mask[8]),
    .ZN(io_pmp_7_mask[9])
  );
  AND2_X1 _6959_ (
    .A1(reg_pmp_7_addr[7]),
    .A2(io_pmp_7_mask[9]),
    .ZN(io_pmp_7_mask[10])
  );
  AND2_X1 _6960_ (
    .A1(reg_pmp_7_addr[8]),
    .A2(io_pmp_7_mask[10]),
    .ZN(io_pmp_7_mask[11])
  );
  AND2_X1 _6961_ (
    .A1(reg_pmp_7_addr[9]),
    .A2(io_pmp_7_mask[11]),
    .ZN(io_pmp_7_mask[12])
  );
  AND2_X1 _6962_ (
    .A1(reg_pmp_7_addr[10]),
    .A2(io_pmp_7_mask[12]),
    .ZN(io_pmp_7_mask[13])
  );
  AND2_X1 _6963_ (
    .A1(reg_pmp_7_addr[11]),
    .A2(io_pmp_7_mask[13]),
    .ZN(io_pmp_7_mask[14])
  );
  AND2_X1 _6964_ (
    .A1(reg_pmp_7_addr[12]),
    .A2(io_pmp_7_mask[14]),
    .ZN(io_pmp_7_mask[15])
  );
  AND2_X1 _6965_ (
    .A1(reg_pmp_7_addr[13]),
    .A2(io_pmp_7_mask[15]),
    .ZN(io_pmp_7_mask[16])
  );
  AND2_X1 _6966_ (
    .A1(reg_pmp_7_addr[14]),
    .A2(io_pmp_7_mask[16]),
    .ZN(io_pmp_7_mask[17])
  );
  AND2_X1 _6967_ (
    .A1(reg_pmp_7_addr[15]),
    .A2(io_pmp_7_mask[17]),
    .ZN(io_pmp_7_mask[18])
  );
  AND2_X1 _6968_ (
    .A1(reg_pmp_7_addr[16]),
    .A2(io_pmp_7_mask[18]),
    .ZN(io_pmp_7_mask[19])
  );
  AND2_X1 _6969_ (
    .A1(reg_pmp_7_addr[17]),
    .A2(io_pmp_7_mask[19]),
    .ZN(io_pmp_7_mask[20])
  );
  AND2_X1 _6970_ (
    .A1(reg_pmp_7_addr[18]),
    .A2(io_pmp_7_mask[20]),
    .ZN(io_pmp_7_mask[21])
  );
  AND2_X1 _6971_ (
    .A1(reg_pmp_7_addr[19]),
    .A2(io_pmp_7_mask[21]),
    .ZN(io_pmp_7_mask[22])
  );
  AND2_X1 _6972_ (
    .A1(reg_pmp_7_addr[20]),
    .A2(io_pmp_7_mask[22]),
    .ZN(io_pmp_7_mask[23])
  );
  AND2_X1 _6973_ (
    .A1(reg_pmp_7_addr[21]),
    .A2(io_pmp_7_mask[23]),
    .ZN(io_pmp_7_mask[24])
  );
  AND2_X1 _6974_ (
    .A1(reg_pmp_7_addr[22]),
    .A2(io_pmp_7_mask[24]),
    .ZN(io_pmp_7_mask[25])
  );
  AND2_X1 _6975_ (
    .A1(reg_pmp_7_addr[23]),
    .A2(io_pmp_7_mask[25]),
    .ZN(io_pmp_7_mask[26])
  );
  AND2_X1 _6976_ (
    .A1(reg_pmp_7_addr[24]),
    .A2(io_pmp_7_mask[26]),
    .ZN(io_pmp_7_mask[27])
  );
  AND2_X1 _6977_ (
    .A1(reg_pmp_7_addr[25]),
    .A2(io_pmp_7_mask[27]),
    .ZN(io_pmp_7_mask[28])
  );
  AND2_X1 _6978_ (
    .A1(reg_pmp_7_addr[26]),
    .A2(io_pmp_7_mask[28]),
    .ZN(io_pmp_7_mask[29])
  );
  AND2_X1 _6979_ (
    .A1(reg_pmp_7_addr[27]),
    .A2(io_pmp_7_mask[29]),
    .ZN(io_pmp_7_mask[30])
  );
  AND2_X1 _6980_ (
    .A1(reg_pmp_7_addr[28]),
    .A2(io_pmp_7_mask[30]),
    .ZN(io_pmp_7_mask[31])
  );
  OR2_X1 _6981_ (
    .A1(io_decode_0_inst[26]),
    .A2(_0666_),
    .ZN(_4318_)
  );
  OR2_X1 _6982_ (
    .A1(_0664_),
    .A2(_4318_),
    .ZN(_4319_)
  );
  INV_X1 _6983_ (
    .A(_4319_),
    .ZN(_4320_)
  );
  OR2_X1 _6984_ (
    .A1(_4312_),
    .A2(_4319_),
    .ZN(_4321_)
  );
  AND2_X1 _6985_ (
    .A1(io_decode_0_inst[21]),
    .A2(io_decode_0_inst[20]),
    .ZN(_4322_)
  );
  INV_X1 _6986_ (
    .A(_4322_),
    .ZN(_4323_)
  );
  AND2_X1 _6987_ (
    .A1(io_decode_0_inst[24]),
    .A2(_4322_),
    .ZN(_4324_)
  );
  OR2_X1 _6988_ (
    .A1(_4321_),
    .A2(_4324_),
    .ZN(_4325_)
  );
  OR2_X1 _6989_ (
    .A1(io_decode_0_inst[21]),
    .A2(_0662_),
    .ZN(_4326_)
  );
  OR2_X1 _6990_ (
    .A1(_4312_),
    .A2(_4326_),
    .ZN(_4327_)
  );
  OR2_X1 _6991_ (
    .A1(_4310_),
    .A2(_4327_),
    .ZN(_4328_)
  );
  OR2_X1 _6992_ (
    .A1(_0666_),
    .A2(_4328_),
    .ZN(_4329_)
  );
  AND2_X1 _6993_ (
    .A1(io_decode_0_inst[30]),
    .A2(_4329_),
    .ZN(_4330_)
  );
  AND2_X1 _6994_ (
    .A1(_4325_),
    .A2(_4330_),
    .ZN(_4331_)
  );
  OR2_X1 _6995_ (
    .A1(_0658_),
    .A2(io_decode_0_inst[23]),
    .ZN(_4332_)
  );
  INV_X1 _6996_ (
    .A(_4332_),
    .ZN(_4333_)
  );
  MUX2_X1 _6997_ (
    .A(io_decode_0_inst[24]),
    .B(_4332_),
    .S(_0662_),
    .Z(_4334_)
  );
  OR2_X1 _6998_ (
    .A1(_0661_),
    .A2(_4334_),
    .ZN(_4335_)
  );
  OR2_X1 _6999_ (
    .A1(io_decode_0_inst[24]),
    .A2(_4313_),
    .ZN(_4336_)
  );
  OR2_X1 _7000_ (
    .A1(_0658_),
    .A2(_0663_),
    .ZN(_4337_)
  );
  OR2_X1 _7001_ (
    .A1(_4326_),
    .A2(_4337_),
    .ZN(_4338_)
  );
  AND2_X1 _7002_ (
    .A1(_4336_),
    .A2(_4338_),
    .ZN(_4339_)
  );
  AND2_X1 _7003_ (
    .A1(_4335_),
    .A2(_4339_),
    .ZN(_4340_)
  );
  OR2_X1 _7004_ (
    .A1(_0664_),
    .A2(_4340_),
    .ZN(_4341_)
  );
  OR2_X1 _7005_ (
    .A1(io_decode_0_inst[21]),
    .A2(io_decode_0_inst[20]),
    .ZN(_4342_)
  );
  INV_X1 _7006_ (
    .A(_4342_),
    .ZN(_4343_)
  );
  OR2_X1 _7007_ (
    .A1(io_decode_0_inst[23]),
    .A2(io_decode_0_inst[24]),
    .ZN(_4344_)
  );
  OR2_X1 _7008_ (
    .A1(_4342_),
    .A2(_4344_),
    .ZN(_4345_)
  );
  AND2_X1 _7009_ (
    .A1(_4341_),
    .A2(_4345_),
    .ZN(_4346_)
  );
  OR2_X1 _7010_ (
    .A1(io_decode_0_inst[26]),
    .A2(_4346_),
    .ZN(_4347_)
  );
  AND2_X1 _7011_ (
    .A1(io_decode_0_inst[22]),
    .A2(io_decode_0_inst[20]),
    .ZN(_4348_)
  );
  OR2_X1 _7012_ (
    .A1(io_decode_0_inst[21]),
    .A2(io_decode_0_inst[23]),
    .ZN(_4349_)
  );
  OR2_X1 _7013_ (
    .A1(_4309_),
    .A2(_4349_),
    .ZN(_4350_)
  );
  OR2_X1 _7014_ (
    .A1(_4348_),
    .A2(_4350_),
    .ZN(_4351_)
  );
  AND2_X1 _7015_ (
    .A1(_4347_),
    .A2(_4351_),
    .ZN(_4352_)
  );
  OR2_X1 _7016_ (
    .A1(io_decode_0_inst[27]),
    .A2(_4352_),
    .ZN(_4353_)
  );
  AND2_X1 _7017_ (
    .A1(io_decode_0_inst[24]),
    .A2(_4320_),
    .ZN(_4354_)
  );
  OR2_X1 _7018_ (
    .A1(_0665_),
    .A2(_4319_),
    .ZN(_4355_)
  );
  OR2_X1 _7019_ (
    .A1(_4326_),
    .A2(_4332_),
    .ZN(_4356_)
  );
  OR2_X1 _7020_ (
    .A1(_4309_),
    .A2(_4317_),
    .ZN(_4357_)
  );
  OR2_X1 _7021_ (
    .A1(_4356_),
    .A2(_4357_),
    .ZN(_4358_)
  );
  OR2_X1 _7022_ (
    .A1(_0664_),
    .A2(_4317_),
    .ZN(_4359_)
  );
  OR2_X1 _7023_ (
    .A1(_0665_),
    .A2(_4359_),
    .ZN(_4360_)
  );
  OR2_X1 _7024_ (
    .A1(io_decode_0_inst[21]),
    .A2(_4332_),
    .ZN(_4361_)
  );
  OR2_X1 _7025_ (
    .A1(_4360_),
    .A2(_4361_),
    .ZN(_4362_)
  );
  AND2_X1 _7026_ (
    .A1(_4358_),
    .A2(_4362_),
    .ZN(_4363_)
  );
  AND2_X1 _7027_ (
    .A1(_4355_),
    .A2(_4363_),
    .ZN(_4364_)
  );
  OR2_X1 _7028_ (
    .A1(io_decode_0_inst[20]),
    .A2(_0663_),
    .ZN(_4365_)
  );
  AND2_X1 _7029_ (
    .A1(io_decode_0_inst[22]),
    .A2(_4323_),
    .ZN(_4366_)
  );
  AND2_X1 _7030_ (
    .A1(_4365_),
    .A2(_4366_),
    .ZN(_4367_)
  );
  OR2_X1 _7031_ (
    .A1(_4360_),
    .A2(_4367_),
    .ZN(_4368_)
  );
  OR2_X1 _7032_ (
    .A1(_4311_),
    .A2(_4316_),
    .ZN(_4369_)
  );
  AND2_X1 _7033_ (
    .A1(_0667_),
    .A2(_4321_),
    .ZN(_4370_)
  );
  AND2_X1 _7034_ (
    .A1(_4369_),
    .A2(_4370_),
    .ZN(_4371_)
  );
  AND2_X1 _7035_ (
    .A1(_4368_),
    .A2(_4371_),
    .ZN(_4372_)
  );
  AND2_X1 _7036_ (
    .A1(_4364_),
    .A2(_4372_),
    .ZN(_4373_)
  );
  AND2_X1 _7037_ (
    .A1(_4353_),
    .A2(_4373_),
    .ZN(_4374_)
  );
  OR2_X1 _7038_ (
    .A1(_4331_),
    .A2(_4374_),
    .ZN(_4375_)
  );
  AND2_X1 _7039_ (
    .A1(_0660_),
    .A2(_4375_),
    .ZN(_4376_)
  );
  OR2_X1 _7040_ (
    .A1(_4332_),
    .A2(_4342_),
    .ZN(_4377_)
  );
  OR2_X1 _7041_ (
    .A1(io_decode_0_inst[25]),
    .A2(_0665_),
    .ZN(_4378_)
  );
  OR2_X1 _7042_ (
    .A1(io_decode_0_inst[26]),
    .A2(_4378_),
    .ZN(_4379_)
  );
  OR2_X1 _7043_ (
    .A1(_4317_),
    .A2(_4378_),
    .ZN(_4380_)
  );
  OR2_X1 _7044_ (
    .A1(_4377_),
    .A2(_4380_),
    .ZN(_4381_)
  );
  AND2_X1 _7045_ (
    .A1(io_decode_0_inst[30]),
    .A2(_4381_),
    .ZN(_4382_)
  );
  OR2_X1 _7046_ (
    .A1(_4312_),
    .A2(_4343_),
    .ZN(_4383_)
  );
  AND2_X1 _7047_ (
    .A1(_4377_),
    .A2(_4383_),
    .ZN(_4384_)
  );
  OR2_X1 _7048_ (
    .A1(_0666_),
    .A2(_4384_),
    .ZN(_4385_)
  );
  OR2_X1 _7049_ (
    .A1(_4312_),
    .A2(_4342_),
    .ZN(_4386_)
  );
  AND2_X1 _7050_ (
    .A1(io_decode_0_inst[22]),
    .A2(_4322_),
    .ZN(_4387_)
  );
  OR2_X1 _7051_ (
    .A1(_0663_),
    .A2(_4387_),
    .ZN(_4388_)
  );
  AND2_X1 _7052_ (
    .A1(_4386_),
    .A2(_4388_),
    .ZN(_4389_)
  );
  AND2_X1 _7053_ (
    .A1(_4385_),
    .A2(_4389_),
    .ZN(_4390_)
  );
  OR2_X1 _7054_ (
    .A1(_4378_),
    .A2(_4390_),
    .ZN(_4391_)
  );
  AND2_X1 _7055_ (
    .A1(_4333_),
    .A2(_4342_),
    .ZN(_4392_)
  );
  OR2_X1 _7056_ (
    .A1(_4312_),
    .A2(_4322_),
    .ZN(_4393_)
  );
  INV_X1 _7057_ (
    .A(_4393_),
    .ZN(_4394_)
  );
  OR2_X1 _7058_ (
    .A1(_4309_),
    .A2(_4394_),
    .ZN(_4395_)
  );
  OR2_X1 _7059_ (
    .A1(_4392_),
    .A2(_4395_),
    .ZN(_4396_)
  );
  OR2_X1 _7060_ (
    .A1(io_decode_0_inst[25]),
    .A2(_4356_),
    .ZN(_4397_)
  );
  OR2_X1 _7061_ (
    .A1(io_decode_0_inst[20]),
    .A2(_4309_),
    .ZN(_4398_)
  );
  OR2_X1 _7062_ (
    .A1(_4312_),
    .A2(_4398_),
    .ZN(_4399_)
  );
  AND2_X1 _7063_ (
    .A1(_4397_),
    .A2(_4399_),
    .ZN(_4400_)
  );
  AND2_X1 _7064_ (
    .A1(_4396_),
    .A2(_4400_),
    .ZN(_4401_)
  );
  AND2_X1 _7065_ (
    .A1(_4391_),
    .A2(_4401_),
    .ZN(_4402_)
  );
  OR2_X1 _7066_ (
    .A1(io_decode_0_inst[26]),
    .A2(_4402_),
    .ZN(_4403_)
  );
  OR2_X1 _7067_ (
    .A1(io_decode_0_inst[26]),
    .A2(io_decode_0_inst[25]),
    .ZN(_4404_)
  );
  OR2_X1 _7068_ (
    .A1(_4332_),
    .A2(_4404_),
    .ZN(_4405_)
  );
  OR2_X1 _7069_ (
    .A1(_0661_),
    .A2(_4405_),
    .ZN(_4406_)
  );
  OR2_X1 _7070_ (
    .A1(_4323_),
    .A2(_4337_),
    .ZN(_4407_)
  );
  OR2_X1 _7071_ (
    .A1(_4379_),
    .A2(_4407_),
    .ZN(_4408_)
  );
  AND2_X1 _7072_ (
    .A1(_4381_),
    .A2(_4408_),
    .ZN(_4409_)
  );
  AND2_X1 _7073_ (
    .A1(_4406_),
    .A2(_4409_),
    .ZN(_4410_)
  );
  AND2_X1 _7074_ (
    .A1(_4403_),
    .A2(_4410_),
    .ZN(_4411_)
  );
  OR2_X1 _7075_ (
    .A1(_4382_),
    .A2(_4411_),
    .ZN(_4412_)
  );
  OR2_X1 _7076_ (
    .A1(_4380_),
    .A2(_4383_),
    .ZN(_4413_)
  );
  AND2_X1 _7077_ (
    .A1(io_decode_0_inst[31]),
    .A2(_4413_),
    .ZN(_4414_)
  );
  AND2_X1 _7078_ (
    .A1(_4412_),
    .A2(_4414_),
    .ZN(_4415_)
  );
  AND2_X1 _7079_ (
    .A1(io_decode_0_inst[29]),
    .A2(io_decode_0_inst[28]),
    .ZN(_4416_)
  );
  INV_X1 _7080_ (
    .A(_4416_),
    .ZN(_4417_)
  );
  AND2_X1 _7081_ (
    .A1(_0660_),
    .A2(io_decode_0_inst[30]),
    .ZN(_4418_)
  );
  AND2_X1 _7082_ (
    .A1(_io_decode_0_read_illegal_T_15),
    .A2(_4416_),
    .ZN(_4419_)
  );
  AND2_X1 _7083_ (
    .A1(_4418_),
    .A2(_4419_),
    .ZN(_4420_)
  );
  AND2_X1 _7084_ (
    .A1(_4354_),
    .A2(_4420_),
    .ZN(_4421_)
  );
  OR2_X1 _7085_ (
    .A1(_4417_),
    .A2(_4421_),
    .ZN(_4422_)
  );
  OR2_X1 _7086_ (
    .A1(_4415_),
    .A2(_4422_),
    .ZN(_4423_)
  );
  OR2_X1 _7087_ (
    .A1(_4376_),
    .A2(_4423_),
    .ZN(io_decode_0_read_illegal)
  );
  AND2_X1 _7088_ (
    .A1(io_decode_0_inst[27]),
    .A2(_io_decode_0_read_illegal_T_15),
    .ZN(_4424_)
  );
  AND2_X1 _7089_ (
    .A1(_4418_),
    .A2(_4424_),
    .ZN(io_decode_0_system_illegal)
  );
  AND2_X1 _7090_ (
    .A1(_2467_),
    .A2(_2511_),
    .ZN(_4425_)
  );
  INV_X1 _7091_ (
    .A(_4425_),
    .ZN(io_eret)
  );
  AND2_X1 _7092_ (
    .A1(_2456_),
    .A2(io_interrupt_cause[1]),
    .ZN(_4426_)
  );
  OR2_X1 _7093_ (
    .A1(reg_singleStepped),
    .A2(_4426_),
    .ZN(_4427_)
  );
  OR2_X1 _7094_ (
    .A1(reg_debug),
    .A2(io_status_cease_r),
    .ZN(_4428_)
  );
  INV_X1 _7095_ (
    .A(_4428_),
    .ZN(_4429_)
  );
  AND2_X1 _7096_ (
    .A1(_4427_),
    .A2(_4429_),
    .ZN(io_interrupt)
  );
  INV_X1 _7097_ (
    .A(large_[16]),
    .ZN(_0622_)
  );
  INV_X1 _7098_ (
    .A(large_[15]),
    .ZN(_0623_)
  );
  INV_X1 _7099_ (
    .A(large_[14]),
    .ZN(_0624_)
  );
  INV_X1 _7100_ (
    .A(large_[13]),
    .ZN(_0625_)
  );
  INV_X1 _7101_ (
    .A(large_1[23]),
    .ZN(_0626_)
  );
  INV_X1 _7102_ (
    .A(large_1[22]),
    .ZN(_0627_)
  );
  INV_X1 _7103_ (
    .A(large_1[20]),
    .ZN(_0628_)
  );
  INV_X1 _7104_ (
    .A(large_1[14]),
    .ZN(_0629_)
  );
  INV_X1 _7105_ (
    .A(large_1[11]),
    .ZN(_0630_)
  );
  INV_X1 _7106_ (
    .A(large_1[10]),
    .ZN(_0631_)
  );
  INV_X1 _7107_ (
    .A(large_1[9]),
    .ZN(_0632_)
  );
  INV_X1 _7108_ (
    .A(large_[50]),
    .ZN(_0633_)
  );
  INV_X1 _7109_ (
    .A(large_[47]),
    .ZN(_0634_)
  );
  INV_X1 _7110_ (
    .A(large_[28]),
    .ZN(_0635_)
  );
  INV_X1 _7111_ (
    .A(small_1[5]),
    .ZN(_0636_)
  );
  INV_X1 _7112_ (
    .A(small_1[4]),
    .ZN(_0637_)
  );
  INV_X1 _7113_ (
    .A(small_1[3]),
    .ZN(_0638_)
  );
  INV_X1 _7114_ (
    .A(small_1[2]),
    .ZN(_0639_)
  );
  INV_X1 _7115_ (
    .A(small_1[1]),
    .ZN(_0640_)
  );
  INV_X1 _7116_ (
    .A(small_1[0]),
    .ZN(_0641_)
  );
  INV_X1 _7117_ (
    .A(large_1[57]),
    .ZN(_0642_)
  );
  INV_X1 _7118_ (
    .A(large_1[56]),
    .ZN(_0643_)
  );
  INV_X1 _7119_ (
    .A(large_1[55]),
    .ZN(_0644_)
  );
  INV_X1 _7120_ (
    .A(large_1[54]),
    .ZN(_0645_)
  );
  INV_X1 _7121_ (
    .A(large_1[53]),
    .ZN(_0646_)
  );
  INV_X1 _7122_ (
    .A(large_1[52]),
    .ZN(_0647_)
  );
  INV_X1 _7123_ (
    .A(large_1[51]),
    .ZN(_0648_)
  );
  INV_X1 _7124_ (
    .A(large_1[50]),
    .ZN(_0649_)
  );
  INV_X1 _7125_ (
    .A(large_1[49]),
    .ZN(_0650_)
  );
  INV_X1 _7126_ (
    .A(large_1[48]),
    .ZN(_0651_)
  );
  INV_X1 _7127_ (
    .A(reg_mcountinhibit[2]),
    .ZN(_0652_)
  );
  INV_X1 _7128_ (
    .A(reg_singleStepped),
    .ZN(_0653_)
  );
  INV_X1 _7129_ (
    .A(reset),
    .ZN(_0654_)
  );
  INV_X1 _7130_ (
    .A(io_rw_cmd[1]),
    .ZN(_0655_)
  );
  INV_X1 _7131_ (
    .A(io_rw_cmd[2]),
    .ZN(_0656_)
  );
  INV_X1 _7132_ (
    .A(io_rw_cmd[0]),
    .ZN(_0657_)
  );
  INV_X1 _7133_ (
    .A(io_decode_0_inst[22]),
    .ZN(_0658_)
  );
  INV_X1 _7134_ (
    .A(io_decode_0_inst[26]),
    .ZN(_0659_)
  );
  INV_X1 _7135_ (
    .A(io_decode_0_inst[31]),
    .ZN(_0660_)
  );
  INV_X1 _7136_ (
    .A(io_decode_0_inst[21]),
    .ZN(_0661_)
  );
  INV_X1 _7137_ (
    .A(io_decode_0_inst[20]),
    .ZN(_0662_)
  );
  INV_X1 _7138_ (
    .A(io_decode_0_inst[23]),
    .ZN(_0663_)
  );
  INV_X1 _7139_ (
    .A(io_decode_0_inst[25]),
    .ZN(_0664_)
  );
  INV_X1 _7140_ (
    .A(io_decode_0_inst[24]),
    .ZN(_0665_)
  );
  INV_X1 _7141_ (
    .A(io_decode_0_inst[27]),
    .ZN(_0666_)
  );
  INV_X1 _7142_ (
    .A(io_decode_0_inst[30]),
    .ZN(_0667_)
  );
  INV_X1 _7143_ (
    .A(io_rw_addr[6]),
    .ZN(_0668_)
  );
  INV_X1 _7144_ (
    .A(io_rw_addr[5]),
    .ZN(_0669_)
  );
  INV_X1 _7145_ (
    .A(io_rw_addr[4]),
    .ZN(_0670_)
  );
  INV_X1 _7146_ (
    .A(io_rw_addr[1]),
    .ZN(_0671_)
  );
  INV_X1 _7147_ (
    .A(io_rw_addr[10]),
    .ZN(_0672_)
  );
  INV_X1 _7148_ (
    .A(io_rw_addr[7]),
    .ZN(_0673_)
  );
  INV_X1 _7149_ (
    .A(io_rw_addr[11]),
    .ZN(_0674_)
  );
  INV_X1 _7150_ (
    .A(io_rw_addr[0]),
    .ZN(_0675_)
  );
  INV_X1 _7151_ (
    .A(reg_mstatus_mie),
    .ZN(_0676_)
  );
  INV_X1 _7152_ (
    .A(io_interrupts_debug),
    .ZN(_0677_)
  );
  INV_X1 _7153_ (
    .A(io_rw_wdata[0]),
    .ZN(_0678_)
  );
  INV_X1 _7154_ (
    .A(io_rw_wdata[1]),
    .ZN(_0679_)
  );
  INV_X1 _7155_ (
    .A(io_rw_wdata[2]),
    .ZN(_0680_)
  );
  INV_X1 _7156_ (
    .A(io_rw_wdata[3]),
    .ZN(_0681_)
  );
  INV_X1 _7157_ (
    .A(io_rw_wdata[4]),
    .ZN(_0682_)
  );
  INV_X1 _7158_ (
    .A(io_rw_wdata[5]),
    .ZN(_0683_)
  );
  INV_X1 _7159_ (
    .A(io_rw_wdata[6]),
    .ZN(_0684_)
  );
  INV_X1 _7160_ (
    .A(io_rw_wdata[7]),
    .ZN(_0685_)
  );
  INV_X1 _7161_ (
    .A(io_rw_wdata[8]),
    .ZN(_0686_)
  );
  INV_X1 _7162_ (
    .A(io_rw_wdata[9]),
    .ZN(_0687_)
  );
  INV_X1 _7163_ (
    .A(io_rw_wdata[10]),
    .ZN(_0688_)
  );
  INV_X1 _7164_ (
    .A(io_rw_wdata[11]),
    .ZN(_0689_)
  );
  INV_X1 _7165_ (
    .A(io_rw_wdata[13]),
    .ZN(_0690_)
  );
  INV_X1 _7166_ (
    .A(io_rw_wdata[14]),
    .ZN(_0691_)
  );
  INV_X1 _7167_ (
    .A(io_rw_wdata[15]),
    .ZN(_0692_)
  );
  INV_X1 _7168_ (
    .A(io_rw_wdata[16]),
    .ZN(_0693_)
  );
  INV_X1 _7169_ (
    .A(io_rw_wdata[17]),
    .ZN(_0694_)
  );
  INV_X1 _7170_ (
    .A(io_rw_wdata[18]),
    .ZN(_0695_)
  );
  INV_X1 _7171_ (
    .A(io_rw_wdata[19]),
    .ZN(_0696_)
  );
  INV_X1 _7172_ (
    .A(io_rw_wdata[20]),
    .ZN(_0697_)
  );
  INV_X1 _7173_ (
    .A(io_rw_wdata[21]),
    .ZN(_0698_)
  );
  INV_X1 _7174_ (
    .A(io_rw_wdata[22]),
    .ZN(_0699_)
  );
  INV_X1 _7175_ (
    .A(io_rw_wdata[23]),
    .ZN(_0700_)
  );
  INV_X1 _7176_ (
    .A(io_rw_wdata[24]),
    .ZN(_0701_)
  );
  INV_X1 _7177_ (
    .A(io_rw_wdata[25]),
    .ZN(_0702_)
  );
  INV_X1 _7178_ (
    .A(io_rw_wdata[26]),
    .ZN(_0703_)
  );
  INV_X1 _7179_ (
    .A(io_rw_wdata[27]),
    .ZN(_0704_)
  );
  INV_X1 _7180_ (
    .A(io_rw_wdata[28]),
    .ZN(_0705_)
  );
  INV_X1 _7181_ (
    .A(io_rw_wdata[29]),
    .ZN(_0706_)
  );
  INV_X1 _7182_ (
    .A(io_rw_wdata[30]),
    .ZN(_0707_)
  );
  INV_X1 _7183_ (
    .A(io_rw_wdata[31]),
    .ZN(_0708_)
  );
  INV_X1 _7184_ (
    .A(io_cause[4]),
    .ZN(_0709_)
  );
  INV_X1 _7185_ (
    .A(io_rw_addr[3]),
    .ZN(_0710_)
  );
  INV_X1 _7186_ (
    .A(_T_15),
    .ZN(_0711_)
  );
  INV_X1 _7187_ (
    .A(_T_18[1]),
    .ZN(_0712_)
  );
  INV_X1 _7188_ (
    .A(_GEN_586[1]),
    .ZN(_0713_)
  );
  INV_X1 _7189_ (
    .A(_T_24[1]),
    .ZN(_0714_)
  );
  INV_X1 _7190_ (
    .A(io_exception),
    .ZN(_0715_)
  );
  OR2_X1 _7191_ (
    .A1(io_rw_addr[2]),
    .A2(io_rw_addr[3]),
    .ZN(_0716_)
  );
  INV_X1 _7192_ (
    .A(_0716_),
    .ZN(_0717_)
  );
  AND2_X1 _7193_ (
    .A1(_0671_),
    .A2(_0717_),
    .ZN(_0718_)
  );
  OR2_X1 _7194_ (
    .A1(io_rw_addr[1]),
    .A2(_0716_),
    .ZN(_0719_)
  );
  AND2_X1 _7195_ (
    .A1(io_rw_addr[0]),
    .A2(_0718_),
    .ZN(_0720_)
  );
  OR2_X1 _7196_ (
    .A1(_0675_),
    .A2(_0719_),
    .ZN(_0721_)
  );
  OR2_X1 _7197_ (
    .A1(io_rw_addr[10]),
    .A2(io_rw_addr[11]),
    .ZN(_0722_)
  );
  INV_X1 _7198_ (
    .A(_0722_),
    .ZN(_0723_)
  );
  AND2_X1 _7199_ (
    .A1(io_rw_addr[8]),
    .A2(io_rw_addr[9]),
    .ZN(_0724_)
  );
  AND2_X1 _7200_ (
    .A1(io_rw_addr[8]),
    .A2(_0723_),
    .ZN(_0725_)
  );
  AND2_X1 _7201_ (
    .A1(_0723_),
    .A2(_0724_),
    .ZN(_0726_)
  );
  AND2_X1 _7202_ (
    .A1(_0668_),
    .A2(io_rw_addr[7]),
    .ZN(_0727_)
  );
  AND2_X1 _7203_ (
    .A1(io_rw_addr[5]),
    .A2(_0670_),
    .ZN(_0728_)
  );
  AND2_X1 _7204_ (
    .A1(_0727_),
    .A2(_0728_),
    .ZN(_0729_)
  );
  AND2_X1 _7205_ (
    .A1(_0726_),
    .A2(_0728_),
    .ZN(_0730_)
  );
  INV_X1 _7206_ (
    .A(_0730_),
    .ZN(_0731_)
  );
  AND2_X1 _7207_ (
    .A1(_0726_),
    .A2(_0729_),
    .ZN(_0732_)
  );
  AND2_X1 _7208_ (
    .A1(_0720_),
    .A2(_0732_),
    .ZN(_0733_)
  );
  AND2_X1 _7209_ (
    .A1(_0655_),
    .A2(_0657_),
    .ZN(_0734_)
  );
  OR2_X1 _7210_ (
    .A1(io_rw_cmd[1]),
    .A2(io_rw_cmd[0]),
    .ZN(_0735_)
  );
  AND2_X1 _7211_ (
    .A1(io_rw_cmd[2]),
    .A2(_0735_),
    .ZN(_0736_)
  );
  OR2_X1 _7212_ (
    .A1(_0656_),
    .A2(_0734_),
    .ZN(_0737_)
  );
  AND2_X1 _7213_ (
    .A1(_0017_),
    .A2(_0733_),
    .ZN(_0738_)
  );
  INV_X1 _7214_ (
    .A(_0738_),
    .ZN(_0739_)
  );
  AND2_X1 _7215_ (
    .A1(_0736_),
    .A2(_0738_),
    .ZN(_0740_)
  );
  OR2_X1 _7216_ (
    .A1(_0737_),
    .A2(_0739_),
    .ZN(_0741_)
  );
  OR2_X1 _7217_ (
    .A1(_0655_),
    .A2(_0657_),
    .ZN(_0742_)
  );
  AND2_X1 _7218_ (
    .A1(io_rw_wdata[16]),
    .A2(_0742_),
    .ZN(_0743_)
  );
  AND2_X1 _7219_ (
    .A1(io_rw_addr[5]),
    .A2(io_rw_addr[4]),
    .ZN(_0744_)
  );
  AND2_X1 _7220_ (
    .A1(_0727_),
    .A2(_0744_),
    .ZN(_0745_)
  );
  AND2_X1 _7221_ (
    .A1(io_rw_addr[10]),
    .A2(_0674_),
    .ZN(_0746_)
  );
  OR2_X1 _7222_ (
    .A1(_0672_),
    .A2(io_rw_addr[11]),
    .ZN(_0747_)
  );
  AND2_X1 _7223_ (
    .A1(_0724_),
    .A2(_0746_),
    .ZN(_0748_)
  );
  AND2_X1 _7224_ (
    .A1(_0745_),
    .A2(_0748_),
    .ZN(_0749_)
  );
  AND2_X1 _7225_ (
    .A1(_0720_),
    .A2(_0749_),
    .ZN(_0750_)
  );
  INV_X1 _7226_ (
    .A(_0750_),
    .ZN(_0751_)
  );
  AND2_X1 _7227_ (
    .A1(reg_dpc[16]),
    .A2(_0750_),
    .ZN(_0752_)
  );
  AND2_X1 _7228_ (
    .A1(_0675_),
    .A2(_0718_),
    .ZN(_0753_)
  );
  AND2_X1 _7229_ (
    .A1(_0732_),
    .A2(_0753_),
    .ZN(_0754_)
  );
  AND2_X1 _7230_ (
    .A1(reg_pmp_2_cfg_r),
    .A2(_0754_),
    .ZN(_0755_)
  );
  OR2_X1 _7231_ (
    .A1(_0752_),
    .A2(_0755_),
    .ZN(_0756_)
  );
  OR2_X1 _7232_ (
    .A1(io_rw_addr[5]),
    .A2(io_rw_addr[4]),
    .ZN(_0757_)
  );
  INV_X1 _7233_ (
    .A(_0757_),
    .ZN(_0758_)
  );
  AND2_X1 _7234_ (
    .A1(io_rw_addr[6]),
    .A2(_0673_),
    .ZN(_0759_)
  );
  AND2_X1 _7235_ (
    .A1(_0758_),
    .A2(_0759_),
    .ZN(_0760_)
  );
  AND2_X1 _7236_ (
    .A1(_0726_),
    .A2(_0760_),
    .ZN(_0761_)
  );
  AND2_X1 _7237_ (
    .A1(io_rw_addr[1]),
    .A2(_0717_),
    .ZN(_0762_)
  );
  AND2_X1 _7238_ (
    .A1(io_rw_addr[0]),
    .A2(_0762_),
    .ZN(_0763_)
  );
  AND2_X1 _7239_ (
    .A1(_0761_),
    .A2(_0763_),
    .ZN(_0764_)
  );
  INV_X1 _7240_ (
    .A(_0764_),
    .ZN(_0765_)
  );
  AND2_X1 _7241_ (
    .A1(reg_mtval[16]),
    .A2(_0764_),
    .ZN(_0766_)
  );
  AND2_X1 _7242_ (
    .A1(_0753_),
    .A2(_0761_),
    .ZN(_0767_)
  );
  AND2_X1 _7243_ (
    .A1(reg_mscratch[16]),
    .A2(_0767_),
    .ZN(_0768_)
  );
  OR2_X1 _7244_ (
    .A1(_0766_),
    .A2(_0768_),
    .ZN(_0769_)
  );
  OR2_X1 _7245_ (
    .A1(_0756_),
    .A2(_0769_),
    .ZN(_0770_)
  );
  AND2_X1 _7246_ (
    .A1(_0668_),
    .A2(_0673_),
    .ZN(_0771_)
  );
  OR2_X1 _7247_ (
    .A1(io_rw_addr[6]),
    .A2(io_rw_addr[7]),
    .ZN(_0772_)
  );
  AND2_X1 _7248_ (
    .A1(_0758_),
    .A2(_0771_),
    .ZN(_0773_)
  );
  OR2_X1 _7249_ (
    .A1(_0757_),
    .A2(_0772_),
    .ZN(_0774_)
  );
  AND2_X1 _7250_ (
    .A1(_0726_),
    .A2(_0773_),
    .ZN(_0775_)
  );
  INV_X1 _7251_ (
    .A(_0775_),
    .ZN(_0776_)
  );
  AND2_X1 _7252_ (
    .A1(io_rw_addr[2]),
    .A2(_0710_),
    .ZN(_0777_)
  );
  AND2_X1 _7253_ (
    .A1(io_rw_addr[0]),
    .A2(_0777_),
    .ZN(_0778_)
  );
  AND2_X1 _7254_ (
    .A1(_0671_),
    .A2(_0778_),
    .ZN(_0779_)
  );
  AND2_X1 _7255_ (
    .A1(_0775_),
    .A2(_0779_),
    .ZN(_0780_)
  );
  INV_X1 _7256_ (
    .A(_0780_),
    .ZN(_0781_)
  );
  AND2_X1 _7257_ (
    .A1(reg_mtvec[16]),
    .A2(_0780_),
    .ZN(_0782_)
  );
  AND2_X1 _7258_ (
    .A1(_0720_),
    .A2(_0761_),
    .ZN(_0783_)
  );
  INV_X1 _7259_ (
    .A(_0783_),
    .ZN(_0784_)
  );
  AND2_X1 _7260_ (
    .A1(reg_mepc[16]),
    .A2(_0783_),
    .ZN(_0785_)
  );
  OR2_X1 _7261_ (
    .A1(_0782_),
    .A2(_0785_),
    .ZN(_0786_)
  );
  AND2_X1 _7262_ (
    .A1(_0726_),
    .A2(_0745_),
    .ZN(_0787_)
  );
  AND2_X1 _7263_ (
    .A1(_0779_),
    .A2(_0787_),
    .ZN(_0788_)
  );
  INV_X1 _7264_ (
    .A(_0788_),
    .ZN(_0789_)
  );
  AND2_X1 _7265_ (
    .A1(reg_pmp_5_addr[16]),
    .A2(_0788_),
    .ZN(_0790_)
  );
  AND2_X1 _7266_ (
    .A1(_0675_),
    .A2(_0762_),
    .ZN(_0791_)
  );
  AND2_X1 _7267_ (
    .A1(_0787_),
    .A2(_0791_),
    .ZN(_0792_)
  );
  INV_X1 _7268_ (
    .A(_0792_),
    .ZN(_0793_)
  );
  AND2_X1 _7269_ (
    .A1(reg_pmp_2_addr[16]),
    .A2(_0792_),
    .ZN(_0794_)
  );
  OR2_X1 _7270_ (
    .A1(_0790_),
    .A2(_0794_),
    .ZN(_0795_)
  );
  OR2_X1 _7271_ (
    .A1(_0786_),
    .A2(_0795_),
    .ZN(_0796_)
  );
  AND2_X1 _7272_ (
    .A1(_0749_),
    .A2(_0762_),
    .ZN(_0797_)
  );
  AND2_X1 _7273_ (
    .A1(reg_dscratch0[16]),
    .A2(_0797_),
    .ZN(_0798_)
  );
  AND2_X1 _7274_ (
    .A1(_0729_),
    .A2(_0748_),
    .ZN(_0799_)
  );
  AND2_X1 _7275_ (
    .A1(_0791_),
    .A2(_0799_),
    .ZN(_0800_)
  );
  AND2_X1 _7276_ (
    .A1(reg_bp_0_address[16]),
    .A2(_0800_),
    .ZN(_0801_)
  );
  OR2_X1 _7277_ (
    .A1(_0798_),
    .A2(_0801_),
    .ZN(_0802_)
  );
  AND2_X1 _7278_ (
    .A1(_0675_),
    .A2(_0777_),
    .ZN(_0803_)
  );
  AND2_X1 _7279_ (
    .A1(_0671_),
    .A2(_0803_),
    .ZN(_0804_)
  );
  AND2_X1 _7280_ (
    .A1(_0787_),
    .A2(_0804_),
    .ZN(_0805_)
  );
  INV_X1 _7281_ (
    .A(_0805_),
    .ZN(_0806_)
  );
  AND2_X1 _7282_ (
    .A1(reg_pmp_4_addr[16]),
    .A2(_0805_),
    .ZN(_0807_)
  );
  AND2_X1 _7283_ (
    .A1(reg_pmp_6_cfg_r),
    .A2(_0733_),
    .ZN(_0808_)
  );
  OR2_X1 _7284_ (
    .A1(_0807_),
    .A2(_0808_),
    .ZN(_0809_)
  );
  OR2_X1 _7285_ (
    .A1(_0802_),
    .A2(_0809_),
    .ZN(_0810_)
  );
  OR2_X1 _7286_ (
    .A1(_0796_),
    .A2(_0810_),
    .ZN(_0811_)
  );
  OR2_X1 _7287_ (
    .A1(_0770_),
    .A2(_0811_),
    .ZN(_0812_)
  );
  AND2_X1 _7288_ (
    .A1(io_rw_addr[1]),
    .A2(_0787_),
    .ZN(_0813_)
  );
  AND2_X1 _7289_ (
    .A1(_0803_),
    .A2(_0813_),
    .ZN(_0814_)
  );
  INV_X1 _7290_ (
    .A(_0814_),
    .ZN(_0815_)
  );
  AND2_X1 _7291_ (
    .A1(reg_pmp_6_addr[16]),
    .A2(_0814_),
    .ZN(_0816_)
  );
  AND2_X1 _7292_ (
    .A1(io_rw_addr[11]),
    .A2(_0724_),
    .ZN(_0817_)
  );
  OR2_X1 _7293_ (
    .A1(io_rw_addr[10]),
    .A2(_0757_),
    .ZN(_0818_)
  );
  INV_X1 _7294_ (
    .A(_0818_),
    .ZN(_0819_)
  );
  AND2_X1 _7295_ (
    .A1(_0817_),
    .A2(_0819_),
    .ZN(_0820_)
  );
  AND2_X1 _7296_ (
    .A1(_0771_),
    .A2(_0820_),
    .ZN(_0821_)
  );
  AND2_X1 _7297_ (
    .A1(_0791_),
    .A2(_0821_),
    .ZN(_0822_)
  );
  AND2_X1 _7298_ (
    .A1(large_[10]),
    .A2(_0822_),
    .ZN(_0823_)
  );
  OR2_X1 _7299_ (
    .A1(_0816_),
    .A2(_0823_),
    .ZN(_0824_)
  );
  AND2_X1 _7300_ (
    .A1(_0672_),
    .A2(_0817_),
    .ZN(_0825_)
  );
  AND2_X1 _7301_ (
    .A1(_0727_),
    .A2(_0820_),
    .ZN(_0826_)
  );
  AND2_X1 _7302_ (
    .A1(_0791_),
    .A2(_0826_),
    .ZN(_0827_)
  );
  INV_X1 _7303_ (
    .A(_0827_),
    .ZN(_0828_)
  );
  AND2_X1 _7304_ (
    .A1(large_[42]),
    .A2(_0827_),
    .ZN(_0829_)
  );
  AND2_X1 _7305_ (
    .A1(_0718_),
    .A2(_0821_),
    .ZN(_0830_)
  );
  AND2_X1 _7306_ (
    .A1(large_1[10]),
    .A2(_0830_),
    .ZN(_0831_)
  );
  OR2_X1 _7307_ (
    .A1(_0829_),
    .A2(_0831_),
    .ZN(_0832_)
  );
  OR2_X1 _7308_ (
    .A1(_0824_),
    .A2(_0832_),
    .ZN(_0833_)
  );
  AND2_X1 _7309_ (
    .A1(_0761_),
    .A2(_0791_),
    .ZN(_0834_)
  );
  INV_X1 _7310_ (
    .A(_0834_),
    .ZN(_0835_)
  );
  AND2_X1 _7311_ (
    .A1(reg_mcause[16]),
    .A2(_0834_),
    .ZN(_0836_)
  );
  AND2_X1 _7312_ (
    .A1(_0753_),
    .A2(_0787_),
    .ZN(_0837_)
  );
  INV_X1 _7313_ (
    .A(_0837_),
    .ZN(_0838_)
  );
  AND2_X1 _7314_ (
    .A1(reg_pmp_0_addr[16]),
    .A2(_0837_),
    .ZN(_0839_)
  );
  OR2_X1 _7315_ (
    .A1(_0836_),
    .A2(_0839_),
    .ZN(_0840_)
  );
  AND2_X1 _7316_ (
    .A1(_0720_),
    .A2(_0787_),
    .ZN(_0841_)
  );
  INV_X1 _7317_ (
    .A(_0841_),
    .ZN(_0842_)
  );
  AND2_X1 _7318_ (
    .A1(reg_pmp_1_addr[16]),
    .A2(_0841_),
    .ZN(_0843_)
  );
  AND2_X1 _7319_ (
    .A1(_0763_),
    .A2(_0787_),
    .ZN(_0844_)
  );
  INV_X1 _7320_ (
    .A(_0844_),
    .ZN(_0845_)
  );
  AND2_X1 _7321_ (
    .A1(reg_pmp_3_addr[16]),
    .A2(_0844_),
    .ZN(_0846_)
  );
  OR2_X1 _7322_ (
    .A1(_0843_),
    .A2(_0846_),
    .ZN(_0847_)
  );
  OR2_X1 _7323_ (
    .A1(_0840_),
    .A2(_0847_),
    .ZN(_0848_)
  );
  AND2_X1 _7324_ (
    .A1(_0778_),
    .A2(_0813_),
    .ZN(_0849_)
  );
  AND2_X1 _7325_ (
    .A1(reg_pmp_7_addr[16]),
    .A2(_0849_),
    .ZN(_0850_)
  );
  AND2_X1 _7326_ (
    .A1(_0718_),
    .A2(_0826_),
    .ZN(_0851_)
  );
  AND2_X1 _7327_ (
    .A1(large_1[42]),
    .A2(_0851_),
    .ZN(_0852_)
  );
  OR2_X1 _7328_ (
    .A1(_0850_),
    .A2(_0852_),
    .ZN(_0853_)
  );
  OR2_X1 _7329_ (
    .A1(_0848_),
    .A2(_0853_),
    .ZN(_0854_)
  );
  OR2_X1 _7330_ (
    .A1(_0833_),
    .A2(_0854_),
    .ZN(_0855_)
  );
  AND2_X1 _7331_ (
    .A1(_0773_),
    .A2(_0825_),
    .ZN(_0856_)
  );
  AND2_X1 _7332_ (
    .A1(_0791_),
    .A2(_0856_),
    .ZN(_0857_)
  );
  INV_X1 _7333_ (
    .A(_0857_),
    .ZN(_0858_)
  );
  AND2_X1 _7334_ (
    .A1(_0718_),
    .A2(_0856_),
    .ZN(_0859_)
  );
  OR2_X1 _7335_ (
    .A1(_0812_),
    .A2(_0855_),
    .ZN(io_rw_rdata[16])
  );
  AND2_X1 _7336_ (
    .A1(io_rw_cmd[1]),
    .A2(_0693_),
    .ZN(_0860_)
  );
  AND2_X1 _7337_ (
    .A1(io_rw_rdata[16]),
    .A2(_0860_),
    .ZN(_0861_)
  );
  OR2_X1 _7338_ (
    .A1(_0743_),
    .A2(_0861_),
    .ZN(_0862_)
  );
  MUX2_X1 _7339_ (
    .A(reg_pmp_6_cfg_r),
    .B(_0862_),
    .S(_0740_),
    .Z(_0019_)
  );
  AND2_X1 _7340_ (
    .A1(io_rw_wdata[18]),
    .A2(_0742_),
    .ZN(_0863_)
  );
  AND2_X1 _7341_ (
    .A1(reg_pmp_2_cfg_x),
    .A2(_0754_),
    .ZN(_0864_)
  );
  AND2_X1 _7342_ (
    .A1(reg_pmp_3_addr[18]),
    .A2(_0844_),
    .ZN(_0865_)
  );
  OR2_X1 _7343_ (
    .A1(_0864_),
    .A2(_0865_),
    .ZN(_0866_)
  );
  AND2_X1 _7344_ (
    .A1(reg_mepc[18]),
    .A2(_0783_),
    .ZN(_0867_)
  );
  AND2_X1 _7345_ (
    .A1(reg_mtval[18]),
    .A2(_0764_),
    .ZN(_0868_)
  );
  OR2_X1 _7346_ (
    .A1(_0867_),
    .A2(_0868_),
    .ZN(_0869_)
  );
  OR2_X1 _7347_ (
    .A1(_0866_),
    .A2(_0869_),
    .ZN(_0870_)
  );
  AND2_X1 _7348_ (
    .A1(reg_mcause[18]),
    .A2(_0834_),
    .ZN(_0871_)
  );
  AND2_X1 _7349_ (
    .A1(reg_pmp_0_addr[18]),
    .A2(_0837_),
    .ZN(_0872_)
  );
  OR2_X1 _7350_ (
    .A1(_0871_),
    .A2(_0872_),
    .ZN(_0873_)
  );
  AND2_X1 _7351_ (
    .A1(reg_dpc[18]),
    .A2(_0750_),
    .ZN(_0874_)
  );
  AND2_X1 _7352_ (
    .A1(reg_pmp_2_addr[18]),
    .A2(_0792_),
    .ZN(_0875_)
  );
  OR2_X1 _7353_ (
    .A1(_0874_),
    .A2(_0875_),
    .ZN(_0876_)
  );
  OR2_X1 _7354_ (
    .A1(_0873_),
    .A2(_0876_),
    .ZN(_0877_)
  );
  AND2_X1 _7355_ (
    .A1(reg_pmp_4_addr[18]),
    .A2(_0805_),
    .ZN(_0878_)
  );
  AND2_X1 _7356_ (
    .A1(reg_mtvec[18]),
    .A2(_0780_),
    .ZN(_0879_)
  );
  OR2_X1 _7357_ (
    .A1(_0878_),
    .A2(_0879_),
    .ZN(_0880_)
  );
  AND2_X1 _7358_ (
    .A1(reg_mscratch[18]),
    .A2(_0767_),
    .ZN(_0881_)
  );
  AND2_X1 _7359_ (
    .A1(reg_pmp_6_cfg_x),
    .A2(_0733_),
    .ZN(_0882_)
  );
  OR2_X1 _7360_ (
    .A1(_0881_),
    .A2(_0882_),
    .ZN(_0883_)
  );
  OR2_X1 _7361_ (
    .A1(_0880_),
    .A2(_0883_),
    .ZN(_0884_)
  );
  OR2_X1 _7362_ (
    .A1(_0877_),
    .A2(_0884_),
    .ZN(_0885_)
  );
  OR2_X1 _7363_ (
    .A1(_0870_),
    .A2(_0885_),
    .ZN(_0886_)
  );
  AND2_X1 _7364_ (
    .A1(large_1[44]),
    .A2(_0851_),
    .ZN(_0887_)
  );
  AND2_X1 _7365_ (
    .A1(large_1[12]),
    .A2(_0830_),
    .ZN(_0888_)
  );
  OR2_X1 _7366_ (
    .A1(_0887_),
    .A2(_0888_),
    .ZN(_0889_)
  );
  AND2_X1 _7367_ (
    .A1(large_[44]),
    .A2(_0827_),
    .ZN(_0890_)
  );
  AND2_X1 _7368_ (
    .A1(large_[12]),
    .A2(_0822_),
    .ZN(_0891_)
  );
  OR2_X1 _7369_ (
    .A1(_0890_),
    .A2(_0891_),
    .ZN(_0892_)
  );
  OR2_X1 _7370_ (
    .A1(_0889_),
    .A2(_0892_),
    .ZN(_0893_)
  );
  AND2_X1 _7371_ (
    .A1(reg_pmp_5_addr[18]),
    .A2(_0788_),
    .ZN(_0894_)
  );
  AND2_X1 _7372_ (
    .A1(reg_bp_0_address[18]),
    .A2(_0800_),
    .ZN(_0895_)
  );
  OR2_X1 _7373_ (
    .A1(_0894_),
    .A2(_0895_),
    .ZN(_0896_)
  );
  AND2_X1 _7374_ (
    .A1(reg_dscratch0[18]),
    .A2(_0797_),
    .ZN(_0897_)
  );
  AND2_X1 _7375_ (
    .A1(reg_pmp_1_addr[18]),
    .A2(_0841_),
    .ZN(_0898_)
  );
  OR2_X1 _7376_ (
    .A1(_0897_),
    .A2(_0898_),
    .ZN(_0899_)
  );
  OR2_X1 _7377_ (
    .A1(_0896_),
    .A2(_0899_),
    .ZN(_0900_)
  );
  AND2_X1 _7378_ (
    .A1(reg_pmp_6_addr[18]),
    .A2(_0814_),
    .ZN(_0901_)
  );
  AND2_X1 _7379_ (
    .A1(reg_pmp_7_addr[18]),
    .A2(_0849_),
    .ZN(_0902_)
  );
  OR2_X1 _7380_ (
    .A1(_0901_),
    .A2(_0902_),
    .ZN(_0903_)
  );
  OR2_X1 _7381_ (
    .A1(_0900_),
    .A2(_0903_),
    .ZN(_0904_)
  );
  OR2_X1 _7382_ (
    .A1(_0893_),
    .A2(_0904_),
    .ZN(_0905_)
  );
  OR2_X1 _7383_ (
    .A1(_0886_),
    .A2(_0905_),
    .ZN(io_rw_rdata[18])
  );
  AND2_X1 _7384_ (
    .A1(io_rw_cmd[1]),
    .A2(_0695_),
    .ZN(_0906_)
  );
  AND2_X1 _7385_ (
    .A1(io_rw_rdata[18]),
    .A2(_0906_),
    .ZN(_0907_)
  );
  OR2_X1 _7386_ (
    .A1(_0863_),
    .A2(_0907_),
    .ZN(_0908_)
  );
  MUX2_X1 _7387_ (
    .A(reg_pmp_6_cfg_x),
    .B(_0908_),
    .S(_0740_),
    .Z(_0020_)
  );
  AND2_X1 _7388_ (
    .A1(io_rw_cmd[2]),
    .A2(_0734_),
    .ZN(_0909_)
  );
  OR2_X1 _7389_ (
    .A1(_0656_),
    .A2(_0735_),
    .ZN(_0910_)
  );
  AND2_X1 _7390_ (
    .A1(_0777_),
    .A2(_0909_),
    .ZN(_0911_)
  );
  AND2_X1 _7391_ (
    .A1(_0775_),
    .A2(_0911_),
    .ZN(_0912_)
  );
  OR2_X1 _7392_ (
    .A1(io_status_cease_r),
    .A2(_0912_),
    .ZN(_0913_)
  );
  AND2_X1 _7393_ (
    .A1(_0654_),
    .A2(_0913_),
    .ZN(_0021_)
  );
  OR2_X1 _7394_ (
    .A1(reg_pmp_6_cfg_a[0]),
    .A2(_0740_),
    .ZN(_0914_)
  );
  AND2_X1 _7395_ (
    .A1(_0654_),
    .A2(_0914_),
    .ZN(_0915_)
  );
  AND2_X1 _7396_ (
    .A1(io_rw_wdata[19]),
    .A2(_0742_),
    .ZN(_0916_)
  );
  AND2_X1 _7397_ (
    .A1(io_rw_cmd[1]),
    .A2(_0696_),
    .ZN(_0917_)
  );
  AND2_X1 _7398_ (
    .A1(reg_bp_0_address[19]),
    .A2(_0800_),
    .ZN(_0918_)
  );
  AND2_X1 _7399_ (
    .A1(reg_pmp_5_addr[19]),
    .A2(_0788_),
    .ZN(_0919_)
  );
  OR2_X1 _7400_ (
    .A1(_0918_),
    .A2(_0919_),
    .ZN(_0920_)
  );
  AND2_X1 _7401_ (
    .A1(reg_pmp_2_cfg_a[0]),
    .A2(_0754_),
    .ZN(_0921_)
  );
  AND2_X1 _7402_ (
    .A1(_0669_),
    .A2(io_rw_addr[4]),
    .ZN(_0922_)
  );
  AND2_X1 _7403_ (
    .A1(io_rw_addr[10]),
    .A2(_0922_),
    .ZN(_0923_)
  );
  AND2_X1 _7404_ (
    .A1(_0771_),
    .A2(_0923_),
    .ZN(_0924_)
  );
  AND2_X1 _7405_ (
    .A1(_0817_),
    .A2(_0924_),
    .ZN(_0925_)
  );
  AND2_X1 _7406_ (
    .A1(_0763_),
    .A2(_0925_),
    .ZN(_0926_)
  );
  OR2_X1 _7407_ (
    .A1(_0921_),
    .A2(_0926_),
    .ZN(_0927_)
  );
  OR2_X1 _7408_ (
    .A1(_0920_),
    .A2(_0927_),
    .ZN(_0928_)
  );
  AND2_X1 _7409_ (
    .A1(reg_mtvec[19]),
    .A2(_0780_),
    .ZN(_0929_)
  );
  AND2_X1 _7410_ (
    .A1(reg_dpc[19]),
    .A2(_0750_),
    .ZN(_0930_)
  );
  OR2_X1 _7411_ (
    .A1(_0929_),
    .A2(_0930_),
    .ZN(_0931_)
  );
  AND2_X1 _7412_ (
    .A1(reg_mepc[19]),
    .A2(_0783_),
    .ZN(_0932_)
  );
  AND2_X1 _7413_ (
    .A1(reg_mcause[19]),
    .A2(_0834_),
    .ZN(_0933_)
  );
  OR2_X1 _7414_ (
    .A1(_0932_),
    .A2(_0933_),
    .ZN(_0934_)
  );
  OR2_X1 _7415_ (
    .A1(_0931_),
    .A2(_0934_),
    .ZN(_0935_)
  );
  OR2_X1 _7416_ (
    .A1(_0928_),
    .A2(_0935_),
    .ZN(_0936_)
  );
  AND2_X1 _7417_ (
    .A1(reg_pmp_2_addr[19]),
    .A2(_0792_),
    .ZN(_0937_)
  );
  AND2_X1 _7418_ (
    .A1(reg_pmp_6_cfg_a[0]),
    .A2(_0733_),
    .ZN(_0938_)
  );
  AND2_X1 _7419_ (
    .A1(reg_pmp_4_addr[19]),
    .A2(_0805_),
    .ZN(_0939_)
  );
  OR2_X1 _7420_ (
    .A1(_0938_),
    .A2(_0939_),
    .ZN(_0940_)
  );
  OR2_X1 _7421_ (
    .A1(_0937_),
    .A2(_0940_),
    .ZN(_0941_)
  );
  AND2_X1 _7422_ (
    .A1(reg_dscratch0[19]),
    .A2(_0797_),
    .ZN(_0942_)
  );
  AND2_X1 _7423_ (
    .A1(reg_pmp_1_addr[19]),
    .A2(_0841_),
    .ZN(_0943_)
  );
  OR2_X1 _7424_ (
    .A1(_0942_),
    .A2(_0943_),
    .ZN(_0944_)
  );
  AND2_X1 _7425_ (
    .A1(reg_mtval[19]),
    .A2(_0764_),
    .ZN(_0945_)
  );
  AND2_X1 _7426_ (
    .A1(reg_pmp_3_addr[19]),
    .A2(_0844_),
    .ZN(_0946_)
  );
  OR2_X1 _7427_ (
    .A1(_0945_),
    .A2(_0946_),
    .ZN(_0947_)
  );
  OR2_X1 _7428_ (
    .A1(_0944_),
    .A2(_0947_),
    .ZN(_0948_)
  );
  OR2_X1 _7429_ (
    .A1(_0941_),
    .A2(_0948_),
    .ZN(_0949_)
  );
  OR2_X1 _7430_ (
    .A1(_0936_),
    .A2(_0949_),
    .ZN(_0950_)
  );
  AND2_X1 _7431_ (
    .A1(large_1[45]),
    .A2(_0851_),
    .ZN(_0951_)
  );
  AND2_X1 _7432_ (
    .A1(reg_pmp_7_addr[19]),
    .A2(_0849_),
    .ZN(_0952_)
  );
  AND2_X1 _7433_ (
    .A1(large_[13]),
    .A2(_0822_),
    .ZN(_0953_)
  );
  OR2_X1 _7434_ (
    .A1(_0952_),
    .A2(_0953_),
    .ZN(_0954_)
  );
  OR2_X1 _7435_ (
    .A1(_0951_),
    .A2(_0954_),
    .ZN(_0955_)
  );
  AND2_X1 _7436_ (
    .A1(large_[45]),
    .A2(_0827_),
    .ZN(_0956_)
  );
  AND2_X1 _7437_ (
    .A1(reg_pmp_0_addr[19]),
    .A2(_0837_),
    .ZN(_0957_)
  );
  AND2_X1 _7438_ (
    .A1(reg_mscratch[19]),
    .A2(_0767_),
    .ZN(_0958_)
  );
  OR2_X1 _7439_ (
    .A1(_0957_),
    .A2(_0958_),
    .ZN(_0959_)
  );
  OR2_X1 _7440_ (
    .A1(_0956_),
    .A2(_0959_),
    .ZN(_0960_)
  );
  AND2_X1 _7441_ (
    .A1(reg_pmp_6_addr[19]),
    .A2(_0814_),
    .ZN(_0961_)
  );
  AND2_X1 _7442_ (
    .A1(large_1[13]),
    .A2(_0830_),
    .ZN(_0962_)
  );
  OR2_X1 _7443_ (
    .A1(_0961_),
    .A2(_0962_),
    .ZN(_0963_)
  );
  OR2_X1 _7444_ (
    .A1(_0960_),
    .A2(_0963_),
    .ZN(_0964_)
  );
  OR2_X1 _7445_ (
    .A1(_0955_),
    .A2(_0964_),
    .ZN(_0965_)
  );
  OR2_X1 _7446_ (
    .A1(_0950_),
    .A2(_0965_),
    .ZN(io_rw_rdata[19])
  );
  AND2_X1 _7447_ (
    .A1(_0917_),
    .A2(io_rw_rdata[19]),
    .ZN(_0966_)
  );
  OR2_X1 _7448_ (
    .A1(_0916_),
    .A2(_0966_),
    .ZN(_0967_)
  );
  OR2_X1 _7449_ (
    .A1(_0741_),
    .A2(_0967_),
    .ZN(_0968_)
  );
  AND2_X1 _7450_ (
    .A1(_0915_),
    .A2(_0968_),
    .ZN(_0022_)
  );
  OR2_X1 _7451_ (
    .A1(reg_pmp_6_cfg_a[1]),
    .A2(_0740_),
    .ZN(_0969_)
  );
  AND2_X1 _7452_ (
    .A1(_0654_),
    .A2(_0969_),
    .ZN(_0970_)
  );
  AND2_X1 _7453_ (
    .A1(io_rw_wdata[20]),
    .A2(_0742_),
    .ZN(_0971_)
  );
  AND2_X1 _7454_ (
    .A1(reg_pmp_4_addr[20]),
    .A2(_0805_),
    .ZN(_0972_)
  );
  AND2_X1 _7455_ (
    .A1(reg_bp_0_address[20]),
    .A2(_0800_),
    .ZN(_0973_)
  );
  OR2_X1 _7456_ (
    .A1(_0972_),
    .A2(_0973_),
    .ZN(_0974_)
  );
  AND2_X1 _7457_ (
    .A1(reg_pmp_2_addr[20]),
    .A2(_0792_),
    .ZN(_0975_)
  );
  AND2_X1 _7458_ (
    .A1(reg_dpc[20]),
    .A2(_0750_),
    .ZN(_0976_)
  );
  OR2_X1 _7459_ (
    .A1(_0975_),
    .A2(_0976_),
    .ZN(_0977_)
  );
  OR2_X1 _7460_ (
    .A1(_0974_),
    .A2(_0977_),
    .ZN(_0978_)
  );
  AND2_X1 _7461_ (
    .A1(reg_pmp_2_cfg_a[1]),
    .A2(_0754_),
    .ZN(_0979_)
  );
  AND2_X1 _7462_ (
    .A1(reg_pmp_5_addr[20]),
    .A2(_0788_),
    .ZN(_0980_)
  );
  OR2_X1 _7463_ (
    .A1(_0979_),
    .A2(_0980_),
    .ZN(_0981_)
  );
  AND2_X1 _7464_ (
    .A1(reg_mepc[20]),
    .A2(_0783_),
    .ZN(_0982_)
  );
  AND2_X1 _7465_ (
    .A1(reg_mscratch[20]),
    .A2(_0767_),
    .ZN(_0983_)
  );
  OR2_X1 _7466_ (
    .A1(_0982_),
    .A2(_0983_),
    .ZN(_0984_)
  );
  OR2_X1 _7467_ (
    .A1(_0981_),
    .A2(_0984_),
    .ZN(_0985_)
  );
  OR2_X1 _7468_ (
    .A1(_0978_),
    .A2(_0985_),
    .ZN(_0986_)
  );
  AND2_X1 _7469_ (
    .A1(reg_pmp_0_addr[20]),
    .A2(_0837_),
    .ZN(_0987_)
  );
  AND2_X1 _7470_ (
    .A1(reg_pmp_3_addr[20]),
    .A2(_0844_),
    .ZN(_0988_)
  );
  AND2_X1 _7471_ (
    .A1(reg_pmp_1_addr[20]),
    .A2(_0841_),
    .ZN(_0989_)
  );
  OR2_X1 _7472_ (
    .A1(_0988_),
    .A2(_0989_),
    .ZN(_0990_)
  );
  OR2_X1 _7473_ (
    .A1(_0987_),
    .A2(_0990_),
    .ZN(_0991_)
  );
  AND2_X1 _7474_ (
    .A1(reg_mtvec[20]),
    .A2(_0780_),
    .ZN(_0992_)
  );
  AND2_X1 _7475_ (
    .A1(reg_mcause[20]),
    .A2(_0834_),
    .ZN(_0993_)
  );
  OR2_X1 _7476_ (
    .A1(_0992_),
    .A2(_0993_),
    .ZN(_0994_)
  );
  AND2_X1 _7477_ (
    .A1(reg_mtval[20]),
    .A2(_0764_),
    .ZN(_0995_)
  );
  AND2_X1 _7478_ (
    .A1(reg_dscratch0[20]),
    .A2(_0797_),
    .ZN(_0996_)
  );
  OR2_X1 _7479_ (
    .A1(_0995_),
    .A2(_0996_),
    .ZN(_0997_)
  );
  OR2_X1 _7480_ (
    .A1(_0994_),
    .A2(_0997_),
    .ZN(_0998_)
  );
  OR2_X1 _7481_ (
    .A1(_0991_),
    .A2(_0998_),
    .ZN(_0999_)
  );
  OR2_X1 _7482_ (
    .A1(_0986_),
    .A2(_0999_),
    .ZN(_1000_)
  );
  AND2_X1 _7483_ (
    .A1(large_1[14]),
    .A2(_0830_),
    .ZN(_1001_)
  );
  AND2_X1 _7484_ (
    .A1(reg_pmp_6_addr[20]),
    .A2(_0814_),
    .ZN(_1002_)
  );
  AND2_X1 _7485_ (
    .A1(large_1[46]),
    .A2(_0851_),
    .ZN(_1003_)
  );
  OR2_X1 _7486_ (
    .A1(_1002_),
    .A2(_1003_),
    .ZN(_1004_)
  );
  OR2_X1 _7487_ (
    .A1(_1001_),
    .A2(_1004_),
    .ZN(_1005_)
  );
  AND2_X1 _7488_ (
    .A1(large_[46]),
    .A2(_0827_),
    .ZN(_1006_)
  );
  AND2_X1 _7489_ (
    .A1(reg_pmp_6_cfg_a[1]),
    .A2(_0733_),
    .ZN(_1007_)
  );
  OR2_X1 _7490_ (
    .A1(_0926_),
    .A2(_1007_),
    .ZN(_1008_)
  );
  OR2_X1 _7491_ (
    .A1(_1006_),
    .A2(_1008_),
    .ZN(_1009_)
  );
  AND2_X1 _7492_ (
    .A1(reg_pmp_7_addr[20]),
    .A2(_0849_),
    .ZN(_1010_)
  );
  AND2_X1 _7493_ (
    .A1(large_[14]),
    .A2(_0822_),
    .ZN(_1011_)
  );
  OR2_X1 _7494_ (
    .A1(_1010_),
    .A2(_1011_),
    .ZN(_1012_)
  );
  OR2_X1 _7495_ (
    .A1(_1009_),
    .A2(_1012_),
    .ZN(_1013_)
  );
  OR2_X1 _7496_ (
    .A1(_1005_),
    .A2(_1013_),
    .ZN(_1014_)
  );
  OR2_X1 _7497_ (
    .A1(_1000_),
    .A2(_1014_),
    .ZN(io_rw_rdata[20])
  );
  AND2_X1 _7498_ (
    .A1(io_rw_cmd[1]),
    .A2(_0697_),
    .ZN(_1015_)
  );
  AND2_X1 _7499_ (
    .A1(io_rw_rdata[20]),
    .A2(_1015_),
    .ZN(_1016_)
  );
  OR2_X1 _7500_ (
    .A1(_0971_),
    .A2(_1016_),
    .ZN(_1017_)
  );
  OR2_X1 _7501_ (
    .A1(_0741_),
    .A2(_1017_),
    .ZN(_1018_)
  );
  AND2_X1 _7502_ (
    .A1(_0970_),
    .A2(_1018_),
    .ZN(_0023_)
  );
  OR2_X1 _7503_ (
    .A1(reg_pmp_6_cfg_l),
    .A2(_0740_),
    .ZN(_1019_)
  );
  AND2_X1 _7504_ (
    .A1(_0654_),
    .A2(_1019_),
    .ZN(_1020_)
  );
  AND2_X1 _7505_ (
    .A1(io_rw_wdata[23]),
    .A2(_0742_),
    .ZN(_1021_)
  );
  AND2_X1 _7506_ (
    .A1(reg_pmp_5_addr[23]),
    .A2(_0788_),
    .ZN(_1022_)
  );
  AND2_X1 _7507_ (
    .A1(reg_bp_0_address[23]),
    .A2(_0800_),
    .ZN(_1023_)
  );
  OR2_X1 _7508_ (
    .A1(_1022_),
    .A2(_1023_),
    .ZN(_1024_)
  );
  AND2_X1 _7509_ (
    .A1(reg_pmp_2_addr[23]),
    .A2(_0792_),
    .ZN(_1025_)
  );
  AND2_X1 _7510_ (
    .A1(reg_pmp_0_addr[23]),
    .A2(_0837_),
    .ZN(_1026_)
  );
  OR2_X1 _7511_ (
    .A1(_1025_),
    .A2(_1026_),
    .ZN(_1027_)
  );
  OR2_X1 _7512_ (
    .A1(_1024_),
    .A2(_1027_),
    .ZN(_1028_)
  );
  AND2_X1 _7513_ (
    .A1(reg_pmp_4_addr[23]),
    .A2(_0805_),
    .ZN(_1029_)
  );
  AND2_X1 _7514_ (
    .A1(reg_mtvec[23]),
    .A2(_0780_),
    .ZN(_1030_)
  );
  OR2_X1 _7515_ (
    .A1(_1029_),
    .A2(_1030_),
    .ZN(_1031_)
  );
  AND2_X1 _7516_ (
    .A1(reg_dpc[23]),
    .A2(_0750_),
    .ZN(_1032_)
  );
  AND2_X1 _7517_ (
    .A1(reg_pmp_1_addr[23]),
    .A2(_0841_),
    .ZN(_1033_)
  );
  OR2_X1 _7518_ (
    .A1(_1032_),
    .A2(_1033_),
    .ZN(_1034_)
  );
  OR2_X1 _7519_ (
    .A1(_1031_),
    .A2(_1034_),
    .ZN(_1035_)
  );
  OR2_X1 _7520_ (
    .A1(_1028_),
    .A2(_1035_),
    .ZN(_1036_)
  );
  AND2_X1 _7521_ (
    .A1(reg_mcause[23]),
    .A2(_0834_),
    .ZN(_1037_)
  );
  AND2_X1 _7522_ (
    .A1(reg_mtval[23]),
    .A2(_0764_),
    .ZN(_1038_)
  );
  AND2_X1 _7523_ (
    .A1(reg_mscratch[23]),
    .A2(_0767_),
    .ZN(_1039_)
  );
  OR2_X1 _7524_ (
    .A1(_1038_),
    .A2(_1039_),
    .ZN(_1040_)
  );
  OR2_X1 _7525_ (
    .A1(_1037_),
    .A2(_1040_),
    .ZN(_1041_)
  );
  AND2_X1 _7526_ (
    .A1(reg_pmp_2_cfg_l),
    .A2(_0754_),
    .ZN(_1042_)
  );
  AND2_X1 _7527_ (
    .A1(reg_pmp_6_cfg_l),
    .A2(_0733_),
    .ZN(_1043_)
  );
  OR2_X1 _7528_ (
    .A1(_1042_),
    .A2(_1043_),
    .ZN(_1044_)
  );
  AND2_X1 _7529_ (
    .A1(reg_dscratch0[23]),
    .A2(_0797_),
    .ZN(_1045_)
  );
  AND2_X1 _7530_ (
    .A1(reg_pmp_3_addr[23]),
    .A2(_0844_),
    .ZN(_1046_)
  );
  OR2_X1 _7531_ (
    .A1(_1045_),
    .A2(_1046_),
    .ZN(_1047_)
  );
  OR2_X1 _7532_ (
    .A1(_1044_),
    .A2(_1047_),
    .ZN(_1048_)
  );
  OR2_X1 _7533_ (
    .A1(_1041_),
    .A2(_1048_),
    .ZN(_1049_)
  );
  OR2_X1 _7534_ (
    .A1(_1036_),
    .A2(_1049_),
    .ZN(_1050_)
  );
  AND2_X1 _7535_ (
    .A1(large_1[17]),
    .A2(_0830_),
    .ZN(_1051_)
  );
  AND2_X1 _7536_ (
    .A1(large_1[49]),
    .A2(_0851_),
    .ZN(_1052_)
  );
  AND2_X1 _7537_ (
    .A1(reg_pmp_6_addr[23]),
    .A2(_0814_),
    .ZN(_1053_)
  );
  OR2_X1 _7538_ (
    .A1(_1052_),
    .A2(_1053_),
    .ZN(_1054_)
  );
  OR2_X1 _7539_ (
    .A1(_1051_),
    .A2(_1054_),
    .ZN(_1055_)
  );
  AND2_X1 _7540_ (
    .A1(reg_pmp_7_addr[23]),
    .A2(_0849_),
    .ZN(_1056_)
  );
  AND2_X1 _7541_ (
    .A1(_0720_),
    .A2(_0775_),
    .ZN(_1057_)
  );
  AND2_X1 _7542_ (
    .A1(_0720_),
    .A2(_0799_),
    .ZN(_1058_)
  );
  INV_X1 _7543_ (
    .A(_1058_),
    .ZN(_1059_)
  );
  OR2_X1 _7544_ (
    .A1(_1057_),
    .A2(_1058_),
    .ZN(_1060_)
  );
  AND2_X1 _7545_ (
    .A1(reg_mepc[23]),
    .A2(_0783_),
    .ZN(_1061_)
  );
  OR2_X1 _7546_ (
    .A1(_1060_),
    .A2(_1061_),
    .ZN(_1062_)
  );
  OR2_X1 _7547_ (
    .A1(_1056_),
    .A2(_1062_),
    .ZN(_1063_)
  );
  AND2_X1 _7548_ (
    .A1(large_[49]),
    .A2(_0827_),
    .ZN(_1064_)
  );
  AND2_X1 _7549_ (
    .A1(large_[17]),
    .A2(_0822_),
    .ZN(_1065_)
  );
  OR2_X1 _7550_ (
    .A1(_1064_),
    .A2(_1065_),
    .ZN(_1066_)
  );
  OR2_X1 _7551_ (
    .A1(_1063_),
    .A2(_1066_),
    .ZN(_1067_)
  );
  OR2_X1 _7552_ (
    .A1(_1055_),
    .A2(_1067_),
    .ZN(_1068_)
  );
  OR2_X1 _7553_ (
    .A1(_1050_),
    .A2(_1068_),
    .ZN(io_rw_rdata[23])
  );
  AND2_X1 _7554_ (
    .A1(io_rw_cmd[1]),
    .A2(_0700_),
    .ZN(_1069_)
  );
  AND2_X1 _7555_ (
    .A1(io_rw_rdata[23]),
    .A2(_1069_),
    .ZN(_1070_)
  );
  OR2_X1 _7556_ (
    .A1(_1021_),
    .A2(_1070_),
    .ZN(_1071_)
  );
  OR2_X1 _7557_ (
    .A1(_0741_),
    .A2(_1071_),
    .ZN(_1072_)
  );
  AND2_X1 _7558_ (
    .A1(_1020_),
    .A2(_1072_),
    .ZN(_0024_)
  );
  AND2_X1 _7559_ (
    .A1(_0015_),
    .A2(_0733_),
    .ZN(_1073_)
  );
  INV_X1 _7560_ (
    .A(_1073_),
    .ZN(_1074_)
  );
  AND2_X1 _7561_ (
    .A1(_0736_),
    .A2(_1073_),
    .ZN(_1075_)
  );
  OR2_X1 _7562_ (
    .A1(_0737_),
    .A2(_1074_),
    .ZN(_1076_)
  );
  AND2_X1 _7563_ (
    .A1(io_rw_wdata[8]),
    .A2(_0742_),
    .ZN(_1077_)
  );
  AND2_X1 _7564_ (
    .A1(reg_pmp_0_addr[8]),
    .A2(_0837_),
    .ZN(_1078_)
  );
  AND2_X1 _7565_ (
    .A1(reg_mtvec[8]),
    .A2(_0780_),
    .ZN(_1079_)
  );
  OR2_X1 _7566_ (
    .A1(_1078_),
    .A2(_1079_),
    .ZN(_1080_)
  );
  AND2_X1 _7567_ (
    .A1(reg_mtval[8]),
    .A2(_0764_),
    .ZN(_1081_)
  );
  AND2_X1 _7568_ (
    .A1(reg_dpc[8]),
    .A2(_0750_),
    .ZN(_1082_)
  );
  OR2_X1 _7569_ (
    .A1(_1081_),
    .A2(_1082_),
    .ZN(_1083_)
  );
  OR2_X1 _7570_ (
    .A1(_1080_),
    .A2(_1083_),
    .ZN(_1084_)
  );
  AND2_X1 _7571_ (
    .A1(reg_bp_0_control_tmatch[1]),
    .A2(_1058_),
    .ZN(_1085_)
  );
  AND2_X1 _7572_ (
    .A1(_0749_),
    .A2(_0753_),
    .ZN(_1086_)
  );
  INV_X1 _7573_ (
    .A(_1086_),
    .ZN(_1087_)
  );
  AND2_X1 _7574_ (
    .A1(reg_dcsr_cause[2]),
    .A2(_1086_),
    .ZN(_1088_)
  );
  OR2_X1 _7575_ (
    .A1(_1085_),
    .A2(_1088_),
    .ZN(_1089_)
  );
  AND2_X1 _7576_ (
    .A1(reg_bp_0_address[8]),
    .A2(_0800_),
    .ZN(_1090_)
  );
  AND2_X1 _7577_ (
    .A1(reg_dscratch0[8]),
    .A2(_0797_),
    .ZN(_1091_)
  );
  OR2_X1 _7578_ (
    .A1(_1090_),
    .A2(_1091_),
    .ZN(_1092_)
  );
  OR2_X1 _7579_ (
    .A1(_1089_),
    .A2(_1092_),
    .ZN(_1093_)
  );
  OR2_X1 _7580_ (
    .A1(_1084_),
    .A2(_1093_),
    .ZN(_1094_)
  );
  AND2_X1 _7581_ (
    .A1(reg_pmp_4_addr[8]),
    .A2(_0805_),
    .ZN(_1095_)
  );
  AND2_X1 _7582_ (
    .A1(reg_mscratch[8]),
    .A2(_0767_),
    .ZN(_1096_)
  );
  AND2_X1 _7583_ (
    .A1(reg_mepc[8]),
    .A2(_0783_),
    .ZN(_1097_)
  );
  OR2_X1 _7584_ (
    .A1(_1096_),
    .A2(_1097_),
    .ZN(_1098_)
  );
  OR2_X1 _7585_ (
    .A1(_1095_),
    .A2(_1098_),
    .ZN(_1099_)
  );
  AND2_X1 _7586_ (
    .A1(reg_pmp_2_addr[8]),
    .A2(_0792_),
    .ZN(_1100_)
  );
  AND2_X1 _7587_ (
    .A1(reg_pmp_5_cfg_r),
    .A2(_0733_),
    .ZN(_1101_)
  );
  OR2_X1 _7588_ (
    .A1(_1100_),
    .A2(_1101_),
    .ZN(_1102_)
  );
  AND2_X1 _7589_ (
    .A1(reg_pmp_1_cfg_r),
    .A2(_0754_),
    .ZN(_1103_)
  );
  AND2_X1 _7590_ (
    .A1(reg_mcause[8]),
    .A2(_0834_),
    .ZN(_1104_)
  );
  OR2_X1 _7591_ (
    .A1(_1103_),
    .A2(_1104_),
    .ZN(_1105_)
  );
  OR2_X1 _7592_ (
    .A1(_1102_),
    .A2(_1105_),
    .ZN(_1106_)
  );
  OR2_X1 _7593_ (
    .A1(_1099_),
    .A2(_1106_),
    .ZN(_1107_)
  );
  OR2_X1 _7594_ (
    .A1(_1094_),
    .A2(_1107_),
    .ZN(_1108_)
  );
  AND2_X1 _7595_ (
    .A1(reg_pmp_7_addr[8]),
    .A2(_0849_),
    .ZN(_1109_)
  );
  AND2_X1 _7596_ (
    .A1(reg_pmp_6_addr[8]),
    .A2(_0814_),
    .ZN(_1110_)
  );
  OR2_X1 _7597_ (
    .A1(_1109_),
    .A2(_1110_),
    .ZN(_1111_)
  );
  AND2_X1 _7598_ (
    .A1(large_[34]),
    .A2(_0827_),
    .ZN(_1112_)
  );
  AND2_X1 _7599_ (
    .A1(large_[2]),
    .A2(_0822_),
    .ZN(_1113_)
  );
  OR2_X1 _7600_ (
    .A1(_1112_),
    .A2(_1113_),
    .ZN(_1114_)
  );
  OR2_X1 _7601_ (
    .A1(_1111_),
    .A2(_1114_),
    .ZN(_1115_)
  );
  AND2_X1 _7602_ (
    .A1(reg_pmp_3_addr[8]),
    .A2(_0844_),
    .ZN(_1116_)
  );
  OR2_X1 _7603_ (
    .A1(_1057_),
    .A2(_1116_),
    .ZN(_1117_)
  );
  AND2_X1 _7604_ (
    .A1(reg_pmp_5_addr[8]),
    .A2(_0788_),
    .ZN(_1118_)
  );
  AND2_X1 _7605_ (
    .A1(reg_pmp_1_addr[8]),
    .A2(_0841_),
    .ZN(_1119_)
  );
  OR2_X1 _7606_ (
    .A1(_1118_),
    .A2(_1119_),
    .ZN(_1120_)
  );
  OR2_X1 _7607_ (
    .A1(_1117_),
    .A2(_1120_),
    .ZN(_1121_)
  );
  AND2_X1 _7608_ (
    .A1(large_1[34]),
    .A2(_0851_),
    .ZN(_1122_)
  );
  AND2_X1 _7609_ (
    .A1(large_1[2]),
    .A2(_0830_),
    .ZN(_1123_)
  );
  OR2_X1 _7610_ (
    .A1(_1122_),
    .A2(_1123_),
    .ZN(_1124_)
  );
  OR2_X1 _7611_ (
    .A1(_1121_),
    .A2(_1124_),
    .ZN(_1125_)
  );
  OR2_X1 _7612_ (
    .A1(_1115_),
    .A2(_1125_),
    .ZN(_1126_)
  );
  OR2_X1 _7613_ (
    .A1(_1108_),
    .A2(_1126_),
    .ZN(io_rw_rdata[8])
  );
  AND2_X1 _7614_ (
    .A1(io_rw_cmd[1]),
    .A2(_0686_),
    .ZN(_1127_)
  );
  AND2_X1 _7615_ (
    .A1(io_rw_rdata[8]),
    .A2(_1127_),
    .ZN(_1128_)
  );
  OR2_X1 _7616_ (
    .A1(_1077_),
    .A2(_1128_),
    .ZN(_1129_)
  );
  MUX2_X1 _7617_ (
    .A(reg_pmp_5_cfg_r),
    .B(_1129_),
    .S(_1075_),
    .Z(_0025_)
  );
  AND2_X1 _7618_ (
    .A1(io_rw_wdata[9]),
    .A2(_0742_),
    .ZN(_1130_)
  );
  AND2_X1 _7619_ (
    .A1(reg_mscratch[9]),
    .A2(_0767_),
    .ZN(_1131_)
  );
  AND2_X1 _7620_ (
    .A1(reg_mtvec[9]),
    .A2(_0780_),
    .ZN(_1132_)
  );
  OR2_X1 _7621_ (
    .A1(_1131_),
    .A2(_1132_),
    .ZN(_1133_)
  );
  AND2_X1 _7622_ (
    .A1(reg_pmp_1_addr[9]),
    .A2(_0841_),
    .ZN(_1134_)
  );
  AND2_X1 _7623_ (
    .A1(reg_pmp_2_addr[9]),
    .A2(_0792_),
    .ZN(_1135_)
  );
  OR2_X1 _7624_ (
    .A1(_1134_),
    .A2(_1135_),
    .ZN(_1136_)
  );
  OR2_X1 _7625_ (
    .A1(_1133_),
    .A2(_1136_),
    .ZN(_1137_)
  );
  AND2_X1 _7626_ (
    .A1(reg_mtval[9]),
    .A2(_0764_),
    .ZN(_1138_)
  );
  AND2_X1 _7627_ (
    .A1(reg_mcause[9]),
    .A2(_0834_),
    .ZN(_1139_)
  );
  OR2_X1 _7628_ (
    .A1(_1138_),
    .A2(_1139_),
    .ZN(_1140_)
  );
  AND2_X1 _7629_ (
    .A1(reg_pmp_0_addr[9]),
    .A2(_0837_),
    .ZN(_1141_)
  );
  AND2_X1 _7630_ (
    .A1(reg_pmp_5_addr[9]),
    .A2(_0788_),
    .ZN(_1142_)
  );
  OR2_X1 _7631_ (
    .A1(_1141_),
    .A2(_1142_),
    .ZN(_1143_)
  );
  OR2_X1 _7632_ (
    .A1(_1140_),
    .A2(_1143_),
    .ZN(_1144_)
  );
  AND2_X1 _7633_ (
    .A1(reg_dscratch0[9]),
    .A2(_0797_),
    .ZN(_1145_)
  );
  AND2_X1 _7634_ (
    .A1(reg_bp_0_address[9]),
    .A2(_0800_),
    .ZN(_1146_)
  );
  OR2_X1 _7635_ (
    .A1(_1145_),
    .A2(_1146_),
    .ZN(_1147_)
  );
  AND2_X1 _7636_ (
    .A1(reg_dpc[9]),
    .A2(_0750_),
    .ZN(_1148_)
  );
  AND2_X1 _7637_ (
    .A1(reg_pmp_4_addr[9]),
    .A2(_0805_),
    .ZN(_1149_)
  );
  OR2_X1 _7638_ (
    .A1(_1148_),
    .A2(_1149_),
    .ZN(_1150_)
  );
  OR2_X1 _7639_ (
    .A1(_1147_),
    .A2(_1150_),
    .ZN(_1151_)
  );
  OR2_X1 _7640_ (
    .A1(_1144_),
    .A2(_1151_),
    .ZN(_1152_)
  );
  OR2_X1 _7641_ (
    .A1(_1137_),
    .A2(_1152_),
    .ZN(_1153_)
  );
  AND2_X1 _7642_ (
    .A1(reg_pmp_7_addr[9]),
    .A2(_0849_),
    .ZN(_1154_)
  );
  AND2_X1 _7643_ (
    .A1(large_1[35]),
    .A2(_0851_),
    .ZN(_1155_)
  );
  OR2_X1 _7644_ (
    .A1(_1154_),
    .A2(_1155_),
    .ZN(_1156_)
  );
  AND2_X1 _7645_ (
    .A1(reg_pmp_6_addr[9]),
    .A2(_0814_),
    .ZN(_1157_)
  );
  AND2_X1 _7646_ (
    .A1(large_1[3]),
    .A2(_0830_),
    .ZN(_1158_)
  );
  OR2_X1 _7647_ (
    .A1(_1157_),
    .A2(_1158_),
    .ZN(_1159_)
  );
  OR2_X1 _7648_ (
    .A1(_1156_),
    .A2(_1159_),
    .ZN(_1160_)
  );
  AND2_X1 _7649_ (
    .A1(reg_pmp_5_cfg_w),
    .A2(_0733_),
    .ZN(_1161_)
  );
  AND2_X1 _7650_ (
    .A1(reg_mepc[9]),
    .A2(_0783_),
    .ZN(_1162_)
  );
  OR2_X1 _7651_ (
    .A1(_1161_),
    .A2(_1162_),
    .ZN(_1163_)
  );
  AND2_X1 _7652_ (
    .A1(reg_pmp_1_cfg_w),
    .A2(_0754_),
    .ZN(_1164_)
  );
  AND2_X1 _7653_ (
    .A1(reg_pmp_3_addr[9]),
    .A2(_0844_),
    .ZN(_1165_)
  );
  OR2_X1 _7654_ (
    .A1(_1164_),
    .A2(_1165_),
    .ZN(_1166_)
  );
  OR2_X1 _7655_ (
    .A1(_1163_),
    .A2(_1166_),
    .ZN(_1167_)
  );
  AND2_X1 _7656_ (
    .A1(large_[35]),
    .A2(_0827_),
    .ZN(_1168_)
  );
  AND2_X1 _7657_ (
    .A1(large_[3]),
    .A2(_0822_),
    .ZN(_1169_)
  );
  OR2_X1 _7658_ (
    .A1(_1168_),
    .A2(_1169_),
    .ZN(_1170_)
  );
  OR2_X1 _7659_ (
    .A1(_1167_),
    .A2(_1170_),
    .ZN(_1171_)
  );
  OR2_X1 _7660_ (
    .A1(_1160_),
    .A2(_1171_),
    .ZN(_1172_)
  );
  OR2_X1 _7661_ (
    .A1(_1153_),
    .A2(_1172_),
    .ZN(io_rw_rdata[9])
  );
  AND2_X1 _7662_ (
    .A1(io_rw_cmd[1]),
    .A2(_0687_),
    .ZN(_1173_)
  );
  AND2_X1 _7663_ (
    .A1(io_rw_rdata[9]),
    .A2(_1173_),
    .ZN(_1174_)
  );
  OR2_X1 _7664_ (
    .A1(_1130_),
    .A2(_1174_),
    .ZN(_1175_)
  );
  AND2_X1 _7665_ (
    .A1(_1129_),
    .A2(_1175_),
    .ZN(_1176_)
  );
  MUX2_X1 _7666_ (
    .A(reg_pmp_5_cfg_w),
    .B(_1176_),
    .S(_1075_),
    .Z(_0026_)
  );
  AND2_X1 _7667_ (
    .A1(reg_pmp_6_cfg_l),
    .A2(reg_pmp_6_cfg_a[0]),
    .ZN(_1177_)
  );
  AND2_X1 _7668_ (
    .A1(_0018_),
    .A2(_1177_),
    .ZN(_1178_)
  );
  OR2_X1 _7669_ (
    .A1(reg_pmp_5_cfg_l),
    .A2(_1178_),
    .ZN(_1179_)
  );
  OR2_X1 _7670_ (
    .A1(_0737_),
    .A2(_1179_),
    .ZN(_1180_)
  );
  OR2_X1 _7671_ (
    .A1(_0789_),
    .A2(_1180_),
    .ZN(_1181_)
  );
  AND2_X1 _7672_ (
    .A1(io_rw_wdata[0]),
    .A2(_0742_),
    .ZN(_1182_)
  );
  AND2_X1 _7673_ (
    .A1(reg_misa[0]),
    .A2(_1057_),
    .ZN(_1183_)
  );
  AND2_X1 _7674_ (
    .A1(reg_pmp_5_addr[0]),
    .A2(_0788_),
    .ZN(_1184_)
  );
  OR2_X1 _7675_ (
    .A1(_1183_),
    .A2(_1184_),
    .ZN(_1185_)
  );
  AND2_X1 _7676_ (
    .A1(reg_mscratch[0]),
    .A2(_0767_),
    .ZN(_1186_)
  );
  AND2_X1 _7677_ (
    .A1(io_hartid),
    .A2(_0777_),
    .ZN(_1187_)
  );
  OR2_X1 _7678_ (
    .A1(_0791_),
    .A2(_1187_),
    .ZN(_1188_)
  );
  AND2_X1 _7679_ (
    .A1(_0925_),
    .A2(_1188_),
    .ZN(_1189_)
  );
  OR2_X1 _7680_ (
    .A1(_1186_),
    .A2(_1189_),
    .ZN(_1190_)
  );
  OR2_X1 _7681_ (
    .A1(_1185_),
    .A2(_1190_),
    .ZN(_1191_)
  );
  AND2_X1 _7682_ (
    .A1(reg_pmp_2_addr[0]),
    .A2(_0792_),
    .ZN(_1192_)
  );
  AND2_X1 _7683_ (
    .A1(reg_pmp_3_addr[0]),
    .A2(_0844_),
    .ZN(_1193_)
  );
  OR2_X1 _7684_ (
    .A1(_1192_),
    .A2(_1193_),
    .ZN(_1194_)
  );
  AND2_X1 _7685_ (
    .A1(reg_dscratch0[0]),
    .A2(_0797_),
    .ZN(_1195_)
  );
  AND2_X1 _7686_ (
    .A1(reg_pmp_1_addr[0]),
    .A2(_0841_),
    .ZN(_1196_)
  );
  OR2_X1 _7687_ (
    .A1(_1195_),
    .A2(_1196_),
    .ZN(_1197_)
  );
  OR2_X1 _7688_ (
    .A1(_1194_),
    .A2(_1197_),
    .ZN(_1198_)
  );
  OR2_X1 _7689_ (
    .A1(_1191_),
    .A2(_1198_),
    .ZN(_1199_)
  );
  AND2_X1 _7690_ (
    .A1(reg_mtvec[0]),
    .A2(_0780_),
    .ZN(_1200_)
  );
  AND2_X1 _7691_ (
    .A1(reg_mcause[0]),
    .A2(_0834_),
    .ZN(_1201_)
  );
  AND2_X1 _7692_ (
    .A1(_0728_),
    .A2(_0771_),
    .ZN(_1202_)
  );
  AND2_X1 _7693_ (
    .A1(_0718_),
    .A2(_1202_),
    .ZN(_1203_)
  );
  AND2_X1 _7694_ (
    .A1(_0726_),
    .A2(_1203_),
    .ZN(_1204_)
  );
  AND2_X1 _7695_ (
    .A1(reg_mcountinhibit[0]),
    .A2(_1204_),
    .ZN(_1205_)
  );
  OR2_X1 _7696_ (
    .A1(_1201_),
    .A2(_1205_),
    .ZN(_1206_)
  );
  OR2_X1 _7697_ (
    .A1(_1200_),
    .A2(_1206_),
    .ZN(_1207_)
  );
  AND2_X1 _7698_ (
    .A1(reg_pmp_0_cfg_r),
    .A2(_0754_),
    .ZN(_1208_)
  );
  AND2_X1 _7699_ (
    .A1(reg_pmp_4_cfg_r),
    .A2(_0733_),
    .ZN(_1209_)
  );
  OR2_X1 _7700_ (
    .A1(_1208_),
    .A2(_1209_),
    .ZN(_1210_)
  );
  AND2_X1 _7701_ (
    .A1(reg_mtval[0]),
    .A2(_0764_),
    .ZN(_1211_)
  );
  AND2_X1 _7702_ (
    .A1(reg_pmp_4_addr[0]),
    .A2(_0805_),
    .ZN(_1212_)
  );
  OR2_X1 _7703_ (
    .A1(_1211_),
    .A2(_1212_),
    .ZN(_1213_)
  );
  OR2_X1 _7704_ (
    .A1(_1210_),
    .A2(_1213_),
    .ZN(_1214_)
  );
  OR2_X1 _7705_ (
    .A1(_1207_),
    .A2(_1214_),
    .ZN(_1215_)
  );
  OR2_X1 _7706_ (
    .A1(_1199_),
    .A2(_1215_),
    .ZN(_1216_)
  );
  AND2_X1 _7707_ (
    .A1(reg_pmp_7_addr[0]),
    .A2(_0849_),
    .ZN(_1217_)
  );
  AND2_X1 _7708_ (
    .A1(small_[0]),
    .A2(_0822_),
    .ZN(_1218_)
  );
  OR2_X1 _7709_ (
    .A1(_1217_),
    .A2(_1218_),
    .ZN(_1219_)
  );
  AND2_X1 _7710_ (
    .A1(reg_pmp_6_addr[0]),
    .A2(_0814_),
    .ZN(_1220_)
  );
  AND2_X1 _7711_ (
    .A1(small_1[0]),
    .A2(_0830_),
    .ZN(_1221_)
  );
  OR2_X1 _7712_ (
    .A1(_1220_),
    .A2(_1221_),
    .ZN(_1222_)
  );
  OR2_X1 _7713_ (
    .A1(_1219_),
    .A2(_1222_),
    .ZN(_1223_)
  );
  AND2_X1 _7714_ (
    .A1(reg_bp_0_address[0]),
    .A2(_0800_),
    .ZN(_1224_)
  );
  OR2_X1 _7715_ (
    .A1(_1086_),
    .A2(_1224_),
    .ZN(_1225_)
  );
  AND2_X1 _7716_ (
    .A1(reg_pmp_0_addr[0]),
    .A2(_0837_),
    .ZN(_1226_)
  );
  AND2_X1 _7717_ (
    .A1(reg_bp_0_control_r),
    .A2(_1058_),
    .ZN(_1227_)
  );
  OR2_X1 _7718_ (
    .A1(_1226_),
    .A2(_1227_),
    .ZN(_1228_)
  );
  OR2_X1 _7719_ (
    .A1(_1225_),
    .A2(_1228_),
    .ZN(_1229_)
  );
  AND2_X1 _7720_ (
    .A1(large_[26]),
    .A2(_0827_),
    .ZN(_1230_)
  );
  AND2_X1 _7721_ (
    .A1(large_1[26]),
    .A2(_0851_),
    .ZN(_1231_)
  );
  OR2_X1 _7722_ (
    .A1(_1230_),
    .A2(_1231_),
    .ZN(_1232_)
  );
  OR2_X1 _7723_ (
    .A1(_1229_),
    .A2(_1232_),
    .ZN(_1233_)
  );
  OR2_X1 _7724_ (
    .A1(_1223_),
    .A2(_1233_),
    .ZN(_1234_)
  );
  AND2_X1 _7725_ (
    .A1(_0718_),
    .A2(_0730_),
    .ZN(_1235_)
  );
  OR2_X1 _7726_ (
    .A1(_0719_),
    .A2(_0731_),
    .ZN(_1236_)
  );
  AND2_X1 _7727_ (
    .A1(_0771_),
    .A2(_1235_),
    .ZN(_1237_)
  );
  OR2_X1 _7728_ (
    .A1(_0772_),
    .A2(_1236_),
    .ZN(_1238_)
  );
  OR2_X1 _7729_ (
    .A1(_1216_),
    .A2(_1234_),
    .ZN(io_rw_rdata[0])
  );
  AND2_X1 _7730_ (
    .A1(io_rw_cmd[1]),
    .A2(_0678_),
    .ZN(_1239_)
  );
  AND2_X1 _7731_ (
    .A1(io_rw_rdata[0]),
    .A2(_1239_),
    .ZN(_1240_)
  );
  OR2_X1 _7732_ (
    .A1(_1182_),
    .A2(_1240_),
    .ZN(_1241_)
  );
  MUX2_X1 _7733_ (
    .A(_1241_),
    .B(reg_pmp_5_addr[0]),
    .S(_1181_),
    .Z(_0027_)
  );
  AND2_X1 _7734_ (
    .A1(io_rw_wdata[1]),
    .A2(_0742_),
    .ZN(_1242_)
  );
  AND2_X1 _7735_ (
    .A1(io_rw_cmd[1]),
    .A2(_0679_),
    .ZN(_1243_)
  );
  AND2_X1 _7736_ (
    .A1(reg_pmp_1_addr[1]),
    .A2(_0841_),
    .ZN(_1244_)
  );
  AND2_X1 _7737_ (
    .A1(reg_pmp_4_addr[1]),
    .A2(_0805_),
    .ZN(_1245_)
  );
  OR2_X1 _7738_ (
    .A1(_1244_),
    .A2(_1245_),
    .ZN(_1246_)
  );
  AND2_X1 _7739_ (
    .A1(reg_pmp_0_addr[1]),
    .A2(_0837_),
    .ZN(_1247_)
  );
  AND2_X1 _7740_ (
    .A1(reg_bp_0_address[1]),
    .A2(_0800_),
    .ZN(_1248_)
  );
  OR2_X1 _7741_ (
    .A1(_1247_),
    .A2(_1248_),
    .ZN(_1249_)
  );
  OR2_X1 _7742_ (
    .A1(_1246_),
    .A2(_1249_),
    .ZN(_1250_)
  );
  AND2_X1 _7743_ (
    .A1(reg_dscratch0[1]),
    .A2(_0797_),
    .ZN(_1251_)
  );
  AND2_X1 _7744_ (
    .A1(_0713_),
    .A2(_0714_),
    .ZN(_1252_)
  );
  AND2_X1 _7745_ (
    .A1(_0750_),
    .A2(_1252_),
    .ZN(_1253_)
  );
  OR2_X1 _7746_ (
    .A1(_1251_),
    .A2(_1253_),
    .ZN(_1254_)
  );
  AND2_X1 _7747_ (
    .A1(reg_pmp_2_addr[1]),
    .A2(_0792_),
    .ZN(_1255_)
  );
  AND2_X1 _7748_ (
    .A1(reg_bp_0_control_w),
    .A2(_1058_),
    .ZN(_1256_)
  );
  OR2_X1 _7749_ (
    .A1(_1255_),
    .A2(_1256_),
    .ZN(_1257_)
  );
  OR2_X1 _7750_ (
    .A1(_1254_),
    .A2(_1257_),
    .ZN(_1258_)
  );
  OR2_X1 _7751_ (
    .A1(_1250_),
    .A2(_1258_),
    .ZN(_1259_)
  );
  AND2_X1 _7752_ (
    .A1(_0712_),
    .A2(_0713_),
    .ZN(_1260_)
  );
  AND2_X1 _7753_ (
    .A1(_0783_),
    .A2(_1260_),
    .ZN(_1261_)
  );
  AND2_X1 _7754_ (
    .A1(reg_mcause[1]),
    .A2(_0834_),
    .ZN(_1262_)
  );
  AND2_X1 _7755_ (
    .A1(reg_mscratch[1]),
    .A2(_0767_),
    .ZN(_1263_)
  );
  OR2_X1 _7756_ (
    .A1(_1262_),
    .A2(_1263_),
    .ZN(_1264_)
  );
  OR2_X1 _7757_ (
    .A1(_1261_),
    .A2(_1264_),
    .ZN(_1265_)
  );
  AND2_X1 _7758_ (
    .A1(reg_pmp_5_addr[1]),
    .A2(_0788_),
    .ZN(_1266_)
  );
  AND2_X1 _7759_ (
    .A1(reg_pmp_4_cfg_w),
    .A2(_0733_),
    .ZN(_1267_)
  );
  OR2_X1 _7760_ (
    .A1(_1266_),
    .A2(_1267_),
    .ZN(_1268_)
  );
  AND2_X1 _7761_ (
    .A1(reg_mtval[1]),
    .A2(_0764_),
    .ZN(_1269_)
  );
  AND2_X1 _7762_ (
    .A1(reg_pmp_3_addr[1]),
    .A2(_0844_),
    .ZN(_1270_)
  );
  OR2_X1 _7763_ (
    .A1(_1269_),
    .A2(_1270_),
    .ZN(_1271_)
  );
  OR2_X1 _7764_ (
    .A1(_1268_),
    .A2(_1271_),
    .ZN(_1272_)
  );
  OR2_X1 _7765_ (
    .A1(_1265_),
    .A2(_1272_),
    .ZN(_1273_)
  );
  OR2_X1 _7766_ (
    .A1(_1259_),
    .A2(_1273_),
    .ZN(_1274_)
  );
  AND2_X1 _7767_ (
    .A1(large_1[27]),
    .A2(_0851_),
    .ZN(_1275_)
  );
  AND2_X1 _7768_ (
    .A1(small_1[1]),
    .A2(_0830_),
    .ZN(_1276_)
  );
  AND2_X1 _7769_ (
    .A1(small_[1]),
    .A2(_0822_),
    .ZN(_1277_)
  );
  OR2_X1 _7770_ (
    .A1(_1276_),
    .A2(_1277_),
    .ZN(_1278_)
  );
  OR2_X1 _7771_ (
    .A1(_1275_),
    .A2(_1278_),
    .ZN(_1279_)
  );
  AND2_X1 _7772_ (
    .A1(reg_pmp_6_addr[1]),
    .A2(_0814_),
    .ZN(_1280_)
  );
  AND2_X1 _7773_ (
    .A1(reg_pmp_0_cfg_w),
    .A2(_0754_),
    .ZN(_1281_)
  );
  OR2_X1 _7774_ (
    .A1(_1086_),
    .A2(_1281_),
    .ZN(_1282_)
  );
  OR2_X1 _7775_ (
    .A1(_1280_),
    .A2(_1282_),
    .ZN(_1283_)
  );
  AND2_X1 _7776_ (
    .A1(large_[27]),
    .A2(_0827_),
    .ZN(_1284_)
  );
  AND2_X1 _7777_ (
    .A1(reg_pmp_7_addr[1]),
    .A2(_0849_),
    .ZN(_1285_)
  );
  OR2_X1 _7778_ (
    .A1(_1284_),
    .A2(_1285_),
    .ZN(_1286_)
  );
  OR2_X1 _7779_ (
    .A1(_1283_),
    .A2(_1286_),
    .ZN(_1287_)
  );
  OR2_X1 _7780_ (
    .A1(_1279_),
    .A2(_1287_),
    .ZN(_1288_)
  );
  OR2_X1 _7781_ (
    .A1(_1274_),
    .A2(_1288_),
    .ZN(io_rw_rdata[1])
  );
  AND2_X1 _7782_ (
    .A1(_1243_),
    .A2(io_rw_rdata[1]),
    .ZN(_1289_)
  );
  OR2_X1 _7783_ (
    .A1(_1242_),
    .A2(_1289_),
    .ZN(_1290_)
  );
  MUX2_X1 _7784_ (
    .A(_1290_),
    .B(reg_pmp_5_addr[1]),
    .S(_1181_),
    .Z(_0028_)
  );
  AND2_X1 _7785_ (
    .A1(io_rw_wdata[2]),
    .A2(_0742_),
    .ZN(_1291_)
  );
  AND2_X1 _7786_ (
    .A1(reg_mepc[2]),
    .A2(_0783_),
    .ZN(_1292_)
  );
  AND2_X1 _7787_ (
    .A1(reg_mscratch[2]),
    .A2(_0767_),
    .ZN(_1293_)
  );
  AND2_X1 _7788_ (
    .A1(reg_dscratch0[2]),
    .A2(_0797_),
    .ZN(_1294_)
  );
  OR2_X1 _7789_ (
    .A1(_1293_),
    .A2(_1294_),
    .ZN(_1295_)
  );
  OR2_X1 _7790_ (
    .A1(_1292_),
    .A2(_1295_),
    .ZN(_1296_)
  );
  AND2_X1 _7791_ (
    .A1(reg_pmp_0_addr[2]),
    .A2(_0837_),
    .ZN(_1297_)
  );
  AND2_X1 _7792_ (
    .A1(reg_mcause[2]),
    .A2(_0834_),
    .ZN(_1298_)
  );
  OR2_X1 _7793_ (
    .A1(_1297_),
    .A2(_1298_),
    .ZN(_1299_)
  );
  AND2_X1 _7794_ (
    .A1(reg_misa[2]),
    .A2(_1057_),
    .ZN(_1300_)
  );
  AND2_X1 _7795_ (
    .A1(reg_mcountinhibit[2]),
    .A2(_1204_),
    .ZN(_1301_)
  );
  OR2_X1 _7796_ (
    .A1(_1300_),
    .A2(_1301_),
    .ZN(_1302_)
  );
  OR2_X1 _7797_ (
    .A1(_1299_),
    .A2(_1302_),
    .ZN(_1303_)
  );
  AND2_X1 _7798_ (
    .A1(reg_bp_0_address[2]),
    .A2(_0800_),
    .ZN(_1304_)
  );
  AND2_X1 _7799_ (
    .A1(reg_dcsr_step),
    .A2(_1086_),
    .ZN(_1305_)
  );
  OR2_X1 _7800_ (
    .A1(_1304_),
    .A2(_1305_),
    .ZN(_1306_)
  );
  AND2_X1 _7801_ (
    .A1(reg_bp_0_control_x),
    .A2(_1058_),
    .ZN(_1307_)
  );
  AND2_X1 _7802_ (
    .A1(reg_mtvec[2]),
    .A2(_read_mtvec_T_4[6]),
    .ZN(_1308_)
  );
  AND2_X1 _7803_ (
    .A1(_0780_),
    .A2(_1308_),
    .ZN(_1309_)
  );
  OR2_X1 _7804_ (
    .A1(_1307_),
    .A2(_1309_),
    .ZN(_1310_)
  );
  OR2_X1 _7805_ (
    .A1(_1306_),
    .A2(_1310_),
    .ZN(_1311_)
  );
  OR2_X1 _7806_ (
    .A1(_1303_),
    .A2(_1311_),
    .ZN(_1312_)
  );
  OR2_X1 _7807_ (
    .A1(_1296_),
    .A2(_1312_),
    .ZN(_1313_)
  );
  AND2_X1 _7808_ (
    .A1(reg_pmp_6_addr[2]),
    .A2(_0814_),
    .ZN(_1314_)
  );
  AND2_X1 _7809_ (
    .A1(reg_pmp_7_addr[2]),
    .A2(_0849_),
    .ZN(_1315_)
  );
  AND2_X1 _7810_ (
    .A1(small_1[2]),
    .A2(_0830_),
    .ZN(_1316_)
  );
  OR2_X1 _7811_ (
    .A1(_1315_),
    .A2(_1316_),
    .ZN(_1317_)
  );
  OR2_X1 _7812_ (
    .A1(_1314_),
    .A2(_1317_),
    .ZN(_1318_)
  );
  AND2_X1 _7813_ (
    .A1(small_[2]),
    .A2(_0822_),
    .ZN(_1319_)
  );
  AND2_X1 _7814_ (
    .A1(reg_pmp_5_addr[2]),
    .A2(_0788_),
    .ZN(_1320_)
  );
  OR2_X1 _7815_ (
    .A1(_0926_),
    .A2(_1320_),
    .ZN(_1321_)
  );
  OR2_X1 _7816_ (
    .A1(_1319_),
    .A2(_1321_),
    .ZN(_1322_)
  );
  AND2_X1 _7817_ (
    .A1(large_[28]),
    .A2(_0827_),
    .ZN(_1323_)
  );
  AND2_X1 _7818_ (
    .A1(large_1[28]),
    .A2(_0851_),
    .ZN(_1324_)
  );
  OR2_X1 _7819_ (
    .A1(_1323_),
    .A2(_1324_),
    .ZN(_1325_)
  );
  OR2_X1 _7820_ (
    .A1(_1322_),
    .A2(_1325_),
    .ZN(_1326_)
  );
  AND2_X1 _7821_ (
    .A1(reg_pmp_3_addr[2]),
    .A2(_0844_),
    .ZN(_1327_)
  );
  AND2_X1 _7822_ (
    .A1(reg_pmp_4_addr[2]),
    .A2(_0805_),
    .ZN(_1328_)
  );
  OR2_X1 _7823_ (
    .A1(_1327_),
    .A2(_1328_),
    .ZN(_1329_)
  );
  AND2_X1 _7824_ (
    .A1(reg_pmp_1_addr[2]),
    .A2(_0841_),
    .ZN(_1330_)
  );
  AND2_X1 _7825_ (
    .A1(reg_mtval[2]),
    .A2(_0764_),
    .ZN(_1331_)
  );
  OR2_X1 _7826_ (
    .A1(_1330_),
    .A2(_1331_),
    .ZN(_1332_)
  );
  OR2_X1 _7827_ (
    .A1(_1329_),
    .A2(_1332_),
    .ZN(_1333_)
  );
  AND2_X1 _7828_ (
    .A1(reg_pmp_4_cfg_x),
    .A2(_0733_),
    .ZN(_1334_)
  );
  AND2_X1 _7829_ (
    .A1(reg_pmp_0_cfg_x),
    .A2(_0754_),
    .ZN(_1335_)
  );
  OR2_X1 _7830_ (
    .A1(_1334_),
    .A2(_1335_),
    .ZN(_1336_)
  );
  AND2_X1 _7831_ (
    .A1(reg_pmp_2_addr[2]),
    .A2(_0792_),
    .ZN(_1337_)
  );
  AND2_X1 _7832_ (
    .A1(reg_dpc[2]),
    .A2(_0750_),
    .ZN(_1338_)
  );
  OR2_X1 _7833_ (
    .A1(_1337_),
    .A2(_1338_),
    .ZN(_1339_)
  );
  OR2_X1 _7834_ (
    .A1(_1336_),
    .A2(_1339_),
    .ZN(_1340_)
  );
  OR2_X1 _7835_ (
    .A1(_1333_),
    .A2(_1340_),
    .ZN(_1341_)
  );
  OR2_X1 _7836_ (
    .A1(_1326_),
    .A2(_1341_),
    .ZN(_1342_)
  );
  OR2_X1 _7837_ (
    .A1(_1318_),
    .A2(_1342_),
    .ZN(_1343_)
  );
  OR2_X1 _7838_ (
    .A1(_1313_),
    .A2(_1343_),
    .ZN(io_rw_rdata[2])
  );
  AND2_X1 _7839_ (
    .A1(io_rw_cmd[1]),
    .A2(_0680_),
    .ZN(_1344_)
  );
  AND2_X1 _7840_ (
    .A1(io_rw_rdata[2]),
    .A2(_1344_),
    .ZN(_1345_)
  );
  OR2_X1 _7841_ (
    .A1(_1291_),
    .A2(_1345_),
    .ZN(_1346_)
  );
  INV_X1 _7842_ (
    .A(_1346_),
    .ZN(_1347_)
  );
  MUX2_X1 _7843_ (
    .A(_1346_),
    .B(reg_pmp_5_addr[2]),
    .S(_1181_),
    .Z(_0029_)
  );
  AND2_X1 _7844_ (
    .A1(io_rw_wdata[3]),
    .A2(_0742_),
    .ZN(_1348_)
  );
  AND2_X1 _7845_ (
    .A1(reg_pmp_4_cfg_a[0]),
    .A2(_0733_),
    .ZN(_1349_)
  );
  AND2_X1 _7846_ (
    .A1(reg_pmp_2_addr[3]),
    .A2(_0792_),
    .ZN(_1350_)
  );
  OR2_X1 _7847_ (
    .A1(_1349_),
    .A2(_1350_),
    .ZN(_1351_)
  );
  AND2_X1 _7848_ (
    .A1(_0775_),
    .A2(_0804_),
    .ZN(_1352_)
  );
  INV_X1 _7849_ (
    .A(_1352_),
    .ZN(_1353_)
  );
  AND2_X1 _7850_ (
    .A1(reg_mie[3]),
    .A2(_1352_),
    .ZN(_1354_)
  );
  AND2_X1 _7851_ (
    .A1(reg_pmp_0_addr[3]),
    .A2(_0837_),
    .ZN(_1355_)
  );
  OR2_X1 _7852_ (
    .A1(_1354_),
    .A2(_1355_),
    .ZN(_1356_)
  );
  OR2_X1 _7853_ (
    .A1(_1351_),
    .A2(_1356_),
    .ZN(_1357_)
  );
  AND2_X1 _7854_ (
    .A1(reg_pmp_4_addr[3]),
    .A2(_0805_),
    .ZN(_1358_)
  );
  AND2_X1 _7855_ (
    .A1(reg_dscratch0[3]),
    .A2(_0797_),
    .ZN(_1359_)
  );
  OR2_X1 _7856_ (
    .A1(_1358_),
    .A2(_1359_),
    .ZN(_1360_)
  );
  AND2_X1 _7857_ (
    .A1(reg_bp_0_address[3]),
    .A2(_0800_),
    .ZN(_1361_)
  );
  AND2_X1 _7858_ (
    .A1(reg_pmp_0_cfg_a[0]),
    .A2(_0754_),
    .ZN(_1362_)
  );
  OR2_X1 _7859_ (
    .A1(_1361_),
    .A2(_1362_),
    .ZN(_1363_)
  );
  OR2_X1 _7860_ (
    .A1(_1360_),
    .A2(_1363_),
    .ZN(_1364_)
  );
  OR2_X1 _7861_ (
    .A1(_1357_),
    .A2(_1364_),
    .ZN(_1365_)
  );
  AND2_X1 _7862_ (
    .A1(reg_mepc[3]),
    .A2(_0783_),
    .ZN(_1366_)
  );
  AND2_X1 _7863_ (
    .A1(_0761_),
    .A2(_0777_),
    .ZN(_1367_)
  );
  AND2_X1 _7864_ (
    .A1(io_interrupts_msip),
    .A2(_1367_),
    .ZN(_1368_)
  );
  OR2_X1 _7865_ (
    .A1(_1366_),
    .A2(_1368_),
    .ZN(_1369_)
  );
  AND2_X1 _7866_ (
    .A1(reg_mscratch[3]),
    .A2(_0767_),
    .ZN(_1370_)
  );
  AND2_X1 _7867_ (
    .A1(reg_mtval[3]),
    .A2(_0764_),
    .ZN(_1371_)
  );
  OR2_X1 _7868_ (
    .A1(_1370_),
    .A2(_1371_),
    .ZN(_1372_)
  );
  OR2_X1 _7869_ (
    .A1(_1369_),
    .A2(_1372_),
    .ZN(_1373_)
  );
  AND2_X1 _7870_ (
    .A1(_0753_),
    .A2(_0775_),
    .ZN(_1374_)
  );
  INV_X1 _7871_ (
    .A(_1374_),
    .ZN(_1375_)
  );
  AND2_X1 _7872_ (
    .A1(reg_mstatus_mie),
    .A2(_1374_),
    .ZN(_1376_)
  );
  AND2_X1 _7873_ (
    .A1(reg_pmp_3_addr[3]),
    .A2(_0844_),
    .ZN(_1377_)
  );
  OR2_X1 _7874_ (
    .A1(_1376_),
    .A2(_1377_),
    .ZN(_1378_)
  );
  AND2_X1 _7875_ (
    .A1(reg_pmp_5_addr[3]),
    .A2(_0788_),
    .ZN(_1379_)
  );
  AND2_X1 _7876_ (
    .A1(reg_mcause[3]),
    .A2(_0834_),
    .ZN(_1380_)
  );
  OR2_X1 _7877_ (
    .A1(_1379_),
    .A2(_1380_),
    .ZN(_1381_)
  );
  OR2_X1 _7878_ (
    .A1(_1378_),
    .A2(_1381_),
    .ZN(_1382_)
  );
  OR2_X1 _7879_ (
    .A1(_1373_),
    .A2(_1382_),
    .ZN(_1383_)
  );
  OR2_X1 _7880_ (
    .A1(_1365_),
    .A2(_1383_),
    .ZN(_1384_)
  );
  AND2_X1 _7881_ (
    .A1(reg_pmp_7_addr[3]),
    .A2(_0849_),
    .ZN(_1385_)
  );
  AND2_X1 _7882_ (
    .A1(reg_pmp_6_addr[3]),
    .A2(_0814_),
    .ZN(_1386_)
  );
  OR2_X1 _7883_ (
    .A1(_1385_),
    .A2(_1386_),
    .ZN(_1387_)
  );
  AND2_X1 _7884_ (
    .A1(large_1[29]),
    .A2(_0851_),
    .ZN(_1388_)
  );
  AND2_X1 _7885_ (
    .A1(small_1[3]),
    .A2(_0830_),
    .ZN(_1389_)
  );
  OR2_X1 _7886_ (
    .A1(_1388_),
    .A2(_1389_),
    .ZN(_1390_)
  );
  OR2_X1 _7887_ (
    .A1(_1387_),
    .A2(_1390_),
    .ZN(_1391_)
  );
  AND2_X1 _7888_ (
    .A1(reg_pmp_1_addr[3]),
    .A2(_0841_),
    .ZN(_1392_)
  );
  AND2_X1 _7889_ (
    .A1(io_rw_addr[6]),
    .A2(io_rw_addr[7]),
    .ZN(_1393_)
  );
  AND2_X1 _7890_ (
    .A1(_0748_),
    .A2(_1393_),
    .ZN(_1394_)
  );
  AND2_X1 _7891_ (
    .A1(reg_custom_0[3]),
    .A2(_1394_),
    .ZN(_1395_)
  );
  OR2_X1 _7892_ (
    .A1(_1392_),
    .A2(_1395_),
    .ZN(_1396_)
  );
  AND2_X1 _7893_ (
    .A1(reg_mtvec[3]),
    .A2(_read_mtvec_T_4[6]),
    .ZN(_1397_)
  );
  AND2_X1 _7894_ (
    .A1(_0780_),
    .A2(_1397_),
    .ZN(_1398_)
  );
  AND2_X1 _7895_ (
    .A1(reg_dpc[3]),
    .A2(_0750_),
    .ZN(_1399_)
  );
  OR2_X1 _7896_ (
    .A1(_1398_),
    .A2(_1399_),
    .ZN(_1400_)
  );
  OR2_X1 _7897_ (
    .A1(_1396_),
    .A2(_1400_),
    .ZN(_1401_)
  );
  AND2_X1 _7898_ (
    .A1(large_[29]),
    .A2(_0827_),
    .ZN(_1402_)
  );
  AND2_X1 _7899_ (
    .A1(small_[3]),
    .A2(_0822_),
    .ZN(_1403_)
  );
  OR2_X1 _7900_ (
    .A1(_1402_),
    .A2(_1403_),
    .ZN(_1404_)
  );
  OR2_X1 _7901_ (
    .A1(_1401_),
    .A2(_1404_),
    .ZN(_1405_)
  );
  OR2_X1 _7902_ (
    .A1(_1391_),
    .A2(_1405_),
    .ZN(_1406_)
  );
  OR2_X1 _7903_ (
    .A1(_1384_),
    .A2(_1406_),
    .ZN(io_rw_rdata[3])
  );
  AND2_X1 _7904_ (
    .A1(io_rw_cmd[1]),
    .A2(_0681_),
    .ZN(_1407_)
  );
  AND2_X1 _7905_ (
    .A1(io_rw_rdata[3]),
    .A2(_1407_),
    .ZN(_1408_)
  );
  OR2_X1 _7906_ (
    .A1(_1348_),
    .A2(_1408_),
    .ZN(_1409_)
  );
  MUX2_X1 _7907_ (
    .A(_1409_),
    .B(reg_pmp_5_addr[3]),
    .S(_1181_),
    .Z(_0030_)
  );
  AND2_X1 _7908_ (
    .A1(io_rw_wdata[4]),
    .A2(_0742_),
    .ZN(_1410_)
  );
  AND2_X1 _7909_ (
    .A1(reg_mscratch[4]),
    .A2(_0767_),
    .ZN(_1411_)
  );
  AND2_X1 _7910_ (
    .A1(reg_mepc[4]),
    .A2(_0783_),
    .ZN(_1412_)
  );
  OR2_X1 _7911_ (
    .A1(_1411_),
    .A2(_1412_),
    .ZN(_1413_)
  );
  AND2_X1 _7912_ (
    .A1(reg_pmp_0_addr[4]),
    .A2(_0837_),
    .ZN(_1414_)
  );
  AND2_X1 _7913_ (
    .A1(reg_pmp_1_addr[4]),
    .A2(_0841_),
    .ZN(_1415_)
  );
  OR2_X1 _7914_ (
    .A1(_1414_),
    .A2(_1415_),
    .ZN(_1416_)
  );
  OR2_X1 _7915_ (
    .A1(_1413_),
    .A2(_1416_),
    .ZN(_1417_)
  );
  AND2_X1 _7916_ (
    .A1(reg_mtvec[4]),
    .A2(_read_mtvec_T_4[6]),
    .ZN(_1418_)
  );
  AND2_X1 _7917_ (
    .A1(_0780_),
    .A2(_1418_),
    .ZN(_1419_)
  );
  AND2_X1 _7918_ (
    .A1(reg_mtval[4]),
    .A2(_0764_),
    .ZN(_1420_)
  );
  OR2_X1 _7919_ (
    .A1(_1419_),
    .A2(_1420_),
    .ZN(_1421_)
  );
  AND2_X1 _7920_ (
    .A1(reg_pmp_5_addr[4]),
    .A2(_0788_),
    .ZN(_1422_)
  );
  AND2_X1 _7921_ (
    .A1(reg_mcause[4]),
    .A2(_0834_),
    .ZN(_1423_)
  );
  OR2_X1 _7922_ (
    .A1(_1422_),
    .A2(_1423_),
    .ZN(_1424_)
  );
  OR2_X1 _7923_ (
    .A1(_1421_),
    .A2(_1424_),
    .ZN(_1425_)
  );
  AND2_X1 _7924_ (
    .A1(reg_pmp_4_addr[4]),
    .A2(_0805_),
    .ZN(_1426_)
  );
  AND2_X1 _7925_ (
    .A1(reg_pmp_0_cfg_a[1]),
    .A2(_0754_),
    .ZN(_1427_)
  );
  OR2_X1 _7926_ (
    .A1(_1426_),
    .A2(_1427_),
    .ZN(_1428_)
  );
  AND2_X1 _7927_ (
    .A1(reg_bp_0_address[4]),
    .A2(_0800_),
    .ZN(_1429_)
  );
  AND2_X1 _7928_ (
    .A1(reg_pmp_4_cfg_a[1]),
    .A2(_0733_),
    .ZN(_1430_)
  );
  OR2_X1 _7929_ (
    .A1(_1429_),
    .A2(_1430_),
    .ZN(_1431_)
  );
  OR2_X1 _7930_ (
    .A1(_1428_),
    .A2(_1431_),
    .ZN(_1432_)
  );
  OR2_X1 _7931_ (
    .A1(_1425_),
    .A2(_1432_),
    .ZN(_1433_)
  );
  OR2_X1 _7932_ (
    .A1(_1417_),
    .A2(_1433_),
    .ZN(_1434_)
  );
  AND2_X1 _7933_ (
    .A1(reg_pmp_6_addr[4]),
    .A2(_0814_),
    .ZN(_1435_)
  );
  AND2_X1 _7934_ (
    .A1(large_1[30]),
    .A2(_0851_),
    .ZN(_1436_)
  );
  OR2_X1 _7935_ (
    .A1(_1435_),
    .A2(_1436_),
    .ZN(_1437_)
  );
  AND2_X1 _7936_ (
    .A1(reg_pmp_7_addr[4]),
    .A2(_0849_),
    .ZN(_1438_)
  );
  AND2_X1 _7937_ (
    .A1(small_1[4]),
    .A2(_0830_),
    .ZN(_1439_)
  );
  OR2_X1 _7938_ (
    .A1(_1438_),
    .A2(_1439_),
    .ZN(_1440_)
  );
  OR2_X1 _7939_ (
    .A1(_1437_),
    .A2(_1440_),
    .ZN(_1441_)
  );
  AND2_X1 _7940_ (
    .A1(reg_pmp_3_addr[4]),
    .A2(_0844_),
    .ZN(_1442_)
  );
  AND2_X1 _7941_ (
    .A1(reg_pmp_2_addr[4]),
    .A2(_0792_),
    .ZN(_1443_)
  );
  OR2_X1 _7942_ (
    .A1(_1442_),
    .A2(_1443_),
    .ZN(_1444_)
  );
  AND2_X1 _7943_ (
    .A1(reg_dpc[4]),
    .A2(_0750_),
    .ZN(_1445_)
  );
  AND2_X1 _7944_ (
    .A1(reg_dscratch0[4]),
    .A2(_0797_),
    .ZN(_1446_)
  );
  OR2_X1 _7945_ (
    .A1(_1445_),
    .A2(_1446_),
    .ZN(_1447_)
  );
  OR2_X1 _7946_ (
    .A1(_1444_),
    .A2(_1447_),
    .ZN(_1448_)
  );
  AND2_X1 _7947_ (
    .A1(large_[30]),
    .A2(_0827_),
    .ZN(_1449_)
  );
  AND2_X1 _7948_ (
    .A1(small_[4]),
    .A2(_0822_),
    .ZN(_1450_)
  );
  OR2_X1 _7949_ (
    .A1(_1449_),
    .A2(_1450_),
    .ZN(_1451_)
  );
  OR2_X1 _7950_ (
    .A1(_1448_),
    .A2(_1451_),
    .ZN(_1452_)
  );
  OR2_X1 _7951_ (
    .A1(_1441_),
    .A2(_1452_),
    .ZN(_1453_)
  );
  OR2_X1 _7952_ (
    .A1(_1434_),
    .A2(_1453_),
    .ZN(io_rw_rdata[4])
  );
  AND2_X1 _7953_ (
    .A1(io_rw_cmd[1]),
    .A2(_0682_),
    .ZN(_1454_)
  );
  AND2_X1 _7954_ (
    .A1(io_rw_rdata[4]),
    .A2(_1454_),
    .ZN(_1455_)
  );
  OR2_X1 _7955_ (
    .A1(_1410_),
    .A2(_1455_),
    .ZN(_1456_)
  );
  MUX2_X1 _7956_ (
    .A(_1456_),
    .B(reg_pmp_5_addr[4]),
    .S(_1181_),
    .Z(_0031_)
  );
  AND2_X1 _7957_ (
    .A1(io_rw_wdata[5]),
    .A2(_0742_),
    .ZN(_1457_)
  );
  AND2_X1 _7958_ (
    .A1(reg_pmp_1_addr[5]),
    .A2(_0841_),
    .ZN(_1458_)
  );
  AND2_X1 _7959_ (
    .A1(reg_pmp_4_addr[5]),
    .A2(_0805_),
    .ZN(_1459_)
  );
  AND2_X1 _7960_ (
    .A1(reg_pmp_2_addr[5]),
    .A2(_0792_),
    .ZN(_1460_)
  );
  AND2_X1 _7961_ (
    .A1(reg_dpc[5]),
    .A2(_0750_),
    .ZN(_1461_)
  );
  AND2_X1 _7962_ (
    .A1(reg_pmp_0_addr[5]),
    .A2(_0837_),
    .ZN(_1462_)
  );
  AND2_X1 _7963_ (
    .A1(reg_bp_0_address[5]),
    .A2(_0800_),
    .ZN(_1463_)
  );
  AND2_X1 _7964_ (
    .A1(reg_mepc[5]),
    .A2(_0783_),
    .ZN(_1464_)
  );
  AND2_X1 _7965_ (
    .A1(reg_mtvec[5]),
    .A2(_read_mtvec_T_4[6]),
    .ZN(_1465_)
  );
  AND2_X1 _7966_ (
    .A1(_0780_),
    .A2(_1465_),
    .ZN(_1466_)
  );
  AND2_X1 _7967_ (
    .A1(reg_pmp_5_addr[5]),
    .A2(_0788_),
    .ZN(_1467_)
  );
  AND2_X1 _7968_ (
    .A1(reg_dscratch0[5]),
    .A2(_0797_),
    .ZN(_1468_)
  );
  AND2_X1 _7969_ (
    .A1(reg_mscratch[5]),
    .A2(_0767_),
    .ZN(_1469_)
  );
  AND2_X1 _7970_ (
    .A1(reg_pmp_3_addr[5]),
    .A2(_0844_),
    .ZN(_1470_)
  );
  AND2_X1 _7971_ (
    .A1(reg_pmp_6_addr[5]),
    .A2(_0814_),
    .ZN(_1471_)
  );
  AND2_X1 _7972_ (
    .A1(reg_pmp_7_addr[5]),
    .A2(_0849_),
    .ZN(_1472_)
  );
  AND2_X1 _7973_ (
    .A1(large_1[31]),
    .A2(_0851_),
    .ZN(_1473_)
  );
  AND2_X1 _7974_ (
    .A1(reg_mtval[5]),
    .A2(_0764_),
    .ZN(_1474_)
  );
  AND2_X1 _7975_ (
    .A1(reg_mcause[5]),
    .A2(_0834_),
    .ZN(_1475_)
  );
  AND2_X1 _7976_ (
    .A1(large_[31]),
    .A2(_0827_),
    .ZN(_1476_)
  );
  OR2_X1 _7977_ (
    .A1(_1458_),
    .A2(_1462_),
    .ZN(_1477_)
  );
  AND2_X1 _7978_ (
    .A1(small_[5]),
    .A2(_0857_),
    .ZN(_1478_)
  );
  AND2_X1 _7979_ (
    .A1(small_1[5]),
    .A2(_0859_),
    .ZN(_1479_)
  );
  OR2_X1 _7980_ (
    .A1(_1460_),
    .A2(_1472_),
    .ZN(_1480_)
  );
  OR2_X1 _7981_ (
    .A1(_1464_),
    .A2(_1475_),
    .ZN(_1481_)
  );
  OR2_X1 _7982_ (
    .A1(_1474_),
    .A2(_1481_),
    .ZN(_1482_)
  );
  OR2_X1 _7983_ (
    .A1(_1480_),
    .A2(_1482_),
    .ZN(_1483_)
  );
  OR2_X1 _7984_ (
    .A1(_1467_),
    .A2(_1477_),
    .ZN(_1484_)
  );
  OR2_X1 _7985_ (
    .A1(_1473_),
    .A2(_1476_),
    .ZN(_1485_)
  );
  OR2_X1 _7986_ (
    .A1(_1484_),
    .A2(_1485_),
    .ZN(_1486_)
  );
  OR2_X1 _7987_ (
    .A1(_1483_),
    .A2(_1486_),
    .ZN(_1487_)
  );
  OR2_X1 _7988_ (
    .A1(_1459_),
    .A2(_1466_),
    .ZN(_1488_)
  );
  OR2_X1 _7989_ (
    .A1(_1471_),
    .A2(_1488_),
    .ZN(_1489_)
  );
  OR2_X1 _7990_ (
    .A1(_1463_),
    .A2(_1469_),
    .ZN(_1490_)
  );
  OR2_X1 _7991_ (
    .A1(_1489_),
    .A2(_1490_),
    .ZN(_1491_)
  );
  OR2_X1 _7992_ (
    .A1(_1461_),
    .A2(_1470_),
    .ZN(_1492_)
  );
  OR2_X1 _7993_ (
    .A1(_1468_),
    .A2(_1478_),
    .ZN(_1493_)
  );
  OR2_X1 _7994_ (
    .A1(_1479_),
    .A2(_1493_),
    .ZN(_1494_)
  );
  OR2_X1 _7995_ (
    .A1(_1492_),
    .A2(_1494_),
    .ZN(_1495_)
  );
  OR2_X1 _7996_ (
    .A1(_1491_),
    .A2(_1495_),
    .ZN(_1496_)
  );
  OR2_X1 _7997_ (
    .A1(_1487_),
    .A2(_1496_),
    .ZN(io_rw_rdata[5])
  );
  AND2_X1 _7998_ (
    .A1(io_rw_cmd[1]),
    .A2(_0683_),
    .ZN(_1497_)
  );
  AND2_X1 _7999_ (
    .A1(io_rw_rdata[5]),
    .A2(_1497_),
    .ZN(_1498_)
  );
  OR2_X1 _8000_ (
    .A1(_1457_),
    .A2(_1498_),
    .ZN(_1499_)
  );
  MUX2_X1 _8001_ (
    .A(_1499_),
    .B(reg_pmp_5_addr[5]),
    .S(_1181_),
    .Z(_0032_)
  );
  AND2_X1 _8002_ (
    .A1(io_rw_wdata[6]),
    .A2(_0742_),
    .ZN(_1500_)
  );
  AND2_X1 _8003_ (
    .A1(reg_pmp_3_addr[6]),
    .A2(_0844_),
    .ZN(_1501_)
  );
  AND2_X1 _8004_ (
    .A1(reg_pmp_2_addr[6]),
    .A2(_0792_),
    .ZN(_1502_)
  );
  AND2_X1 _8005_ (
    .A1(reg_dcsr_cause[0]),
    .A2(_1086_),
    .ZN(_1503_)
  );
  AND2_X1 _8006_ (
    .A1(reg_mepc[6]),
    .A2(_0783_),
    .ZN(_1504_)
  );
  AND2_X1 _8007_ (
    .A1(reg_pmp_5_addr[6]),
    .A2(_0788_),
    .ZN(_1505_)
  );
  AND2_X1 _8008_ (
    .A1(reg_dpc[6]),
    .A2(_0750_),
    .ZN(_1506_)
  );
  AND2_X1 _8009_ (
    .A1(reg_pmp_1_addr[6]),
    .A2(_0841_),
    .ZN(_1507_)
  );
  AND2_X1 _8010_ (
    .A1(reg_pmp_0_addr[6]),
    .A2(_0837_),
    .ZN(_1508_)
  );
  AND2_X1 _8011_ (
    .A1(reg_pmp_4_addr[6]),
    .A2(_0805_),
    .ZN(_1509_)
  );
  AND2_X1 _8012_ (
    .A1(reg_mcause[6]),
    .A2(_0834_),
    .ZN(_1510_)
  );
  AND2_X1 _8013_ (
    .A1(reg_mtval[6]),
    .A2(_0764_),
    .ZN(_1511_)
  );
  AND2_X1 _8014_ (
    .A1(reg_mscratch[6]),
    .A2(_0767_),
    .ZN(_1512_)
  );
  AND2_X1 _8015_ (
    .A1(large_[32]),
    .A2(_0827_),
    .ZN(_1513_)
  );
  AND2_X1 _8016_ (
    .A1(large_1[32]),
    .A2(_0851_),
    .ZN(_1514_)
  );
  AND2_X1 _8017_ (
    .A1(reg_dscratch0[6]),
    .A2(_0797_),
    .ZN(_1515_)
  );
  AND2_X1 _8018_ (
    .A1(reg_bp_0_address[6]),
    .A2(_0800_),
    .ZN(_1516_)
  );
  AND2_X1 _8019_ (
    .A1(reg_mtvec[6]),
    .A2(_read_mtvec_T_4[6]),
    .ZN(_1517_)
  );
  AND2_X1 _8020_ (
    .A1(_0780_),
    .A2(_1517_),
    .ZN(_1518_)
  );
  AND2_X1 _8021_ (
    .A1(reg_pmp_6_addr[6]),
    .A2(_0814_),
    .ZN(_1519_)
  );
  AND2_X1 _8022_ (
    .A1(reg_pmp_7_addr[6]),
    .A2(_0849_),
    .ZN(_1520_)
  );
  OR2_X1 _8023_ (
    .A1(_1502_),
    .A2(_1508_),
    .ZN(_1521_)
  );
  AND2_X1 _8024_ (
    .A1(large_[0]),
    .A2(_0857_),
    .ZN(_1522_)
  );
  AND2_X1 _8025_ (
    .A1(large_1[0]),
    .A2(_0859_),
    .ZN(_1523_)
  );
  OR2_X1 _8026_ (
    .A1(_1505_),
    .A2(_1509_),
    .ZN(_1524_)
  );
  OR2_X1 _8027_ (
    .A1(_1503_),
    .A2(_1524_),
    .ZN(_1525_)
  );
  OR2_X1 _8028_ (
    .A1(_1506_),
    .A2(_1515_),
    .ZN(_1526_)
  );
  OR2_X1 _8029_ (
    .A1(_1504_),
    .A2(_1511_),
    .ZN(_1527_)
  );
  OR2_X1 _8030_ (
    .A1(_1526_),
    .A2(_1527_),
    .ZN(_1528_)
  );
  OR2_X1 _8031_ (
    .A1(_1525_),
    .A2(_1528_),
    .ZN(_1529_)
  );
  OR2_X1 _8032_ (
    .A1(_1510_),
    .A2(_1519_),
    .ZN(_1530_)
  );
  OR2_X1 _8033_ (
    .A1(_1507_),
    .A2(_1530_),
    .ZN(_1531_)
  );
  OR2_X1 _8034_ (
    .A1(_1529_),
    .A2(_1531_),
    .ZN(_1532_)
  );
  OR2_X1 _8035_ (
    .A1(_1058_),
    .A2(_1516_),
    .ZN(_1533_)
  );
  OR2_X1 _8036_ (
    .A1(_1520_),
    .A2(_1533_),
    .ZN(_1534_)
  );
  OR2_X1 _8037_ (
    .A1(_1512_),
    .A2(_1513_),
    .ZN(_1535_)
  );
  OR2_X1 _8038_ (
    .A1(_1534_),
    .A2(_1535_),
    .ZN(_1536_)
  );
  OR2_X1 _8039_ (
    .A1(_1522_),
    .A2(_1523_),
    .ZN(_1537_)
  );
  OR2_X1 _8040_ (
    .A1(_1501_),
    .A2(_1518_),
    .ZN(_1538_)
  );
  OR2_X1 _8041_ (
    .A1(_1537_),
    .A2(_1538_),
    .ZN(_1539_)
  );
  OR2_X1 _8042_ (
    .A1(_1514_),
    .A2(_1521_),
    .ZN(_1540_)
  );
  OR2_X1 _8043_ (
    .A1(_1539_),
    .A2(_1540_),
    .ZN(_1541_)
  );
  OR2_X1 _8044_ (
    .A1(_1536_),
    .A2(_1541_),
    .ZN(_1542_)
  );
  OR2_X1 _8045_ (
    .A1(_1532_),
    .A2(_1542_),
    .ZN(io_rw_rdata[6])
  );
  AND2_X1 _8046_ (
    .A1(io_rw_cmd[1]),
    .A2(_0684_),
    .ZN(_1543_)
  );
  AND2_X1 _8047_ (
    .A1(io_rw_rdata[6]),
    .A2(_1543_),
    .ZN(_1544_)
  );
  OR2_X1 _8048_ (
    .A1(_1500_),
    .A2(_1544_),
    .ZN(_1545_)
  );
  MUX2_X1 _8049_ (
    .A(_1545_),
    .B(reg_pmp_5_addr[6]),
    .S(_1181_),
    .Z(_0033_)
  );
  AND2_X1 _8050_ (
    .A1(io_rw_wdata[7]),
    .A2(_0742_),
    .ZN(_1546_)
  );
  AND2_X1 _8051_ (
    .A1(reg_pmp_0_cfg_l),
    .A2(_0754_),
    .ZN(_1547_)
  );
  AND2_X1 _8052_ (
    .A1(reg_mscratch[7]),
    .A2(_0767_),
    .ZN(_1548_)
  );
  AND2_X1 _8053_ (
    .A1(reg_pmp_4_cfg_l),
    .A2(_0733_),
    .ZN(_1549_)
  );
  AND2_X1 _8054_ (
    .A1(reg_mie[7]),
    .A2(_1352_),
    .ZN(_1550_)
  );
  AND2_X1 _8055_ (
    .A1(reg_dpc[7]),
    .A2(_0750_),
    .ZN(_1551_)
  );
  AND2_X1 _8056_ (
    .A1(reg_bp_0_control_tmatch[0]),
    .A2(_1058_),
    .ZN(_1552_)
  );
  AND2_X1 _8057_ (
    .A1(reg_mtvec[7]),
    .A2(_0780_),
    .ZN(_1553_)
  );
  AND2_X1 _8058_ (
    .A1(reg_pmp_5_addr[7]),
    .A2(_0788_),
    .ZN(_1554_)
  );
  AND2_X1 _8059_ (
    .A1(reg_mtval[7]),
    .A2(_0764_),
    .ZN(_1555_)
  );
  AND2_X1 _8060_ (
    .A1(reg_dscratch0[7]),
    .A2(_0797_),
    .ZN(_1556_)
  );
  AND2_X1 _8061_ (
    .A1(reg_pmp_2_addr[7]),
    .A2(_0792_),
    .ZN(_1557_)
  );
  AND2_X1 _8062_ (
    .A1(reg_pmp_7_addr[7]),
    .A2(_0849_),
    .ZN(_1558_)
  );
  AND2_X1 _8063_ (
    .A1(large_1[33]),
    .A2(_0851_),
    .ZN(_1559_)
  );
  AND2_X1 _8064_ (
    .A1(large_[33]),
    .A2(_0827_),
    .ZN(_1560_)
  );
  AND2_X1 _8065_ (
    .A1(reg_pmp_4_addr[7]),
    .A2(_0805_),
    .ZN(_1561_)
  );
  AND2_X1 _8066_ (
    .A1(reg_pmp_1_addr[7]),
    .A2(_0841_),
    .ZN(_1562_)
  );
  AND2_X1 _8067_ (
    .A1(reg_pmp_6_addr[7]),
    .A2(_0814_),
    .ZN(_1563_)
  );
  AND2_X1 _8068_ (
    .A1(io_interrupts_mtip),
    .A2(_1367_),
    .ZN(_1564_)
  );
  AND2_X1 _8069_ (
    .A1(reg_mcause[7]),
    .A2(_0834_),
    .ZN(_1565_)
  );
  AND2_X1 _8070_ (
    .A1(reg_mstatus_mpie),
    .A2(_1374_),
    .ZN(_1566_)
  );
  AND2_X1 _8071_ (
    .A1(reg_pmp_0_addr[7]),
    .A2(_0837_),
    .ZN(_1567_)
  );
  AND2_X1 _8072_ (
    .A1(reg_dcsr_cause[1]),
    .A2(_1086_),
    .ZN(_1568_)
  );
  AND2_X1 _8073_ (
    .A1(reg_mepc[7]),
    .A2(_0783_),
    .ZN(_1569_)
  );
  AND2_X1 _8074_ (
    .A1(reg_pmp_3_addr[7]),
    .A2(_0844_),
    .ZN(_1570_)
  );
  AND2_X1 _8075_ (
    .A1(reg_bp_0_address[7]),
    .A2(_0800_),
    .ZN(_1571_)
  );
  OR2_X1 _8076_ (
    .A1(_1548_),
    .A2(_1553_),
    .ZN(_1572_)
  );
  AND2_X1 _8077_ (
    .A1(large_1[1]),
    .A2(_0859_),
    .ZN(_1573_)
  );
  OR2_X1 _8078_ (
    .A1(_1555_),
    .A2(_1573_),
    .ZN(_1574_)
  );
  OR2_X1 _8079_ (
    .A1(_1572_),
    .A2(_1574_),
    .ZN(_1575_)
  );
  AND2_X1 _8080_ (
    .A1(large_[1]),
    .A2(_0857_),
    .ZN(_1576_)
  );
  OR2_X1 _8081_ (
    .A1(_1557_),
    .A2(_1562_),
    .ZN(_1577_)
  );
  OR2_X1 _8082_ (
    .A1(_1560_),
    .A2(_1577_),
    .ZN(_1578_)
  );
  OR2_X1 _8083_ (
    .A1(_1550_),
    .A2(_1566_),
    .ZN(_1579_)
  );
  OR2_X1 _8084_ (
    .A1(_1547_),
    .A2(_1549_),
    .ZN(_1580_)
  );
  OR2_X1 _8085_ (
    .A1(_1563_),
    .A2(_1580_),
    .ZN(_1581_)
  );
  OR2_X1 _8086_ (
    .A1(_1561_),
    .A2(_1570_),
    .ZN(_1582_)
  );
  OR2_X1 _8087_ (
    .A1(_1552_),
    .A2(_1582_),
    .ZN(_1583_)
  );
  OR2_X1 _8088_ (
    .A1(_1564_),
    .A2(_1579_),
    .ZN(_1584_)
  );
  OR2_X1 _8089_ (
    .A1(_1554_),
    .A2(_1567_),
    .ZN(_1585_)
  );
  OR2_X1 _8090_ (
    .A1(_1559_),
    .A2(_1585_),
    .ZN(_1586_)
  );
  OR2_X1 _8091_ (
    .A1(_1584_),
    .A2(_1586_),
    .ZN(_1587_)
  );
  OR2_X1 _8092_ (
    .A1(_1583_),
    .A2(_1587_),
    .ZN(_1588_)
  );
  OR2_X1 _8093_ (
    .A1(_1565_),
    .A2(_1568_),
    .ZN(_1589_)
  );
  OR2_X1 _8094_ (
    .A1(_1576_),
    .A2(_1589_),
    .ZN(_1590_)
  );
  OR2_X1 _8095_ (
    .A1(_1556_),
    .A2(_1571_),
    .ZN(_1591_)
  );
  OR2_X1 _8096_ (
    .A1(_1590_),
    .A2(_1591_),
    .ZN(_1592_)
  );
  OR2_X1 _8097_ (
    .A1(_1551_),
    .A2(_1569_),
    .ZN(_1593_)
  );
  OR2_X1 _8098_ (
    .A1(_1575_),
    .A2(_1593_),
    .ZN(_1594_)
  );
  OR2_X1 _8099_ (
    .A1(_1592_),
    .A2(_1594_),
    .ZN(_1595_)
  );
  OR2_X1 _8100_ (
    .A1(_1558_),
    .A2(_1578_),
    .ZN(_1596_)
  );
  OR2_X1 _8101_ (
    .A1(_1581_),
    .A2(_1596_),
    .ZN(_1597_)
  );
  OR2_X1 _8102_ (
    .A1(_1595_),
    .A2(_1597_),
    .ZN(_1598_)
  );
  OR2_X1 _8103_ (
    .A1(_1588_),
    .A2(_1598_),
    .ZN(io_rw_rdata[7])
  );
  AND2_X1 _8104_ (
    .A1(io_rw_cmd[1]),
    .A2(_0685_),
    .ZN(_1599_)
  );
  AND2_X1 _8105_ (
    .A1(io_rw_rdata[7]),
    .A2(_1599_),
    .ZN(_1600_)
  );
  OR2_X1 _8106_ (
    .A1(_1546_),
    .A2(_1600_),
    .ZN(_1601_)
  );
  MUX2_X1 _8107_ (
    .A(_1601_),
    .B(reg_pmp_5_addr[7]),
    .S(_1181_),
    .Z(_0034_)
  );
  MUX2_X1 _8108_ (
    .A(_1129_),
    .B(reg_pmp_5_addr[8]),
    .S(_1181_),
    .Z(_0035_)
  );
  MUX2_X1 _8109_ (
    .A(_1175_),
    .B(reg_pmp_5_addr[9]),
    .S(_1181_),
    .Z(_0036_)
  );
  AND2_X1 _8110_ (
    .A1(io_rw_wdata[10]),
    .A2(_0742_),
    .ZN(_1602_)
  );
  AND2_X1 _8111_ (
    .A1(reg_dscratch0[10]),
    .A2(_0797_),
    .ZN(_1603_)
  );
  AND2_X1 _8112_ (
    .A1(reg_pmp_1_addr[10]),
    .A2(_0841_),
    .ZN(_1604_)
  );
  OR2_X1 _8113_ (
    .A1(_1603_),
    .A2(_1604_),
    .ZN(_1605_)
  );
  AND2_X1 _8114_ (
    .A1(reg_bp_0_address[10]),
    .A2(_0800_),
    .ZN(_1606_)
  );
  AND2_X1 _8115_ (
    .A1(reg_pmp_5_addr[10]),
    .A2(_0788_),
    .ZN(_1607_)
  );
  OR2_X1 _8116_ (
    .A1(_1606_),
    .A2(_1607_),
    .ZN(_1608_)
  );
  OR2_X1 _8117_ (
    .A1(_1605_),
    .A2(_1608_),
    .ZN(_1609_)
  );
  AND2_X1 _8118_ (
    .A1(reg_mepc[10]),
    .A2(_0783_),
    .ZN(_1610_)
  );
  AND2_X1 _8119_ (
    .A1(reg_pmp_0_addr[10]),
    .A2(_0837_),
    .ZN(_1611_)
  );
  OR2_X1 _8120_ (
    .A1(_1610_),
    .A2(_1611_),
    .ZN(_1612_)
  );
  AND2_X1 _8121_ (
    .A1(reg_pmp_1_cfg_x),
    .A2(_0754_),
    .ZN(_1613_)
  );
  AND2_X1 _8122_ (
    .A1(reg_pmp_3_addr[10]),
    .A2(_0844_),
    .ZN(_1614_)
  );
  OR2_X1 _8123_ (
    .A1(_1613_),
    .A2(_1614_),
    .ZN(_1615_)
  );
  OR2_X1 _8124_ (
    .A1(_1612_),
    .A2(_1615_),
    .ZN(_1616_)
  );
  AND2_X1 _8125_ (
    .A1(reg_mtvec[10]),
    .A2(_0780_),
    .ZN(_1617_)
  );
  AND2_X1 _8126_ (
    .A1(reg_mtval[10]),
    .A2(_0764_),
    .ZN(_1618_)
  );
  OR2_X1 _8127_ (
    .A1(_1617_),
    .A2(_1618_),
    .ZN(_1619_)
  );
  AND2_X1 _8128_ (
    .A1(reg_pmp_5_cfg_x),
    .A2(_0733_),
    .ZN(_1620_)
  );
  AND2_X1 _8129_ (
    .A1(reg_mcause[10]),
    .A2(_0834_),
    .ZN(_1621_)
  );
  OR2_X1 _8130_ (
    .A1(_1620_),
    .A2(_1621_),
    .ZN(_1622_)
  );
  OR2_X1 _8131_ (
    .A1(_1619_),
    .A2(_1622_),
    .ZN(_1623_)
  );
  OR2_X1 _8132_ (
    .A1(_1616_),
    .A2(_1623_),
    .ZN(_1624_)
  );
  OR2_X1 _8133_ (
    .A1(_1609_),
    .A2(_1624_),
    .ZN(_1625_)
  );
  AND2_X1 _8134_ (
    .A1(reg_pmp_7_addr[10]),
    .A2(_0849_),
    .ZN(_1626_)
  );
  AND2_X1 _8135_ (
    .A1(large_[36]),
    .A2(_0827_),
    .ZN(_1627_)
  );
  OR2_X1 _8136_ (
    .A1(_1626_),
    .A2(_1627_),
    .ZN(_1628_)
  );
  AND2_X1 _8137_ (
    .A1(large_1[36]),
    .A2(_0851_),
    .ZN(_1629_)
  );
  AND2_X1 _8138_ (
    .A1(large_[4]),
    .A2(_0822_),
    .ZN(_1630_)
  );
  OR2_X1 _8139_ (
    .A1(_1629_),
    .A2(_1630_),
    .ZN(_1631_)
  );
  OR2_X1 _8140_ (
    .A1(_1628_),
    .A2(_1631_),
    .ZN(_1632_)
  );
  AND2_X1 _8141_ (
    .A1(reg_dpc[10]),
    .A2(_0750_),
    .ZN(_1633_)
  );
  AND2_X1 _8142_ (
    .A1(reg_mscratch[10]),
    .A2(_0767_),
    .ZN(_1634_)
  );
  OR2_X1 _8143_ (
    .A1(_1633_),
    .A2(_1634_),
    .ZN(_1635_)
  );
  AND2_X1 _8144_ (
    .A1(reg_pmp_4_addr[10]),
    .A2(_0805_),
    .ZN(_1636_)
  );
  AND2_X1 _8145_ (
    .A1(reg_pmp_2_addr[10]),
    .A2(_0792_),
    .ZN(_1637_)
  );
  OR2_X1 _8146_ (
    .A1(_1636_),
    .A2(_1637_),
    .ZN(_1638_)
  );
  OR2_X1 _8147_ (
    .A1(_1635_),
    .A2(_1638_),
    .ZN(_1639_)
  );
  AND2_X1 _8148_ (
    .A1(reg_pmp_6_addr[10]),
    .A2(_0814_),
    .ZN(_1640_)
  );
  AND2_X1 _8149_ (
    .A1(large_1[4]),
    .A2(_0830_),
    .ZN(_1641_)
  );
  OR2_X1 _8150_ (
    .A1(_1640_),
    .A2(_1641_),
    .ZN(_1642_)
  );
  OR2_X1 _8151_ (
    .A1(_1639_),
    .A2(_1642_),
    .ZN(_1643_)
  );
  OR2_X1 _8152_ (
    .A1(_1632_),
    .A2(_1643_),
    .ZN(_1644_)
  );
  OR2_X1 _8153_ (
    .A1(_1625_),
    .A2(_1644_),
    .ZN(io_rw_rdata[10])
  );
  AND2_X1 _8154_ (
    .A1(io_rw_cmd[1]),
    .A2(_0688_),
    .ZN(_1645_)
  );
  AND2_X1 _8155_ (
    .A1(io_rw_rdata[10]),
    .A2(_1645_),
    .ZN(_1646_)
  );
  OR2_X1 _8156_ (
    .A1(_1602_),
    .A2(_1646_),
    .ZN(_1647_)
  );
  MUX2_X1 _8157_ (
    .A(_1647_),
    .B(reg_pmp_5_addr[10]),
    .S(_1181_),
    .Z(_0037_)
  );
  AND2_X1 _8158_ (
    .A1(io_rw_wdata[11]),
    .A2(_0742_),
    .ZN(_1648_)
  );
  AND2_X1 _8159_ (
    .A1(reg_mtval[11]),
    .A2(_0764_),
    .ZN(_1649_)
  );
  AND2_X1 _8160_ (
    .A1(reg_mscratch[11]),
    .A2(_0767_),
    .ZN(_1650_)
  );
  OR2_X1 _8161_ (
    .A1(_1649_),
    .A2(_1650_),
    .ZN(_1651_)
  );
  AND2_X1 _8162_ (
    .A1(reg_mtvec[11]),
    .A2(_0780_),
    .ZN(_1652_)
  );
  AND2_X1 _8163_ (
    .A1(reg_mepc[11]),
    .A2(_0783_),
    .ZN(_1653_)
  );
  OR2_X1 _8164_ (
    .A1(_1652_),
    .A2(_1653_),
    .ZN(_1654_)
  );
  OR2_X1 _8165_ (
    .A1(_1651_),
    .A2(_1654_),
    .ZN(_1655_)
  );
  AND2_X1 _8166_ (
    .A1(reg_pmp_5_addr[11]),
    .A2(_0788_),
    .ZN(_1656_)
  );
  AND2_X1 _8167_ (
    .A1(reg_pmp_4_addr[11]),
    .A2(_0805_),
    .ZN(_1657_)
  );
  OR2_X1 _8168_ (
    .A1(_1656_),
    .A2(_1657_),
    .ZN(_1658_)
  );
  AND2_X1 _8169_ (
    .A1(reg_mcause[11]),
    .A2(_0834_),
    .ZN(_1659_)
  );
  AND2_X1 _8170_ (
    .A1(reg_dscratch0[11]),
    .A2(_0797_),
    .ZN(_1660_)
  );
  OR2_X1 _8171_ (
    .A1(_1659_),
    .A2(_1660_),
    .ZN(_1661_)
  );
  OR2_X1 _8172_ (
    .A1(_1658_),
    .A2(_1661_),
    .ZN(_1662_)
  );
  OR2_X1 _8173_ (
    .A1(_1655_),
    .A2(_1662_),
    .ZN(_1663_)
  );
  AND2_X1 _8174_ (
    .A1(reg_bp_0_address[11]),
    .A2(_0800_),
    .ZN(_1664_)
  );
  AND2_X1 _8175_ (
    .A1(reg_pmp_1_cfg_a[0]),
    .A2(_0754_),
    .ZN(_1665_)
  );
  AND2_X1 _8176_ (
    .A1(reg_pmp_5_cfg_a[0]),
    .A2(_0733_),
    .ZN(_1666_)
  );
  OR2_X1 _8177_ (
    .A1(_1665_),
    .A2(_1666_),
    .ZN(_1667_)
  );
  OR2_X1 _8178_ (
    .A1(_1664_),
    .A2(_1667_),
    .ZN(_1668_)
  );
  AND2_X1 _8179_ (
    .A1(io_interrupts_meip),
    .A2(_1367_),
    .ZN(_1669_)
  );
  AND2_X1 _8180_ (
    .A1(reg_pmp_2_addr[11]),
    .A2(_0792_),
    .ZN(_1670_)
  );
  OR2_X1 _8181_ (
    .A1(_1669_),
    .A2(_1670_),
    .ZN(_1671_)
  );
  AND2_X1 _8182_ (
    .A1(reg_dpc[11]),
    .A2(_0750_),
    .ZN(_1672_)
  );
  AND2_X1 _8183_ (
    .A1(reg_pmp_1_addr[11]),
    .A2(_0841_),
    .ZN(_1673_)
  );
  OR2_X1 _8184_ (
    .A1(_1672_),
    .A2(_1673_),
    .ZN(_1674_)
  );
  OR2_X1 _8185_ (
    .A1(_1671_),
    .A2(_1674_),
    .ZN(_1675_)
  );
  OR2_X1 _8186_ (
    .A1(_1668_),
    .A2(_1675_),
    .ZN(_1676_)
  );
  OR2_X1 _8187_ (
    .A1(_1663_),
    .A2(_1676_),
    .ZN(_1677_)
  );
  AND2_X1 _8188_ (
    .A1(reg_pmp_7_addr[11]),
    .A2(_0849_),
    .ZN(_1678_)
  );
  AND2_X1 _8189_ (
    .A1(large_1[37]),
    .A2(_0851_),
    .ZN(_1679_)
  );
  OR2_X1 _8190_ (
    .A1(_1678_),
    .A2(_1679_),
    .ZN(_1680_)
  );
  AND2_X1 _8191_ (
    .A1(large_[37]),
    .A2(_0827_),
    .ZN(_1681_)
  );
  AND2_X1 _8192_ (
    .A1(large_1[5]),
    .A2(_0830_),
    .ZN(_1682_)
  );
  OR2_X1 _8193_ (
    .A1(_1681_),
    .A2(_1682_),
    .ZN(_1683_)
  );
  OR2_X1 _8194_ (
    .A1(_1680_),
    .A2(_1683_),
    .ZN(_1684_)
  );
  AND2_X1 _8195_ (
    .A1(reg_pmp_0_addr[11]),
    .A2(_0837_),
    .ZN(_1685_)
  );
  OR2_X1 _8196_ (
    .A1(_1374_),
    .A2(_1685_),
    .ZN(_1686_)
  );
  AND2_X1 _8197_ (
    .A1(reg_mie[11]),
    .A2(_1352_),
    .ZN(_1687_)
  );
  AND2_X1 _8198_ (
    .A1(reg_pmp_3_addr[11]),
    .A2(_0844_),
    .ZN(_1688_)
  );
  OR2_X1 _8199_ (
    .A1(_1687_),
    .A2(_1688_),
    .ZN(_1689_)
  );
  OR2_X1 _8200_ (
    .A1(_1686_),
    .A2(_1689_),
    .ZN(_1690_)
  );
  AND2_X1 _8201_ (
    .A1(reg_pmp_6_addr[11]),
    .A2(_0814_),
    .ZN(_1691_)
  );
  AND2_X1 _8202_ (
    .A1(large_[5]),
    .A2(_0822_),
    .ZN(_1692_)
  );
  OR2_X1 _8203_ (
    .A1(_1691_),
    .A2(_1692_),
    .ZN(_1693_)
  );
  OR2_X1 _8204_ (
    .A1(_1690_),
    .A2(_1693_),
    .ZN(_1694_)
  );
  OR2_X1 _8205_ (
    .A1(_1684_),
    .A2(_1694_),
    .ZN(_1695_)
  );
  OR2_X1 _8206_ (
    .A1(_1677_),
    .A2(_1695_),
    .ZN(io_rw_rdata[11])
  );
  AND2_X1 _8207_ (
    .A1(io_rw_cmd[1]),
    .A2(_0689_),
    .ZN(_1696_)
  );
  AND2_X1 _8208_ (
    .A1(io_rw_rdata[11]),
    .A2(_1696_),
    .ZN(_1697_)
  );
  OR2_X1 _8209_ (
    .A1(_1648_),
    .A2(_1697_),
    .ZN(_1698_)
  );
  MUX2_X1 _8210_ (
    .A(_1698_),
    .B(reg_pmp_5_addr[11]),
    .S(_1181_),
    .Z(_0038_)
  );
  AND2_X1 _8211_ (
    .A1(reg_pmp_1_addr[12]),
    .A2(_0841_),
    .ZN(_1699_)
  );
  AND2_X1 _8212_ (
    .A1(reg_mepc[12]),
    .A2(_0783_),
    .ZN(_1700_)
  );
  OR2_X1 _8213_ (
    .A1(_1699_),
    .A2(_1700_),
    .ZN(_1701_)
  );
  AND2_X1 _8214_ (
    .A1(reg_dscratch0[12]),
    .A2(_0797_),
    .ZN(_1702_)
  );
  AND2_X1 _8215_ (
    .A1(reg_dpc[12]),
    .A2(_0750_),
    .ZN(_1703_)
  );
  OR2_X1 _8216_ (
    .A1(_1702_),
    .A2(_1703_),
    .ZN(_1704_)
  );
  OR2_X1 _8217_ (
    .A1(_1701_),
    .A2(_1704_),
    .ZN(_1705_)
  );
  AND2_X1 _8218_ (
    .A1(reg_pmp_2_addr[12]),
    .A2(_0792_),
    .ZN(_1706_)
  );
  AND2_X1 _8219_ (
    .A1(reg_pmp_0_addr[12]),
    .A2(_0837_),
    .ZN(_1707_)
  );
  OR2_X1 _8220_ (
    .A1(_1706_),
    .A2(_1707_),
    .ZN(_1708_)
  );
  AND2_X1 _8221_ (
    .A1(reg_pmp_5_addr[12]),
    .A2(_0788_),
    .ZN(_1709_)
  );
  AND2_X1 _8222_ (
    .A1(reg_pmp_4_addr[12]),
    .A2(_0805_),
    .ZN(_1710_)
  );
  OR2_X1 _8223_ (
    .A1(_1709_),
    .A2(_1710_),
    .ZN(_1711_)
  );
  OR2_X1 _8224_ (
    .A1(_1708_),
    .A2(_1711_),
    .ZN(_1712_)
  );
  OR2_X1 _8225_ (
    .A1(_1705_),
    .A2(_1712_),
    .ZN(_1713_)
  );
  AND2_X1 _8226_ (
    .A1(reg_mtval[12]),
    .A2(_0764_),
    .ZN(_1714_)
  );
  AND2_X1 _8227_ (
    .A1(reg_mcause[12]),
    .A2(_0834_),
    .ZN(_1715_)
  );
  OR2_X1 _8228_ (
    .A1(_1714_),
    .A2(_1715_),
    .ZN(_1716_)
  );
  AND2_X1 _8229_ (
    .A1(reg_mscratch[12]),
    .A2(_0767_),
    .ZN(_1717_)
  );
  AND2_X1 _8230_ (
    .A1(reg_mtvec[12]),
    .A2(_0780_),
    .ZN(_1718_)
  );
  OR2_X1 _8231_ (
    .A1(_1717_),
    .A2(_1718_),
    .ZN(_1719_)
  );
  OR2_X1 _8232_ (
    .A1(_1716_),
    .A2(_1719_),
    .ZN(_1720_)
  );
  AND2_X1 _8233_ (
    .A1(reg_bp_0_control_action),
    .A2(_1058_),
    .ZN(_1721_)
  );
  AND2_X1 _8234_ (
    .A1(reg_pmp_3_addr[12]),
    .A2(_0844_),
    .ZN(_1722_)
  );
  OR2_X1 _8235_ (
    .A1(_1721_),
    .A2(_1722_),
    .ZN(_1723_)
  );
  AND2_X1 _8236_ (
    .A1(reg_misa[12]),
    .A2(_1057_),
    .ZN(_1724_)
  );
  AND2_X1 _8237_ (
    .A1(reg_pmp_5_cfg_a[1]),
    .A2(_0733_),
    .ZN(_1725_)
  );
  OR2_X1 _8238_ (
    .A1(_1724_),
    .A2(_1725_),
    .ZN(_1726_)
  );
  OR2_X1 _8239_ (
    .A1(_1723_),
    .A2(_1726_),
    .ZN(_1727_)
  );
  OR2_X1 _8240_ (
    .A1(_1720_),
    .A2(_1727_),
    .ZN(_1728_)
  );
  OR2_X1 _8241_ (
    .A1(_1713_),
    .A2(_1728_),
    .ZN(_1729_)
  );
  AND2_X1 _8242_ (
    .A1(reg_pmp_7_addr[12]),
    .A2(_0849_),
    .ZN(_1730_)
  );
  AND2_X1 _8243_ (
    .A1(large_[6]),
    .A2(_0822_),
    .ZN(_1731_)
  );
  OR2_X1 _8244_ (
    .A1(_1730_),
    .A2(_1731_),
    .ZN(_1732_)
  );
  AND2_X1 _8245_ (
    .A1(large_1[38]),
    .A2(_0851_),
    .ZN(_1733_)
  );
  AND2_X1 _8246_ (
    .A1(reg_pmp_6_addr[12]),
    .A2(_0814_),
    .ZN(_1734_)
  );
  OR2_X1 _8247_ (
    .A1(_1733_),
    .A2(_1734_),
    .ZN(_1735_)
  );
  OR2_X1 _8248_ (
    .A1(_1732_),
    .A2(_1735_),
    .ZN(_1736_)
  );
  OR2_X1 _8249_ (
    .A1(_0926_),
    .A2(_1374_),
    .ZN(_1737_)
  );
  AND2_X1 _8250_ (
    .A1(reg_bp_0_address[12]),
    .A2(_0800_),
    .ZN(_1738_)
  );
  AND2_X1 _8251_ (
    .A1(reg_pmp_1_cfg_a[1]),
    .A2(_0754_),
    .ZN(_1739_)
  );
  OR2_X1 _8252_ (
    .A1(_1738_),
    .A2(_1739_),
    .ZN(_1740_)
  );
  OR2_X1 _8253_ (
    .A1(_1737_),
    .A2(_1740_),
    .ZN(_1741_)
  );
  AND2_X1 _8254_ (
    .A1(large_[38]),
    .A2(_0827_),
    .ZN(_1742_)
  );
  AND2_X1 _8255_ (
    .A1(large_1[6]),
    .A2(_0830_),
    .ZN(_1743_)
  );
  OR2_X1 _8256_ (
    .A1(_1742_),
    .A2(_1743_),
    .ZN(_1744_)
  );
  OR2_X1 _8257_ (
    .A1(_1741_),
    .A2(_1744_),
    .ZN(_1745_)
  );
  OR2_X1 _8258_ (
    .A1(_1736_),
    .A2(_1745_),
    .ZN(_1746_)
  );
  OR2_X1 _8259_ (
    .A1(_1729_),
    .A2(_1746_),
    .ZN(io_rw_rdata[12])
  );
  AND2_X1 _8260_ (
    .A1(io_rw_cmd[1]),
    .A2(io_rw_rdata[12]),
    .ZN(_1747_)
  );
  MUX2_X1 _8261_ (
    .A(_1747_),
    .B(_0742_),
    .S(io_rw_wdata[12]),
    .Z(_1748_)
  );
  MUX2_X1 _8262_ (
    .A(_1748_),
    .B(reg_pmp_5_addr[12]),
    .S(_1181_),
    .Z(_0039_)
  );
  AND2_X1 _8263_ (
    .A1(io_rw_wdata[13]),
    .A2(_0742_),
    .ZN(_1749_)
  );
  AND2_X1 _8264_ (
    .A1(reg_pmp_3_addr[13]),
    .A2(_0844_),
    .ZN(_1750_)
  );
  AND2_X1 _8265_ (
    .A1(reg_mepc[13]),
    .A2(_0783_),
    .ZN(_1751_)
  );
  OR2_X1 _8266_ (
    .A1(_1750_),
    .A2(_1751_),
    .ZN(_1752_)
  );
  AND2_X1 _8267_ (
    .A1(reg_mtval[13]),
    .A2(_0764_),
    .ZN(_1753_)
  );
  AND2_X1 _8268_ (
    .A1(reg_pmp_4_addr[13]),
    .A2(_0805_),
    .ZN(_1754_)
  );
  OR2_X1 _8269_ (
    .A1(_1753_),
    .A2(_1754_),
    .ZN(_1755_)
  );
  OR2_X1 _8270_ (
    .A1(_1752_),
    .A2(_1755_),
    .ZN(_1756_)
  );
  AND2_X1 _8271_ (
    .A1(reg_dscratch0[13]),
    .A2(_0797_),
    .ZN(_1757_)
  );
  AND2_X1 _8272_ (
    .A1(reg_pmp_1_addr[13]),
    .A2(_0841_),
    .ZN(_1758_)
  );
  OR2_X1 _8273_ (
    .A1(_1757_),
    .A2(_1758_),
    .ZN(_1759_)
  );
  AND2_X1 _8274_ (
    .A1(reg_mscratch[13]),
    .A2(_0767_),
    .ZN(_1760_)
  );
  AND2_X1 _8275_ (
    .A1(reg_mtvec[13]),
    .A2(_0780_),
    .ZN(_1761_)
  );
  OR2_X1 _8276_ (
    .A1(_1760_),
    .A2(_1761_),
    .ZN(_1762_)
  );
  OR2_X1 _8277_ (
    .A1(_1759_),
    .A2(_1762_),
    .ZN(_1763_)
  );
  AND2_X1 _8278_ (
    .A1(reg_bp_0_address[13]),
    .A2(_0800_),
    .ZN(_1764_)
  );
  AND2_X1 _8279_ (
    .A1(reg_pmp_5_addr[13]),
    .A2(_0788_),
    .ZN(_1765_)
  );
  OR2_X1 _8280_ (
    .A1(_1764_),
    .A2(_1765_),
    .ZN(_1766_)
  );
  AND2_X1 _8281_ (
    .A1(reg_pmp_0_addr[13]),
    .A2(_0837_),
    .ZN(_1767_)
  );
  AND2_X1 _8282_ (
    .A1(reg_dpc[13]),
    .A2(_0750_),
    .ZN(_1768_)
  );
  OR2_X1 _8283_ (
    .A1(_1767_),
    .A2(_1768_),
    .ZN(_1769_)
  );
  OR2_X1 _8284_ (
    .A1(_1766_),
    .A2(_1769_),
    .ZN(_1770_)
  );
  OR2_X1 _8285_ (
    .A1(_1763_),
    .A2(_1770_),
    .ZN(_1771_)
  );
  OR2_X1 _8286_ (
    .A1(_1756_),
    .A2(_1771_),
    .ZN(_1772_)
  );
  AND2_X1 _8287_ (
    .A1(reg_pmp_7_addr[13]),
    .A2(_0849_),
    .ZN(_1773_)
  );
  AND2_X1 _8288_ (
    .A1(large_[39]),
    .A2(_0827_),
    .ZN(_1774_)
  );
  AND2_X1 _8289_ (
    .A1(large_1[7]),
    .A2(_0830_),
    .ZN(_1775_)
  );
  OR2_X1 _8290_ (
    .A1(_1774_),
    .A2(_1775_),
    .ZN(_1776_)
  );
  OR2_X1 _8291_ (
    .A1(_1773_),
    .A2(_1776_),
    .ZN(_1777_)
  );
  AND2_X1 _8292_ (
    .A1(large_1[39]),
    .A2(_0851_),
    .ZN(_1778_)
  );
  AND2_X1 _8293_ (
    .A1(reg_pmp_2_addr[13]),
    .A2(_0792_),
    .ZN(_1779_)
  );
  AND2_X1 _8294_ (
    .A1(reg_mcause[13]),
    .A2(_0834_),
    .ZN(_1780_)
  );
  OR2_X1 _8295_ (
    .A1(_1779_),
    .A2(_1780_),
    .ZN(_1781_)
  );
  OR2_X1 _8296_ (
    .A1(_1778_),
    .A2(_1781_),
    .ZN(_1782_)
  );
  AND2_X1 _8297_ (
    .A1(reg_pmp_6_addr[13]),
    .A2(_0814_),
    .ZN(_1783_)
  );
  AND2_X1 _8298_ (
    .A1(large_[7]),
    .A2(_0822_),
    .ZN(_1784_)
  );
  OR2_X1 _8299_ (
    .A1(_1783_),
    .A2(_1784_),
    .ZN(_1785_)
  );
  OR2_X1 _8300_ (
    .A1(_1782_),
    .A2(_1785_),
    .ZN(_1786_)
  );
  OR2_X1 _8301_ (
    .A1(_1777_),
    .A2(_1786_),
    .ZN(_1787_)
  );
  OR2_X1 _8302_ (
    .A1(_1772_),
    .A2(_1787_),
    .ZN(io_rw_rdata[13])
  );
  AND2_X1 _8303_ (
    .A1(io_rw_cmd[1]),
    .A2(_0690_),
    .ZN(_1788_)
  );
  AND2_X1 _8304_ (
    .A1(io_rw_rdata[13]),
    .A2(_1788_),
    .ZN(_1789_)
  );
  OR2_X1 _8305_ (
    .A1(_1749_),
    .A2(_1789_),
    .ZN(_1790_)
  );
  MUX2_X1 _8306_ (
    .A(_1790_),
    .B(reg_pmp_5_addr[13]),
    .S(_1181_),
    .Z(_0040_)
  );
  AND2_X1 _8307_ (
    .A1(io_rw_wdata[14]),
    .A2(_0742_),
    .ZN(_1791_)
  );
  AND2_X1 _8308_ (
    .A1(reg_pmp_0_addr[14]),
    .A2(_0837_),
    .ZN(_1792_)
  );
  AND2_X1 _8309_ (
    .A1(reg_dscratch0[14]),
    .A2(_0797_),
    .ZN(_1793_)
  );
  OR2_X1 _8310_ (
    .A1(_1792_),
    .A2(_1793_),
    .ZN(_1794_)
  );
  AND2_X1 _8311_ (
    .A1(reg_pmp_3_addr[14]),
    .A2(_0844_),
    .ZN(_1795_)
  );
  AND2_X1 _8312_ (
    .A1(reg_mtvec[14]),
    .A2(_0780_),
    .ZN(_1796_)
  );
  OR2_X1 _8313_ (
    .A1(_1795_),
    .A2(_1796_),
    .ZN(_1797_)
  );
  OR2_X1 _8314_ (
    .A1(_1794_),
    .A2(_1797_),
    .ZN(_1798_)
  );
  AND2_X1 _8315_ (
    .A1(reg_dpc[14]),
    .A2(_0750_),
    .ZN(_1799_)
  );
  AND2_X1 _8316_ (
    .A1(reg_bp_0_address[14]),
    .A2(_0800_),
    .ZN(_1800_)
  );
  OR2_X1 _8317_ (
    .A1(_1799_),
    .A2(_1800_),
    .ZN(_1801_)
  );
  AND2_X1 _8318_ (
    .A1(reg_pmp_5_addr[14]),
    .A2(_0788_),
    .ZN(_1802_)
  );
  AND2_X1 _8319_ (
    .A1(reg_pmp_1_addr[14]),
    .A2(_0841_),
    .ZN(_1803_)
  );
  OR2_X1 _8320_ (
    .A1(_1802_),
    .A2(_1803_),
    .ZN(_1804_)
  );
  OR2_X1 _8321_ (
    .A1(_1801_),
    .A2(_1804_),
    .ZN(_1805_)
  );
  AND2_X1 _8322_ (
    .A1(reg_mscratch[14]),
    .A2(_0767_),
    .ZN(_1806_)
  );
  AND2_X1 _8323_ (
    .A1(reg_mcause[14]),
    .A2(_0834_),
    .ZN(_1807_)
  );
  OR2_X1 _8324_ (
    .A1(_1806_),
    .A2(_1807_),
    .ZN(_1808_)
  );
  AND2_X1 _8325_ (
    .A1(reg_mepc[14]),
    .A2(_0783_),
    .ZN(_1809_)
  );
  AND2_X1 _8326_ (
    .A1(reg_mtval[14]),
    .A2(_0764_),
    .ZN(_1810_)
  );
  OR2_X1 _8327_ (
    .A1(_1809_),
    .A2(_1810_),
    .ZN(_1811_)
  );
  OR2_X1 _8328_ (
    .A1(_1808_),
    .A2(_1811_),
    .ZN(_1812_)
  );
  OR2_X1 _8329_ (
    .A1(_1805_),
    .A2(_1812_),
    .ZN(_1813_)
  );
  OR2_X1 _8330_ (
    .A1(_1798_),
    .A2(_1813_),
    .ZN(_1814_)
  );
  AND2_X1 _8331_ (
    .A1(large_1[8]),
    .A2(_0830_),
    .ZN(_1815_)
  );
  AND2_X1 _8332_ (
    .A1(reg_pmp_6_addr[14]),
    .A2(_0814_),
    .ZN(_1816_)
  );
  AND2_X1 _8333_ (
    .A1(reg_pmp_7_addr[14]),
    .A2(_0849_),
    .ZN(_1817_)
  );
  OR2_X1 _8334_ (
    .A1(_1816_),
    .A2(_1817_),
    .ZN(_1818_)
  );
  OR2_X1 _8335_ (
    .A1(_1815_),
    .A2(_1818_),
    .ZN(_1819_)
  );
  AND2_X1 _8336_ (
    .A1(large_[8]),
    .A2(_0822_),
    .ZN(_1820_)
  );
  AND2_X1 _8337_ (
    .A1(reg_pmp_4_addr[14]),
    .A2(_0805_),
    .ZN(_1821_)
  );
  AND2_X1 _8338_ (
    .A1(reg_pmp_2_addr[14]),
    .A2(_0792_),
    .ZN(_1822_)
  );
  OR2_X1 _8339_ (
    .A1(_1821_),
    .A2(_1822_),
    .ZN(_1823_)
  );
  OR2_X1 _8340_ (
    .A1(_1820_),
    .A2(_1823_),
    .ZN(_1824_)
  );
  AND2_X1 _8341_ (
    .A1(large_1[40]),
    .A2(_0851_),
    .ZN(_1825_)
  );
  AND2_X1 _8342_ (
    .A1(large_[40]),
    .A2(_0827_),
    .ZN(_1826_)
  );
  OR2_X1 _8343_ (
    .A1(_1825_),
    .A2(_1826_),
    .ZN(_1827_)
  );
  OR2_X1 _8344_ (
    .A1(_1824_),
    .A2(_1827_),
    .ZN(_1828_)
  );
  OR2_X1 _8345_ (
    .A1(_1819_),
    .A2(_1828_),
    .ZN(_1829_)
  );
  OR2_X1 _8346_ (
    .A1(_1814_),
    .A2(_1829_),
    .ZN(io_rw_rdata[14])
  );
  AND2_X1 _8347_ (
    .A1(io_rw_cmd[1]),
    .A2(_0691_),
    .ZN(_1830_)
  );
  AND2_X1 _8348_ (
    .A1(io_rw_rdata[14]),
    .A2(_1830_),
    .ZN(_1831_)
  );
  OR2_X1 _8349_ (
    .A1(_1791_),
    .A2(_1831_),
    .ZN(_1832_)
  );
  MUX2_X1 _8350_ (
    .A(_1832_),
    .B(reg_pmp_5_addr[14]),
    .S(_1181_),
    .Z(_0041_)
  );
  AND2_X1 _8351_ (
    .A1(io_rw_wdata[15]),
    .A2(_0742_),
    .ZN(_1833_)
  );
  AND2_X1 _8352_ (
    .A1(reg_pmp_5_cfg_l),
    .A2(_0733_),
    .ZN(_1834_)
  );
  AND2_X1 _8353_ (
    .A1(reg_pmp_1_cfg_l),
    .A2(_0754_),
    .ZN(_1835_)
  );
  OR2_X1 _8354_ (
    .A1(_1834_),
    .A2(_1835_),
    .ZN(_1836_)
  );
  AND2_X1 _8355_ (
    .A1(reg_pmp_2_addr[15]),
    .A2(_0792_),
    .ZN(_1837_)
  );
  AND2_X1 _8356_ (
    .A1(reg_bp_0_address[15]),
    .A2(_0800_),
    .ZN(_1838_)
  );
  OR2_X1 _8357_ (
    .A1(_1837_),
    .A2(_1838_),
    .ZN(_1839_)
  );
  OR2_X1 _8358_ (
    .A1(_1836_),
    .A2(_1839_),
    .ZN(_1840_)
  );
  AND2_X1 _8359_ (
    .A1(reg_pmp_1_addr[15]),
    .A2(_0841_),
    .ZN(_1841_)
  );
  AND2_X1 _8360_ (
    .A1(reg_pmp_3_addr[15]),
    .A2(_0844_),
    .ZN(_1842_)
  );
  OR2_X1 _8361_ (
    .A1(_1841_),
    .A2(_1842_),
    .ZN(_1843_)
  );
  AND2_X1 _8362_ (
    .A1(reg_dcsr_ebreakm),
    .A2(_1086_),
    .ZN(_1844_)
  );
  AND2_X1 _8363_ (
    .A1(reg_pmp_5_addr[15]),
    .A2(_0788_),
    .ZN(_1845_)
  );
  OR2_X1 _8364_ (
    .A1(_1844_),
    .A2(_1845_),
    .ZN(_1846_)
  );
  OR2_X1 _8365_ (
    .A1(_1843_),
    .A2(_1846_),
    .ZN(_1847_)
  );
  OR2_X1 _8366_ (
    .A1(_1840_),
    .A2(_1847_),
    .ZN(_1848_)
  );
  AND2_X1 _8367_ (
    .A1(reg_mtvec[15]),
    .A2(_0780_),
    .ZN(_1849_)
  );
  AND2_X1 _8368_ (
    .A1(reg_dscratch0[15]),
    .A2(_0797_),
    .ZN(_1850_)
  );
  AND2_X1 _8369_ (
    .A1(reg_mtval[15]),
    .A2(_0764_),
    .ZN(_1851_)
  );
  OR2_X1 _8370_ (
    .A1(_1850_),
    .A2(_1851_),
    .ZN(_1852_)
  );
  OR2_X1 _8371_ (
    .A1(_1849_),
    .A2(_1852_),
    .ZN(_1853_)
  );
  AND2_X1 _8372_ (
    .A1(reg_dpc[15]),
    .A2(_0750_),
    .ZN(_1854_)
  );
  AND2_X1 _8373_ (
    .A1(reg_mepc[15]),
    .A2(_0783_),
    .ZN(_1855_)
  );
  OR2_X1 _8374_ (
    .A1(_1854_),
    .A2(_1855_),
    .ZN(_1856_)
  );
  AND2_X1 _8375_ (
    .A1(reg_mscratch[15]),
    .A2(_0767_),
    .ZN(_1857_)
  );
  AND2_X1 _8376_ (
    .A1(reg_mcause[15]),
    .A2(_0834_),
    .ZN(_1858_)
  );
  OR2_X1 _8377_ (
    .A1(_1857_),
    .A2(_1858_),
    .ZN(_1859_)
  );
  OR2_X1 _8378_ (
    .A1(_1856_),
    .A2(_1859_),
    .ZN(_1860_)
  );
  OR2_X1 _8379_ (
    .A1(_1853_),
    .A2(_1860_),
    .ZN(_1861_)
  );
  OR2_X1 _8380_ (
    .A1(_1848_),
    .A2(_1861_),
    .ZN(_1862_)
  );
  AND2_X1 _8381_ (
    .A1(large_1[9]),
    .A2(_0830_),
    .ZN(_1863_)
  );
  AND2_X1 _8382_ (
    .A1(large_1[41]),
    .A2(_0851_),
    .ZN(_1864_)
  );
  AND2_X1 _8383_ (
    .A1(large_[9]),
    .A2(_0822_),
    .ZN(_1865_)
  );
  OR2_X1 _8384_ (
    .A1(_1864_),
    .A2(_1865_),
    .ZN(_1866_)
  );
  OR2_X1 _8385_ (
    .A1(_1863_),
    .A2(_1866_),
    .ZN(_1867_)
  );
  AND2_X1 _8386_ (
    .A1(reg_pmp_6_addr[15]),
    .A2(_0814_),
    .ZN(_1868_)
  );
  AND2_X1 _8387_ (
    .A1(reg_pmp_4_addr[15]),
    .A2(_0805_),
    .ZN(_1869_)
  );
  AND2_X1 _8388_ (
    .A1(reg_pmp_0_addr[15]),
    .A2(_0837_),
    .ZN(_1870_)
  );
  OR2_X1 _8389_ (
    .A1(_1869_),
    .A2(_1870_),
    .ZN(_1871_)
  );
  OR2_X1 _8390_ (
    .A1(_1868_),
    .A2(_1871_),
    .ZN(_1872_)
  );
  AND2_X1 _8391_ (
    .A1(reg_pmp_7_addr[15]),
    .A2(_0849_),
    .ZN(_1873_)
  );
  AND2_X1 _8392_ (
    .A1(large_[41]),
    .A2(_0827_),
    .ZN(_1874_)
  );
  OR2_X1 _8393_ (
    .A1(_1873_),
    .A2(_1874_),
    .ZN(_1875_)
  );
  OR2_X1 _8394_ (
    .A1(_1872_),
    .A2(_1875_),
    .ZN(_1876_)
  );
  OR2_X1 _8395_ (
    .A1(_1867_),
    .A2(_1876_),
    .ZN(_1877_)
  );
  OR2_X1 _8396_ (
    .A1(_1862_),
    .A2(_1877_),
    .ZN(io_rw_rdata[15])
  );
  AND2_X1 _8397_ (
    .A1(io_rw_cmd[1]),
    .A2(_0692_),
    .ZN(_1878_)
  );
  AND2_X1 _8398_ (
    .A1(io_rw_rdata[15]),
    .A2(_1878_),
    .ZN(_1879_)
  );
  OR2_X1 _8399_ (
    .A1(_1833_),
    .A2(_1879_),
    .ZN(_1880_)
  );
  MUX2_X1 _8400_ (
    .A(_1880_),
    .B(reg_pmp_5_addr[15]),
    .S(_1181_),
    .Z(_0042_)
  );
  MUX2_X1 _8401_ (
    .A(_0862_),
    .B(reg_pmp_5_addr[16]),
    .S(_1181_),
    .Z(_0043_)
  );
  AND2_X1 _8402_ (
    .A1(io_rw_wdata[17]),
    .A2(_0742_),
    .ZN(_1881_)
  );
  AND2_X1 _8403_ (
    .A1(reg_mcause[17]),
    .A2(_0834_),
    .ZN(_1882_)
  );
  AND2_X1 _8404_ (
    .A1(reg_mscratch[17]),
    .A2(_0767_),
    .ZN(_1883_)
  );
  OR2_X1 _8405_ (
    .A1(_1882_),
    .A2(_1883_),
    .ZN(_1884_)
  );
  AND2_X1 _8406_ (
    .A1(reg_mtvec[17]),
    .A2(_0780_),
    .ZN(_1885_)
  );
  AND2_X1 _8407_ (
    .A1(reg_mepc[17]),
    .A2(_0783_),
    .ZN(_1886_)
  );
  OR2_X1 _8408_ (
    .A1(_1885_),
    .A2(_1886_),
    .ZN(_1887_)
  );
  OR2_X1 _8409_ (
    .A1(_1884_),
    .A2(_1887_),
    .ZN(_1888_)
  );
  AND2_X1 _8410_ (
    .A1(reg_mtval[17]),
    .A2(_0764_),
    .ZN(_1889_)
  );
  AND2_X1 _8411_ (
    .A1(reg_dpc[17]),
    .A2(_0750_),
    .ZN(_1890_)
  );
  OR2_X1 _8412_ (
    .A1(_1889_),
    .A2(_1890_),
    .ZN(_1891_)
  );
  AND2_X1 _8413_ (
    .A1(reg_pmp_4_addr[17]),
    .A2(_0805_),
    .ZN(_1892_)
  );
  AND2_X1 _8414_ (
    .A1(reg_pmp_6_cfg_w),
    .A2(_0733_),
    .ZN(_1893_)
  );
  OR2_X1 _8415_ (
    .A1(_1892_),
    .A2(_1893_),
    .ZN(_1894_)
  );
  OR2_X1 _8416_ (
    .A1(_1891_),
    .A2(_1894_),
    .ZN(_1895_)
  );
  AND2_X1 _8417_ (
    .A1(reg_bp_0_address[17]),
    .A2(_0800_),
    .ZN(_1896_)
  );
  AND2_X1 _8418_ (
    .A1(reg_pmp_5_addr[17]),
    .A2(_0788_),
    .ZN(_1897_)
  );
  OR2_X1 _8419_ (
    .A1(_1896_),
    .A2(_1897_),
    .ZN(_1898_)
  );
  AND2_X1 _8420_ (
    .A1(reg_pmp_2_cfg_w),
    .A2(_0754_),
    .ZN(_1899_)
  );
  AND2_X1 _8421_ (
    .A1(reg_dscratch0[17]),
    .A2(_0797_),
    .ZN(_1900_)
  );
  OR2_X1 _8422_ (
    .A1(_1899_),
    .A2(_1900_),
    .ZN(_1901_)
  );
  OR2_X1 _8423_ (
    .A1(_1898_),
    .A2(_1901_),
    .ZN(_1902_)
  );
  OR2_X1 _8424_ (
    .A1(_1895_),
    .A2(_1902_),
    .ZN(_1903_)
  );
  OR2_X1 _8425_ (
    .A1(_1888_),
    .A2(_1903_),
    .ZN(_1904_)
  );
  AND2_X1 _8426_ (
    .A1(reg_pmp_7_addr[17]),
    .A2(_0849_),
    .ZN(_1905_)
  );
  AND2_X1 _8427_ (
    .A1(large_[11]),
    .A2(_0822_),
    .ZN(_1906_)
  );
  OR2_X1 _8428_ (
    .A1(_1905_),
    .A2(_1906_),
    .ZN(_1907_)
  );
  AND2_X1 _8429_ (
    .A1(reg_pmp_6_addr[17]),
    .A2(_0814_),
    .ZN(_1908_)
  );
  AND2_X1 _8430_ (
    .A1(large_1[11]),
    .A2(_0830_),
    .ZN(_1909_)
  );
  OR2_X1 _8431_ (
    .A1(_1908_),
    .A2(_1909_),
    .ZN(_1910_)
  );
  OR2_X1 _8432_ (
    .A1(_1907_),
    .A2(_1910_),
    .ZN(_1911_)
  );
  AND2_X1 _8433_ (
    .A1(reg_pmp_3_addr[17]),
    .A2(_0844_),
    .ZN(_1912_)
  );
  AND2_X1 _8434_ (
    .A1(reg_pmp_1_addr[17]),
    .A2(_0841_),
    .ZN(_1913_)
  );
  OR2_X1 _8435_ (
    .A1(_1912_),
    .A2(_1913_),
    .ZN(_1914_)
  );
  AND2_X1 _8436_ (
    .A1(reg_pmp_0_addr[17]),
    .A2(_0837_),
    .ZN(_1915_)
  );
  AND2_X1 _8437_ (
    .A1(reg_pmp_2_addr[17]),
    .A2(_0792_),
    .ZN(_1916_)
  );
  OR2_X1 _8438_ (
    .A1(_1915_),
    .A2(_1916_),
    .ZN(_1917_)
  );
  OR2_X1 _8439_ (
    .A1(_1914_),
    .A2(_1917_),
    .ZN(_1918_)
  );
  AND2_X1 _8440_ (
    .A1(large_[43]),
    .A2(_0827_),
    .ZN(_1919_)
  );
  AND2_X1 _8441_ (
    .A1(large_1[43]),
    .A2(_0851_),
    .ZN(_1920_)
  );
  OR2_X1 _8442_ (
    .A1(_1919_),
    .A2(_1920_),
    .ZN(_1921_)
  );
  OR2_X1 _8443_ (
    .A1(_1918_),
    .A2(_1921_),
    .ZN(_1922_)
  );
  OR2_X1 _8444_ (
    .A1(_1911_),
    .A2(_1922_),
    .ZN(_1923_)
  );
  OR2_X1 _8445_ (
    .A1(_1904_),
    .A2(_1923_),
    .ZN(io_rw_rdata[17])
  );
  AND2_X1 _8446_ (
    .A1(io_rw_cmd[1]),
    .A2(_0694_),
    .ZN(_1924_)
  );
  AND2_X1 _8447_ (
    .A1(io_rw_rdata[17]),
    .A2(_1924_),
    .ZN(_1925_)
  );
  OR2_X1 _8448_ (
    .A1(_1881_),
    .A2(_1925_),
    .ZN(_1926_)
  );
  MUX2_X1 _8449_ (
    .A(_1926_),
    .B(reg_pmp_5_addr[17]),
    .S(_1181_),
    .Z(_0044_)
  );
  MUX2_X1 _8450_ (
    .A(_0908_),
    .B(reg_pmp_5_addr[18]),
    .S(_1181_),
    .Z(_0045_)
  );
  MUX2_X1 _8451_ (
    .A(_0967_),
    .B(reg_pmp_5_addr[19]),
    .S(_1181_),
    .Z(_0046_)
  );
  MUX2_X1 _8452_ (
    .A(_1017_),
    .B(reg_pmp_5_addr[20]),
    .S(_1181_),
    .Z(_0047_)
  );
  AND2_X1 _8453_ (
    .A1(io_rw_wdata[21]),
    .A2(_0742_),
    .ZN(_1927_)
  );
  AND2_X1 _8454_ (
    .A1(reg_dpc[21]),
    .A2(_0750_),
    .ZN(_1928_)
  );
  AND2_X1 _8455_ (
    .A1(reg_bp_0_address[21]),
    .A2(_0800_),
    .ZN(_1929_)
  );
  OR2_X1 _8456_ (
    .A1(_1928_),
    .A2(_1929_),
    .ZN(_1930_)
  );
  AND2_X1 _8457_ (
    .A1(reg_pmp_2_addr[21]),
    .A2(_0792_),
    .ZN(_1931_)
  );
  AND2_X1 _8458_ (
    .A1(reg_dscratch0[21]),
    .A2(_0797_),
    .ZN(_1932_)
  );
  OR2_X1 _8459_ (
    .A1(_1931_),
    .A2(_1932_),
    .ZN(_1933_)
  );
  OR2_X1 _8460_ (
    .A1(_1930_),
    .A2(_1933_),
    .ZN(_1934_)
  );
  AND2_X1 _8461_ (
    .A1(reg_pmp_5_addr[21]),
    .A2(_0788_),
    .ZN(_1935_)
  );
  AND2_X1 _8462_ (
    .A1(reg_pmp_1_addr[21]),
    .A2(_0841_),
    .ZN(_1936_)
  );
  OR2_X1 _8463_ (
    .A1(_1935_),
    .A2(_1936_),
    .ZN(_1937_)
  );
  AND2_X1 _8464_ (
    .A1(reg_mepc[21]),
    .A2(_0783_),
    .ZN(_1938_)
  );
  AND2_X1 _8465_ (
    .A1(reg_mtval[21]),
    .A2(_0764_),
    .ZN(_1939_)
  );
  OR2_X1 _8466_ (
    .A1(_1938_),
    .A2(_1939_),
    .ZN(_1940_)
  );
  OR2_X1 _8467_ (
    .A1(_1937_),
    .A2(_1940_),
    .ZN(_1941_)
  );
  AND2_X1 _8468_ (
    .A1(reg_pmp_4_addr[21]),
    .A2(_0805_),
    .ZN(_1942_)
  );
  AND2_X1 _8469_ (
    .A1(reg_mtvec[21]),
    .A2(_0780_),
    .ZN(_1943_)
  );
  OR2_X1 _8470_ (
    .A1(_1942_),
    .A2(_1943_),
    .ZN(_1944_)
  );
  AND2_X1 _8471_ (
    .A1(reg_pmp_0_addr[21]),
    .A2(_0837_),
    .ZN(_1945_)
  );
  AND2_X1 _8472_ (
    .A1(reg_mcause[21]),
    .A2(_0834_),
    .ZN(_1946_)
  );
  OR2_X1 _8473_ (
    .A1(_1945_),
    .A2(_1946_),
    .ZN(_1947_)
  );
  OR2_X1 _8474_ (
    .A1(_1944_),
    .A2(_1947_),
    .ZN(_1948_)
  );
  OR2_X1 _8475_ (
    .A1(_1941_),
    .A2(_1948_),
    .ZN(_1949_)
  );
  OR2_X1 _8476_ (
    .A1(_1934_),
    .A2(_1949_),
    .ZN(_1950_)
  );
  AND2_X1 _8477_ (
    .A1(large_1[47]),
    .A2(_0851_),
    .ZN(_1951_)
  );
  AND2_X1 _8478_ (
    .A1(reg_pmp_7_addr[21]),
    .A2(_0849_),
    .ZN(_1952_)
  );
  AND2_X1 _8479_ (
    .A1(large_[47]),
    .A2(_0827_),
    .ZN(_1953_)
  );
  OR2_X1 _8480_ (
    .A1(_1952_),
    .A2(_1953_),
    .ZN(_1954_)
  );
  OR2_X1 _8481_ (
    .A1(_1951_),
    .A2(_1954_),
    .ZN(_1955_)
  );
  AND2_X1 _8482_ (
    .A1(large_[15]),
    .A2(_0822_),
    .ZN(_1956_)
  );
  AND2_X1 _8483_ (
    .A1(reg_mscratch[21]),
    .A2(_0767_),
    .ZN(_1957_)
  );
  AND2_X1 _8484_ (
    .A1(reg_pmp_3_addr[21]),
    .A2(_0844_),
    .ZN(_1958_)
  );
  OR2_X1 _8485_ (
    .A1(_1957_),
    .A2(_1958_),
    .ZN(_1959_)
  );
  OR2_X1 _8486_ (
    .A1(_1956_),
    .A2(_1959_),
    .ZN(_1960_)
  );
  AND2_X1 _8487_ (
    .A1(reg_pmp_6_addr[21]),
    .A2(_0814_),
    .ZN(_1961_)
  );
  AND2_X1 _8488_ (
    .A1(large_1[15]),
    .A2(_0830_),
    .ZN(_1962_)
  );
  OR2_X1 _8489_ (
    .A1(_1961_),
    .A2(_1962_),
    .ZN(_1963_)
  );
  OR2_X1 _8490_ (
    .A1(_1960_),
    .A2(_1963_),
    .ZN(_1964_)
  );
  OR2_X1 _8491_ (
    .A1(_1955_),
    .A2(_1964_),
    .ZN(_1965_)
  );
  OR2_X1 _8492_ (
    .A1(_1950_),
    .A2(_1965_),
    .ZN(io_rw_rdata[21])
  );
  AND2_X1 _8493_ (
    .A1(io_rw_cmd[1]),
    .A2(_0698_),
    .ZN(_1966_)
  );
  AND2_X1 _8494_ (
    .A1(io_rw_rdata[21]),
    .A2(_1966_),
    .ZN(_1967_)
  );
  OR2_X1 _8495_ (
    .A1(_1927_),
    .A2(_1967_),
    .ZN(_1968_)
  );
  MUX2_X1 _8496_ (
    .A(_1968_),
    .B(reg_pmp_5_addr[21]),
    .S(_1181_),
    .Z(_0048_)
  );
  AND2_X1 _8497_ (
    .A1(io_rw_wdata[22]),
    .A2(_0742_),
    .ZN(_1969_)
  );
  AND2_X1 _8498_ (
    .A1(reg_pmp_1_addr[22]),
    .A2(_0841_),
    .ZN(_1970_)
  );
  AND2_X1 _8499_ (
    .A1(reg_pmp_5_addr[22]),
    .A2(_0788_),
    .ZN(_1971_)
  );
  AND2_X1 _8500_ (
    .A1(reg_pmp_2_addr[22]),
    .A2(_0792_),
    .ZN(_1972_)
  );
  AND2_X1 _8501_ (
    .A1(reg_dscratch0[22]),
    .A2(_0797_),
    .ZN(_1973_)
  );
  AND2_X1 _8502_ (
    .A1(reg_mtvec[22]),
    .A2(_0780_),
    .ZN(_1974_)
  );
  AND2_X1 _8503_ (
    .A1(reg_pmp_4_addr[22]),
    .A2(_0805_),
    .ZN(_1975_)
  );
  OR2_X1 _8504_ (
    .A1(_1974_),
    .A2(_1975_),
    .ZN(_1976_)
  );
  AND2_X1 _8505_ (
    .A1(reg_mscratch[22]),
    .A2(_0767_),
    .ZN(_1977_)
  );
  AND2_X1 _8506_ (
    .A1(reg_bp_0_address[22]),
    .A2(_0800_),
    .ZN(_1978_)
  );
  AND2_X1 _8507_ (
    .A1(reg_pmp_3_addr[22]),
    .A2(_0844_),
    .ZN(_1979_)
  );
  AND2_X1 _8508_ (
    .A1(reg_dpc[22]),
    .A2(_0750_),
    .ZN(_1980_)
  );
  AND2_X1 _8509_ (
    .A1(reg_pmp_0_addr[22]),
    .A2(_0837_),
    .ZN(_1981_)
  );
  AND2_X1 _8510_ (
    .A1(reg_mepc[22]),
    .A2(_0783_),
    .ZN(_1982_)
  );
  AND2_X1 _8511_ (
    .A1(reg_pmp_7_addr[22]),
    .A2(_0849_),
    .ZN(_1983_)
  );
  AND2_X1 _8512_ (
    .A1(reg_pmp_6_addr[22]),
    .A2(_0814_),
    .ZN(_1984_)
  );
  AND2_X1 _8513_ (
    .A1(large_[48]),
    .A2(_0827_),
    .ZN(_1985_)
  );
  AND2_X1 _8514_ (
    .A1(large_1[48]),
    .A2(_0851_),
    .ZN(_1986_)
  );
  AND2_X1 _8515_ (
    .A1(reg_mtval[22]),
    .A2(_0764_),
    .ZN(_1987_)
  );
  AND2_X1 _8516_ (
    .A1(reg_mcause[22]),
    .A2(_0834_),
    .ZN(_1988_)
  );
  OR2_X1 _8517_ (
    .A1(_1977_),
    .A2(_1987_),
    .ZN(_1989_)
  );
  OR2_X1 _8518_ (
    .A1(_1988_),
    .A2(_1989_),
    .ZN(_1990_)
  );
  OR2_X1 _8519_ (
    .A1(_1970_),
    .A2(_1981_),
    .ZN(_1991_)
  );
  AND2_X1 _8520_ (
    .A1(large_[16]),
    .A2(_0857_),
    .ZN(_1992_)
  );
  AND2_X1 _8521_ (
    .A1(large_1[16]),
    .A2(_0859_),
    .ZN(_1993_)
  );
  OR2_X1 _8522_ (
    .A1(_1972_),
    .A2(_1984_),
    .ZN(_1994_)
  );
  OR2_X1 _8523_ (
    .A1(_1990_),
    .A2(_1994_),
    .ZN(_1995_)
  );
  OR2_X1 _8524_ (
    .A1(_1979_),
    .A2(_1991_),
    .ZN(_1996_)
  );
  OR2_X1 _8525_ (
    .A1(_1985_),
    .A2(_1986_),
    .ZN(_1997_)
  );
  OR2_X1 _8526_ (
    .A1(_1996_),
    .A2(_1997_),
    .ZN(_1998_)
  );
  OR2_X1 _8527_ (
    .A1(_1995_),
    .A2(_1998_),
    .ZN(_1999_)
  );
  OR2_X1 _8528_ (
    .A1(_1976_),
    .A2(_1983_),
    .ZN(_2000_)
  );
  OR2_X1 _8529_ (
    .A1(_1978_),
    .A2(_1982_),
    .ZN(_2001_)
  );
  OR2_X1 _8530_ (
    .A1(_2000_),
    .A2(_2001_),
    .ZN(_2002_)
  );
  OR2_X1 _8531_ (
    .A1(_1971_),
    .A2(_1973_),
    .ZN(_2003_)
  );
  OR2_X1 _8532_ (
    .A1(_1980_),
    .A2(_1992_),
    .ZN(_2004_)
  );
  OR2_X1 _8533_ (
    .A1(_1993_),
    .A2(_2004_),
    .ZN(_2005_)
  );
  OR2_X1 _8534_ (
    .A1(_2003_),
    .A2(_2005_),
    .ZN(_2006_)
  );
  OR2_X1 _8535_ (
    .A1(_2002_),
    .A2(_2006_),
    .ZN(_2007_)
  );
  OR2_X1 _8536_ (
    .A1(_1999_),
    .A2(_2007_),
    .ZN(io_rw_rdata[22])
  );
  AND2_X1 _8537_ (
    .A1(io_rw_cmd[1]),
    .A2(_0699_),
    .ZN(_2008_)
  );
  AND2_X1 _8538_ (
    .A1(io_rw_rdata[22]),
    .A2(_2008_),
    .ZN(_2009_)
  );
  OR2_X1 _8539_ (
    .A1(_1969_),
    .A2(_2009_),
    .ZN(_2010_)
  );
  MUX2_X1 _8540_ (
    .A(_2010_),
    .B(reg_pmp_5_addr[22]),
    .S(_1181_),
    .Z(_0049_)
  );
  MUX2_X1 _8541_ (
    .A(_1071_),
    .B(reg_pmp_5_addr[23]),
    .S(_1181_),
    .Z(_0050_)
  );
  AND2_X1 _8542_ (
    .A1(io_rw_wdata[24]),
    .A2(_0742_),
    .ZN(_2011_)
  );
  AND2_X1 _8543_ (
    .A1(reg_mcause[24]),
    .A2(_0834_),
    .ZN(_2012_)
  );
  AND2_X1 _8544_ (
    .A1(reg_pmp_1_addr[24]),
    .A2(_0841_),
    .ZN(_2013_)
  );
  OR2_X1 _8545_ (
    .A1(_2012_),
    .A2(_2013_),
    .ZN(_2014_)
  );
  AND2_X1 _8546_ (
    .A1(reg_mtvec[24]),
    .A2(_0780_),
    .ZN(_2015_)
  );
  AND2_X1 _8547_ (
    .A1(reg_mscratch[24]),
    .A2(_0767_),
    .ZN(_2016_)
  );
  OR2_X1 _8548_ (
    .A1(_2015_),
    .A2(_2016_),
    .ZN(_2017_)
  );
  OR2_X1 _8549_ (
    .A1(_2014_),
    .A2(_2017_),
    .ZN(_2018_)
  );
  AND2_X1 _8550_ (
    .A1(reg_mtval[24]),
    .A2(_0764_),
    .ZN(_2019_)
  );
  AND2_X1 _8551_ (
    .A1(reg_pmp_0_addr[24]),
    .A2(_0837_),
    .ZN(_2020_)
  );
  OR2_X1 _8552_ (
    .A1(_2019_),
    .A2(_2020_),
    .ZN(_2021_)
  );
  AND2_X1 _8553_ (
    .A1(reg_pmp_2_addr[24]),
    .A2(_0792_),
    .ZN(_2022_)
  );
  AND2_X1 _8554_ (
    .A1(reg_dscratch0[24]),
    .A2(_0797_),
    .ZN(_2023_)
  );
  OR2_X1 _8555_ (
    .A1(_2022_),
    .A2(_2023_),
    .ZN(_2024_)
  );
  OR2_X1 _8556_ (
    .A1(_2021_),
    .A2(_2024_),
    .ZN(_2025_)
  );
  AND2_X1 _8557_ (
    .A1(reg_mepc[24]),
    .A2(_0783_),
    .ZN(_2026_)
  );
  AND2_X1 _8558_ (
    .A1(reg_pmp_4_addr[24]),
    .A2(_0805_),
    .ZN(_2027_)
  );
  OR2_X1 _8559_ (
    .A1(_2026_),
    .A2(_2027_),
    .ZN(_2028_)
  );
  AND2_X1 _8560_ (
    .A1(reg_pmp_5_addr[24]),
    .A2(_0788_),
    .ZN(_2029_)
  );
  AND2_X1 _8561_ (
    .A1(reg_dpc[24]),
    .A2(_0750_),
    .ZN(_2030_)
  );
  OR2_X1 _8562_ (
    .A1(_2029_),
    .A2(_2030_),
    .ZN(_2031_)
  );
  OR2_X1 _8563_ (
    .A1(_2028_),
    .A2(_2031_),
    .ZN(_2032_)
  );
  OR2_X1 _8564_ (
    .A1(_2025_),
    .A2(_2032_),
    .ZN(_2033_)
  );
  OR2_X1 _8565_ (
    .A1(_2018_),
    .A2(_2033_),
    .ZN(_2034_)
  );
  AND2_X1 _8566_ (
    .A1(large_[18]),
    .A2(_0822_),
    .ZN(_2035_)
  );
  AND2_X1 _8567_ (
    .A1(large_1[18]),
    .A2(_0830_),
    .ZN(_2036_)
  );
  OR2_X1 _8568_ (
    .A1(_2035_),
    .A2(_2036_),
    .ZN(_2037_)
  );
  AND2_X1 _8569_ (
    .A1(reg_pmp_6_addr[24]),
    .A2(_0814_),
    .ZN(_2038_)
  );
  AND2_X1 _8570_ (
    .A1(reg_pmp_7_addr[24]),
    .A2(_0849_),
    .ZN(_2039_)
  );
  OR2_X1 _8571_ (
    .A1(_2038_),
    .A2(_2039_),
    .ZN(_2040_)
  );
  OR2_X1 _8572_ (
    .A1(_2037_),
    .A2(_2040_),
    .ZN(_2041_)
  );
  AND2_X1 _8573_ (
    .A1(large_1[50]),
    .A2(_0851_),
    .ZN(_2042_)
  );
  AND2_X1 _8574_ (
    .A1(large_[50]),
    .A2(_0827_),
    .ZN(_2043_)
  );
  OR2_X1 _8575_ (
    .A1(_2042_),
    .A2(_2043_),
    .ZN(_2044_)
  );
  AND2_X1 _8576_ (
    .A1(reg_pmp_3_cfg_r),
    .A2(_0754_),
    .ZN(_2045_)
  );
  AND2_X1 _8577_ (
    .A1(reg_bp_0_address[24]),
    .A2(_0800_),
    .ZN(_2046_)
  );
  OR2_X1 _8578_ (
    .A1(_2045_),
    .A2(_2046_),
    .ZN(_2047_)
  );
  AND2_X1 _8579_ (
    .A1(reg_pmp_7_cfg_r),
    .A2(_0733_),
    .ZN(_2048_)
  );
  AND2_X1 _8580_ (
    .A1(reg_pmp_3_addr[24]),
    .A2(_0844_),
    .ZN(_2049_)
  );
  OR2_X1 _8581_ (
    .A1(_2048_),
    .A2(_2049_),
    .ZN(_2050_)
  );
  OR2_X1 _8582_ (
    .A1(_2047_),
    .A2(_2050_),
    .ZN(_2051_)
  );
  OR2_X1 _8583_ (
    .A1(_2044_),
    .A2(_2051_),
    .ZN(_2052_)
  );
  OR2_X1 _8584_ (
    .A1(_2041_),
    .A2(_2052_),
    .ZN(_2053_)
  );
  OR2_X1 _8585_ (
    .A1(_2034_),
    .A2(_2053_),
    .ZN(io_rw_rdata[24])
  );
  AND2_X1 _8586_ (
    .A1(io_rw_cmd[1]),
    .A2(_0701_),
    .ZN(_2054_)
  );
  AND2_X1 _8587_ (
    .A1(io_rw_rdata[24]),
    .A2(_2054_),
    .ZN(_2055_)
  );
  OR2_X1 _8588_ (
    .A1(_2011_),
    .A2(_2055_),
    .ZN(_2056_)
  );
  MUX2_X1 _8589_ (
    .A(_2056_),
    .B(reg_pmp_5_addr[24]),
    .S(_1181_),
    .Z(_0051_)
  );
  AND2_X1 _8590_ (
    .A1(io_rw_wdata[25]),
    .A2(_0742_),
    .ZN(_2057_)
  );
  AND2_X1 _8591_ (
    .A1(reg_pmp_7_cfg_w),
    .A2(_0733_),
    .ZN(_2058_)
  );
  AND2_X1 _8592_ (
    .A1(reg_pmp_4_addr[25]),
    .A2(_0805_),
    .ZN(_2059_)
  );
  OR2_X1 _8593_ (
    .A1(_2058_),
    .A2(_2059_),
    .ZN(_2060_)
  );
  AND2_X1 _8594_ (
    .A1(reg_mtvec[25]),
    .A2(_0780_),
    .ZN(_2061_)
  );
  AND2_X1 _8595_ (
    .A1(reg_pmp_5_addr[25]),
    .A2(_0788_),
    .ZN(_2062_)
  );
  OR2_X1 _8596_ (
    .A1(_2061_),
    .A2(_2062_),
    .ZN(_2063_)
  );
  OR2_X1 _8597_ (
    .A1(_2060_),
    .A2(_2063_),
    .ZN(_2064_)
  );
  AND2_X1 _8598_ (
    .A1(reg_mepc[25]),
    .A2(_0783_),
    .ZN(_2065_)
  );
  AND2_X1 _8599_ (
    .A1(reg_pmp_3_addr[25]),
    .A2(_0844_),
    .ZN(_2066_)
  );
  OR2_X1 _8600_ (
    .A1(_2065_),
    .A2(_2066_),
    .ZN(_2067_)
  );
  AND2_X1 _8601_ (
    .A1(reg_mtval[25]),
    .A2(_0764_),
    .ZN(_2068_)
  );
  AND2_X1 _8602_ (
    .A1(reg_pmp_0_addr[25]),
    .A2(_0837_),
    .ZN(_2069_)
  );
  OR2_X1 _8603_ (
    .A1(_2068_),
    .A2(_2069_),
    .ZN(_2070_)
  );
  OR2_X1 _8604_ (
    .A1(_2067_),
    .A2(_2070_),
    .ZN(_2071_)
  );
  AND2_X1 _8605_ (
    .A1(reg_dscratch0[25]),
    .A2(_0797_),
    .ZN(_2072_)
  );
  AND2_X1 _8606_ (
    .A1(reg_pmp_1_addr[25]),
    .A2(_0841_),
    .ZN(_2073_)
  );
  OR2_X1 _8607_ (
    .A1(_2072_),
    .A2(_2073_),
    .ZN(_2074_)
  );
  AND2_X1 _8608_ (
    .A1(reg_mcause[25]),
    .A2(_0834_),
    .ZN(_2075_)
  );
  AND2_X1 _8609_ (
    .A1(reg_bp_0_address[25]),
    .A2(_0800_),
    .ZN(_2076_)
  );
  OR2_X1 _8610_ (
    .A1(_2075_),
    .A2(_2076_),
    .ZN(_2077_)
  );
  OR2_X1 _8611_ (
    .A1(_2074_),
    .A2(_2077_),
    .ZN(_2078_)
  );
  OR2_X1 _8612_ (
    .A1(_2071_),
    .A2(_2078_),
    .ZN(_2079_)
  );
  OR2_X1 _8613_ (
    .A1(_2064_),
    .A2(_2079_),
    .ZN(_2080_)
  );
  AND2_X1 _8614_ (
    .A1(reg_pmp_6_addr[25]),
    .A2(_0814_),
    .ZN(_2081_)
  );
  AND2_X1 _8615_ (
    .A1(large_[19]),
    .A2(_0822_),
    .ZN(_2082_)
  );
  OR2_X1 _8616_ (
    .A1(_2081_),
    .A2(_2082_),
    .ZN(_2083_)
  );
  AND2_X1 _8617_ (
    .A1(reg_pmp_7_addr[25]),
    .A2(_0849_),
    .ZN(_2084_)
  );
  AND2_X1 _8618_ (
    .A1(large_1[51]),
    .A2(_0851_),
    .ZN(_2085_)
  );
  OR2_X1 _8619_ (
    .A1(_2084_),
    .A2(_2085_),
    .ZN(_2086_)
  );
  OR2_X1 _8620_ (
    .A1(_2083_),
    .A2(_2086_),
    .ZN(_2087_)
  );
  AND2_X1 _8621_ (
    .A1(reg_mscratch[25]),
    .A2(_0767_),
    .ZN(_2088_)
  );
  AND2_X1 _8622_ (
    .A1(reg_pmp_2_addr[25]),
    .A2(_0792_),
    .ZN(_2089_)
  );
  OR2_X1 _8623_ (
    .A1(_2088_),
    .A2(_2089_),
    .ZN(_2090_)
  );
  AND2_X1 _8624_ (
    .A1(reg_dpc[25]),
    .A2(_0750_),
    .ZN(_2091_)
  );
  AND2_X1 _8625_ (
    .A1(reg_pmp_3_cfg_w),
    .A2(_0754_),
    .ZN(_2092_)
  );
  OR2_X1 _8626_ (
    .A1(_2091_),
    .A2(_2092_),
    .ZN(_2093_)
  );
  OR2_X1 _8627_ (
    .A1(_2090_),
    .A2(_2093_),
    .ZN(_2094_)
  );
  AND2_X1 _8628_ (
    .A1(large_[51]),
    .A2(_0827_),
    .ZN(_2095_)
  );
  AND2_X1 _8629_ (
    .A1(large_1[19]),
    .A2(_0830_),
    .ZN(_2096_)
  );
  OR2_X1 _8630_ (
    .A1(_2095_),
    .A2(_2096_),
    .ZN(_2097_)
  );
  OR2_X1 _8631_ (
    .A1(_2094_),
    .A2(_2097_),
    .ZN(_2098_)
  );
  OR2_X1 _8632_ (
    .A1(_2087_),
    .A2(_2098_),
    .ZN(_2099_)
  );
  OR2_X1 _8633_ (
    .A1(_2080_),
    .A2(_2099_),
    .ZN(io_rw_rdata[25])
  );
  AND2_X1 _8634_ (
    .A1(io_rw_cmd[1]),
    .A2(_0702_),
    .ZN(_2100_)
  );
  AND2_X1 _8635_ (
    .A1(io_rw_rdata[25]),
    .A2(_2100_),
    .ZN(_2101_)
  );
  OR2_X1 _8636_ (
    .A1(_2057_),
    .A2(_2101_),
    .ZN(_2102_)
  );
  MUX2_X1 _8637_ (
    .A(_2102_),
    .B(reg_pmp_5_addr[25]),
    .S(_1181_),
    .Z(_0052_)
  );
  AND2_X1 _8638_ (
    .A1(io_rw_wdata[26]),
    .A2(_0742_),
    .ZN(_2103_)
  );
  AND2_X1 _8639_ (
    .A1(reg_pmp_3_addr[26]),
    .A2(_0844_),
    .ZN(_2104_)
  );
  AND2_X1 _8640_ (
    .A1(reg_mtval[26]),
    .A2(_0764_),
    .ZN(_2105_)
  );
  OR2_X1 _8641_ (
    .A1(_2104_),
    .A2(_2105_),
    .ZN(_2106_)
  );
  AND2_X1 _8642_ (
    .A1(reg_pmp_1_addr[26]),
    .A2(_0841_),
    .ZN(_2107_)
  );
  AND2_X1 _8643_ (
    .A1(reg_pmp_7_cfg_x),
    .A2(_0733_),
    .ZN(_2108_)
  );
  OR2_X1 _8644_ (
    .A1(_2107_),
    .A2(_2108_),
    .ZN(_2109_)
  );
  OR2_X1 _8645_ (
    .A1(_2106_),
    .A2(_2109_),
    .ZN(_2110_)
  );
  AND2_X1 _8646_ (
    .A1(reg_mscratch[26]),
    .A2(_0767_),
    .ZN(_2111_)
  );
  AND2_X1 _8647_ (
    .A1(reg_pmp_2_addr[26]),
    .A2(_0792_),
    .ZN(_2112_)
  );
  OR2_X1 _8648_ (
    .A1(_2111_),
    .A2(_2112_),
    .ZN(_2113_)
  );
  AND2_X1 _8649_ (
    .A1(reg_pmp_3_cfg_x),
    .A2(_0754_),
    .ZN(_2114_)
  );
  AND2_X1 _8650_ (
    .A1(reg_mtvec[26]),
    .A2(_0780_),
    .ZN(_2115_)
  );
  OR2_X1 _8651_ (
    .A1(_2114_),
    .A2(_2115_),
    .ZN(_2116_)
  );
  OR2_X1 _8652_ (
    .A1(_2113_),
    .A2(_2116_),
    .ZN(_2117_)
  );
  AND2_X1 _8653_ (
    .A1(reg_pmp_4_addr[26]),
    .A2(_0805_),
    .ZN(_2118_)
  );
  AND2_X1 _8654_ (
    .A1(reg_pmp_0_addr[26]),
    .A2(_0837_),
    .ZN(_2119_)
  );
  OR2_X1 _8655_ (
    .A1(_2118_),
    .A2(_2119_),
    .ZN(_2120_)
  );
  AND2_X1 _8656_ (
    .A1(reg_bp_0_address[26]),
    .A2(_0800_),
    .ZN(_2121_)
  );
  AND2_X1 _8657_ (
    .A1(reg_mepc[26]),
    .A2(_0783_),
    .ZN(_2122_)
  );
  OR2_X1 _8658_ (
    .A1(_2121_),
    .A2(_2122_),
    .ZN(_2123_)
  );
  OR2_X1 _8659_ (
    .A1(_2120_),
    .A2(_2123_),
    .ZN(_2124_)
  );
  OR2_X1 _8660_ (
    .A1(_2117_),
    .A2(_2124_),
    .ZN(_2125_)
  );
  OR2_X1 _8661_ (
    .A1(_2110_),
    .A2(_2125_),
    .ZN(_2126_)
  );
  AND2_X1 _8662_ (
    .A1(large_1[52]),
    .A2(_0851_),
    .ZN(_2127_)
  );
  AND2_X1 _8663_ (
    .A1(large_1[20]),
    .A2(_0830_),
    .ZN(_2128_)
  );
  OR2_X1 _8664_ (
    .A1(_2127_),
    .A2(_2128_),
    .ZN(_2129_)
  );
  AND2_X1 _8665_ (
    .A1(large_[52]),
    .A2(_0827_),
    .ZN(_2130_)
  );
  AND2_X1 _8666_ (
    .A1(large_[20]),
    .A2(_0822_),
    .ZN(_2131_)
  );
  OR2_X1 _8667_ (
    .A1(_2130_),
    .A2(_2131_),
    .ZN(_2132_)
  );
  OR2_X1 _8668_ (
    .A1(_2129_),
    .A2(_2132_),
    .ZN(_2133_)
  );
  AND2_X1 _8669_ (
    .A1(reg_mcause[26]),
    .A2(_0834_),
    .ZN(_2134_)
  );
  AND2_X1 _8670_ (
    .A1(reg_dscratch0[26]),
    .A2(_0797_),
    .ZN(_2135_)
  );
  OR2_X1 _8671_ (
    .A1(_2134_),
    .A2(_2135_),
    .ZN(_2136_)
  );
  AND2_X1 _8672_ (
    .A1(reg_pmp_5_addr[26]),
    .A2(_0788_),
    .ZN(_2137_)
  );
  AND2_X1 _8673_ (
    .A1(reg_dpc[26]),
    .A2(_0750_),
    .ZN(_2138_)
  );
  OR2_X1 _8674_ (
    .A1(_2137_),
    .A2(_2138_),
    .ZN(_2139_)
  );
  OR2_X1 _8675_ (
    .A1(_2136_),
    .A2(_2139_),
    .ZN(_2140_)
  );
  AND2_X1 _8676_ (
    .A1(reg_pmp_6_addr[26]),
    .A2(_0814_),
    .ZN(_2141_)
  );
  AND2_X1 _8677_ (
    .A1(reg_pmp_7_addr[26]),
    .A2(_0849_),
    .ZN(_2142_)
  );
  OR2_X1 _8678_ (
    .A1(_2141_),
    .A2(_2142_),
    .ZN(_2143_)
  );
  OR2_X1 _8679_ (
    .A1(_2140_),
    .A2(_2143_),
    .ZN(_2144_)
  );
  OR2_X1 _8680_ (
    .A1(_2133_),
    .A2(_2144_),
    .ZN(_2145_)
  );
  OR2_X1 _8681_ (
    .A1(_2126_),
    .A2(_2145_),
    .ZN(io_rw_rdata[26])
  );
  AND2_X1 _8682_ (
    .A1(io_rw_cmd[1]),
    .A2(_0703_),
    .ZN(_2146_)
  );
  AND2_X1 _8683_ (
    .A1(io_rw_rdata[26]),
    .A2(_2146_),
    .ZN(_2147_)
  );
  OR2_X1 _8684_ (
    .A1(_2103_),
    .A2(_2147_),
    .ZN(_2148_)
  );
  MUX2_X1 _8685_ (
    .A(_2148_),
    .B(reg_pmp_5_addr[26]),
    .S(_1181_),
    .Z(_0053_)
  );
  AND2_X1 _8686_ (
    .A1(reg_bp_0_control_dmode),
    .A2(_1058_),
    .ZN(_2149_)
  );
  AND2_X1 _8687_ (
    .A1(reg_bp_0_address[27]),
    .A2(_0800_),
    .ZN(_2150_)
  );
  OR2_X1 _8688_ (
    .A1(_2149_),
    .A2(_2150_),
    .ZN(_2151_)
  );
  AND2_X1 _8689_ (
    .A1(reg_pmp_3_cfg_a[0]),
    .A2(_0754_),
    .ZN(_2152_)
  );
  AND2_X1 _8690_ (
    .A1(reg_mtval[27]),
    .A2(_0764_),
    .ZN(_2153_)
  );
  OR2_X1 _8691_ (
    .A1(_2152_),
    .A2(_2153_),
    .ZN(_2154_)
  );
  OR2_X1 _8692_ (
    .A1(_2151_),
    .A2(_2154_),
    .ZN(_2155_)
  );
  AND2_X1 _8693_ (
    .A1(reg_dpc[27]),
    .A2(_0750_),
    .ZN(_2156_)
  );
  AND2_X1 _8694_ (
    .A1(reg_pmp_4_addr[27]),
    .A2(_0805_),
    .ZN(_2157_)
  );
  OR2_X1 _8695_ (
    .A1(_2156_),
    .A2(_2157_),
    .ZN(_2158_)
  );
  AND2_X1 _8696_ (
    .A1(reg_pmp_5_addr[27]),
    .A2(_0788_),
    .ZN(_2159_)
  );
  AND2_X1 _8697_ (
    .A1(reg_pmp_0_addr[27]),
    .A2(_0837_),
    .ZN(_2160_)
  );
  OR2_X1 _8698_ (
    .A1(_2159_),
    .A2(_2160_),
    .ZN(_2161_)
  );
  OR2_X1 _8699_ (
    .A1(_2158_),
    .A2(_2161_),
    .ZN(_2162_)
  );
  OR2_X1 _8700_ (
    .A1(_2155_),
    .A2(_2162_),
    .ZN(_2163_)
  );
  AND2_X1 _8701_ (
    .A1(reg_pmp_3_addr[27]),
    .A2(_0844_),
    .ZN(_2164_)
  );
  AND2_X1 _8702_ (
    .A1(reg_pmp_1_addr[27]),
    .A2(_0841_),
    .ZN(_2165_)
  );
  AND2_X1 _8703_ (
    .A1(reg_mepc[27]),
    .A2(_0783_),
    .ZN(_2166_)
  );
  OR2_X1 _8704_ (
    .A1(_2165_),
    .A2(_2166_),
    .ZN(_2167_)
  );
  OR2_X1 _8705_ (
    .A1(_2164_),
    .A2(_2167_),
    .ZN(_2168_)
  );
  AND2_X1 _8706_ (
    .A1(reg_mtvec[27]),
    .A2(_0780_),
    .ZN(_2169_)
  );
  AND2_X1 _8707_ (
    .A1(reg_mscratch[27]),
    .A2(_0767_),
    .ZN(_2170_)
  );
  OR2_X1 _8708_ (
    .A1(_2169_),
    .A2(_2170_),
    .ZN(_2171_)
  );
  AND2_X1 _8709_ (
    .A1(reg_pmp_2_addr[27]),
    .A2(_0792_),
    .ZN(_2172_)
  );
  AND2_X1 _8710_ (
    .A1(reg_mcause[27]),
    .A2(_0834_),
    .ZN(_2173_)
  );
  OR2_X1 _8711_ (
    .A1(_2172_),
    .A2(_2173_),
    .ZN(_2174_)
  );
  OR2_X1 _8712_ (
    .A1(_2171_),
    .A2(_2174_),
    .ZN(_2175_)
  );
  OR2_X1 _8713_ (
    .A1(_2168_),
    .A2(_2175_),
    .ZN(_2176_)
  );
  OR2_X1 _8714_ (
    .A1(_2163_),
    .A2(_2176_),
    .ZN(_2177_)
  );
  AND2_X1 _8715_ (
    .A1(large_1[21]),
    .A2(_0830_),
    .ZN(_2178_)
  );
  AND2_X1 _8716_ (
    .A1(large_[53]),
    .A2(_0827_),
    .ZN(_2179_)
  );
  AND2_X1 _8717_ (
    .A1(large_1[53]),
    .A2(_0851_),
    .ZN(_2180_)
  );
  OR2_X1 _8718_ (
    .A1(_2179_),
    .A2(_2180_),
    .ZN(_2181_)
  );
  OR2_X1 _8719_ (
    .A1(_2178_),
    .A2(_2181_),
    .ZN(_2182_)
  );
  AND2_X1 _8720_ (
    .A1(large_[21]),
    .A2(_0822_),
    .ZN(_2183_)
  );
  AND2_X1 _8721_ (
    .A1(reg_dscratch0[27]),
    .A2(_0797_),
    .ZN(_2184_)
  );
  AND2_X1 _8722_ (
    .A1(reg_pmp_7_cfg_a[0]),
    .A2(_0733_),
    .ZN(_2185_)
  );
  OR2_X1 _8723_ (
    .A1(_2184_),
    .A2(_2185_),
    .ZN(_2186_)
  );
  OR2_X1 _8724_ (
    .A1(_2183_),
    .A2(_2186_),
    .ZN(_2187_)
  );
  AND2_X1 _8725_ (
    .A1(reg_pmp_7_addr[27]),
    .A2(_0849_),
    .ZN(_2188_)
  );
  AND2_X1 _8726_ (
    .A1(reg_pmp_6_addr[27]),
    .A2(_0814_),
    .ZN(_2189_)
  );
  OR2_X1 _8727_ (
    .A1(_2188_),
    .A2(_2189_),
    .ZN(_2190_)
  );
  OR2_X1 _8728_ (
    .A1(_2187_),
    .A2(_2190_),
    .ZN(_2191_)
  );
  OR2_X1 _8729_ (
    .A1(_2182_),
    .A2(_2191_),
    .ZN(_2192_)
  );
  OR2_X1 _8730_ (
    .A1(_2177_),
    .A2(_2192_),
    .ZN(io_rw_rdata[27])
  );
  AND2_X1 _8731_ (
    .A1(io_rw_cmd[1]),
    .A2(io_rw_rdata[27]),
    .ZN(_2193_)
  );
  OR2_X1 _8732_ (
    .A1(_0704_),
    .A2(_0742_),
    .ZN(_2194_)
  );
  MUX2_X1 _8733_ (
    .A(_0742_),
    .B(_2193_),
    .S(_0704_),
    .Z(_2195_)
  );
  MUX2_X1 _8734_ (
    .A(_2195_),
    .B(reg_pmp_5_addr[27]),
    .S(_1181_),
    .Z(_0054_)
  );
  AND2_X1 _8735_ (
    .A1(io_rw_wdata[28]),
    .A2(_0742_),
    .ZN(_2196_)
  );
  AND2_X1 _8736_ (
    .A1(reg_dscratch0[28]),
    .A2(_0797_),
    .ZN(_2197_)
  );
  AND2_X1 _8737_ (
    .A1(reg_mtval[28]),
    .A2(_0764_),
    .ZN(_2198_)
  );
  AND2_X1 _8738_ (
    .A1(reg_mtvec[28]),
    .A2(_0780_),
    .ZN(_2199_)
  );
  AND2_X1 _8739_ (
    .A1(reg_pmp_2_addr[28]),
    .A2(_0792_),
    .ZN(_2200_)
  );
  AND2_X1 _8740_ (
    .A1(reg_pmp_7_cfg_a[1]),
    .A2(_0733_),
    .ZN(_2201_)
  );
  AND2_X1 _8741_ (
    .A1(reg_pmp_3_addr[28]),
    .A2(_0844_),
    .ZN(_2202_)
  );
  AND2_X1 _8742_ (
    .A1(reg_dpc[28]),
    .A2(_0750_),
    .ZN(_2203_)
  );
  AND2_X1 _8743_ (
    .A1(reg_pmp_3_cfg_a[1]),
    .A2(_0754_),
    .ZN(_2204_)
  );
  AND2_X1 _8744_ (
    .A1(reg_mepc[28]),
    .A2(_0783_),
    .ZN(_2205_)
  );
  AND2_X1 _8745_ (
    .A1(reg_mscratch[28]),
    .A2(_0767_),
    .ZN(_2206_)
  );
  OR2_X1 _8746_ (
    .A1(_2205_),
    .A2(_2206_),
    .ZN(_2207_)
  );
  AND2_X1 _8747_ (
    .A1(reg_pmp_4_addr[28]),
    .A2(_0805_),
    .ZN(_2208_)
  );
  AND2_X1 _8748_ (
    .A1(reg_bp_0_address[28]),
    .A2(_0800_),
    .ZN(_2209_)
  );
  AND2_X1 _8749_ (
    .A1(large_1[54]),
    .A2(_0851_),
    .ZN(_2210_)
  );
  AND2_X1 _8750_ (
    .A1(large_[54]),
    .A2(_0827_),
    .ZN(_2211_)
  );
  AND2_X1 _8751_ (
    .A1(reg_pmp_5_addr[28]),
    .A2(_0788_),
    .ZN(_2212_)
  );
  AND2_X1 _8752_ (
    .A1(reg_mcause[28]),
    .A2(_0834_),
    .ZN(_2213_)
  );
  AND2_X1 _8753_ (
    .A1(reg_pmp_1_addr[28]),
    .A2(_0841_),
    .ZN(_2214_)
  );
  AND2_X1 _8754_ (
    .A1(reg_pmp_0_addr[28]),
    .A2(_0837_),
    .ZN(_2215_)
  );
  AND2_X1 _8755_ (
    .A1(reg_pmp_7_addr[28]),
    .A2(_0849_),
    .ZN(_2216_)
  );
  AND2_X1 _8756_ (
    .A1(reg_pmp_6_addr[28]),
    .A2(_0814_),
    .ZN(_2217_)
  );
  OR2_X1 _8757_ (
    .A1(_2200_),
    .A2(_2202_),
    .ZN(_2218_)
  );
  OR2_X1 _8758_ (
    .A1(_2211_),
    .A2(_2218_),
    .ZN(_2219_)
  );
  OR2_X1 _8759_ (
    .A1(_2198_),
    .A2(_2199_),
    .ZN(_2220_)
  );
  OR2_X1 _8760_ (
    .A1(_2213_),
    .A2(_2215_),
    .ZN(_2221_)
  );
  OR2_X1 _8761_ (
    .A1(_2220_),
    .A2(_2221_),
    .ZN(_2222_)
  );
  OR2_X1 _8762_ (
    .A1(_2219_),
    .A2(_2222_),
    .ZN(_2223_)
  );
  OR2_X1 _8763_ (
    .A1(_2201_),
    .A2(_2204_),
    .ZN(_2224_)
  );
  OR2_X1 _8764_ (
    .A1(_2217_),
    .A2(_2224_),
    .ZN(_2225_)
  );
  AND2_X1 _8765_ (
    .A1(large_1[22]),
    .A2(_0859_),
    .ZN(_2226_)
  );
  OR2_X1 _8766_ (
    .A1(_2208_),
    .A2(_2226_),
    .ZN(_2227_)
  );
  AND2_X1 _8767_ (
    .A1(large_[22]),
    .A2(_0857_),
    .ZN(_2228_)
  );
  OR2_X1 _8768_ (
    .A1(_2212_),
    .A2(_2228_),
    .ZN(_2229_)
  );
  OR2_X1 _8769_ (
    .A1(_2227_),
    .A2(_2229_),
    .ZN(_2230_)
  );
  OR2_X1 _8770_ (
    .A1(_2225_),
    .A2(_2230_),
    .ZN(_2231_)
  );
  OR2_X1 _8771_ (
    .A1(_2223_),
    .A2(_2231_),
    .ZN(_2232_)
  );
  OR2_X1 _8772_ (
    .A1(_2207_),
    .A2(_2214_),
    .ZN(_2233_)
  );
  OR2_X1 _8773_ (
    .A1(_2210_),
    .A2(_2233_),
    .ZN(_2234_)
  );
  OR2_X1 _8774_ (
    .A1(_2203_),
    .A2(_2209_),
    .ZN(_2235_)
  );
  OR2_X1 _8775_ (
    .A1(_2216_),
    .A2(_2235_),
    .ZN(_2236_)
  );
  OR2_X1 _8776_ (
    .A1(_2197_),
    .A2(_2236_),
    .ZN(_2237_)
  );
  OR2_X1 _8777_ (
    .A1(_2234_),
    .A2(_2237_),
    .ZN(_2238_)
  );
  OR2_X1 _8778_ (
    .A1(_2232_),
    .A2(_2238_),
    .ZN(io_rw_rdata[28])
  );
  AND2_X1 _8779_ (
    .A1(io_rw_cmd[1]),
    .A2(_0705_),
    .ZN(_2239_)
  );
  AND2_X1 _8780_ (
    .A1(io_rw_rdata[28]),
    .A2(_2239_),
    .ZN(_2240_)
  );
  OR2_X1 _8781_ (
    .A1(_2196_),
    .A2(_2240_),
    .ZN(_2241_)
  );
  MUX2_X1 _8782_ (
    .A(_2241_),
    .B(reg_pmp_5_addr[28]),
    .S(_1181_),
    .Z(_0055_)
  );
  AND2_X1 _8783_ (
    .A1(io_rw_wdata[29]),
    .A2(_0742_),
    .ZN(_2242_)
  );
  AND2_X1 _8784_ (
    .A1(reg_pmp_1_addr[29]),
    .A2(_0841_),
    .ZN(_2243_)
  );
  AND2_X1 _8785_ (
    .A1(reg_pmp_3_addr[29]),
    .A2(_0844_),
    .ZN(_2244_)
  );
  OR2_X1 _8786_ (
    .A1(_2243_),
    .A2(_2244_),
    .ZN(_2245_)
  );
  AND2_X1 _8787_ (
    .A1(reg_mtvec[29]),
    .A2(_0780_),
    .ZN(_2246_)
  );
  AND2_X1 _8788_ (
    .A1(reg_pmp_2_addr[29]),
    .A2(_0792_),
    .ZN(_2247_)
  );
  OR2_X1 _8789_ (
    .A1(_2246_),
    .A2(_2247_),
    .ZN(_2248_)
  );
  OR2_X1 _8790_ (
    .A1(_2245_),
    .A2(_2248_),
    .ZN(_2249_)
  );
  AND2_X1 _8791_ (
    .A1(reg_mscratch[29]),
    .A2(_0767_),
    .ZN(_2250_)
  );
  AND2_X1 _8792_ (
    .A1(reg_mepc[29]),
    .A2(_0783_),
    .ZN(_2251_)
  );
  OR2_X1 _8793_ (
    .A1(_2250_),
    .A2(_2251_),
    .ZN(_2252_)
  );
  AND2_X1 _8794_ (
    .A1(reg_pmp_0_addr[29]),
    .A2(_0837_),
    .ZN(_2253_)
  );
  AND2_X1 _8795_ (
    .A1(reg_pmp_4_addr[29]),
    .A2(_0805_),
    .ZN(_2254_)
  );
  OR2_X1 _8796_ (
    .A1(_2253_),
    .A2(_2254_),
    .ZN(_2255_)
  );
  OR2_X1 _8797_ (
    .A1(_2252_),
    .A2(_2255_),
    .ZN(_2256_)
  );
  AND2_X1 _8798_ (
    .A1(reg_dscratch0[29]),
    .A2(_0797_),
    .ZN(_2257_)
  );
  AND2_X1 _8799_ (
    .A1(reg_mtval[29]),
    .A2(_0764_),
    .ZN(_2258_)
  );
  OR2_X1 _8800_ (
    .A1(_2257_),
    .A2(_2258_),
    .ZN(_2259_)
  );
  AND2_X1 _8801_ (
    .A1(reg_mcause[29]),
    .A2(_0834_),
    .ZN(_2260_)
  );
  AND2_X1 _8802_ (
    .A1(reg_pmp_5_addr[29]),
    .A2(_0788_),
    .ZN(_2261_)
  );
  OR2_X1 _8803_ (
    .A1(_2260_),
    .A2(_2261_),
    .ZN(_2262_)
  );
  OR2_X1 _8804_ (
    .A1(_2259_),
    .A2(_2262_),
    .ZN(_2263_)
  );
  OR2_X1 _8805_ (
    .A1(_2256_),
    .A2(_2263_),
    .ZN(_2264_)
  );
  OR2_X1 _8806_ (
    .A1(_2249_),
    .A2(_2264_),
    .ZN(_2265_)
  );
  AND2_X1 _8807_ (
    .A1(large_[55]),
    .A2(_0827_),
    .ZN(_2266_)
  );
  AND2_X1 _8808_ (
    .A1(large_[23]),
    .A2(_0822_),
    .ZN(_2267_)
  );
  OR2_X1 _8809_ (
    .A1(_2266_),
    .A2(_2267_),
    .ZN(_2268_)
  );
  AND2_X1 _8810_ (
    .A1(large_1[55]),
    .A2(_0851_),
    .ZN(_2269_)
  );
  AND2_X1 _8811_ (
    .A1(large_1[23]),
    .A2(_0830_),
    .ZN(_2270_)
  );
  OR2_X1 _8812_ (
    .A1(_2269_),
    .A2(_2270_),
    .ZN(_2271_)
  );
  OR2_X1 _8813_ (
    .A1(_2268_),
    .A2(_2271_),
    .ZN(_2272_)
  );
  OR2_X1 _8814_ (
    .A1(_0926_),
    .A2(_1058_),
    .ZN(_2273_)
  );
  AND2_X1 _8815_ (
    .A1(reg_dpc[29]),
    .A2(_0750_),
    .ZN(_2274_)
  );
  AND2_X1 _8816_ (
    .A1(reg_bp_0_address[29]),
    .A2(_0800_),
    .ZN(_2275_)
  );
  OR2_X1 _8817_ (
    .A1(_2274_),
    .A2(_2275_),
    .ZN(_2276_)
  );
  OR2_X1 _8818_ (
    .A1(_2273_),
    .A2(_2276_),
    .ZN(_2277_)
  );
  AND2_X1 _8819_ (
    .A1(reg_pmp_6_addr[29]),
    .A2(_0814_),
    .ZN(_2278_)
  );
  AND2_X1 _8820_ (
    .A1(reg_pmp_7_addr[29]),
    .A2(_0849_),
    .ZN(_2279_)
  );
  OR2_X1 _8821_ (
    .A1(_2278_),
    .A2(_2279_),
    .ZN(_2280_)
  );
  OR2_X1 _8822_ (
    .A1(_2277_),
    .A2(_2280_),
    .ZN(_2281_)
  );
  OR2_X1 _8823_ (
    .A1(_2272_),
    .A2(_2281_),
    .ZN(_2282_)
  );
  OR2_X1 _8824_ (
    .A1(_2265_),
    .A2(_2282_),
    .ZN(io_rw_rdata[29])
  );
  AND2_X1 _8825_ (
    .A1(io_rw_cmd[1]),
    .A2(_0706_),
    .ZN(_2283_)
  );
  AND2_X1 _8826_ (
    .A1(io_rw_rdata[29]),
    .A2(_2283_),
    .ZN(_2284_)
  );
  OR2_X1 _8827_ (
    .A1(_2242_),
    .A2(_2284_),
    .ZN(_2285_)
  );
  MUX2_X1 _8828_ (
    .A(_2285_),
    .B(reg_pmp_5_addr[29]),
    .S(_1181_),
    .Z(_0056_)
  );
  AND2_X1 _8829_ (
    .A1(_0006_),
    .A2(_0754_),
    .ZN(_2286_)
  );
  INV_X1 _8830_ (
    .A(_2286_),
    .ZN(_2287_)
  );
  AND2_X1 _8831_ (
    .A1(_0736_),
    .A2(_2286_),
    .ZN(_2288_)
  );
  OR2_X1 _8832_ (
    .A1(_0737_),
    .A2(_2287_),
    .ZN(_2289_)
  );
  AND2_X1 _8833_ (
    .A1(_1241_),
    .A2(_1290_),
    .ZN(_2290_)
  );
  MUX2_X1 _8834_ (
    .A(reg_pmp_0_cfg_w),
    .B(_2290_),
    .S(_2288_),
    .Z(_0057_)
  );
  OR2_X1 _8835_ (
    .A1(reg_pmp_5_cfg_a[0]),
    .A2(_1075_),
    .ZN(_2291_)
  );
  AND2_X1 _8836_ (
    .A1(_0654_),
    .A2(_2291_),
    .ZN(_2292_)
  );
  OR2_X1 _8837_ (
    .A1(_1076_),
    .A2(_1698_),
    .ZN(_2293_)
  );
  AND2_X1 _8838_ (
    .A1(_2292_),
    .A2(_2293_),
    .ZN(_0058_)
  );
  OR2_X1 _8839_ (
    .A1(reg_pmp_5_cfg_a[1]),
    .A2(_1075_),
    .ZN(_2294_)
  );
  AND2_X1 _8840_ (
    .A1(_0654_),
    .A2(_2294_),
    .ZN(_2295_)
  );
  OR2_X1 _8841_ (
    .A1(_1076_),
    .A2(_1748_),
    .ZN(_2296_)
  );
  AND2_X1 _8842_ (
    .A1(_2295_),
    .A2(_2296_),
    .ZN(_0059_)
  );
  OR2_X1 _8843_ (
    .A1(reg_pmp_5_cfg_l),
    .A2(_1075_),
    .ZN(_2297_)
  );
  AND2_X1 _8844_ (
    .A1(_0654_),
    .A2(_2297_),
    .ZN(_2298_)
  );
  OR2_X1 _8845_ (
    .A1(_1076_),
    .A2(_1880_),
    .ZN(_2299_)
  );
  AND2_X1 _8846_ (
    .A1(_2298_),
    .A2(_2299_),
    .ZN(_0060_)
  );
  AND2_X1 _8847_ (
    .A1(reg_pmp_5_cfg_l),
    .A2(reg_pmp_5_cfg_a[0]),
    .ZN(_2300_)
  );
  AND2_X1 _8848_ (
    .A1(_0016_),
    .A2(_2300_),
    .ZN(_2301_)
  );
  OR2_X1 _8849_ (
    .A1(reg_pmp_4_cfg_l),
    .A2(_2301_),
    .ZN(_2302_)
  );
  OR2_X1 _8850_ (
    .A1(_0737_),
    .A2(_2302_),
    .ZN(_2303_)
  );
  OR2_X1 _8851_ (
    .A1(_0806_),
    .A2(_2303_),
    .ZN(_2304_)
  );
  MUX2_X1 _8852_ (
    .A(_1241_),
    .B(reg_pmp_4_addr[0]),
    .S(_2304_),
    .Z(_0061_)
  );
  MUX2_X1 _8853_ (
    .A(_1290_),
    .B(reg_pmp_4_addr[1]),
    .S(_2304_),
    .Z(_0062_)
  );
  MUX2_X1 _8854_ (
    .A(_1346_),
    .B(reg_pmp_4_addr[2]),
    .S(_2304_),
    .Z(_0063_)
  );
  MUX2_X1 _8855_ (
    .A(_1409_),
    .B(reg_pmp_4_addr[3]),
    .S(_2304_),
    .Z(_0064_)
  );
  MUX2_X1 _8856_ (
    .A(_1456_),
    .B(reg_pmp_4_addr[4]),
    .S(_2304_),
    .Z(_0065_)
  );
  MUX2_X1 _8857_ (
    .A(_1499_),
    .B(reg_pmp_4_addr[5]),
    .S(_2304_),
    .Z(_0066_)
  );
  MUX2_X1 _8858_ (
    .A(_1545_),
    .B(reg_pmp_4_addr[6]),
    .S(_2304_),
    .Z(_0067_)
  );
  MUX2_X1 _8859_ (
    .A(_1601_),
    .B(reg_pmp_4_addr[7]),
    .S(_2304_),
    .Z(_0068_)
  );
  MUX2_X1 _8860_ (
    .A(_1129_),
    .B(reg_pmp_4_addr[8]),
    .S(_2304_),
    .Z(_0069_)
  );
  MUX2_X1 _8861_ (
    .A(_1175_),
    .B(reg_pmp_4_addr[9]),
    .S(_2304_),
    .Z(_0070_)
  );
  MUX2_X1 _8862_ (
    .A(_1647_),
    .B(reg_pmp_4_addr[10]),
    .S(_2304_),
    .Z(_0071_)
  );
  MUX2_X1 _8863_ (
    .A(_1698_),
    .B(reg_pmp_4_addr[11]),
    .S(_2304_),
    .Z(_0072_)
  );
  MUX2_X1 _8864_ (
    .A(_1748_),
    .B(reg_pmp_4_addr[12]),
    .S(_2304_),
    .Z(_0073_)
  );
  MUX2_X1 _8865_ (
    .A(_1790_),
    .B(reg_pmp_4_addr[13]),
    .S(_2304_),
    .Z(_0074_)
  );
  MUX2_X1 _8866_ (
    .A(_1832_),
    .B(reg_pmp_4_addr[14]),
    .S(_2304_),
    .Z(_0075_)
  );
  MUX2_X1 _8867_ (
    .A(_1880_),
    .B(reg_pmp_4_addr[15]),
    .S(_2304_),
    .Z(_0076_)
  );
  MUX2_X1 _8868_ (
    .A(_0862_),
    .B(reg_pmp_4_addr[16]),
    .S(_2304_),
    .Z(_0077_)
  );
  MUX2_X1 _8869_ (
    .A(_1926_),
    .B(reg_pmp_4_addr[17]),
    .S(_2304_),
    .Z(_0078_)
  );
  MUX2_X1 _8870_ (
    .A(_0908_),
    .B(reg_pmp_4_addr[18]),
    .S(_2304_),
    .Z(_0079_)
  );
  MUX2_X1 _8871_ (
    .A(_0967_),
    .B(reg_pmp_4_addr[19]),
    .S(_2304_),
    .Z(_0080_)
  );
  MUX2_X1 _8872_ (
    .A(_1017_),
    .B(reg_pmp_4_addr[20]),
    .S(_2304_),
    .Z(_0081_)
  );
  MUX2_X1 _8873_ (
    .A(_1968_),
    .B(reg_pmp_4_addr[21]),
    .S(_2304_),
    .Z(_0082_)
  );
  MUX2_X1 _8874_ (
    .A(_2010_),
    .B(reg_pmp_4_addr[22]),
    .S(_2304_),
    .Z(_0083_)
  );
  MUX2_X1 _8875_ (
    .A(_1071_),
    .B(reg_pmp_4_addr[23]),
    .S(_2304_),
    .Z(_0084_)
  );
  MUX2_X1 _8876_ (
    .A(_2056_),
    .B(reg_pmp_4_addr[24]),
    .S(_2304_),
    .Z(_0085_)
  );
  MUX2_X1 _8877_ (
    .A(_2102_),
    .B(reg_pmp_4_addr[25]),
    .S(_2304_),
    .Z(_0086_)
  );
  MUX2_X1 _8878_ (
    .A(_2148_),
    .B(reg_pmp_4_addr[26]),
    .S(_2304_),
    .Z(_0087_)
  );
  MUX2_X1 _8879_ (
    .A(_2195_),
    .B(reg_pmp_4_addr[27]),
    .S(_2304_),
    .Z(_0088_)
  );
  MUX2_X1 _8880_ (
    .A(_2241_),
    .B(reg_pmp_4_addr[28]),
    .S(_2304_),
    .Z(_0089_)
  );
  MUX2_X1 _8881_ (
    .A(_2285_),
    .B(reg_pmp_4_addr[29]),
    .S(_2304_),
    .Z(_0090_)
  );
  AND2_X1 _8882_ (
    .A1(_0013_),
    .A2(_0733_),
    .ZN(_2305_)
  );
  INV_X1 _8883_ (
    .A(_2305_),
    .ZN(_2306_)
  );
  AND2_X1 _8884_ (
    .A1(_0736_),
    .A2(_2305_),
    .ZN(_2307_)
  );
  OR2_X1 _8885_ (
    .A1(_0737_),
    .A2(_2306_),
    .ZN(_2308_)
  );
  MUX2_X1 _8886_ (
    .A(reg_pmp_4_cfg_w),
    .B(_2290_),
    .S(_2307_),
    .Z(_0091_)
  );
  MUX2_X1 _8887_ (
    .A(reg_pmp_4_cfg_x),
    .B(_1346_),
    .S(_2307_),
    .Z(_0092_)
  );
  OR2_X1 _8888_ (
    .A1(reg_pmp_4_cfg_a[0]),
    .A2(_2307_),
    .ZN(_2309_)
  );
  AND2_X1 _8889_ (
    .A1(_0654_),
    .A2(_2309_),
    .ZN(_2310_)
  );
  OR2_X1 _8890_ (
    .A1(_1409_),
    .A2(_2308_),
    .ZN(_2311_)
  );
  AND2_X1 _8891_ (
    .A1(_2310_),
    .A2(_2311_),
    .ZN(_0093_)
  );
  OR2_X1 _8892_ (
    .A1(reg_pmp_4_cfg_a[1]),
    .A2(_2307_),
    .ZN(_2312_)
  );
  AND2_X1 _8893_ (
    .A1(_0654_),
    .A2(_2312_),
    .ZN(_2313_)
  );
  OR2_X1 _8894_ (
    .A1(_1456_),
    .A2(_2308_),
    .ZN(_2314_)
  );
  AND2_X1 _8895_ (
    .A1(_2313_),
    .A2(_2314_),
    .ZN(_0094_)
  );
  OR2_X1 _8896_ (
    .A1(reg_pmp_4_cfg_l),
    .A2(_2307_),
    .ZN(_2315_)
  );
  AND2_X1 _8897_ (
    .A1(_0654_),
    .A2(_2315_),
    .ZN(_2316_)
  );
  OR2_X1 _8898_ (
    .A1(_1601_),
    .A2(_2308_),
    .ZN(_2317_)
  );
  AND2_X1 _8899_ (
    .A1(_2316_),
    .A2(_2317_),
    .ZN(_0095_)
  );
  AND2_X1 _8900_ (
    .A1(_0011_),
    .A2(_0754_),
    .ZN(_2318_)
  );
  INV_X1 _8901_ (
    .A(_2318_),
    .ZN(_2319_)
  );
  AND2_X1 _8902_ (
    .A1(_0736_),
    .A2(_2318_),
    .ZN(_2320_)
  );
  OR2_X1 _8903_ (
    .A1(_0737_),
    .A2(_2319_),
    .ZN(_2321_)
  );
  AND2_X1 _8904_ (
    .A1(_2056_),
    .A2(_2102_),
    .ZN(_2322_)
  );
  MUX2_X1 _8905_ (
    .A(reg_pmp_3_cfg_w),
    .B(_2322_),
    .S(_2320_),
    .Z(_0096_)
  );
  MUX2_X1 _8906_ (
    .A(reg_pmp_3_cfg_x),
    .B(_2148_),
    .S(_2320_),
    .Z(_0097_)
  );
  MUX2_X1 _8907_ (
    .A(reg_pmp_3_cfg_r),
    .B(_2056_),
    .S(_2320_),
    .Z(_0098_)
  );
  AND2_X1 _8908_ (
    .A1(_0009_),
    .A2(_0754_),
    .ZN(_2323_)
  );
  INV_X1 _8909_ (
    .A(_2323_),
    .ZN(_2324_)
  );
  AND2_X1 _8910_ (
    .A1(_0736_),
    .A2(_2323_),
    .ZN(_2325_)
  );
  OR2_X1 _8911_ (
    .A1(_0737_),
    .A2(_2324_),
    .ZN(_2326_)
  );
  AND2_X1 _8912_ (
    .A1(_0862_),
    .A2(_1926_),
    .ZN(_2327_)
  );
  MUX2_X1 _8913_ (
    .A(reg_pmp_2_cfg_w),
    .B(_2327_),
    .S(_2325_),
    .Z(_0099_)
  );
  OR2_X1 _8914_ (
    .A1(reg_pmp_3_cfg_a[0]),
    .A2(_2320_),
    .ZN(_2328_)
  );
  AND2_X1 _8915_ (
    .A1(_0654_),
    .A2(_2328_),
    .ZN(_2329_)
  );
  OR2_X1 _8916_ (
    .A1(_2195_),
    .A2(_2321_),
    .ZN(_2330_)
  );
  AND2_X1 _8917_ (
    .A1(_2329_),
    .A2(_2330_),
    .ZN(_0100_)
  );
  OR2_X1 _8918_ (
    .A1(reg_pmp_3_cfg_a[1]),
    .A2(_2320_),
    .ZN(_2331_)
  );
  AND2_X1 _8919_ (
    .A1(_0654_),
    .A2(_2331_),
    .ZN(_2332_)
  );
  OR2_X1 _8920_ (
    .A1(_2241_),
    .A2(_2321_),
    .ZN(_2333_)
  );
  AND2_X1 _8921_ (
    .A1(_2332_),
    .A2(_2333_),
    .ZN(_0101_)
  );
  OR2_X1 _8922_ (
    .A1(reg_pmp_3_cfg_l),
    .A2(_2320_),
    .ZN(_2334_)
  );
  AND2_X1 _8923_ (
    .A1(_0654_),
    .A2(_2334_),
    .ZN(_2335_)
  );
  AND2_X1 _8924_ (
    .A1(io_rw_wdata[31]),
    .A2(_0742_),
    .ZN(_2336_)
  );
  AND2_X1 _8925_ (
    .A1(large_1[57]),
    .A2(_0851_),
    .ZN(_2337_)
  );
  AND2_X1 _8926_ (
    .A1(large_[57]),
    .A2(_0827_),
    .ZN(_2338_)
  );
  AND2_X1 _8927_ (
    .A1(large_1[25]),
    .A2(_0830_),
    .ZN(_2339_)
  );
  OR2_X1 _8928_ (
    .A1(_2338_),
    .A2(_2339_),
    .ZN(_2340_)
  );
  OR2_X1 _8929_ (
    .A1(_2337_),
    .A2(_2340_),
    .ZN(_2341_)
  );
  AND2_X1 _8930_ (
    .A1(reg_pmp_7_cfg_l),
    .A2(_0733_),
    .ZN(_2342_)
  );
  AND2_X1 _8931_ (
    .A1(reg_pmp_3_cfg_l),
    .A2(_0754_),
    .ZN(_2343_)
  );
  OR2_X1 _8932_ (
    .A1(_2342_),
    .A2(_2343_),
    .ZN(_2344_)
  );
  AND2_X1 _8933_ (
    .A1(reg_bp_0_address[31]),
    .A2(_0800_),
    .ZN(_2345_)
  );
  AND2_X1 _8934_ (
    .A1(reg_mepc[31]),
    .A2(_0783_),
    .ZN(_2346_)
  );
  OR2_X1 _8935_ (
    .A1(_2345_),
    .A2(_2346_),
    .ZN(_2347_)
  );
  OR2_X1 _8936_ (
    .A1(_2344_),
    .A2(_2347_),
    .ZN(_2348_)
  );
  AND2_X1 _8937_ (
    .A1(reg_mcause[31]),
    .A2(_0834_),
    .ZN(_2349_)
  );
  AND2_X1 _8938_ (
    .A1(reg_dpc[31]),
    .A2(_0750_),
    .ZN(_2350_)
  );
  OR2_X1 _8939_ (
    .A1(_2349_),
    .A2(_2350_),
    .ZN(_2351_)
  );
  AND2_X1 _8940_ (
    .A1(reg_dscratch0[31]),
    .A2(_0797_),
    .ZN(_2352_)
  );
  AND2_X1 _8941_ (
    .A1(reg_mtvec[31]),
    .A2(_0780_),
    .ZN(_2353_)
  );
  OR2_X1 _8942_ (
    .A1(_2352_),
    .A2(_2353_),
    .ZN(_2354_)
  );
  OR2_X1 _8943_ (
    .A1(_2351_),
    .A2(_2354_),
    .ZN(_2355_)
  );
  AND2_X1 _8944_ (
    .A1(large_[25]),
    .A2(_0822_),
    .ZN(_2356_)
  );
  AND2_X1 _8945_ (
    .A1(reg_mtval[31]),
    .A2(_0764_),
    .ZN(_2357_)
  );
  AND2_X1 _8946_ (
    .A1(reg_mscratch[31]),
    .A2(_0767_),
    .ZN(_2358_)
  );
  OR2_X1 _8947_ (
    .A1(_2357_),
    .A2(_2358_),
    .ZN(_2359_)
  );
  OR2_X1 _8948_ (
    .A1(_2356_),
    .A2(_2359_),
    .ZN(_2360_)
  );
  OR2_X1 _8949_ (
    .A1(_2355_),
    .A2(_2360_),
    .ZN(_2361_)
  );
  OR2_X1 _8950_ (
    .A1(_2348_),
    .A2(_2361_),
    .ZN(_2362_)
  );
  OR2_X1 _8951_ (
    .A1(_2341_),
    .A2(_2362_),
    .ZN(io_rw_rdata[31])
  );
  AND2_X1 _8952_ (
    .A1(io_rw_cmd[1]),
    .A2(_0708_),
    .ZN(_2363_)
  );
  AND2_X1 _8953_ (
    .A1(io_rw_rdata[31]),
    .A2(_2363_),
    .ZN(_2364_)
  );
  OR2_X1 _8954_ (
    .A1(_2336_),
    .A2(_2364_),
    .ZN(_2365_)
  );
  OR2_X1 _8955_ (
    .A1(_2321_),
    .A2(_2365_),
    .ZN(_2366_)
  );
  AND2_X1 _8956_ (
    .A1(_2335_),
    .A2(_2366_),
    .ZN(_0102_)
  );
  AND2_X1 _8957_ (
    .A1(reg_pmp_3_cfg_l),
    .A2(reg_pmp_3_cfg_a[0]),
    .ZN(_2367_)
  );
  AND2_X1 _8958_ (
    .A1(_0012_),
    .A2(_2367_),
    .ZN(_2368_)
  );
  OR2_X1 _8959_ (
    .A1(reg_pmp_2_cfg_l),
    .A2(_2368_),
    .ZN(_2369_)
  );
  OR2_X1 _8960_ (
    .A1(_0737_),
    .A2(_2369_),
    .ZN(_2370_)
  );
  OR2_X1 _8961_ (
    .A1(_0793_),
    .A2(_2370_),
    .ZN(_2371_)
  );
  MUX2_X1 _8962_ (
    .A(_1241_),
    .B(reg_pmp_2_addr[0]),
    .S(_2371_),
    .Z(_0103_)
  );
  MUX2_X1 _8963_ (
    .A(_1290_),
    .B(reg_pmp_2_addr[1]),
    .S(_2371_),
    .Z(_0104_)
  );
  MUX2_X1 _8964_ (
    .A(_1346_),
    .B(reg_pmp_2_addr[2]),
    .S(_2371_),
    .Z(_0105_)
  );
  MUX2_X1 _8965_ (
    .A(_1409_),
    .B(reg_pmp_2_addr[3]),
    .S(_2371_),
    .Z(_0106_)
  );
  MUX2_X1 _8966_ (
    .A(_1456_),
    .B(reg_pmp_2_addr[4]),
    .S(_2371_),
    .Z(_0107_)
  );
  MUX2_X1 _8967_ (
    .A(_1499_),
    .B(reg_pmp_2_addr[5]),
    .S(_2371_),
    .Z(_0108_)
  );
  MUX2_X1 _8968_ (
    .A(_1545_),
    .B(reg_pmp_2_addr[6]),
    .S(_2371_),
    .Z(_0109_)
  );
  MUX2_X1 _8969_ (
    .A(_1601_),
    .B(reg_pmp_2_addr[7]),
    .S(_2371_),
    .Z(_0110_)
  );
  MUX2_X1 _8970_ (
    .A(_1129_),
    .B(reg_pmp_2_addr[8]),
    .S(_2371_),
    .Z(_0111_)
  );
  MUX2_X1 _8971_ (
    .A(_1175_),
    .B(reg_pmp_2_addr[9]),
    .S(_2371_),
    .Z(_0112_)
  );
  MUX2_X1 _8972_ (
    .A(_1647_),
    .B(reg_pmp_2_addr[10]),
    .S(_2371_),
    .Z(_0113_)
  );
  MUX2_X1 _8973_ (
    .A(_1698_),
    .B(reg_pmp_2_addr[11]),
    .S(_2371_),
    .Z(_0114_)
  );
  MUX2_X1 _8974_ (
    .A(_1748_),
    .B(reg_pmp_2_addr[12]),
    .S(_2371_),
    .Z(_0115_)
  );
  MUX2_X1 _8975_ (
    .A(_1790_),
    .B(reg_pmp_2_addr[13]),
    .S(_2371_),
    .Z(_0116_)
  );
  MUX2_X1 _8976_ (
    .A(_1832_),
    .B(reg_pmp_2_addr[14]),
    .S(_2371_),
    .Z(_0117_)
  );
  MUX2_X1 _8977_ (
    .A(_1880_),
    .B(reg_pmp_2_addr[15]),
    .S(_2371_),
    .Z(_0118_)
  );
  MUX2_X1 _8978_ (
    .A(_0862_),
    .B(reg_pmp_2_addr[16]),
    .S(_2371_),
    .Z(_0119_)
  );
  MUX2_X1 _8979_ (
    .A(_1926_),
    .B(reg_pmp_2_addr[17]),
    .S(_2371_),
    .Z(_0120_)
  );
  MUX2_X1 _8980_ (
    .A(_0908_),
    .B(reg_pmp_2_addr[18]),
    .S(_2371_),
    .Z(_0121_)
  );
  MUX2_X1 _8981_ (
    .A(_0967_),
    .B(reg_pmp_2_addr[19]),
    .S(_2371_),
    .Z(_0122_)
  );
  MUX2_X1 _8982_ (
    .A(_1017_),
    .B(reg_pmp_2_addr[20]),
    .S(_2371_),
    .Z(_0123_)
  );
  MUX2_X1 _8983_ (
    .A(_1968_),
    .B(reg_pmp_2_addr[21]),
    .S(_2371_),
    .Z(_0124_)
  );
  MUX2_X1 _8984_ (
    .A(_2010_),
    .B(reg_pmp_2_addr[22]),
    .S(_2371_),
    .Z(_0125_)
  );
  MUX2_X1 _8985_ (
    .A(_1071_),
    .B(reg_pmp_2_addr[23]),
    .S(_2371_),
    .Z(_0126_)
  );
  MUX2_X1 _8986_ (
    .A(_2056_),
    .B(reg_pmp_2_addr[24]),
    .S(_2371_),
    .Z(_0127_)
  );
  MUX2_X1 _8987_ (
    .A(_2102_),
    .B(reg_pmp_2_addr[25]),
    .S(_2371_),
    .Z(_0128_)
  );
  MUX2_X1 _8988_ (
    .A(_2148_),
    .B(reg_pmp_2_addr[26]),
    .S(_2371_),
    .Z(_0129_)
  );
  MUX2_X1 _8989_ (
    .A(_2195_),
    .B(reg_pmp_2_addr[27]),
    .S(_2371_),
    .Z(_0130_)
  );
  MUX2_X1 _8990_ (
    .A(_2241_),
    .B(reg_pmp_2_addr[28]),
    .S(_2371_),
    .Z(_0131_)
  );
  MUX2_X1 _8991_ (
    .A(_2285_),
    .B(reg_pmp_2_addr[29]),
    .S(_2371_),
    .Z(_0132_)
  );
  AND2_X1 _8992_ (
    .A1(_0007_),
    .A2(_0754_),
    .ZN(_2372_)
  );
  INV_X1 _8993_ (
    .A(_2372_),
    .ZN(_2373_)
  );
  AND2_X1 _8994_ (
    .A1(_0736_),
    .A2(_2372_),
    .ZN(_2374_)
  );
  OR2_X1 _8995_ (
    .A1(_0737_),
    .A2(_2373_),
    .ZN(_2375_)
  );
  MUX2_X1 _8996_ (
    .A(reg_pmp_1_cfg_w),
    .B(_1176_),
    .S(_2374_),
    .Z(_0133_)
  );
  MUX2_X1 _8997_ (
    .A(reg_pmp_2_cfg_r),
    .B(_0862_),
    .S(_2325_),
    .Z(_0134_)
  );
  AND2_X1 _8998_ (
    .A1(reg_pmp_4_cfg_l),
    .A2(reg_pmp_4_cfg_a[0]),
    .ZN(_2376_)
  );
  AND2_X1 _8999_ (
    .A1(_0014_),
    .A2(_2376_),
    .ZN(_2377_)
  );
  OR2_X1 _9000_ (
    .A1(reg_pmp_3_cfg_l),
    .A2(_2377_),
    .ZN(_2378_)
  );
  OR2_X1 _9001_ (
    .A1(_0737_),
    .A2(_2378_),
    .ZN(_2379_)
  );
  OR2_X1 _9002_ (
    .A1(_0845_),
    .A2(_2379_),
    .ZN(_2380_)
  );
  MUX2_X1 _9003_ (
    .A(_1241_),
    .B(reg_pmp_3_addr[0]),
    .S(_2380_),
    .Z(_0135_)
  );
  MUX2_X1 _9004_ (
    .A(_1290_),
    .B(reg_pmp_3_addr[1]),
    .S(_2380_),
    .Z(_0136_)
  );
  MUX2_X1 _9005_ (
    .A(_1346_),
    .B(reg_pmp_3_addr[2]),
    .S(_2380_),
    .Z(_0137_)
  );
  MUX2_X1 _9006_ (
    .A(_1409_),
    .B(reg_pmp_3_addr[3]),
    .S(_2380_),
    .Z(_0138_)
  );
  MUX2_X1 _9007_ (
    .A(_1456_),
    .B(reg_pmp_3_addr[4]),
    .S(_2380_),
    .Z(_0139_)
  );
  MUX2_X1 _9008_ (
    .A(_1499_),
    .B(reg_pmp_3_addr[5]),
    .S(_2380_),
    .Z(_0140_)
  );
  MUX2_X1 _9009_ (
    .A(_1545_),
    .B(reg_pmp_3_addr[6]),
    .S(_2380_),
    .Z(_0141_)
  );
  MUX2_X1 _9010_ (
    .A(_1601_),
    .B(reg_pmp_3_addr[7]),
    .S(_2380_),
    .Z(_0142_)
  );
  MUX2_X1 _9011_ (
    .A(_1129_),
    .B(reg_pmp_3_addr[8]),
    .S(_2380_),
    .Z(_0143_)
  );
  MUX2_X1 _9012_ (
    .A(_1175_),
    .B(reg_pmp_3_addr[9]),
    .S(_2380_),
    .Z(_0144_)
  );
  MUX2_X1 _9013_ (
    .A(_1647_),
    .B(reg_pmp_3_addr[10]),
    .S(_2380_),
    .Z(_0145_)
  );
  MUX2_X1 _9014_ (
    .A(_1698_),
    .B(reg_pmp_3_addr[11]),
    .S(_2380_),
    .Z(_0146_)
  );
  MUX2_X1 _9015_ (
    .A(_1748_),
    .B(reg_pmp_3_addr[12]),
    .S(_2380_),
    .Z(_0147_)
  );
  MUX2_X1 _9016_ (
    .A(_1790_),
    .B(reg_pmp_3_addr[13]),
    .S(_2380_),
    .Z(_0148_)
  );
  MUX2_X1 _9017_ (
    .A(_1832_),
    .B(reg_pmp_3_addr[14]),
    .S(_2380_),
    .Z(_0149_)
  );
  MUX2_X1 _9018_ (
    .A(_1880_),
    .B(reg_pmp_3_addr[15]),
    .S(_2380_),
    .Z(_0150_)
  );
  MUX2_X1 _9019_ (
    .A(_0862_),
    .B(reg_pmp_3_addr[16]),
    .S(_2380_),
    .Z(_0151_)
  );
  MUX2_X1 _9020_ (
    .A(_1926_),
    .B(reg_pmp_3_addr[17]),
    .S(_2380_),
    .Z(_0152_)
  );
  MUX2_X1 _9021_ (
    .A(_0908_),
    .B(reg_pmp_3_addr[18]),
    .S(_2380_),
    .Z(_0153_)
  );
  MUX2_X1 _9022_ (
    .A(_0967_),
    .B(reg_pmp_3_addr[19]),
    .S(_2380_),
    .Z(_0154_)
  );
  MUX2_X1 _9023_ (
    .A(_1017_),
    .B(reg_pmp_3_addr[20]),
    .S(_2380_),
    .Z(_0155_)
  );
  MUX2_X1 _9024_ (
    .A(_1968_),
    .B(reg_pmp_3_addr[21]),
    .S(_2380_),
    .Z(_0156_)
  );
  MUX2_X1 _9025_ (
    .A(_2010_),
    .B(reg_pmp_3_addr[22]),
    .S(_2380_),
    .Z(_0157_)
  );
  MUX2_X1 _9026_ (
    .A(_1071_),
    .B(reg_pmp_3_addr[23]),
    .S(_2380_),
    .Z(_0158_)
  );
  MUX2_X1 _9027_ (
    .A(_2056_),
    .B(reg_pmp_3_addr[24]),
    .S(_2380_),
    .Z(_0159_)
  );
  MUX2_X1 _9028_ (
    .A(_2102_),
    .B(reg_pmp_3_addr[25]),
    .S(_2380_),
    .Z(_0160_)
  );
  MUX2_X1 _9029_ (
    .A(_2148_),
    .B(reg_pmp_3_addr[26]),
    .S(_2380_),
    .Z(_0161_)
  );
  MUX2_X1 _9030_ (
    .A(_2195_),
    .B(reg_pmp_3_addr[27]),
    .S(_2380_),
    .Z(_0162_)
  );
  MUX2_X1 _9031_ (
    .A(_2241_),
    .B(reg_pmp_3_addr[28]),
    .S(_2380_),
    .Z(_0163_)
  );
  MUX2_X1 _9032_ (
    .A(_2285_),
    .B(reg_pmp_3_addr[29]),
    .S(_2380_),
    .Z(_0164_)
  );
  OR2_X1 _9033_ (
    .A1(reg_pmp_2_cfg_a[0]),
    .A2(_2325_),
    .ZN(_2381_)
  );
  AND2_X1 _9034_ (
    .A1(_0654_),
    .A2(_2381_),
    .ZN(_2382_)
  );
  OR2_X1 _9035_ (
    .A1(_0967_),
    .A2(_2326_),
    .ZN(_2383_)
  );
  AND2_X1 _9036_ (
    .A1(_2382_),
    .A2(_2383_),
    .ZN(_0165_)
  );
  OR2_X1 _9037_ (
    .A1(reg_pmp_2_cfg_a[1]),
    .A2(_2325_),
    .ZN(_2384_)
  );
  AND2_X1 _9038_ (
    .A1(_0654_),
    .A2(_2384_),
    .ZN(_2385_)
  );
  OR2_X1 _9039_ (
    .A1(_1017_),
    .A2(_2326_),
    .ZN(_2386_)
  );
  AND2_X1 _9040_ (
    .A1(_2385_),
    .A2(_2386_),
    .ZN(_0166_)
  );
  OR2_X1 _9041_ (
    .A1(reg_pmp_2_cfg_l),
    .A2(_2325_),
    .ZN(_2387_)
  );
  AND2_X1 _9042_ (
    .A1(_0654_),
    .A2(_2387_),
    .ZN(_2388_)
  );
  OR2_X1 _9043_ (
    .A1(_1071_),
    .A2(_2326_),
    .ZN(_2389_)
  );
  AND2_X1 _9044_ (
    .A1(_2388_),
    .A2(_2389_),
    .ZN(_0167_)
  );
  MUX2_X1 _9045_ (
    .A(reg_pmp_1_cfg_r),
    .B(_1129_),
    .S(_2374_),
    .Z(_0168_)
  );
  MUX2_X1 _9046_ (
    .A(reg_pmp_4_cfg_r),
    .B(_1241_),
    .S(_2307_),
    .Z(_0169_)
  );
  MUX2_X1 _9047_ (
    .A(reg_pmp_1_cfg_x),
    .B(_1647_),
    .S(_2374_),
    .Z(_0170_)
  );
  MUX2_X1 _9048_ (
    .A(reg_pmp_2_cfg_x),
    .B(_0908_),
    .S(_2325_),
    .Z(_0171_)
  );
  OR2_X1 _9049_ (
    .A1(reg_pmp_1_cfg_a[0]),
    .A2(_2374_),
    .ZN(_2390_)
  );
  AND2_X1 _9050_ (
    .A1(_0654_),
    .A2(_2390_),
    .ZN(_2391_)
  );
  OR2_X1 _9051_ (
    .A1(_1698_),
    .A2(_2375_),
    .ZN(_2392_)
  );
  AND2_X1 _9052_ (
    .A1(_2391_),
    .A2(_2392_),
    .ZN(_0172_)
  );
  OR2_X1 _9053_ (
    .A1(reg_pmp_1_cfg_a[1]),
    .A2(_2374_),
    .ZN(_2393_)
  );
  AND2_X1 _9054_ (
    .A1(_0654_),
    .A2(_2393_),
    .ZN(_2394_)
  );
  OR2_X1 _9055_ (
    .A1(_1748_),
    .A2(_2375_),
    .ZN(_2395_)
  );
  AND2_X1 _9056_ (
    .A1(_2394_),
    .A2(_2395_),
    .ZN(_0173_)
  );
  OR2_X1 _9057_ (
    .A1(reg_pmp_1_cfg_l),
    .A2(_2374_),
    .ZN(_2396_)
  );
  AND2_X1 _9058_ (
    .A1(_0654_),
    .A2(_2396_),
    .ZN(_2397_)
  );
  OR2_X1 _9059_ (
    .A1(_1880_),
    .A2(_2375_),
    .ZN(_2398_)
  );
  AND2_X1 _9060_ (
    .A1(_2397_),
    .A2(_2398_),
    .ZN(_0174_)
  );
  MUX2_X1 _9061_ (
    .A(reg_pmp_0_cfg_r),
    .B(_1241_),
    .S(_2288_),
    .Z(_0175_)
  );
  AND2_X1 _9062_ (
    .A1(reg_pmp_1_cfg_l),
    .A2(reg_pmp_1_cfg_a[0]),
    .ZN(_2399_)
  );
  AND2_X1 _9063_ (
    .A1(_0008_),
    .A2(_2399_),
    .ZN(_2400_)
  );
  OR2_X1 _9064_ (
    .A1(reg_pmp_0_cfg_l),
    .A2(_2400_),
    .ZN(_2401_)
  );
  OR2_X1 _9065_ (
    .A1(_0737_),
    .A2(_2401_),
    .ZN(_2402_)
  );
  OR2_X1 _9066_ (
    .A1(_0838_),
    .A2(_2402_),
    .ZN(_2403_)
  );
  MUX2_X1 _9067_ (
    .A(_1241_),
    .B(reg_pmp_0_addr[0]),
    .S(_2403_),
    .Z(_0176_)
  );
  MUX2_X1 _9068_ (
    .A(_1290_),
    .B(reg_pmp_0_addr[1]),
    .S(_2403_),
    .Z(_0177_)
  );
  MUX2_X1 _9069_ (
    .A(_1346_),
    .B(reg_pmp_0_addr[2]),
    .S(_2403_),
    .Z(_0178_)
  );
  MUX2_X1 _9070_ (
    .A(_1409_),
    .B(reg_pmp_0_addr[3]),
    .S(_2403_),
    .Z(_0179_)
  );
  MUX2_X1 _9071_ (
    .A(_1456_),
    .B(reg_pmp_0_addr[4]),
    .S(_2403_),
    .Z(_0180_)
  );
  MUX2_X1 _9072_ (
    .A(_1499_),
    .B(reg_pmp_0_addr[5]),
    .S(_2403_),
    .Z(_0181_)
  );
  MUX2_X1 _9073_ (
    .A(_1545_),
    .B(reg_pmp_0_addr[6]),
    .S(_2403_),
    .Z(_0182_)
  );
  MUX2_X1 _9074_ (
    .A(_1601_),
    .B(reg_pmp_0_addr[7]),
    .S(_2403_),
    .Z(_0183_)
  );
  MUX2_X1 _9075_ (
    .A(_1129_),
    .B(reg_pmp_0_addr[8]),
    .S(_2403_),
    .Z(_0184_)
  );
  MUX2_X1 _9076_ (
    .A(_1175_),
    .B(reg_pmp_0_addr[9]),
    .S(_2403_),
    .Z(_0185_)
  );
  MUX2_X1 _9077_ (
    .A(_1647_),
    .B(reg_pmp_0_addr[10]),
    .S(_2403_),
    .Z(_0186_)
  );
  MUX2_X1 _9078_ (
    .A(_1698_),
    .B(reg_pmp_0_addr[11]),
    .S(_2403_),
    .Z(_0187_)
  );
  MUX2_X1 _9079_ (
    .A(_1748_),
    .B(reg_pmp_0_addr[12]),
    .S(_2403_),
    .Z(_0188_)
  );
  MUX2_X1 _9080_ (
    .A(_1790_),
    .B(reg_pmp_0_addr[13]),
    .S(_2403_),
    .Z(_0189_)
  );
  MUX2_X1 _9081_ (
    .A(_1832_),
    .B(reg_pmp_0_addr[14]),
    .S(_2403_),
    .Z(_0190_)
  );
  MUX2_X1 _9082_ (
    .A(_1880_),
    .B(reg_pmp_0_addr[15]),
    .S(_2403_),
    .Z(_0191_)
  );
  MUX2_X1 _9083_ (
    .A(_0862_),
    .B(reg_pmp_0_addr[16]),
    .S(_2403_),
    .Z(_0192_)
  );
  MUX2_X1 _9084_ (
    .A(_1926_),
    .B(reg_pmp_0_addr[17]),
    .S(_2403_),
    .Z(_0193_)
  );
  MUX2_X1 _9085_ (
    .A(_0908_),
    .B(reg_pmp_0_addr[18]),
    .S(_2403_),
    .Z(_0194_)
  );
  MUX2_X1 _9086_ (
    .A(_0967_),
    .B(reg_pmp_0_addr[19]),
    .S(_2403_),
    .Z(_0195_)
  );
  MUX2_X1 _9087_ (
    .A(_1017_),
    .B(reg_pmp_0_addr[20]),
    .S(_2403_),
    .Z(_0196_)
  );
  MUX2_X1 _9088_ (
    .A(_1968_),
    .B(reg_pmp_0_addr[21]),
    .S(_2403_),
    .Z(_0197_)
  );
  MUX2_X1 _9089_ (
    .A(_2010_),
    .B(reg_pmp_0_addr[22]),
    .S(_2403_),
    .Z(_0198_)
  );
  MUX2_X1 _9090_ (
    .A(_1071_),
    .B(reg_pmp_0_addr[23]),
    .S(_2403_),
    .Z(_0199_)
  );
  MUX2_X1 _9091_ (
    .A(_2056_),
    .B(reg_pmp_0_addr[24]),
    .S(_2403_),
    .Z(_0200_)
  );
  MUX2_X1 _9092_ (
    .A(_2102_),
    .B(reg_pmp_0_addr[25]),
    .S(_2403_),
    .Z(_0201_)
  );
  MUX2_X1 _9093_ (
    .A(_2148_),
    .B(reg_pmp_0_addr[26]),
    .S(_2403_),
    .Z(_0202_)
  );
  MUX2_X1 _9094_ (
    .A(_2195_),
    .B(reg_pmp_0_addr[27]),
    .S(_2403_),
    .Z(_0203_)
  );
  MUX2_X1 _9095_ (
    .A(_2241_),
    .B(reg_pmp_0_addr[28]),
    .S(_2403_),
    .Z(_0204_)
  );
  MUX2_X1 _9096_ (
    .A(_2285_),
    .B(reg_pmp_0_addr[29]),
    .S(_2403_),
    .Z(_0205_)
  );
  MUX2_X1 _9097_ (
    .A(reg_pmp_0_cfg_x),
    .B(_1346_),
    .S(_2288_),
    .Z(_0206_)
  );
  OR2_X1 _9098_ (
    .A1(reg_debug),
    .A2(_0005_),
    .ZN(_2404_)
  );
  AND2_X1 _9099_ (
    .A1(_0736_),
    .A2(_2404_),
    .ZN(_2405_)
  );
  INV_X1 _9100_ (
    .A(_2405_),
    .ZN(_2406_)
  );
  AND2_X1 _9101_ (
    .A1(_0800_),
    .A2(_2405_),
    .ZN(_2407_)
  );
  MUX2_X1 _9102_ (
    .A(reg_bp_0_address[0]),
    .B(_1241_),
    .S(_2407_),
    .Z(_0207_)
  );
  MUX2_X1 _9103_ (
    .A(reg_bp_0_address[1]),
    .B(_1290_),
    .S(_2407_),
    .Z(_0208_)
  );
  MUX2_X1 _9104_ (
    .A(reg_bp_0_address[2]),
    .B(_1346_),
    .S(_2407_),
    .Z(_0209_)
  );
  MUX2_X1 _9105_ (
    .A(reg_bp_0_address[3]),
    .B(_1409_),
    .S(_2407_),
    .Z(_0210_)
  );
  MUX2_X1 _9106_ (
    .A(reg_bp_0_address[4]),
    .B(_1456_),
    .S(_2407_),
    .Z(_0211_)
  );
  MUX2_X1 _9107_ (
    .A(reg_bp_0_address[5]),
    .B(_1499_),
    .S(_2407_),
    .Z(_0212_)
  );
  MUX2_X1 _9108_ (
    .A(reg_bp_0_address[6]),
    .B(_1545_),
    .S(_2407_),
    .Z(_0213_)
  );
  MUX2_X1 _9109_ (
    .A(reg_bp_0_address[7]),
    .B(_1601_),
    .S(_2407_),
    .Z(_0214_)
  );
  MUX2_X1 _9110_ (
    .A(reg_bp_0_address[8]),
    .B(_1129_),
    .S(_2407_),
    .Z(_0215_)
  );
  MUX2_X1 _9111_ (
    .A(reg_bp_0_address[9]),
    .B(_1175_),
    .S(_2407_),
    .Z(_0216_)
  );
  MUX2_X1 _9112_ (
    .A(reg_bp_0_address[10]),
    .B(_1647_),
    .S(_2407_),
    .Z(_0217_)
  );
  MUX2_X1 _9113_ (
    .A(reg_bp_0_address[11]),
    .B(_1698_),
    .S(_2407_),
    .Z(_0218_)
  );
  MUX2_X1 _9114_ (
    .A(reg_bp_0_address[12]),
    .B(_1748_),
    .S(_2407_),
    .Z(_0219_)
  );
  MUX2_X1 _9115_ (
    .A(reg_bp_0_address[13]),
    .B(_1790_),
    .S(_2407_),
    .Z(_0220_)
  );
  MUX2_X1 _9116_ (
    .A(reg_bp_0_address[14]),
    .B(_1832_),
    .S(_2407_),
    .Z(_0221_)
  );
  MUX2_X1 _9117_ (
    .A(reg_bp_0_address[15]),
    .B(_1880_),
    .S(_2407_),
    .Z(_0222_)
  );
  MUX2_X1 _9118_ (
    .A(reg_bp_0_address[16]),
    .B(_0862_),
    .S(_2407_),
    .Z(_0223_)
  );
  MUX2_X1 _9119_ (
    .A(reg_bp_0_address[17]),
    .B(_1926_),
    .S(_2407_),
    .Z(_0224_)
  );
  MUX2_X1 _9120_ (
    .A(reg_bp_0_address[18]),
    .B(_0908_),
    .S(_2407_),
    .Z(_0225_)
  );
  MUX2_X1 _9121_ (
    .A(reg_bp_0_address[19]),
    .B(_0967_),
    .S(_2407_),
    .Z(_0226_)
  );
  MUX2_X1 _9122_ (
    .A(reg_bp_0_address[20]),
    .B(_1017_),
    .S(_2407_),
    .Z(_0227_)
  );
  MUX2_X1 _9123_ (
    .A(reg_bp_0_address[21]),
    .B(_1968_),
    .S(_2407_),
    .Z(_0228_)
  );
  MUX2_X1 _9124_ (
    .A(reg_bp_0_address[22]),
    .B(_2010_),
    .S(_2407_),
    .Z(_0229_)
  );
  MUX2_X1 _9125_ (
    .A(reg_bp_0_address[23]),
    .B(_1071_),
    .S(_2407_),
    .Z(_0230_)
  );
  MUX2_X1 _9126_ (
    .A(reg_bp_0_address[24]),
    .B(_2056_),
    .S(_2407_),
    .Z(_0231_)
  );
  MUX2_X1 _9127_ (
    .A(reg_bp_0_address[25]),
    .B(_2102_),
    .S(_2407_),
    .Z(_0232_)
  );
  MUX2_X1 _9128_ (
    .A(reg_bp_0_address[26]),
    .B(_2148_),
    .S(_2407_),
    .Z(_0233_)
  );
  MUX2_X1 _9129_ (
    .A(reg_bp_0_address[27]),
    .B(_2195_),
    .S(_2407_),
    .Z(_0234_)
  );
  MUX2_X1 _9130_ (
    .A(reg_bp_0_address[28]),
    .B(_2241_),
    .S(_2407_),
    .Z(_0235_)
  );
  MUX2_X1 _9131_ (
    .A(reg_bp_0_address[29]),
    .B(_2285_),
    .S(_2407_),
    .Z(_0236_)
  );
  AND2_X1 _9132_ (
    .A1(io_rw_wdata[30]),
    .A2(_0742_),
    .ZN(_2408_)
  );
  AND2_X1 _9133_ (
    .A1(large_[56]),
    .A2(_0827_),
    .ZN(_2409_)
  );
  AND2_X1 _9134_ (
    .A1(large_1[56]),
    .A2(_0851_),
    .ZN(_2410_)
  );
  AND2_X1 _9135_ (
    .A1(reg_dscratch0[30]),
    .A2(_0797_),
    .ZN(_2411_)
  );
  AND2_X1 _9136_ (
    .A1(reg_mtval[30]),
    .A2(_0764_),
    .ZN(_2412_)
  );
  AND2_X1 _9137_ (
    .A1(reg_bp_0_address[30]),
    .A2(_0800_),
    .ZN(_2413_)
  );
  AND2_X1 _9138_ (
    .A1(reg_mepc[30]),
    .A2(_0783_),
    .ZN(_2414_)
  );
  AND2_X1 _9139_ (
    .A1(reg_dpc[30]),
    .A2(_0750_),
    .ZN(_2415_)
  );
  AND2_X1 _9140_ (
    .A1(reg_mtvec[30]),
    .A2(_0780_),
    .ZN(_2416_)
  );
  AND2_X1 _9141_ (
    .A1(reg_mcause[30]),
    .A2(_0834_),
    .ZN(_2417_)
  );
  AND2_X1 _9142_ (
    .A1(reg_mscratch[30]),
    .A2(_0767_),
    .ZN(_2418_)
  );
  OR2_X1 _9143_ (
    .A1(_1057_),
    .A2(_1086_),
    .ZN(_2419_)
  );
  OR2_X1 _9144_ (
    .A1(_2411_),
    .A2(_2415_),
    .ZN(_2420_)
  );
  OR2_X1 _9145_ (
    .A1(_2413_),
    .A2(_2420_),
    .ZN(_2421_)
  );
  AND2_X1 _9146_ (
    .A1(large_[24]),
    .A2(_0857_),
    .ZN(_2422_)
  );
  OR2_X1 _9147_ (
    .A1(_2412_),
    .A2(_2414_),
    .ZN(_2423_)
  );
  OR2_X1 _9148_ (
    .A1(_2422_),
    .A2(_2423_),
    .ZN(_2424_)
  );
  OR2_X1 _9149_ (
    .A1(_2409_),
    .A2(_2424_),
    .ZN(_2425_)
  );
  OR2_X1 _9150_ (
    .A1(_2421_),
    .A2(_2425_),
    .ZN(_2426_)
  );
  AND2_X1 _9151_ (
    .A1(large_1[24]),
    .A2(_0859_),
    .ZN(_2427_)
  );
  OR2_X1 _9152_ (
    .A1(_2417_),
    .A2(_2418_),
    .ZN(_2428_)
  );
  OR2_X1 _9153_ (
    .A1(_2427_),
    .A2(_2428_),
    .ZN(_2429_)
  );
  OR2_X1 _9154_ (
    .A1(_2416_),
    .A2(_2429_),
    .ZN(_2430_)
  );
  OR2_X1 _9155_ (
    .A1(_2410_),
    .A2(_2419_),
    .ZN(_2431_)
  );
  OR2_X1 _9156_ (
    .A1(_2430_),
    .A2(_2431_),
    .ZN(_2432_)
  );
  OR2_X1 _9157_ (
    .A1(_2426_),
    .A2(_2432_),
    .ZN(io_rw_rdata[30])
  );
  AND2_X1 _9158_ (
    .A1(io_rw_cmd[1]),
    .A2(_0707_),
    .ZN(_2433_)
  );
  AND2_X1 _9159_ (
    .A1(io_rw_rdata[30]),
    .A2(_2433_),
    .ZN(_2434_)
  );
  OR2_X1 _9160_ (
    .A1(_2408_),
    .A2(_2434_),
    .ZN(_2435_)
  );
  MUX2_X1 _9161_ (
    .A(reg_bp_0_address[30]),
    .B(_2435_),
    .S(_2407_),
    .Z(_0237_)
  );
  MUX2_X1 _9162_ (
    .A(reg_bp_0_address[31]),
    .B(_2365_),
    .S(_2407_),
    .Z(_0238_)
  );
  OR2_X1 _9163_ (
    .A1(reg_pmp_0_cfg_a[0]),
    .A2(_2288_),
    .ZN(_2436_)
  );
  AND2_X1 _9164_ (
    .A1(_0654_),
    .A2(_2436_),
    .ZN(_2437_)
  );
  OR2_X1 _9165_ (
    .A1(_1409_),
    .A2(_2289_),
    .ZN(_2438_)
  );
  AND2_X1 _9166_ (
    .A1(_2437_),
    .A2(_2438_),
    .ZN(_0239_)
  );
  OR2_X1 _9167_ (
    .A1(reg_pmp_0_cfg_a[1]),
    .A2(_2288_),
    .ZN(_2439_)
  );
  AND2_X1 _9168_ (
    .A1(_0654_),
    .A2(_2439_),
    .ZN(_2440_)
  );
  OR2_X1 _9169_ (
    .A1(_1456_),
    .A2(_2289_),
    .ZN(_2441_)
  );
  AND2_X1 _9170_ (
    .A1(_2440_),
    .A2(_2441_),
    .ZN(_0240_)
  );
  OR2_X1 _9171_ (
    .A1(reg_pmp_0_cfg_l),
    .A2(_2288_),
    .ZN(_2442_)
  );
  AND2_X1 _9172_ (
    .A1(_0654_),
    .A2(_2442_),
    .ZN(_2443_)
  );
  OR2_X1 _9173_ (
    .A1(_1601_),
    .A2(_2289_),
    .ZN(_2444_)
  );
  AND2_X1 _9174_ (
    .A1(_2443_),
    .A2(_2444_),
    .ZN(_0241_)
  );
  AND2_X1 _9175_ (
    .A1(_1058_),
    .A2(_2405_),
    .ZN(_2445_)
  );
  OR2_X1 _9176_ (
    .A1(_1059_),
    .A2(_2406_),
    .ZN(_2446_)
  );
  MUX2_X1 _9177_ (
    .A(reg_bp_0_control_tmatch[0]),
    .B(_1601_),
    .S(_2445_),
    .Z(_0242_)
  );
  MUX2_X1 _9178_ (
    .A(reg_bp_0_control_tmatch[1]),
    .B(_1129_),
    .S(_2445_),
    .Z(_0243_)
  );
  OR2_X1 _9179_ (
    .A1(_1241_),
    .A2(_2446_),
    .ZN(_2447_)
  );
  OR2_X1 _9180_ (
    .A1(reg_bp_0_control_r),
    .A2(_2445_),
    .ZN(_2448_)
  );
  AND2_X1 _9181_ (
    .A1(_0654_),
    .A2(_2448_),
    .ZN(_2449_)
  );
  AND2_X1 _9182_ (
    .A1(_2447_),
    .A2(_2449_),
    .ZN(_0244_)
  );
  OR2_X1 _9183_ (
    .A1(_1290_),
    .A2(_2446_),
    .ZN(_2450_)
  );
  OR2_X1 _9184_ (
    .A1(reg_bp_0_control_w),
    .A2(_2445_),
    .ZN(_2451_)
  );
  AND2_X1 _9185_ (
    .A1(_0654_),
    .A2(_2451_),
    .ZN(_2452_)
  );
  AND2_X1 _9186_ (
    .A1(_2450_),
    .A2(_2452_),
    .ZN(_0245_)
  );
  OR2_X1 _9187_ (
    .A1(_1346_),
    .A2(_2446_),
    .ZN(_2453_)
  );
  OR2_X1 _9188_ (
    .A1(reg_bp_0_control_x),
    .A2(_2445_),
    .ZN(_2454_)
  );
  AND2_X1 _9189_ (
    .A1(_0654_),
    .A2(_2454_),
    .ZN(_2455_)
  );
  AND2_X1 _9190_ (
    .A1(_2453_),
    .A2(_2455_),
    .ZN(_0246_)
  );
  AND2_X1 _9191_ (
    .A1(reg_dcsr_step),
    .A2(_io_decode_0_read_illegal_T_15),
    .ZN(io_singleStep)
  );
  INV_X1 _9192_ (
    .A(io_singleStep),
    .ZN(_2456_)
  );
  OR2_X1 _9193_ (
    .A1(io_rw_addr[8]),
    .A2(io_rw_addr[9]),
    .ZN(_2457_)
  );
  OR2_X1 _9194_ (
    .A1(_0722_),
    .A2(_2457_),
    .ZN(_2458_)
  );
  OR2_X1 _9195_ (
    .A1(_0774_),
    .A2(_2458_),
    .ZN(_2459_)
  );
  INV_X1 _9196_ (
    .A(_2459_),
    .ZN(_2460_)
  );
  AND2_X1 _9197_ (
    .A1(_0753_),
    .A2(_2460_),
    .ZN(_2461_)
  );
  AND2_X1 _9198_ (
    .A1(_0909_),
    .A2(_2461_),
    .ZN(_2462_)
  );
  INV_X1 _9199_ (
    .A(_2462_),
    .ZN(_2463_)
  );
  OR2_X1 _9200_ (
    .A1(_0721_),
    .A2(_2459_),
    .ZN(_2464_)
  );
  OR2_X1 _9201_ (
    .A1(_0910_),
    .A2(_2464_),
    .ZN(_2465_)
  );
  INV_X1 _9202_ (
    .A(_2465_),
    .ZN(_2466_)
  );
  AND2_X1 _9203_ (
    .A1(_2463_),
    .A2(_2465_),
    .ZN(_2467_)
  );
  INV_X1 _9204_ (
    .A(_2467_),
    .ZN(_2468_)
  );
  AND2_X1 _9205_ (
    .A1(_0715_),
    .A2(_2467_),
    .ZN(_2469_)
  );
  INV_X1 _9206_ (
    .A(_2469_),
    .ZN(io_trace_0_exception)
  );
  OR2_X1 _9207_ (
    .A1(io_retire),
    .A2(io_trace_0_exception),
    .ZN(io_trace_0_valid)
  );
  OR2_X1 _9208_ (
    .A1(reg_singleStepped),
    .A2(io_trace_0_valid),
    .ZN(_2470_)
  );
  AND2_X1 _9209_ (
    .A1(io_singleStep),
    .A2(_2470_),
    .ZN(_0247_)
  );
  AND2_X1 _9210_ (
    .A1(reg_bp_0_control_action),
    .A2(_2446_),
    .ZN(_2471_)
  );
  AND2_X1 _9211_ (
    .A1(reg_bp_0_control_dmode),
    .A2(io_rw_cmd[1]),
    .ZN(_2472_)
  );
  OR2_X1 _9212_ (
    .A1(io_rw_wdata[27]),
    .A2(_2472_),
    .ZN(_2473_)
  );
  AND2_X1 _9213_ (
    .A1(reg_debug),
    .A2(_2194_),
    .ZN(_2474_)
  );
  AND2_X1 _9214_ (
    .A1(_2473_),
    .A2(_2474_),
    .ZN(_2475_)
  );
  AND2_X1 _9215_ (
    .A1(_2445_),
    .A2(_2475_),
    .ZN(_2476_)
  );
  AND2_X1 _9216_ (
    .A1(reg_bp_0_control_action),
    .A2(io_rw_cmd[1]),
    .ZN(_2477_)
  );
  MUX2_X1 _9217_ (
    .A(_2477_),
    .B(_0742_),
    .S(io_rw_wdata[12]),
    .Z(_2478_)
  );
  AND2_X1 _9218_ (
    .A1(_2476_),
    .A2(_2478_),
    .ZN(_2479_)
  );
  OR2_X1 _9219_ (
    .A1(_2471_),
    .A2(_2479_),
    .ZN(_2480_)
  );
  AND2_X1 _9220_ (
    .A1(_0654_),
    .A2(_2480_),
    .ZN(_0248_)
  );
  MUX2_X1 _9221_ (
    .A(reg_bp_0_control_dmode),
    .B(_2475_),
    .S(_2445_),
    .Z(_2481_)
  );
  AND2_X1 _9222_ (
    .A1(_0654_),
    .A2(_2481_),
    .ZN(_0249_)
  );
  AND2_X1 _9223_ (
    .A1(_0736_),
    .A2(_0797_),
    .ZN(_2482_)
  );
  MUX2_X1 _9224_ (
    .A(reg_dscratch0[0]),
    .B(_1241_),
    .S(_2482_),
    .Z(_0250_)
  );
  MUX2_X1 _9225_ (
    .A(reg_dscratch0[1]),
    .B(_1290_),
    .S(_2482_),
    .Z(_0251_)
  );
  MUX2_X1 _9226_ (
    .A(reg_dscratch0[2]),
    .B(_1346_),
    .S(_2482_),
    .Z(_0252_)
  );
  MUX2_X1 _9227_ (
    .A(reg_dscratch0[3]),
    .B(_1409_),
    .S(_2482_),
    .Z(_0253_)
  );
  MUX2_X1 _9228_ (
    .A(reg_dscratch0[4]),
    .B(_1456_),
    .S(_2482_),
    .Z(_0254_)
  );
  MUX2_X1 _9229_ (
    .A(reg_dscratch0[5]),
    .B(_1499_),
    .S(_2482_),
    .Z(_0255_)
  );
  MUX2_X1 _9230_ (
    .A(reg_dscratch0[6]),
    .B(_1545_),
    .S(_2482_),
    .Z(_0256_)
  );
  MUX2_X1 _9231_ (
    .A(reg_dscratch0[7]),
    .B(_1601_),
    .S(_2482_),
    .Z(_0257_)
  );
  MUX2_X1 _9232_ (
    .A(reg_dscratch0[8]),
    .B(_1129_),
    .S(_2482_),
    .Z(_0258_)
  );
  MUX2_X1 _9233_ (
    .A(reg_dscratch0[9]),
    .B(_1175_),
    .S(_2482_),
    .Z(_0259_)
  );
  MUX2_X1 _9234_ (
    .A(reg_dscratch0[10]),
    .B(_1647_),
    .S(_2482_),
    .Z(_0260_)
  );
  MUX2_X1 _9235_ (
    .A(reg_dscratch0[11]),
    .B(_1698_),
    .S(_2482_),
    .Z(_0261_)
  );
  MUX2_X1 _9236_ (
    .A(reg_dscratch0[12]),
    .B(_1748_),
    .S(_2482_),
    .Z(_0262_)
  );
  MUX2_X1 _9237_ (
    .A(reg_dscratch0[13]),
    .B(_1790_),
    .S(_2482_),
    .Z(_0263_)
  );
  MUX2_X1 _9238_ (
    .A(reg_dscratch0[14]),
    .B(_1832_),
    .S(_2482_),
    .Z(_0264_)
  );
  MUX2_X1 _9239_ (
    .A(reg_dscratch0[15]),
    .B(_1880_),
    .S(_2482_),
    .Z(_0265_)
  );
  MUX2_X1 _9240_ (
    .A(reg_dscratch0[16]),
    .B(_0862_),
    .S(_2482_),
    .Z(_0266_)
  );
  MUX2_X1 _9241_ (
    .A(reg_dscratch0[17]),
    .B(_1926_),
    .S(_2482_),
    .Z(_0267_)
  );
  MUX2_X1 _9242_ (
    .A(reg_dscratch0[18]),
    .B(_0908_),
    .S(_2482_),
    .Z(_0268_)
  );
  MUX2_X1 _9243_ (
    .A(reg_dscratch0[19]),
    .B(_0967_),
    .S(_2482_),
    .Z(_0269_)
  );
  MUX2_X1 _9244_ (
    .A(reg_dscratch0[20]),
    .B(_1017_),
    .S(_2482_),
    .Z(_0270_)
  );
  MUX2_X1 _9245_ (
    .A(reg_dscratch0[21]),
    .B(_1968_),
    .S(_2482_),
    .Z(_0271_)
  );
  MUX2_X1 _9246_ (
    .A(reg_dscratch0[22]),
    .B(_2010_),
    .S(_2482_),
    .Z(_0272_)
  );
  MUX2_X1 _9247_ (
    .A(reg_dscratch0[23]),
    .B(_1071_),
    .S(_2482_),
    .Z(_0273_)
  );
  MUX2_X1 _9248_ (
    .A(reg_dscratch0[24]),
    .B(_2056_),
    .S(_2482_),
    .Z(_0274_)
  );
  MUX2_X1 _9249_ (
    .A(reg_dscratch0[25]),
    .B(_2102_),
    .S(_2482_),
    .Z(_0275_)
  );
  MUX2_X1 _9250_ (
    .A(reg_dscratch0[26]),
    .B(_2148_),
    .S(_2482_),
    .Z(_0276_)
  );
  MUX2_X1 _9251_ (
    .A(reg_dscratch0[27]),
    .B(_2195_),
    .S(_2482_),
    .Z(_0277_)
  );
  MUX2_X1 _9252_ (
    .A(reg_dscratch0[28]),
    .B(_2241_),
    .S(_2482_),
    .Z(_0278_)
  );
  MUX2_X1 _9253_ (
    .A(reg_dscratch0[29]),
    .B(_2285_),
    .S(_2482_),
    .Z(_0279_)
  );
  MUX2_X1 _9254_ (
    .A(reg_dscratch0[30]),
    .B(_2435_),
    .S(_2482_),
    .Z(_0280_)
  );
  MUX2_X1 _9255_ (
    .A(reg_dscratch0[31]),
    .B(_2365_),
    .S(_2482_),
    .Z(_0281_)
  );
  AND2_X1 _9256_ (
    .A1(io_cause[5]),
    .A2(_2467_),
    .ZN(_2483_)
  );
  INV_X1 _9257_ (
    .A(_2483_),
    .ZN(_2484_)
  );
  AND2_X1 _9258_ (
    .A1(io_cause[7]),
    .A2(_2467_),
    .ZN(_2485_)
  );
  AND2_X1 _9259_ (
    .A1(io_cause[6]),
    .A2(_2467_),
    .ZN(_2486_)
  );
  OR2_X1 _9260_ (
    .A1(_2485_),
    .A2(_2486_),
    .ZN(_2487_)
  );
  INV_X1 _9261_ (
    .A(_2487_),
    .ZN(_2488_)
  );
  AND2_X1 _9262_ (
    .A1(_2484_),
    .A2(_2488_),
    .ZN(_2489_)
  );
  OR2_X1 _9263_ (
    .A1(io_cause[0]),
    .A2(_2468_),
    .ZN(_2490_)
  );
  INV_X1 _9264_ (
    .A(_2490_),
    .ZN(_2491_)
  );
  AND2_X1 _9265_ (
    .A1(io_cause[2]),
    .A2(_2467_),
    .ZN(_2492_)
  );
  AND2_X1 _9266_ (
    .A1(io_cause[3]),
    .A2(_2465_),
    .ZN(_2493_)
  );
  AND2_X1 _9267_ (
    .A1(io_cause[1]),
    .A2(_0709_),
    .ZN(_2494_)
  );
  AND2_X1 _9268_ (
    .A1(_2493_),
    .A2(_2494_),
    .ZN(_2495_)
  );
  AND2_X1 _9269_ (
    .A1(_2492_),
    .A2(_2495_),
    .ZN(_2496_)
  );
  OR2_X1 _9270_ (
    .A1(_2462_),
    .A2(_2493_),
    .ZN(_2497_)
  );
  AND2_X1 _9271_ (
    .A1(_2491_),
    .A2(_2496_),
    .ZN(_2498_)
  );
  AND2_X1 _9272_ (
    .A1(_2489_),
    .A2(_2498_),
    .ZN(_2499_)
  );
  INV_X1 _9273_ (
    .A(_2499_),
    .ZN(_2500_)
  );
  OR2_X1 _9274_ (
    .A1(reg_singleStepped),
    .A2(reg_debug),
    .ZN(_2501_)
  );
  AND2_X1 _9275_ (
    .A1(reg_dcsr_ebreakm),
    .A2(_2466_),
    .ZN(_2502_)
  );
  OR2_X1 _9276_ (
    .A1(_2501_),
    .A2(_2502_),
    .ZN(_2503_)
  );
  INV_X1 _9277_ (
    .A(_2503_),
    .ZN(_2504_)
  );
  AND2_X1 _9278_ (
    .A1(_2500_),
    .A2(_2504_),
    .ZN(_2505_)
  );
  OR2_X1 _9279_ (
    .A1(_2499_),
    .A2(_2503_),
    .ZN(_2506_)
  );
  OR2_X1 _9280_ (
    .A1(_2469_),
    .A2(_2506_),
    .ZN(_2507_)
  );
  OR2_X1 _9281_ (
    .A1(reg_debug),
    .A2(io_trace_0_exception),
    .ZN(_2508_)
  );
  OR2_X1 _9282_ (
    .A1(_0716_),
    .A2(_0776_),
    .ZN(_2509_)
  );
  AND2_X1 _9283_ (
    .A1(_0747_),
    .A2(_2509_),
    .ZN(_2510_)
  );
  OR2_X1 _9284_ (
    .A1(_0910_),
    .A2(_2510_),
    .ZN(_2511_)
  );
  INV_X1 _9285_ (
    .A(_2511_),
    .ZN(_2512_)
  );
  AND2_X1 _9286_ (
    .A1(io_rw_addr[10]),
    .A2(io_rw_addr[7]),
    .ZN(_2513_)
  );
  INV_X1 _9287_ (
    .A(_2513_),
    .ZN(_2514_)
  );
  AND2_X1 _9288_ (
    .A1(_2512_),
    .A2(_2513_),
    .ZN(_2515_)
  );
  OR2_X1 _9289_ (
    .A1(reset),
    .A2(_2515_),
    .ZN(_2516_)
  );
  INV_X1 _9290_ (
    .A(_2516_),
    .ZN(_2517_)
  );
  AND2_X1 _9291_ (
    .A1(_2508_),
    .A2(_2517_),
    .ZN(_2518_)
  );
  AND2_X1 _9292_ (
    .A1(_2507_),
    .A2(_2518_),
    .ZN(_0282_)
  );
  AND2_X1 _9293_ (
    .A1(_2512_),
    .A2(_2514_),
    .ZN(_2519_)
  );
  INV_X1 _9294_ (
    .A(_2519_),
    .ZN(_2520_)
  );
  AND2_X1 _9295_ (
    .A1(reg_mstatus_mie),
    .A2(_2520_),
    .ZN(_2521_)
  );
  AND2_X1 _9296_ (
    .A1(_2507_),
    .A2(_2521_),
    .ZN(_2522_)
  );
  AND2_X1 _9297_ (
    .A1(_0736_),
    .A2(_1374_),
    .ZN(_2523_)
  );
  OR2_X1 _9298_ (
    .A1(_0737_),
    .A2(_1375_),
    .ZN(_2524_)
  );
  AND2_X1 _9299_ (
    .A1(reg_mstatus_mpie),
    .A2(_2519_),
    .ZN(_2525_)
  );
  OR2_X1 _9300_ (
    .A1(_2519_),
    .A2(_2523_),
    .ZN(_2526_)
  );
  OR2_X1 _9301_ (
    .A1(_2523_),
    .A2(_2525_),
    .ZN(_2527_)
  );
  OR2_X1 _9302_ (
    .A1(_2522_),
    .A2(_2527_),
    .ZN(_2528_)
  );
  OR2_X1 _9303_ (
    .A1(_1409_),
    .A2(_2524_),
    .ZN(_2529_)
  );
  AND2_X1 _9304_ (
    .A1(_0654_),
    .A2(_2529_),
    .ZN(_2530_)
  );
  AND2_X1 _9305_ (
    .A1(_2528_),
    .A2(_2530_),
    .ZN(_0283_)
  );
  AND2_X1 _9306_ (
    .A1(_0736_),
    .A2(_1086_),
    .ZN(_2531_)
  );
  OR2_X1 _9307_ (
    .A1(_0737_),
    .A2(_1087_),
    .ZN(_2532_)
  );
  OR2_X1 _9308_ (
    .A1(_1346_),
    .A2(_2532_),
    .ZN(_2533_)
  );
  OR2_X1 _9309_ (
    .A1(reg_dcsr_step),
    .A2(_2531_),
    .ZN(_2534_)
  );
  AND2_X1 _9310_ (
    .A1(_0654_),
    .A2(_2534_),
    .ZN(_2535_)
  );
  AND2_X1 _9311_ (
    .A1(_2533_),
    .A2(_2535_),
    .ZN(_0284_)
  );
  AND2_X1 _9312_ (
    .A1(_io_decode_0_read_illegal_T_15),
    .A2(io_trace_0_exception),
    .ZN(_2536_)
  );
  AND2_X1 _9313_ (
    .A1(_2506_),
    .A2(_2536_),
    .ZN(_2537_)
  );
  INV_X1 _9314_ (
    .A(_2537_),
    .ZN(_2538_)
  );
  AND2_X1 _9315_ (
    .A1(io_cause[31]),
    .A2(_2467_),
    .ZN(_2539_)
  );
  OR2_X1 _9316_ (
    .A1(_2500_),
    .A2(_2539_),
    .ZN(_2540_)
  );
  AND2_X1 _9317_ (
    .A1(_0653_),
    .A2(_2540_),
    .ZN(_2541_)
  );
  MUX2_X1 _9318_ (
    .A(reg_dcsr_cause[0]),
    .B(_2541_),
    .S(_2537_),
    .Z(_2542_)
  );
  AND2_X1 _9319_ (
    .A1(_0654_),
    .A2(_2542_),
    .ZN(_0285_)
  );
  AND2_X1 _9320_ (
    .A1(reg_dcsr_cause[1]),
    .A2(_2538_),
    .ZN(_2543_)
  );
  AND2_X1 _9321_ (
    .A1(_2499_),
    .A2(_2536_),
    .ZN(_2544_)
  );
  AND2_X1 _9322_ (
    .A1(_0653_),
    .A2(_2544_),
    .ZN(_2545_)
  );
  OR2_X1 _9323_ (
    .A1(_2543_),
    .A2(_2545_),
    .ZN(_2546_)
  );
  AND2_X1 _9324_ (
    .A1(_0654_),
    .A2(_2546_),
    .ZN(_0286_)
  );
  MUX2_X1 _9325_ (
    .A(reg_dcsr_cause[2]),
    .B(reg_singleStepped),
    .S(_2537_),
    .Z(_2547_)
  );
  AND2_X1 _9326_ (
    .A1(_0654_),
    .A2(_2547_),
    .ZN(_0287_)
  );
  OR2_X1 _9327_ (
    .A1(_1880_),
    .A2(_2532_),
    .ZN(_2548_)
  );
  OR2_X1 _9328_ (
    .A1(reg_dcsr_ebreakm),
    .A2(_2531_),
    .ZN(_2549_)
  );
  AND2_X1 _9329_ (
    .A1(_0654_),
    .A2(_2549_),
    .ZN(_2550_)
  );
  AND2_X1 _9330_ (
    .A1(_2548_),
    .A2(_2550_),
    .ZN(_0288_)
  );
  MUX2_X1 _9331_ (
    .A(reg_mstatus_mie),
    .B(reg_mstatus_mpie),
    .S(_2507_),
    .Z(_2551_)
  );
  OR2_X1 _9332_ (
    .A1(_2526_),
    .A2(_2551_),
    .ZN(_2552_)
  );
  OR2_X1 _9333_ (
    .A1(_1601_),
    .A2(_2524_),
    .ZN(_2553_)
  );
  AND2_X1 _9334_ (
    .A1(_0654_),
    .A2(_2553_),
    .ZN(_2554_)
  );
  AND2_X1 _9335_ (
    .A1(_2552_),
    .A2(_2554_),
    .ZN(_0289_)
  );
  AND2_X1 _9336_ (
    .A1(_0736_),
    .A2(_1237_),
    .ZN(_2555_)
  );
  OR2_X1 _9337_ (
    .A1(_0737_),
    .A2(_1238_),
    .ZN(_2556_)
  );
  OR2_X1 _9338_ (
    .A1(reg_mcountinhibit[0]),
    .A2(_2555_),
    .ZN(_2557_)
  );
  AND2_X1 _9339_ (
    .A1(_0654_),
    .A2(_2557_),
    .ZN(_2558_)
  );
  OR2_X1 _9340_ (
    .A1(_1241_),
    .A2(_2556_),
    .ZN(_2559_)
  );
  AND2_X1 _9341_ (
    .A1(_2558_),
    .A2(_2559_),
    .ZN(_0290_)
  );
  OR2_X1 _9342_ (
    .A1(reg_mcountinhibit[2]),
    .A2(_2555_),
    .ZN(_2560_)
  );
  AND2_X1 _9343_ (
    .A1(_0654_),
    .A2(_2560_),
    .ZN(_2561_)
  );
  OR2_X1 _9344_ (
    .A1(_1346_),
    .A2(_2556_),
    .ZN(_2562_)
  );
  AND2_X1 _9345_ (
    .A1(_2561_),
    .A2(_2562_),
    .ZN(_0291_)
  );
  OR2_X1 _9346_ (
    .A1(reg_dcsr_step),
    .A2(io_rw_addr[9]),
    .ZN(_2563_)
  );
  INV_X1 _9347_ (
    .A(_2563_),
    .ZN(_2564_)
  );
  AND2_X1 _9348_ (
    .A1(_io_decode_0_read_illegal_T_15),
    .A2(_2564_),
    .ZN(_2565_)
  );
  AND2_X1 _9349_ (
    .A1(_0909_),
    .A2(_2565_),
    .ZN(_2566_)
  );
  AND2_X1 _9350_ (
    .A1(_0725_),
    .A2(_2566_),
    .ZN(_2567_)
  );
  OR2_X1 _9351_ (
    .A1(reg_wfi),
    .A2(_2567_),
    .ZN(_2568_)
  );
  OR2_X1 _9352_ (
    .A1(reset),
    .A2(io_interrupts_debug),
    .ZN(_2569_)
  );
  AND2_X1 _9353_ (
    .A1(reg_mie[7]),
    .A2(io_interrupts_mtip),
    .ZN(_2570_)
  );
  AND2_X1 _9354_ (
    .A1(reg_mie[3]),
    .A2(io_interrupts_msip),
    .ZN(_2571_)
  );
  AND2_X1 _9355_ (
    .A1(reg_mie[11]),
    .A2(io_interrupts_meip),
    .ZN(_2572_)
  );
  OR2_X1 _9356_ (
    .A1(_2571_),
    .A2(_2572_),
    .ZN(_2573_)
  );
  INV_X1 _9357_ (
    .A(_2573_),
    .ZN(_2574_)
  );
  OR2_X1 _9358_ (
    .A1(_2570_),
    .A2(_2573_),
    .ZN(_2575_)
  );
  OR2_X1 _9359_ (
    .A1(_2569_),
    .A2(_2575_),
    .ZN(_2576_)
  );
  INV_X1 _9360_ (
    .A(_2576_),
    .ZN(_2577_)
  );
  AND2_X1 _9361_ (
    .A1(_2568_),
    .A2(_2577_),
    .ZN(_2578_)
  );
  AND2_X1 _9362_ (
    .A1(_2469_),
    .A2(_2578_),
    .ZN(_0292_)
  );
  MUX2_X1 _9363_ (
    .A(io_gva),
    .B(reg_mstatus_gva),
    .S(_2507_),
    .Z(_2579_)
  );
  AND2_X1 _9364_ (
    .A1(_0654_),
    .A2(_2579_),
    .ZN(_0293_)
  );
  AND2_X1 _9365_ (
    .A1(large_1[17]),
    .A2(large_1[16]),
    .ZN(_2580_)
  );
  AND2_X1 _9366_ (
    .A1(large_1[21]),
    .A2(large_1[15]),
    .ZN(_2581_)
  );
  AND2_X1 _9367_ (
    .A1(large_1[20]),
    .A2(_2581_),
    .ZN(_2582_)
  );
  AND2_X1 _9368_ (
    .A1(large_1[19]),
    .A2(large_1[18]),
    .ZN(_2583_)
  );
  AND2_X1 _9369_ (
    .A1(_2580_),
    .A2(_2583_),
    .ZN(_2584_)
  );
  AND2_X1 _9370_ (
    .A1(_2582_),
    .A2(_2584_),
    .ZN(_2585_)
  );
  AND2_X1 _9371_ (
    .A1(large_1[22]),
    .A2(_2585_),
    .ZN(_2586_)
  );
  INV_X1 _9372_ (
    .A(_2586_),
    .ZN(_2587_)
  );
  AND2_X1 _9373_ (
    .A1(large_1[23]),
    .A2(_2586_),
    .ZN(_2588_)
  );
  OR2_X1 _9374_ (
    .A1(_0626_),
    .A2(_2587_),
    .ZN(_2589_)
  );
  AND2_X1 _9375_ (
    .A1(large_1[13]),
    .A2(large_1[12]),
    .ZN(_2590_)
  );
  INV_X1 _9376_ (
    .A(_2590_),
    .ZN(_2591_)
  );
  AND2_X1 _9377_ (
    .A1(large_1[14]),
    .A2(_2590_),
    .ZN(_2592_)
  );
  OR2_X1 _9378_ (
    .A1(_0629_),
    .A2(_2591_),
    .ZN(_2593_)
  );
  AND2_X1 _9379_ (
    .A1(large_1[8]),
    .A2(large_1[7]),
    .ZN(_2594_)
  );
  INV_X1 _9380_ (
    .A(_2594_),
    .ZN(_2595_)
  );
  AND2_X1 _9381_ (
    .A1(large_1[9]),
    .A2(_2594_),
    .ZN(_2596_)
  );
  OR2_X1 _9382_ (
    .A1(_0632_),
    .A2(_2595_),
    .ZN(_2597_)
  );
  AND2_X1 _9383_ (
    .A1(large_1[4]),
    .A2(large_1[3]),
    .ZN(_2598_)
  );
  AND2_X1 _9384_ (
    .A1(large_1[3]),
    .A2(large_1[2]),
    .ZN(_2599_)
  );
  AND2_X1 _9385_ (
    .A1(large_1[5]),
    .A2(large_1[4]),
    .ZN(_2600_)
  );
  AND2_X1 _9386_ (
    .A1(_2599_),
    .A2(_2600_),
    .ZN(_2601_)
  );
  AND2_X1 _9387_ (
    .A1(large_1[6]),
    .A2(_2601_),
    .ZN(_2602_)
  );
  OR2_X1 _9388_ (
    .A1(reg_wfi),
    .A2(io_status_cease_r),
    .ZN(io_csr_stall)
  );
  INV_X1 _9389_ (
    .A(io_csr_stall),
    .ZN(_2603_)
  );
  AND2_X1 _9390_ (
    .A1(small_1[0]),
    .A2(_2603_),
    .ZN(_2604_)
  );
  OR2_X1 _9391_ (
    .A1(_0641_),
    .A2(io_csr_stall),
    .ZN(_2605_)
  );
  AND2_X1 _9392_ (
    .A1(small_1[1]),
    .A2(_2604_),
    .ZN(_2606_)
  );
  OR2_X1 _9393_ (
    .A1(_0640_),
    .A2(_2605_),
    .ZN(_2607_)
  );
  AND2_X1 _9394_ (
    .A1(small_1[2]),
    .A2(_2606_),
    .ZN(_2608_)
  );
  OR2_X1 _9395_ (
    .A1(_0639_),
    .A2(_2607_),
    .ZN(_2609_)
  );
  AND2_X1 _9396_ (
    .A1(small_1[3]),
    .A2(_2608_),
    .ZN(_2610_)
  );
  OR2_X1 _9397_ (
    .A1(_0638_),
    .A2(_2609_),
    .ZN(_2611_)
  );
  AND2_X1 _9398_ (
    .A1(small_1[4]),
    .A2(_2610_),
    .ZN(_2612_)
  );
  OR2_X1 _9399_ (
    .A1(_0637_),
    .A2(_2611_),
    .ZN(_2613_)
  );
  AND2_X1 _9400_ (
    .A1(small_1[5]),
    .A2(_T_15),
    .ZN(_2614_)
  );
  AND2_X1 _9401_ (
    .A1(_2612_),
    .A2(_2614_),
    .ZN(_2615_)
  );
  AND2_X1 _9402_ (
    .A1(large_1[0]),
    .A2(_2615_),
    .ZN(_2616_)
  );
  AND2_X1 _9403_ (
    .A1(large_1[1]),
    .A2(_2616_),
    .ZN(_2617_)
  );
  AND2_X1 _9404_ (
    .A1(_2602_),
    .A2(_2617_),
    .ZN(_2618_)
  );
  AND2_X1 _9405_ (
    .A1(_2596_),
    .A2(_2618_),
    .ZN(_2619_)
  );
  AND2_X1 _9406_ (
    .A1(large_1[10]),
    .A2(_2619_),
    .ZN(_2620_)
  );
  AND2_X1 _9407_ (
    .A1(large_1[11]),
    .A2(_2620_),
    .ZN(_2621_)
  );
  AND2_X1 _9408_ (
    .A1(_2592_),
    .A2(_2621_),
    .ZN(_2622_)
  );
  AND2_X1 _9409_ (
    .A1(_2588_),
    .A2(_2622_),
    .ZN(_2623_)
  );
  AND2_X1 _9410_ (
    .A1(small_1[5]),
    .A2(_2612_),
    .ZN(_2624_)
  );
  OR2_X1 _9411_ (
    .A1(_0636_),
    .A2(_2613_),
    .ZN(_2625_)
  );
  AND2_X1 _9412_ (
    .A1(_T_15),
    .A2(_2624_),
    .ZN(_2626_)
  );
  OR2_X1 _9413_ (
    .A1(_0711_),
    .A2(_2625_),
    .ZN(_2627_)
  );
  AND2_X1 _9414_ (
    .A1(large_1[0]),
    .A2(_2626_),
    .ZN(_2628_)
  );
  AND2_X1 _9415_ (
    .A1(large_1[1]),
    .A2(_2628_),
    .ZN(_2629_)
  );
  AND2_X1 _9416_ (
    .A1(_2602_),
    .A2(_2629_),
    .ZN(_2630_)
  );
  AND2_X1 _9417_ (
    .A1(_2596_),
    .A2(_2630_),
    .ZN(_2631_)
  );
  AND2_X1 _9418_ (
    .A1(large_1[10]),
    .A2(_2631_),
    .ZN(_2632_)
  );
  AND2_X1 _9419_ (
    .A1(large_1[11]),
    .A2(_2632_),
    .ZN(_2633_)
  );
  AND2_X1 _9420_ (
    .A1(_2592_),
    .A2(_2633_),
    .ZN(_2634_)
  );
  AND2_X1 _9421_ (
    .A1(large_1[25]),
    .A2(large_1[24]),
    .ZN(_2635_)
  );
  AND2_X1 _9422_ (
    .A1(large_1[1]),
    .A2(large_1[0]),
    .ZN(_2636_)
  );
  AND2_X1 _9423_ (
    .A1(_2599_),
    .A2(_2636_),
    .ZN(_2637_)
  );
  INV_X1 _9424_ (
    .A(_2637_),
    .ZN(_2638_)
  );
  AND2_X1 _9425_ (
    .A1(large_1[6]),
    .A2(_2600_),
    .ZN(_2639_)
  );
  INV_X1 _9426_ (
    .A(_2639_),
    .ZN(_2640_)
  );
  AND2_X1 _9427_ (
    .A1(_2626_),
    .A2(_2639_),
    .ZN(_2641_)
  );
  OR2_X1 _9428_ (
    .A1(_2627_),
    .A2(_2640_),
    .ZN(_2642_)
  );
  AND2_X1 _9429_ (
    .A1(_2637_),
    .A2(_2641_),
    .ZN(_2643_)
  );
  OR2_X1 _9430_ (
    .A1(_2638_),
    .A2(_2642_),
    .ZN(_2644_)
  );
  AND2_X1 _9431_ (
    .A1(_2596_),
    .A2(_2643_),
    .ZN(_2645_)
  );
  OR2_X1 _9432_ (
    .A1(_2597_),
    .A2(_2644_),
    .ZN(_2646_)
  );
  AND2_X1 _9433_ (
    .A1(large_1[10]),
    .A2(_2645_),
    .ZN(_2647_)
  );
  OR2_X1 _9434_ (
    .A1(_0631_),
    .A2(_2646_),
    .ZN(_2648_)
  );
  AND2_X1 _9435_ (
    .A1(large_1[11]),
    .A2(_2647_),
    .ZN(_2649_)
  );
  OR2_X1 _9436_ (
    .A1(_0630_),
    .A2(_2648_),
    .ZN(_2650_)
  );
  AND2_X1 _9437_ (
    .A1(_2592_),
    .A2(_2649_),
    .ZN(_2651_)
  );
  OR2_X1 _9438_ (
    .A1(_2593_),
    .A2(_2650_),
    .ZN(_2652_)
  );
  AND2_X1 _9439_ (
    .A1(_2588_),
    .A2(_2651_),
    .ZN(_2653_)
  );
  OR2_X1 _9440_ (
    .A1(_2589_),
    .A2(_2652_),
    .ZN(_2654_)
  );
  AND2_X1 _9441_ (
    .A1(large_1[24]),
    .A2(_2653_),
    .ZN(_2655_)
  );
  INV_X1 _9442_ (
    .A(_2655_),
    .ZN(_2656_)
  );
  AND2_X1 _9443_ (
    .A1(large_1[25]),
    .A2(_2655_),
    .ZN(_2657_)
  );
  INV_X1 _9444_ (
    .A(_2657_),
    .ZN(_2658_)
  );
  OR2_X1 _9445_ (
    .A1(large_1[26]),
    .A2(_2657_),
    .ZN(_2659_)
  );
  AND2_X1 _9446_ (
    .A1(_0736_),
    .A2(_0851_),
    .ZN(_2660_)
  );
  INV_X1 _9447_ (
    .A(_2660_),
    .ZN(_2661_)
  );
  AND2_X1 _9448_ (
    .A1(_0736_),
    .A2(_0830_),
    .ZN(_2662_)
  );
  OR2_X1 _9449_ (
    .A1(_0737_),
    .A2(_0851_),
    .ZN(_2663_)
  );
  OR2_X1 _9450_ (
    .A1(_0830_),
    .A2(_2663_),
    .ZN(_2664_)
  );
  INV_X1 _9451_ (
    .A(_2664_),
    .ZN(_2665_)
  );
  OR2_X1 _9452_ (
    .A1(_0737_),
    .A2(_2665_),
    .ZN(_2666_)
  );
  AND2_X1 _9453_ (
    .A1(_0736_),
    .A2(_0859_),
    .ZN(_2667_)
  );
  INV_X1 _9454_ (
    .A(_2667_),
    .ZN(_2668_)
  );
  AND2_X1 _9455_ (
    .A1(_2661_),
    .A2(_2668_),
    .ZN(_2669_)
  );
  OR2_X1 _9456_ (
    .A1(_2660_),
    .A2(_2667_),
    .ZN(_2670_)
  );
  AND2_X1 _9457_ (
    .A1(large_1[26]),
    .A2(_2657_),
    .ZN(_2671_)
  );
  INV_X1 _9458_ (
    .A(_2671_),
    .ZN(_2672_)
  );
  AND2_X1 _9459_ (
    .A1(_2669_),
    .A2(_2672_),
    .ZN(_2673_)
  );
  AND2_X1 _9460_ (
    .A1(_2659_),
    .A2(_2673_),
    .ZN(_2674_)
  );
  AND2_X1 _9461_ (
    .A1(_1241_),
    .A2(_2660_),
    .ZN(_2675_)
  );
  AND2_X1 _9462_ (
    .A1(large_1[26]),
    .A2(_2662_),
    .ZN(_2676_)
  );
  OR2_X1 _9463_ (
    .A1(_2675_),
    .A2(_2676_),
    .ZN(_2677_)
  );
  OR2_X1 _9464_ (
    .A1(_2674_),
    .A2(_2677_),
    .ZN(_2678_)
  );
  AND2_X1 _9465_ (
    .A1(_0654_),
    .A2(_2678_),
    .ZN(_0294_)
  );
  AND2_X1 _9466_ (
    .A1(large_1[27]),
    .A2(large_1[26]),
    .ZN(_2679_)
  );
  AND2_X1 _9467_ (
    .A1(_2635_),
    .A2(_2679_),
    .ZN(_2680_)
  );
  AND2_X1 _9468_ (
    .A1(_2653_),
    .A2(_2680_),
    .ZN(_2681_)
  );
  XOR2_X1 _9469_ (
    .A(large_1[27]),
    .B(_2671_),
    .Z(_2682_)
  );
  AND2_X1 _9470_ (
    .A1(_2669_),
    .A2(_2682_),
    .ZN(_2683_)
  );
  AND2_X1 _9471_ (
    .A1(_1290_),
    .A2(_2660_),
    .ZN(_2684_)
  );
  AND2_X1 _9472_ (
    .A1(large_1[27]),
    .A2(_2662_),
    .ZN(_2685_)
  );
  OR2_X1 _9473_ (
    .A1(_2684_),
    .A2(_2685_),
    .ZN(_2686_)
  );
  OR2_X1 _9474_ (
    .A1(_2683_),
    .A2(_2686_),
    .ZN(_2687_)
  );
  AND2_X1 _9475_ (
    .A1(_0654_),
    .A2(_2687_),
    .ZN(_0295_)
  );
  OR2_X1 _9476_ (
    .A1(large_1[28]),
    .A2(_2681_),
    .ZN(_2688_)
  );
  AND2_X1 _9477_ (
    .A1(_2669_),
    .A2(_2688_),
    .ZN(_2689_)
  );
  AND2_X1 _9478_ (
    .A1(large_1[28]),
    .A2(_2681_),
    .ZN(_2690_)
  );
  INV_X1 _9479_ (
    .A(_2690_),
    .ZN(_2691_)
  );
  AND2_X1 _9480_ (
    .A1(_2689_),
    .A2(_2691_),
    .ZN(_2692_)
  );
  AND2_X1 _9481_ (
    .A1(_1346_),
    .A2(_2660_),
    .ZN(_2693_)
  );
  AND2_X1 _9482_ (
    .A1(large_1[28]),
    .A2(_2662_),
    .ZN(_2694_)
  );
  OR2_X1 _9483_ (
    .A1(_2693_),
    .A2(_2694_),
    .ZN(_2695_)
  );
  OR2_X1 _9484_ (
    .A1(_2692_),
    .A2(_2695_),
    .ZN(_2696_)
  );
  AND2_X1 _9485_ (
    .A1(_0654_),
    .A2(_2696_),
    .ZN(_0296_)
  );
  OR2_X1 _9486_ (
    .A1(large_1[29]),
    .A2(_2690_),
    .ZN(_2697_)
  );
  AND2_X1 _9487_ (
    .A1(large_1[29]),
    .A2(large_1[28]),
    .ZN(_2698_)
  );
  AND2_X1 _9488_ (
    .A1(large_1[29]),
    .A2(_2690_),
    .ZN(_2699_)
  );
  INV_X1 _9489_ (
    .A(_2699_),
    .ZN(_2700_)
  );
  AND2_X1 _9490_ (
    .A1(_2669_),
    .A2(_2700_),
    .ZN(_2701_)
  );
  AND2_X1 _9491_ (
    .A1(_2697_),
    .A2(_2701_),
    .ZN(_2702_)
  );
  AND2_X1 _9492_ (
    .A1(_1409_),
    .A2(_2660_),
    .ZN(_2703_)
  );
  AND2_X1 _9493_ (
    .A1(large_1[29]),
    .A2(_2667_),
    .ZN(_2704_)
  );
  OR2_X1 _9494_ (
    .A1(_2703_),
    .A2(_2704_),
    .ZN(_2705_)
  );
  OR2_X1 _9495_ (
    .A1(_2702_),
    .A2(_2705_),
    .ZN(_2706_)
  );
  AND2_X1 _9496_ (
    .A1(_0654_),
    .A2(_2706_),
    .ZN(_0297_)
  );
  AND2_X1 _9497_ (
    .A1(large_1[30]),
    .A2(_2699_),
    .ZN(_2707_)
  );
  XOR2_X1 _9498_ (
    .A(large_1[30]),
    .B(_2699_),
    .Z(_2708_)
  );
  AND2_X1 _9499_ (
    .A1(_2669_),
    .A2(_2708_),
    .ZN(_2709_)
  );
  AND2_X1 _9500_ (
    .A1(_1456_),
    .A2(_2660_),
    .ZN(_2710_)
  );
  AND2_X1 _9501_ (
    .A1(large_1[30]),
    .A2(_2662_),
    .ZN(_2711_)
  );
  OR2_X1 _9502_ (
    .A1(_2710_),
    .A2(_2711_),
    .ZN(_2712_)
  );
  OR2_X1 _9503_ (
    .A1(_2709_),
    .A2(_2712_),
    .ZN(_2713_)
  );
  AND2_X1 _9504_ (
    .A1(_0654_),
    .A2(_2713_),
    .ZN(_0298_)
  );
  OR2_X1 _9505_ (
    .A1(large_1[31]),
    .A2(_2707_),
    .ZN(_2714_)
  );
  AND2_X1 _9506_ (
    .A1(large_1[31]),
    .A2(large_1[30]),
    .ZN(_2715_)
  );
  AND2_X1 _9507_ (
    .A1(large_1[31]),
    .A2(_2707_),
    .ZN(_2716_)
  );
  OR2_X1 _9508_ (
    .A1(_2670_),
    .A2(_2716_),
    .ZN(_2717_)
  );
  INV_X1 _9509_ (
    .A(_2717_),
    .ZN(_2718_)
  );
  AND2_X1 _9510_ (
    .A1(_2714_),
    .A2(_2718_),
    .ZN(_2719_)
  );
  AND2_X1 _9511_ (
    .A1(_1499_),
    .A2(_2660_),
    .ZN(_2720_)
  );
  AND2_X1 _9512_ (
    .A1(large_1[31]),
    .A2(_2662_),
    .ZN(_2721_)
  );
  OR2_X1 _9513_ (
    .A1(_2720_),
    .A2(_2721_),
    .ZN(_2722_)
  );
  OR2_X1 _9514_ (
    .A1(_2719_),
    .A2(_2722_),
    .ZN(_2723_)
  );
  AND2_X1 _9515_ (
    .A1(_0654_),
    .A2(_2723_),
    .ZN(_0299_)
  );
  AND2_X1 _9516_ (
    .A1(_2698_),
    .A2(_2715_),
    .ZN(_2724_)
  );
  AND2_X1 _9517_ (
    .A1(_2681_),
    .A2(_2724_),
    .ZN(_2725_)
  );
  AND2_X1 _9518_ (
    .A1(large_1[32]),
    .A2(_2725_),
    .ZN(_2726_)
  );
  XOR2_X1 _9519_ (
    .A(large_1[32]),
    .B(_2725_),
    .Z(_2727_)
  );
  AND2_X1 _9520_ (
    .A1(_2669_),
    .A2(_2727_),
    .ZN(_2728_)
  );
  AND2_X1 _9521_ (
    .A1(_1545_),
    .A2(_2660_),
    .ZN(_2729_)
  );
  AND2_X1 _9522_ (
    .A1(large_1[32]),
    .A2(_2662_),
    .ZN(_2730_)
  );
  OR2_X1 _9523_ (
    .A1(_2729_),
    .A2(_2730_),
    .ZN(_2731_)
  );
  OR2_X1 _9524_ (
    .A1(_2728_),
    .A2(_2731_),
    .ZN(_2732_)
  );
  AND2_X1 _9525_ (
    .A1(_0654_),
    .A2(_2732_),
    .ZN(_0300_)
  );
  OR2_X1 _9526_ (
    .A1(large_1[33]),
    .A2(_2726_),
    .ZN(_2733_)
  );
  AND2_X1 _9527_ (
    .A1(large_1[33]),
    .A2(_2726_),
    .ZN(_2734_)
  );
  INV_X1 _9528_ (
    .A(_2734_),
    .ZN(_2735_)
  );
  AND2_X1 _9529_ (
    .A1(_2669_),
    .A2(_2735_),
    .ZN(_2736_)
  );
  AND2_X1 _9530_ (
    .A1(_2733_),
    .A2(_2736_),
    .ZN(_2737_)
  );
  AND2_X1 _9531_ (
    .A1(_1601_),
    .A2(_2660_),
    .ZN(_2738_)
  );
  AND2_X1 _9532_ (
    .A1(large_1[33]),
    .A2(_2667_),
    .ZN(_2739_)
  );
  OR2_X1 _9533_ (
    .A1(_2738_),
    .A2(_2739_),
    .ZN(_2740_)
  );
  OR2_X1 _9534_ (
    .A1(_2737_),
    .A2(_2740_),
    .ZN(_2741_)
  );
  AND2_X1 _9535_ (
    .A1(_0654_),
    .A2(_2741_),
    .ZN(_0301_)
  );
  OR2_X1 _9536_ (
    .A1(large_1[34]),
    .A2(_2734_),
    .ZN(_2742_)
  );
  AND2_X1 _9537_ (
    .A1(large_1[34]),
    .A2(large_1[33]),
    .ZN(_2743_)
  );
  AND2_X1 _9538_ (
    .A1(_2726_),
    .A2(_2743_),
    .ZN(_2744_)
  );
  INV_X1 _9539_ (
    .A(_2744_),
    .ZN(_2745_)
  );
  AND2_X1 _9540_ (
    .A1(_2742_),
    .A2(_2745_),
    .ZN(_2746_)
  );
  AND2_X1 _9541_ (
    .A1(_2669_),
    .A2(_2746_),
    .ZN(_2747_)
  );
  AND2_X1 _9542_ (
    .A1(_1129_),
    .A2(_2660_),
    .ZN(_2748_)
  );
  AND2_X1 _9543_ (
    .A1(large_1[34]),
    .A2(_2662_),
    .ZN(_2749_)
  );
  OR2_X1 _9544_ (
    .A1(_2748_),
    .A2(_2749_),
    .ZN(_2750_)
  );
  OR2_X1 _9545_ (
    .A1(_2747_),
    .A2(_2750_),
    .ZN(_2751_)
  );
  AND2_X1 _9546_ (
    .A1(_0654_),
    .A2(_2751_),
    .ZN(_0302_)
  );
  OR2_X1 _9547_ (
    .A1(large_1[35]),
    .A2(_2744_),
    .ZN(_2752_)
  );
  AND2_X1 _9548_ (
    .A1(large_1[35]),
    .A2(_2743_),
    .ZN(_2753_)
  );
  AND2_X1 _9549_ (
    .A1(_2726_),
    .A2(_2753_),
    .ZN(_2754_)
  );
  INV_X1 _9550_ (
    .A(_2754_),
    .ZN(_2755_)
  );
  AND2_X1 _9551_ (
    .A1(_2669_),
    .A2(_2755_),
    .ZN(_2756_)
  );
  AND2_X1 _9552_ (
    .A1(_2752_),
    .A2(_2756_),
    .ZN(_2757_)
  );
  AND2_X1 _9553_ (
    .A1(_1175_),
    .A2(_2660_),
    .ZN(_2758_)
  );
  AND2_X1 _9554_ (
    .A1(large_1[35]),
    .A2(_2662_),
    .ZN(_2759_)
  );
  OR2_X1 _9555_ (
    .A1(_2758_),
    .A2(_2759_),
    .ZN(_2760_)
  );
  OR2_X1 _9556_ (
    .A1(_2757_),
    .A2(_2760_),
    .ZN(_2761_)
  );
  AND2_X1 _9557_ (
    .A1(_0654_),
    .A2(_2761_),
    .ZN(_0303_)
  );
  AND2_X1 _9558_ (
    .A1(large_1[36]),
    .A2(_2754_),
    .ZN(_2762_)
  );
  XOR2_X1 _9559_ (
    .A(large_1[36]),
    .B(_2754_),
    .Z(_2763_)
  );
  AND2_X1 _9560_ (
    .A1(_2669_),
    .A2(_2763_),
    .ZN(_2764_)
  );
  AND2_X1 _9561_ (
    .A1(_1647_),
    .A2(_2660_),
    .ZN(_2765_)
  );
  AND2_X1 _9562_ (
    .A1(large_1[36]),
    .A2(_2662_),
    .ZN(_2766_)
  );
  OR2_X1 _9563_ (
    .A1(_2765_),
    .A2(_2766_),
    .ZN(_2767_)
  );
  OR2_X1 _9564_ (
    .A1(_2764_),
    .A2(_2767_),
    .ZN(_2768_)
  );
  AND2_X1 _9565_ (
    .A1(_0654_),
    .A2(_2768_),
    .ZN(_0304_)
  );
  OR2_X1 _9566_ (
    .A1(large_1[37]),
    .A2(_2762_),
    .ZN(_2769_)
  );
  AND2_X1 _9567_ (
    .A1(large_1[37]),
    .A2(_2762_),
    .ZN(_2770_)
  );
  INV_X1 _9568_ (
    .A(_2770_),
    .ZN(_2771_)
  );
  AND2_X1 _9569_ (
    .A1(_2669_),
    .A2(_2771_),
    .ZN(_2772_)
  );
  AND2_X1 _9570_ (
    .A1(_2769_),
    .A2(_2772_),
    .ZN(_2773_)
  );
  AND2_X1 _9571_ (
    .A1(_1698_),
    .A2(_2660_),
    .ZN(_2774_)
  );
  AND2_X1 _9572_ (
    .A1(large_1[37]),
    .A2(_2662_),
    .ZN(_2775_)
  );
  OR2_X1 _9573_ (
    .A1(_2774_),
    .A2(_2775_),
    .ZN(_2776_)
  );
  OR2_X1 _9574_ (
    .A1(_2773_),
    .A2(_2776_),
    .ZN(_2777_)
  );
  AND2_X1 _9575_ (
    .A1(_0654_),
    .A2(_2777_),
    .ZN(_0305_)
  );
  OR2_X1 _9576_ (
    .A1(large_1[38]),
    .A2(_2770_),
    .ZN(_2778_)
  );
  AND2_X1 _9577_ (
    .A1(large_1[38]),
    .A2(large_1[37]),
    .ZN(_2779_)
  );
  AND2_X1 _9578_ (
    .A1(large_1[36]),
    .A2(_2779_),
    .ZN(_2780_)
  );
  AND2_X1 _9579_ (
    .A1(_2754_),
    .A2(_2780_),
    .ZN(_2781_)
  );
  INV_X1 _9580_ (
    .A(_2781_),
    .ZN(_2782_)
  );
  AND2_X1 _9581_ (
    .A1(_2778_),
    .A2(_2782_),
    .ZN(_2783_)
  );
  AND2_X1 _9582_ (
    .A1(_2669_),
    .A2(_2783_),
    .ZN(_2784_)
  );
  AND2_X1 _9583_ (
    .A1(_1748_),
    .A2(_2660_),
    .ZN(_2785_)
  );
  AND2_X1 _9584_ (
    .A1(large_1[38]),
    .A2(_2662_),
    .ZN(_2786_)
  );
  OR2_X1 _9585_ (
    .A1(_2785_),
    .A2(_2786_),
    .ZN(_2787_)
  );
  OR2_X1 _9586_ (
    .A1(_2784_),
    .A2(_2787_),
    .ZN(_2788_)
  );
  AND2_X1 _9587_ (
    .A1(_0654_),
    .A2(_2788_),
    .ZN(_0306_)
  );
  OR2_X1 _9588_ (
    .A1(large_1[39]),
    .A2(_2781_),
    .ZN(_2789_)
  );
  AND2_X1 _9589_ (
    .A1(large_1[39]),
    .A2(_2781_),
    .ZN(_2790_)
  );
  INV_X1 _9590_ (
    .A(_2790_),
    .ZN(_2791_)
  );
  AND2_X1 _9591_ (
    .A1(_2669_),
    .A2(_2791_),
    .ZN(_2792_)
  );
  AND2_X1 _9592_ (
    .A1(_2789_),
    .A2(_2792_),
    .ZN(_2793_)
  );
  AND2_X1 _9593_ (
    .A1(_1790_),
    .A2(_2660_),
    .ZN(_2794_)
  );
  AND2_X1 _9594_ (
    .A1(large_1[39]),
    .A2(_2662_),
    .ZN(_2795_)
  );
  OR2_X1 _9595_ (
    .A1(_2794_),
    .A2(_2795_),
    .ZN(_2796_)
  );
  OR2_X1 _9596_ (
    .A1(_2793_),
    .A2(_2796_),
    .ZN(_2797_)
  );
  AND2_X1 _9597_ (
    .A1(_0654_),
    .A2(_2797_),
    .ZN(_0307_)
  );
  AND2_X1 _9598_ (
    .A1(_2680_),
    .A2(_2715_),
    .ZN(_2798_)
  );
  AND2_X1 _9599_ (
    .A1(large_1[39]),
    .A2(large_1[32]),
    .ZN(_2799_)
  );
  AND2_X1 _9600_ (
    .A1(_2698_),
    .A2(_2799_),
    .ZN(_2800_)
  );
  AND2_X1 _9601_ (
    .A1(_2753_),
    .A2(_2800_),
    .ZN(_2801_)
  );
  AND2_X1 _9602_ (
    .A1(_2780_),
    .A2(_2801_),
    .ZN(_2802_)
  );
  AND2_X1 _9603_ (
    .A1(_2798_),
    .A2(_2802_),
    .ZN(_2803_)
  );
  AND2_X1 _9604_ (
    .A1(_2623_),
    .A2(_2803_),
    .ZN(_2804_)
  );
  AND2_X1 _9605_ (
    .A1(_2680_),
    .A2(_2799_),
    .ZN(_2805_)
  );
  AND2_X1 _9606_ (
    .A1(_2724_),
    .A2(_2753_),
    .ZN(_2806_)
  );
  AND2_X1 _9607_ (
    .A1(_2780_),
    .A2(_2805_),
    .ZN(_2807_)
  );
  AND2_X1 _9608_ (
    .A1(_2806_),
    .A2(_2807_),
    .ZN(_2808_)
  );
  INV_X1 _9609_ (
    .A(_2808_),
    .ZN(_2809_)
  );
  AND2_X1 _9610_ (
    .A1(_2653_),
    .A2(_2808_),
    .ZN(_2810_)
  );
  OR2_X1 _9611_ (
    .A1(_2654_),
    .A2(_2809_),
    .ZN(_2811_)
  );
  AND2_X1 _9612_ (
    .A1(large_1[40]),
    .A2(_2810_),
    .ZN(_2812_)
  );
  XOR2_X1 _9613_ (
    .A(large_1[40]),
    .B(_2810_),
    .Z(_2813_)
  );
  AND2_X1 _9614_ (
    .A1(_2669_),
    .A2(_2813_),
    .ZN(_2814_)
  );
  AND2_X1 _9615_ (
    .A1(_1832_),
    .A2(_2660_),
    .ZN(_2815_)
  );
  AND2_X1 _9616_ (
    .A1(large_1[40]),
    .A2(_2662_),
    .ZN(_2816_)
  );
  OR2_X1 _9617_ (
    .A1(_2815_),
    .A2(_2816_),
    .ZN(_2817_)
  );
  OR2_X1 _9618_ (
    .A1(_2814_),
    .A2(_2817_),
    .ZN(_2818_)
  );
  AND2_X1 _9619_ (
    .A1(_0654_),
    .A2(_2818_),
    .ZN(_0308_)
  );
  OR2_X1 _9620_ (
    .A1(large_1[41]),
    .A2(_2812_),
    .ZN(_2819_)
  );
  AND2_X1 _9621_ (
    .A1(large_1[41]),
    .A2(large_1[40]),
    .ZN(_2820_)
  );
  AND2_X1 _9622_ (
    .A1(large_1[41]),
    .A2(_2812_),
    .ZN(_2821_)
  );
  INV_X1 _9623_ (
    .A(_2821_),
    .ZN(_2822_)
  );
  AND2_X1 _9624_ (
    .A1(_2669_),
    .A2(_2822_),
    .ZN(_2823_)
  );
  AND2_X1 _9625_ (
    .A1(_2819_),
    .A2(_2823_),
    .ZN(_2824_)
  );
  AND2_X1 _9626_ (
    .A1(_1880_),
    .A2(_2660_),
    .ZN(_2825_)
  );
  AND2_X1 _9627_ (
    .A1(large_1[41]),
    .A2(_2662_),
    .ZN(_2826_)
  );
  OR2_X1 _9628_ (
    .A1(_2825_),
    .A2(_2826_),
    .ZN(_2827_)
  );
  OR2_X1 _9629_ (
    .A1(_2824_),
    .A2(_2827_),
    .ZN(_2828_)
  );
  AND2_X1 _9630_ (
    .A1(_0654_),
    .A2(_2828_),
    .ZN(_0309_)
  );
  AND2_X1 _9631_ (
    .A1(large_1[42]),
    .A2(_2821_),
    .ZN(_2829_)
  );
  XOR2_X1 _9632_ (
    .A(large_1[42]),
    .B(_2821_),
    .Z(_2830_)
  );
  AND2_X1 _9633_ (
    .A1(_2669_),
    .A2(_2830_),
    .ZN(_2831_)
  );
  AND2_X1 _9634_ (
    .A1(_0862_),
    .A2(_2660_),
    .ZN(_2832_)
  );
  AND2_X1 _9635_ (
    .A1(large_1[42]),
    .A2(_2662_),
    .ZN(_2833_)
  );
  OR2_X1 _9636_ (
    .A1(_2832_),
    .A2(_2833_),
    .ZN(_2834_)
  );
  OR2_X1 _9637_ (
    .A1(_2831_),
    .A2(_2834_),
    .ZN(_2835_)
  );
  AND2_X1 _9638_ (
    .A1(_0654_),
    .A2(_2835_),
    .ZN(_0310_)
  );
  OR2_X1 _9639_ (
    .A1(large_1[43]),
    .A2(_2829_),
    .ZN(_2836_)
  );
  AND2_X1 _9640_ (
    .A1(large_1[43]),
    .A2(large_1[42]),
    .ZN(_2837_)
  );
  AND2_X1 _9641_ (
    .A1(large_1[43]),
    .A2(_2829_),
    .ZN(_2838_)
  );
  INV_X1 _9642_ (
    .A(_2838_),
    .ZN(_2839_)
  );
  AND2_X1 _9643_ (
    .A1(_2669_),
    .A2(_2839_),
    .ZN(_2840_)
  );
  AND2_X1 _9644_ (
    .A1(_2836_),
    .A2(_2840_),
    .ZN(_2841_)
  );
  AND2_X1 _9645_ (
    .A1(_1926_),
    .A2(_2660_),
    .ZN(_2842_)
  );
  AND2_X1 _9646_ (
    .A1(large_1[43]),
    .A2(_2667_),
    .ZN(_2843_)
  );
  OR2_X1 _9647_ (
    .A1(_2842_),
    .A2(_2843_),
    .ZN(_2844_)
  );
  OR2_X1 _9648_ (
    .A1(_2841_),
    .A2(_2844_),
    .ZN(_2845_)
  );
  AND2_X1 _9649_ (
    .A1(_0654_),
    .A2(_2845_),
    .ZN(_0311_)
  );
  AND2_X1 _9650_ (
    .A1(_2820_),
    .A2(_2837_),
    .ZN(_2846_)
  );
  INV_X1 _9651_ (
    .A(_2846_),
    .ZN(_2847_)
  );
  AND2_X1 _9652_ (
    .A1(_2810_),
    .A2(_2846_),
    .ZN(_2848_)
  );
  AND2_X1 _9653_ (
    .A1(large_1[44]),
    .A2(_2848_),
    .ZN(_2849_)
  );
  XOR2_X1 _9654_ (
    .A(large_1[44]),
    .B(_2848_),
    .Z(_2850_)
  );
  AND2_X1 _9655_ (
    .A1(_2669_),
    .A2(_2850_),
    .ZN(_2851_)
  );
  AND2_X1 _9656_ (
    .A1(_0908_),
    .A2(_2660_),
    .ZN(_2852_)
  );
  AND2_X1 _9657_ (
    .A1(large_1[44]),
    .A2(_2662_),
    .ZN(_2853_)
  );
  OR2_X1 _9658_ (
    .A1(_2852_),
    .A2(_2853_),
    .ZN(_2854_)
  );
  OR2_X1 _9659_ (
    .A1(_2851_),
    .A2(_2854_),
    .ZN(_2855_)
  );
  AND2_X1 _9660_ (
    .A1(_0654_),
    .A2(_2855_),
    .ZN(_0312_)
  );
  OR2_X1 _9661_ (
    .A1(large_1[45]),
    .A2(_2849_),
    .ZN(_2856_)
  );
  AND2_X1 _9662_ (
    .A1(large_1[45]),
    .A2(large_1[44]),
    .ZN(_2857_)
  );
  AND2_X1 _9663_ (
    .A1(large_1[45]),
    .A2(_2849_),
    .ZN(_2858_)
  );
  INV_X1 _9664_ (
    .A(_2858_),
    .ZN(_2859_)
  );
  AND2_X1 _9665_ (
    .A1(_2669_),
    .A2(_2859_),
    .ZN(_2860_)
  );
  AND2_X1 _9666_ (
    .A1(_2856_),
    .A2(_2860_),
    .ZN(_2861_)
  );
  AND2_X1 _9667_ (
    .A1(_0967_),
    .A2(_2660_),
    .ZN(_2862_)
  );
  AND2_X1 _9668_ (
    .A1(large_1[45]),
    .A2(_2662_),
    .ZN(_2863_)
  );
  OR2_X1 _9669_ (
    .A1(_2862_),
    .A2(_2863_),
    .ZN(_2864_)
  );
  OR2_X1 _9670_ (
    .A1(_2861_),
    .A2(_2864_),
    .ZN(_2865_)
  );
  AND2_X1 _9671_ (
    .A1(_0654_),
    .A2(_2865_),
    .ZN(_0313_)
  );
  AND2_X1 _9672_ (
    .A1(large_1[46]),
    .A2(_2858_),
    .ZN(_2866_)
  );
  XOR2_X1 _9673_ (
    .A(large_1[46]),
    .B(_2858_),
    .Z(_2867_)
  );
  AND2_X1 _9674_ (
    .A1(_2669_),
    .A2(_2867_),
    .ZN(_2868_)
  );
  AND2_X1 _9675_ (
    .A1(_1017_),
    .A2(_2660_),
    .ZN(_2869_)
  );
  AND2_X1 _9676_ (
    .A1(large_1[46]),
    .A2(_2662_),
    .ZN(_2870_)
  );
  OR2_X1 _9677_ (
    .A1(_2869_),
    .A2(_2870_),
    .ZN(_2871_)
  );
  OR2_X1 _9678_ (
    .A1(_2868_),
    .A2(_2871_),
    .ZN(_2872_)
  );
  AND2_X1 _9679_ (
    .A1(_0654_),
    .A2(_2872_),
    .ZN(_0314_)
  );
  OR2_X1 _9680_ (
    .A1(large_1[47]),
    .A2(_2866_),
    .ZN(_2873_)
  );
  AND2_X1 _9681_ (
    .A1(large_1[47]),
    .A2(large_1[46]),
    .ZN(_2874_)
  );
  AND2_X1 _9682_ (
    .A1(_2857_),
    .A2(_2874_),
    .ZN(_2875_)
  );
  INV_X1 _9683_ (
    .A(_2875_),
    .ZN(_2876_)
  );
  AND2_X1 _9684_ (
    .A1(large_1[47]),
    .A2(_2866_),
    .ZN(_2877_)
  );
  INV_X1 _9685_ (
    .A(_2877_),
    .ZN(_2878_)
  );
  AND2_X1 _9686_ (
    .A1(_2669_),
    .A2(_2878_),
    .ZN(_2879_)
  );
  AND2_X1 _9687_ (
    .A1(_2873_),
    .A2(_2879_),
    .ZN(_2880_)
  );
  AND2_X1 _9688_ (
    .A1(_1968_),
    .A2(_2660_),
    .ZN(_2881_)
  );
  AND2_X1 _9689_ (
    .A1(large_1[47]),
    .A2(_2662_),
    .ZN(_2882_)
  );
  OR2_X1 _9690_ (
    .A1(_2881_),
    .A2(_2882_),
    .ZN(_2883_)
  );
  OR2_X1 _9691_ (
    .A1(_2880_),
    .A2(_2883_),
    .ZN(_2884_)
  );
  AND2_X1 _9692_ (
    .A1(_0654_),
    .A2(_2884_),
    .ZN(_0315_)
  );
  AND2_X1 _9693_ (
    .A1(_2846_),
    .A2(_2875_),
    .ZN(_2885_)
  );
  OR2_X1 _9694_ (
    .A1(_2847_),
    .A2(_2876_),
    .ZN(_2886_)
  );
  AND2_X1 _9695_ (
    .A1(_2804_),
    .A2(_2885_),
    .ZN(_2887_)
  );
  AND2_X1 _9696_ (
    .A1(large_1[48]),
    .A2(_2887_),
    .ZN(_2888_)
  );
  AND2_X1 _9697_ (
    .A1(_2810_),
    .A2(_2885_),
    .ZN(_2889_)
  );
  OR2_X1 _9698_ (
    .A1(_2811_),
    .A2(_2886_),
    .ZN(_2890_)
  );
  AND2_X1 _9699_ (
    .A1(large_1[48]),
    .A2(_2889_),
    .ZN(_2891_)
  );
  OR2_X1 _9700_ (
    .A1(_0651_),
    .A2(_2890_),
    .ZN(_2892_)
  );
  XOR2_X1 _9701_ (
    .A(_0651_),
    .B(_2890_),
    .Z(_2893_)
  );
  AND2_X1 _9702_ (
    .A1(_2669_),
    .A2(_2893_),
    .ZN(_2894_)
  );
  AND2_X1 _9703_ (
    .A1(_2010_),
    .A2(_2660_),
    .ZN(_2895_)
  );
  AND2_X1 _9704_ (
    .A1(large_1[48]),
    .A2(_2662_),
    .ZN(_2896_)
  );
  OR2_X1 _9705_ (
    .A1(_2895_),
    .A2(_2896_),
    .ZN(_2897_)
  );
  OR2_X1 _9706_ (
    .A1(_2894_),
    .A2(_2897_),
    .ZN(_2898_)
  );
  AND2_X1 _9707_ (
    .A1(_0654_),
    .A2(_2898_),
    .ZN(_0316_)
  );
  OR2_X1 _9708_ (
    .A1(large_1[49]),
    .A2(_2891_),
    .ZN(_2899_)
  );
  AND2_X1 _9709_ (
    .A1(large_1[49]),
    .A2(_2891_),
    .ZN(_2900_)
  );
  OR2_X1 _9710_ (
    .A1(_2670_),
    .A2(_2900_),
    .ZN(_2901_)
  );
  INV_X1 _9711_ (
    .A(_2901_),
    .ZN(_2902_)
  );
  AND2_X1 _9712_ (
    .A1(_2899_),
    .A2(_2902_),
    .ZN(_2903_)
  );
  AND2_X1 _9713_ (
    .A1(_1071_),
    .A2(_2660_),
    .ZN(_2904_)
  );
  AND2_X1 _9714_ (
    .A1(large_1[49]),
    .A2(_2662_),
    .ZN(_2905_)
  );
  OR2_X1 _9715_ (
    .A1(_2904_),
    .A2(_2905_),
    .ZN(_2906_)
  );
  OR2_X1 _9716_ (
    .A1(_2903_),
    .A2(_2906_),
    .ZN(_2907_)
  );
  AND2_X1 _9717_ (
    .A1(_0654_),
    .A2(_2907_),
    .ZN(_0317_)
  );
  OR2_X1 _9718_ (
    .A1(large_1[50]),
    .A2(_2900_),
    .ZN(_2908_)
  );
  AND2_X1 _9719_ (
    .A1(large_1[50]),
    .A2(large_1[49]),
    .ZN(_2909_)
  );
  OR2_X1 _9720_ (
    .A1(_0649_),
    .A2(_0650_),
    .ZN(_2910_)
  );
  AND2_X1 _9721_ (
    .A1(_2888_),
    .A2(_2909_),
    .ZN(_2911_)
  );
  AND2_X1 _9722_ (
    .A1(_2891_),
    .A2(_2909_),
    .ZN(_2912_)
  );
  OR2_X1 _9723_ (
    .A1(_2892_),
    .A2(_2910_),
    .ZN(_2913_)
  );
  AND2_X1 _9724_ (
    .A1(_2908_),
    .A2(_2913_),
    .ZN(_2914_)
  );
  AND2_X1 _9725_ (
    .A1(_2669_),
    .A2(_2914_),
    .ZN(_2915_)
  );
  AND2_X1 _9726_ (
    .A1(_2056_),
    .A2(_2660_),
    .ZN(_2916_)
  );
  AND2_X1 _9727_ (
    .A1(large_1[50]),
    .A2(_2662_),
    .ZN(_2917_)
  );
  OR2_X1 _9728_ (
    .A1(_2916_),
    .A2(_2917_),
    .ZN(_2918_)
  );
  OR2_X1 _9729_ (
    .A1(_2915_),
    .A2(_2918_),
    .ZN(_2919_)
  );
  AND2_X1 _9730_ (
    .A1(_0654_),
    .A2(_2919_),
    .ZN(_0318_)
  );
  OR2_X1 _9731_ (
    .A1(large_1[51]),
    .A2(_2911_),
    .ZN(_2920_)
  );
  AND2_X1 _9732_ (
    .A1(large_1[51]),
    .A2(_2911_),
    .ZN(_2921_)
  );
  AND2_X1 _9733_ (
    .A1(large_1[51]),
    .A2(_2912_),
    .ZN(_2922_)
  );
  OR2_X1 _9734_ (
    .A1(_0648_),
    .A2(_2913_),
    .ZN(_2923_)
  );
  OR2_X1 _9735_ (
    .A1(_2670_),
    .A2(_2922_),
    .ZN(_2924_)
  );
  INV_X1 _9736_ (
    .A(_2924_),
    .ZN(_2925_)
  );
  AND2_X1 _9737_ (
    .A1(_2920_),
    .A2(_2925_),
    .ZN(_2926_)
  );
  AND2_X1 _9738_ (
    .A1(_2102_),
    .A2(_2660_),
    .ZN(_2927_)
  );
  AND2_X1 _9739_ (
    .A1(large_1[51]),
    .A2(_2667_),
    .ZN(_2928_)
  );
  OR2_X1 _9740_ (
    .A1(_2927_),
    .A2(_2928_),
    .ZN(_2929_)
  );
  OR2_X1 _9741_ (
    .A1(_2926_),
    .A2(_2929_),
    .ZN(_2930_)
  );
  AND2_X1 _9742_ (
    .A1(_0654_),
    .A2(_2930_),
    .ZN(_0319_)
  );
  AND2_X1 _9743_ (
    .A1(large_1[52]),
    .A2(_2921_),
    .ZN(_2931_)
  );
  AND2_X1 _9744_ (
    .A1(large_1[52]),
    .A2(_2922_),
    .ZN(_2932_)
  );
  OR2_X1 _9745_ (
    .A1(_0647_),
    .A2(_2923_),
    .ZN(_2933_)
  );
  XOR2_X1 _9746_ (
    .A(_0647_),
    .B(_2923_),
    .Z(_2934_)
  );
  AND2_X1 _9747_ (
    .A1(_2669_),
    .A2(_2934_),
    .ZN(_2935_)
  );
  AND2_X1 _9748_ (
    .A1(_2148_),
    .A2(_2660_),
    .ZN(_2936_)
  );
  AND2_X1 _9749_ (
    .A1(large_1[52]),
    .A2(_2662_),
    .ZN(_2937_)
  );
  OR2_X1 _9750_ (
    .A1(_2936_),
    .A2(_2937_),
    .ZN(_2938_)
  );
  OR2_X1 _9751_ (
    .A1(_2935_),
    .A2(_2938_),
    .ZN(_2939_)
  );
  AND2_X1 _9752_ (
    .A1(_0654_),
    .A2(_2939_),
    .ZN(_0320_)
  );
  OR2_X1 _9753_ (
    .A1(large_1[53]),
    .A2(_2931_),
    .ZN(_2940_)
  );
  AND2_X1 _9754_ (
    .A1(large_1[53]),
    .A2(_2931_),
    .ZN(_2941_)
  );
  AND2_X1 _9755_ (
    .A1(large_1[53]),
    .A2(_2932_),
    .ZN(_2942_)
  );
  OR2_X1 _9756_ (
    .A1(_0646_),
    .A2(_2933_),
    .ZN(_2943_)
  );
  OR2_X1 _9757_ (
    .A1(_2670_),
    .A2(_2942_),
    .ZN(_2944_)
  );
  INV_X1 _9758_ (
    .A(_2944_),
    .ZN(_2945_)
  );
  AND2_X1 _9759_ (
    .A1(_2940_),
    .A2(_2945_),
    .ZN(_2946_)
  );
  AND2_X1 _9760_ (
    .A1(_2195_),
    .A2(_2660_),
    .ZN(_2947_)
  );
  AND2_X1 _9761_ (
    .A1(large_1[53]),
    .A2(_2662_),
    .ZN(_2948_)
  );
  OR2_X1 _9762_ (
    .A1(_2947_),
    .A2(_2948_),
    .ZN(_2949_)
  );
  OR2_X1 _9763_ (
    .A1(_2946_),
    .A2(_2949_),
    .ZN(_2950_)
  );
  AND2_X1 _9764_ (
    .A1(_0654_),
    .A2(_2950_),
    .ZN(_0321_)
  );
  AND2_X1 _9765_ (
    .A1(large_1[54]),
    .A2(_2941_),
    .ZN(_2951_)
  );
  OR2_X1 _9766_ (
    .A1(_0645_),
    .A2(_2943_),
    .ZN(_2952_)
  );
  XOR2_X1 _9767_ (
    .A(_0645_),
    .B(_2943_),
    .Z(_2953_)
  );
  AND2_X1 _9768_ (
    .A1(_2669_),
    .A2(_2953_),
    .ZN(_2954_)
  );
  AND2_X1 _9769_ (
    .A1(_2241_),
    .A2(_2660_),
    .ZN(_2955_)
  );
  AND2_X1 _9770_ (
    .A1(large_1[54]),
    .A2(_2662_),
    .ZN(_2956_)
  );
  OR2_X1 _9771_ (
    .A1(_2955_),
    .A2(_2956_),
    .ZN(_2957_)
  );
  OR2_X1 _9772_ (
    .A1(_2954_),
    .A2(_2957_),
    .ZN(_2958_)
  );
  AND2_X1 _9773_ (
    .A1(_0654_),
    .A2(_2958_),
    .ZN(_0322_)
  );
  OR2_X1 _9774_ (
    .A1(large_1[55]),
    .A2(_2951_),
    .ZN(_2959_)
  );
  AND2_X1 _9775_ (
    .A1(large_1[55]),
    .A2(_2951_),
    .ZN(_2960_)
  );
  OR2_X1 _9776_ (
    .A1(_0644_),
    .A2(_2952_),
    .ZN(_2961_)
  );
  AND2_X1 _9777_ (
    .A1(_2669_),
    .A2(_2961_),
    .ZN(_2962_)
  );
  AND2_X1 _9778_ (
    .A1(_2959_),
    .A2(_2962_),
    .ZN(_2963_)
  );
  AND2_X1 _9779_ (
    .A1(_2285_),
    .A2(_2660_),
    .ZN(_2964_)
  );
  AND2_X1 _9780_ (
    .A1(large_1[55]),
    .A2(_2662_),
    .ZN(_2965_)
  );
  OR2_X1 _9781_ (
    .A1(_2964_),
    .A2(_2965_),
    .ZN(_2966_)
  );
  OR2_X1 _9782_ (
    .A1(_2963_),
    .A2(_2966_),
    .ZN(_2967_)
  );
  AND2_X1 _9783_ (
    .A1(_0654_),
    .A2(_2967_),
    .ZN(_0323_)
  );
  OR2_X1 _9784_ (
    .A1(large_1[56]),
    .A2(_2960_),
    .ZN(_2968_)
  );
  OR2_X1 _9785_ (
    .A1(_0643_),
    .A2(_2961_),
    .ZN(_2969_)
  );
  AND2_X1 _9786_ (
    .A1(_2669_),
    .A2(_2969_),
    .ZN(_2970_)
  );
  AND2_X1 _9787_ (
    .A1(_2968_),
    .A2(_2970_),
    .ZN(_2971_)
  );
  AND2_X1 _9788_ (
    .A1(_2435_),
    .A2(_2660_),
    .ZN(_2972_)
  );
  AND2_X1 _9789_ (
    .A1(large_1[56]),
    .A2(_2662_),
    .ZN(_2973_)
  );
  OR2_X1 _9790_ (
    .A1(_2972_),
    .A2(_2973_),
    .ZN(_2974_)
  );
  OR2_X1 _9791_ (
    .A1(_2971_),
    .A2(_2974_),
    .ZN(_2975_)
  );
  AND2_X1 _9792_ (
    .A1(_0654_),
    .A2(_2975_),
    .ZN(_0324_)
  );
  XOR2_X1 _9793_ (
    .A(_0642_),
    .B(_2969_),
    .Z(_2976_)
  );
  AND2_X1 _9794_ (
    .A1(_2669_),
    .A2(_2976_),
    .ZN(_2977_)
  );
  AND2_X1 _9795_ (
    .A1(_2365_),
    .A2(_2660_),
    .ZN(_2978_)
  );
  AND2_X1 _9796_ (
    .A1(large_1[57]),
    .A2(_2667_),
    .ZN(_2979_)
  );
  OR2_X1 _9797_ (
    .A1(_2978_),
    .A2(_2979_),
    .ZN(_2980_)
  );
  OR2_X1 _9798_ (
    .A1(_2977_),
    .A2(_2980_),
    .ZN(_2981_)
  );
  AND2_X1 _9799_ (
    .A1(_0654_),
    .A2(_2981_),
    .ZN(_0325_)
  );
  OR2_X1 _9800_ (
    .A1(reg_mcountinhibit[0]),
    .A2(io_csr_stall),
    .ZN(_2982_)
  );
  XOR2_X1 _9801_ (
    .A(_0641_),
    .B(_2982_),
    .Z(_2983_)
  );
  AND2_X1 _9802_ (
    .A1(_2665_),
    .A2(_2983_),
    .ZN(_2984_)
  );
  AND2_X1 _9803_ (
    .A1(small_1[0]),
    .A2(_2660_),
    .ZN(_2985_)
  );
  AND2_X1 _9804_ (
    .A1(_0737_),
    .A2(_2983_),
    .ZN(_2986_)
  );
  OR2_X1 _9805_ (
    .A1(_2985_),
    .A2(_2986_),
    .ZN(_2987_)
  );
  OR2_X1 _9806_ (
    .A1(_2984_),
    .A2(_2987_),
    .ZN(_2988_)
  );
  AND2_X1 _9807_ (
    .A1(_1241_),
    .A2(_2667_),
    .ZN(_2989_)
  );
  OR2_X1 _9808_ (
    .A1(_2988_),
    .A2(_2989_),
    .ZN(_2990_)
  );
  AND2_X1 _9809_ (
    .A1(_0654_),
    .A2(_2990_),
    .ZN(_0326_)
  );
  AND2_X1 _9810_ (
    .A1(small_1[1]),
    .A2(_2660_),
    .ZN(_2991_)
  );
  OR2_X1 _9811_ (
    .A1(reg_mcountinhibit[0]),
    .A2(_2605_),
    .ZN(_2992_)
  );
  XOR2_X1 _9812_ (
    .A(_0640_),
    .B(_2992_),
    .Z(_2993_)
  );
  AND2_X1 _9813_ (
    .A1(_2666_),
    .A2(_2993_),
    .ZN(_2994_)
  );
  OR2_X1 _9814_ (
    .A1(_2991_),
    .A2(_2994_),
    .ZN(_2995_)
  );
  AND2_X1 _9815_ (
    .A1(_1290_),
    .A2(_2662_),
    .ZN(_2996_)
  );
  OR2_X1 _9816_ (
    .A1(_2995_),
    .A2(_2996_),
    .ZN(_2997_)
  );
  AND2_X1 _9817_ (
    .A1(_0654_),
    .A2(_2997_),
    .ZN(_0327_)
  );
  AND2_X1 _9818_ (
    .A1(small_1[2]),
    .A2(_2660_),
    .ZN(_2998_)
  );
  OR2_X1 _9819_ (
    .A1(reg_mcountinhibit[0]),
    .A2(_2607_),
    .ZN(_2999_)
  );
  XOR2_X1 _9820_ (
    .A(_0639_),
    .B(_2999_),
    .Z(_3000_)
  );
  AND2_X1 _9821_ (
    .A1(_2666_),
    .A2(_3000_),
    .ZN(_3001_)
  );
  OR2_X1 _9822_ (
    .A1(_2998_),
    .A2(_3001_),
    .ZN(_3002_)
  );
  AND2_X1 _9823_ (
    .A1(_1346_),
    .A2(_2667_),
    .ZN(_3003_)
  );
  OR2_X1 _9824_ (
    .A1(_3002_),
    .A2(_3003_),
    .ZN(_3004_)
  );
  AND2_X1 _9825_ (
    .A1(_0654_),
    .A2(_3004_),
    .ZN(_0328_)
  );
  AND2_X1 _9826_ (
    .A1(small_1[3]),
    .A2(_2660_),
    .ZN(_3005_)
  );
  OR2_X1 _9827_ (
    .A1(reg_mcountinhibit[0]),
    .A2(_2609_),
    .ZN(_3006_)
  );
  XOR2_X1 _9828_ (
    .A(_0638_),
    .B(_3006_),
    .Z(_3007_)
  );
  AND2_X1 _9829_ (
    .A1(_2669_),
    .A2(_3007_),
    .ZN(_3008_)
  );
  OR2_X1 _9830_ (
    .A1(_3005_),
    .A2(_3008_),
    .ZN(_3009_)
  );
  AND2_X1 _9831_ (
    .A1(_1409_),
    .A2(_2662_),
    .ZN(_3010_)
  );
  OR2_X1 _9832_ (
    .A1(_3009_),
    .A2(_3010_),
    .ZN(_3011_)
  );
  AND2_X1 _9833_ (
    .A1(_0654_),
    .A2(_3011_),
    .ZN(_0329_)
  );
  OR2_X1 _9834_ (
    .A1(reg_mcountinhibit[0]),
    .A2(_2611_),
    .ZN(_3012_)
  );
  OR2_X1 _9835_ (
    .A1(_0637_),
    .A2(_3012_),
    .ZN(_3013_)
  );
  XOR2_X1 _9836_ (
    .A(_0637_),
    .B(_3012_),
    .Z(_3014_)
  );
  AND2_X1 _9837_ (
    .A1(_2669_),
    .A2(_3014_),
    .ZN(_3015_)
  );
  AND2_X1 _9838_ (
    .A1(small_1[4]),
    .A2(_2660_),
    .ZN(_3016_)
  );
  OR2_X1 _9839_ (
    .A1(_3015_),
    .A2(_3016_),
    .ZN(_3017_)
  );
  AND2_X1 _9840_ (
    .A1(_1456_),
    .A2(_2662_),
    .ZN(_3018_)
  );
  OR2_X1 _9841_ (
    .A1(_3017_),
    .A2(_3018_),
    .ZN(_3019_)
  );
  AND2_X1 _9842_ (
    .A1(_0654_),
    .A2(_3019_),
    .ZN(_0330_)
  );
  AND2_X1 _9843_ (
    .A1(_1499_),
    .A2(_2662_),
    .ZN(_3020_)
  );
  AND2_X1 _9844_ (
    .A1(small_1[5]),
    .A2(_2660_),
    .ZN(_3021_)
  );
  XOR2_X1 _9845_ (
    .A(_0636_),
    .B(_3013_),
    .Z(_3022_)
  );
  AND2_X1 _9846_ (
    .A1(_2669_),
    .A2(_3022_),
    .ZN(_3023_)
  );
  OR2_X1 _9847_ (
    .A1(_3021_),
    .A2(_3023_),
    .ZN(_3024_)
  );
  OR2_X1 _9848_ (
    .A1(_3020_),
    .A2(_3024_),
    .ZN(_3025_)
  );
  AND2_X1 _9849_ (
    .A1(_0654_),
    .A2(_3025_),
    .ZN(_0331_)
  );
  AND2_X1 _9850_ (
    .A1(_0736_),
    .A2(_0767_),
    .ZN(_3026_)
  );
  MUX2_X1 _9851_ (
    .A(reg_mscratch[0]),
    .B(_1241_),
    .S(_3026_),
    .Z(_0332_)
  );
  MUX2_X1 _9852_ (
    .A(reg_mscratch[1]),
    .B(_1290_),
    .S(_3026_),
    .Z(_0333_)
  );
  MUX2_X1 _9853_ (
    .A(reg_mscratch[2]),
    .B(_1346_),
    .S(_3026_),
    .Z(_0334_)
  );
  MUX2_X1 _9854_ (
    .A(reg_mscratch[3]),
    .B(_1409_),
    .S(_3026_),
    .Z(_0335_)
  );
  MUX2_X1 _9855_ (
    .A(reg_mscratch[4]),
    .B(_1456_),
    .S(_3026_),
    .Z(_0336_)
  );
  MUX2_X1 _9856_ (
    .A(reg_mscratch[5]),
    .B(_1499_),
    .S(_3026_),
    .Z(_0337_)
  );
  MUX2_X1 _9857_ (
    .A(reg_mscratch[6]),
    .B(_1545_),
    .S(_3026_),
    .Z(_0338_)
  );
  MUX2_X1 _9858_ (
    .A(reg_mscratch[7]),
    .B(_1601_),
    .S(_3026_),
    .Z(_0339_)
  );
  MUX2_X1 _9859_ (
    .A(reg_mscratch[8]),
    .B(_1129_),
    .S(_3026_),
    .Z(_0340_)
  );
  MUX2_X1 _9860_ (
    .A(reg_mscratch[9]),
    .B(_1175_),
    .S(_3026_),
    .Z(_0341_)
  );
  MUX2_X1 _9861_ (
    .A(reg_mscratch[10]),
    .B(_1647_),
    .S(_3026_),
    .Z(_0342_)
  );
  MUX2_X1 _9862_ (
    .A(reg_mscratch[11]),
    .B(_1698_),
    .S(_3026_),
    .Z(_0343_)
  );
  MUX2_X1 _9863_ (
    .A(reg_mscratch[12]),
    .B(_1748_),
    .S(_3026_),
    .Z(_0344_)
  );
  MUX2_X1 _9864_ (
    .A(reg_mscratch[13]),
    .B(_1790_),
    .S(_3026_),
    .Z(_0345_)
  );
  MUX2_X1 _9865_ (
    .A(reg_mscratch[14]),
    .B(_1832_),
    .S(_3026_),
    .Z(_0346_)
  );
  MUX2_X1 _9866_ (
    .A(reg_mscratch[15]),
    .B(_1880_),
    .S(_3026_),
    .Z(_0347_)
  );
  MUX2_X1 _9867_ (
    .A(reg_mscratch[16]),
    .B(_0862_),
    .S(_3026_),
    .Z(_0348_)
  );
  MUX2_X1 _9868_ (
    .A(reg_mscratch[17]),
    .B(_1926_),
    .S(_3026_),
    .Z(_0349_)
  );
  MUX2_X1 _9869_ (
    .A(reg_mscratch[18]),
    .B(_0908_),
    .S(_3026_),
    .Z(_0350_)
  );
  MUX2_X1 _9870_ (
    .A(reg_mscratch[19]),
    .B(_0967_),
    .S(_3026_),
    .Z(_0351_)
  );
  MUX2_X1 _9871_ (
    .A(reg_mscratch[20]),
    .B(_1017_),
    .S(_3026_),
    .Z(_0352_)
  );
  MUX2_X1 _9872_ (
    .A(reg_mscratch[21]),
    .B(_1968_),
    .S(_3026_),
    .Z(_0353_)
  );
  MUX2_X1 _9873_ (
    .A(reg_mscratch[22]),
    .B(_2010_),
    .S(_3026_),
    .Z(_0354_)
  );
  MUX2_X1 _9874_ (
    .A(reg_mscratch[23]),
    .B(_1071_),
    .S(_3026_),
    .Z(_0355_)
  );
  MUX2_X1 _9875_ (
    .A(reg_mscratch[24]),
    .B(_2056_),
    .S(_3026_),
    .Z(_0356_)
  );
  MUX2_X1 _9876_ (
    .A(reg_mscratch[25]),
    .B(_2102_),
    .S(_3026_),
    .Z(_0357_)
  );
  MUX2_X1 _9877_ (
    .A(reg_mscratch[26]),
    .B(_2148_),
    .S(_3026_),
    .Z(_0358_)
  );
  MUX2_X1 _9878_ (
    .A(reg_mscratch[27]),
    .B(_2195_),
    .S(_3026_),
    .Z(_0359_)
  );
  MUX2_X1 _9879_ (
    .A(reg_mscratch[28]),
    .B(_2241_),
    .S(_3026_),
    .Z(_0360_)
  );
  MUX2_X1 _9880_ (
    .A(reg_mscratch[29]),
    .B(_2285_),
    .S(_3026_),
    .Z(_0361_)
  );
  MUX2_X1 _9881_ (
    .A(reg_mscratch[30]),
    .B(_2435_),
    .S(_3026_),
    .Z(_0362_)
  );
  MUX2_X1 _9882_ (
    .A(reg_mscratch[31]),
    .B(_2365_),
    .S(_3026_),
    .Z(_0363_)
  );
  MUX2_X1 _9883_ (
    .A(reg_pmp_5_cfg_x),
    .B(_1647_),
    .S(_1075_),
    .Z(_0364_)
  );
  AND2_X1 _9884_ (
    .A1(reg_pmp_2_cfg_l),
    .A2(reg_pmp_2_cfg_a[0]),
    .ZN(_3027_)
  );
  AND2_X1 _9885_ (
    .A1(_0010_),
    .A2(_3027_),
    .ZN(_3028_)
  );
  OR2_X1 _9886_ (
    .A1(reg_pmp_1_cfg_l),
    .A2(_3028_),
    .ZN(_3029_)
  );
  OR2_X1 _9887_ (
    .A1(_0737_),
    .A2(_3029_),
    .ZN(_3030_)
  );
  OR2_X1 _9888_ (
    .A1(_0842_),
    .A2(_3030_),
    .ZN(_3031_)
  );
  MUX2_X1 _9889_ (
    .A(_1241_),
    .B(reg_pmp_1_addr[0]),
    .S(_3031_),
    .Z(_0365_)
  );
  MUX2_X1 _9890_ (
    .A(_1290_),
    .B(reg_pmp_1_addr[1]),
    .S(_3031_),
    .Z(_0366_)
  );
  MUX2_X1 _9891_ (
    .A(_1346_),
    .B(reg_pmp_1_addr[2]),
    .S(_3031_),
    .Z(_0367_)
  );
  MUX2_X1 _9892_ (
    .A(_1409_),
    .B(reg_pmp_1_addr[3]),
    .S(_3031_),
    .Z(_0368_)
  );
  MUX2_X1 _9893_ (
    .A(_1456_),
    .B(reg_pmp_1_addr[4]),
    .S(_3031_),
    .Z(_0369_)
  );
  MUX2_X1 _9894_ (
    .A(_1499_),
    .B(reg_pmp_1_addr[5]),
    .S(_3031_),
    .Z(_0370_)
  );
  MUX2_X1 _9895_ (
    .A(_1545_),
    .B(reg_pmp_1_addr[6]),
    .S(_3031_),
    .Z(_0371_)
  );
  MUX2_X1 _9896_ (
    .A(_1601_),
    .B(reg_pmp_1_addr[7]),
    .S(_3031_),
    .Z(_0372_)
  );
  MUX2_X1 _9897_ (
    .A(_1129_),
    .B(reg_pmp_1_addr[8]),
    .S(_3031_),
    .Z(_0373_)
  );
  MUX2_X1 _9898_ (
    .A(_1175_),
    .B(reg_pmp_1_addr[9]),
    .S(_3031_),
    .Z(_0374_)
  );
  MUX2_X1 _9899_ (
    .A(_1647_),
    .B(reg_pmp_1_addr[10]),
    .S(_3031_),
    .Z(_0375_)
  );
  MUX2_X1 _9900_ (
    .A(_1698_),
    .B(reg_pmp_1_addr[11]),
    .S(_3031_),
    .Z(_0376_)
  );
  MUX2_X1 _9901_ (
    .A(_1748_),
    .B(reg_pmp_1_addr[12]),
    .S(_3031_),
    .Z(_0377_)
  );
  MUX2_X1 _9902_ (
    .A(_1790_),
    .B(reg_pmp_1_addr[13]),
    .S(_3031_),
    .Z(_0378_)
  );
  MUX2_X1 _9903_ (
    .A(_1832_),
    .B(reg_pmp_1_addr[14]),
    .S(_3031_),
    .Z(_0379_)
  );
  MUX2_X1 _9904_ (
    .A(_1880_),
    .B(reg_pmp_1_addr[15]),
    .S(_3031_),
    .Z(_0380_)
  );
  MUX2_X1 _9905_ (
    .A(_0862_),
    .B(reg_pmp_1_addr[16]),
    .S(_3031_),
    .Z(_0381_)
  );
  MUX2_X1 _9906_ (
    .A(_1926_),
    .B(reg_pmp_1_addr[17]),
    .S(_3031_),
    .Z(_0382_)
  );
  MUX2_X1 _9907_ (
    .A(_0908_),
    .B(reg_pmp_1_addr[18]),
    .S(_3031_),
    .Z(_0383_)
  );
  MUX2_X1 _9908_ (
    .A(_0967_),
    .B(reg_pmp_1_addr[19]),
    .S(_3031_),
    .Z(_0384_)
  );
  MUX2_X1 _9909_ (
    .A(_1017_),
    .B(reg_pmp_1_addr[20]),
    .S(_3031_),
    .Z(_0385_)
  );
  MUX2_X1 _9910_ (
    .A(_1968_),
    .B(reg_pmp_1_addr[21]),
    .S(_3031_),
    .Z(_0386_)
  );
  MUX2_X1 _9911_ (
    .A(_2010_),
    .B(reg_pmp_1_addr[22]),
    .S(_3031_),
    .Z(_0387_)
  );
  MUX2_X1 _9912_ (
    .A(_1071_),
    .B(reg_pmp_1_addr[23]),
    .S(_3031_),
    .Z(_0388_)
  );
  MUX2_X1 _9913_ (
    .A(_2056_),
    .B(reg_pmp_1_addr[24]),
    .S(_3031_),
    .Z(_0389_)
  );
  MUX2_X1 _9914_ (
    .A(_2102_),
    .B(reg_pmp_1_addr[25]),
    .S(_3031_),
    .Z(_0390_)
  );
  MUX2_X1 _9915_ (
    .A(_2148_),
    .B(reg_pmp_1_addr[26]),
    .S(_3031_),
    .Z(_0391_)
  );
  DFF_X1 \io_status_cease_r$_SDFF_PP0_  (
    .CK(clock),
    .D(_0021_),
    .Q(io_status_cease_r),
    .QN(_5008_)
  );
  DFF_X1 \large_1[0]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0569_),
    .Q(large_1[0]),
    .QN(_large_r_T_3[0])
  );
  DFF_X1 \large_1[10]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0579_),
    .Q(large_1[10]),
    .QN(_4471_)
  );
  DFF_X1 \large_1[11]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0580_),
    .Q(large_1[11]),
    .QN(_4470_)
  );
  DFF_X1 \large_1[12]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0581_),
    .Q(large_1[12]),
    .QN(_4469_)
  );
  DFF_X1 \large_1[13]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0582_),
    .Q(large_1[13]),
    .QN(_4468_)
  );
  DFF_X1 \large_1[14]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0583_),
    .Q(large_1[14]),
    .QN(_4467_)
  );
  DFF_X1 \large_1[15]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0584_),
    .Q(large_1[15]),
    .QN(_4466_)
  );
  DFF_X1 \large_1[16]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0585_),
    .Q(large_1[16]),
    .QN(_4465_)
  );
  DFF_X1 \large_1[17]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0586_),
    .Q(large_1[17]),
    .QN(_4464_)
  );
  DFF_X1 \large_1[18]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0587_),
    .Q(large_1[18]),
    .QN(_4463_)
  );
  DFF_X1 \large_1[19]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0588_),
    .Q(large_1[19]),
    .QN(_4462_)
  );
  DFF_X1 \large_1[1]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0570_),
    .Q(large_1[1]),
    .QN(_4480_)
  );
  DFF_X1 \large_1[20]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0589_),
    .Q(large_1[20]),
    .QN(_4461_)
  );
  DFF_X1 \large_1[21]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0590_),
    .Q(large_1[21]),
    .QN(_4460_)
  );
  DFF_X1 \large_1[22]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0591_),
    .Q(large_1[22]),
    .QN(_4459_)
  );
  DFF_X1 \large_1[23]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0592_),
    .Q(large_1[23]),
    .QN(_4458_)
  );
  DFF_X1 \large_1[24]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0593_),
    .Q(large_1[24]),
    .QN(_4457_)
  );
  DFF_X1 \large_1[25]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0594_),
    .Q(large_1[25]),
    .QN(_4456_)
  );
  DFF_X1 \large_1[26]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0294_),
    .Q(large_1[26]),
    .QN(_4751_)
  );
  DFF_X1 \large_1[27]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0295_),
    .Q(large_1[27]),
    .QN(_4750_)
  );
  DFF_X1 \large_1[28]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0296_),
    .Q(large_1[28]),
    .QN(_4749_)
  );
  DFF_X1 \large_1[29]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0297_),
    .Q(large_1[29]),
    .QN(_4748_)
  );
  DFF_X1 \large_1[2]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0571_),
    .Q(large_1[2]),
    .QN(_4479_)
  );
  DFF_X1 \large_1[30]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0298_),
    .Q(large_1[30]),
    .QN(_4747_)
  );
  DFF_X1 \large_1[31]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0299_),
    .Q(large_1[31]),
    .QN(_4746_)
  );
  DFF_X1 \large_1[32]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0300_),
    .Q(large_1[32]),
    .QN(_4745_)
  );
  DFF_X1 \large_1[33]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0301_),
    .Q(large_1[33]),
    .QN(_4744_)
  );
  DFF_X1 \large_1[34]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0302_),
    .Q(large_1[34]),
    .QN(_4743_)
  );
  DFF_X1 \large_1[35]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0303_),
    .Q(large_1[35]),
    .QN(_4742_)
  );
  DFF_X1 \large_1[36]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0304_),
    .Q(large_1[36]),
    .QN(_4741_)
  );
  DFF_X1 \large_1[37]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0305_),
    .Q(large_1[37]),
    .QN(_4740_)
  );
  DFF_X1 \large_1[38]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0306_),
    .Q(large_1[38]),
    .QN(_4739_)
  );
  DFF_X1 \large_1[39]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0307_),
    .Q(large_1[39]),
    .QN(_4738_)
  );
  DFF_X1 \large_1[3]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0572_),
    .Q(large_1[3]),
    .QN(_4478_)
  );
  DFF_X1 \large_1[40]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0308_),
    .Q(large_1[40]),
    .QN(_4737_)
  );
  DFF_X1 \large_1[41]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0309_),
    .Q(large_1[41]),
    .QN(_4736_)
  );
  DFF_X1 \large_1[42]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0310_),
    .Q(large_1[42]),
    .QN(_4735_)
  );
  DFF_X1 \large_1[43]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0311_),
    .Q(large_1[43]),
    .QN(_4734_)
  );
  DFF_X1 \large_1[44]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0312_),
    .Q(large_1[44]),
    .QN(_4733_)
  );
  DFF_X1 \large_1[45]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0313_),
    .Q(large_1[45]),
    .QN(_4732_)
  );
  DFF_X1 \large_1[46]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0314_),
    .Q(large_1[46]),
    .QN(_4731_)
  );
  DFF_X1 \large_1[47]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0315_),
    .Q(large_1[47]),
    .QN(_4730_)
  );
  DFF_X1 \large_1[48]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0316_),
    .Q(large_1[48]),
    .QN(_4729_)
  );
  DFF_X1 \large_1[49]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0317_),
    .Q(large_1[49]),
    .QN(_4728_)
  );
  DFF_X1 \large_1[4]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0573_),
    .Q(large_1[4]),
    .QN(_4477_)
  );
  DFF_X1 \large_1[50]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0318_),
    .Q(large_1[50]),
    .QN(_4727_)
  );
  DFF_X1 \large_1[51]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0319_),
    .Q(large_1[51]),
    .QN(_4726_)
  );
  DFF_X1 \large_1[52]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0320_),
    .Q(large_1[52]),
    .QN(_4725_)
  );
  DFF_X1 \large_1[53]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0321_),
    .Q(large_1[53]),
    .QN(_4724_)
  );
  DFF_X1 \large_1[54]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0322_),
    .Q(large_1[54]),
    .QN(_4723_)
  );
  DFF_X1 \large_1[55]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0323_),
    .Q(large_1[55]),
    .QN(_4722_)
  );
  DFF_X1 \large_1[56]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0324_),
    .Q(large_1[56]),
    .QN(_4721_)
  );
  DFF_X1 \large_1[57]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0325_),
    .Q(large_1[57]),
    .QN(_4720_)
  );
  DFF_X1 \large_1[5]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0574_),
    .Q(large_1[5]),
    .QN(_4476_)
  );
  DFF_X1 \large_1[6]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0575_),
    .Q(large_1[6]),
    .QN(_4475_)
  );
  DFF_X1 \large_1[7]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0576_),
    .Q(large_1[7]),
    .QN(_4474_)
  );
  DFF_X1 \large_1[8]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0577_),
    .Q(large_1[8]),
    .QN(_4473_)
  );
  DFF_X1 \large_1[9]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0578_),
    .Q(large_1[9]),
    .QN(_4472_)
  );
  DFF_X1 \large_[0]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0595_),
    .Q(large_[0]),
    .QN(_large_r_T_1[0])
  );
  DFF_X1 \large_[10]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0605_),
    .Q(large_[10]),
    .QN(_4446_)
  );
  DFF_X1 \large_[11]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0606_),
    .Q(large_[11]),
    .QN(_4445_)
  );
  DFF_X1 \large_[12]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0607_),
    .Q(large_[12]),
    .QN(_4444_)
  );
  DFF_X1 \large_[13]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0608_),
    .Q(large_[13]),
    .QN(_4443_)
  );
  DFF_X1 \large_[14]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0609_),
    .Q(large_[14]),
    .QN(_4442_)
  );
  DFF_X1 \large_[15]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0610_),
    .Q(large_[15]),
    .QN(_4441_)
  );
  DFF_X1 \large_[16]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0611_),
    .Q(large_[16]),
    .QN(_4440_)
  );
  DFF_X1 \large_[17]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0612_),
    .Q(large_[17]),
    .QN(_4439_)
  );
  DFF_X1 \large_[18]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0613_),
    .Q(large_[18]),
    .QN(_4438_)
  );
  DFF_X1 \large_[19]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0614_),
    .Q(large_[19]),
    .QN(_4437_)
  );
  DFF_X1 \large_[1]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0596_),
    .Q(large_[1]),
    .QN(_4455_)
  );
  DFF_X1 \large_[20]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0615_),
    .Q(large_[20]),
    .QN(_4436_)
  );
  DFF_X1 \large_[21]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0616_),
    .Q(large_[21]),
    .QN(_4435_)
  );
  DFF_X1 \large_[22]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0617_),
    .Q(large_[22]),
    .QN(_4434_)
  );
  DFF_X1 \large_[23]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0618_),
    .Q(large_[23]),
    .QN(_4433_)
  );
  DFF_X1 \large_[24]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0619_),
    .Q(large_[24]),
    .QN(_4432_)
  );
  DFF_X1 \large_[25]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0620_),
    .Q(large_[25]),
    .QN(_4431_)
  );
  DFF_X1 \large_[26]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0429_),
    .Q(large_[26]),
    .QN(_4617_)
  );
  DFF_X1 \large_[27]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0430_),
    .Q(large_[27]),
    .QN(_4616_)
  );
  DFF_X1 \large_[28]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0431_),
    .Q(large_[28]),
    .QN(_4615_)
  );
  DFF_X1 \large_[29]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0432_),
    .Q(large_[29]),
    .QN(_4614_)
  );
  DFF_X1 \large_[2]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0597_),
    .Q(large_[2]),
    .QN(_4454_)
  );
  DFF_X1 \large_[30]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0433_),
    .Q(large_[30]),
    .QN(_4613_)
  );
  DFF_X1 \large_[31]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0434_),
    .Q(large_[31]),
    .QN(_4612_)
  );
  DFF_X1 \large_[32]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0435_),
    .Q(large_[32]),
    .QN(_4611_)
  );
  DFF_X1 \large_[33]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0436_),
    .Q(large_[33]),
    .QN(_4610_)
  );
  DFF_X1 \large_[34]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0437_),
    .Q(large_[34]),
    .QN(_4609_)
  );
  DFF_X1 \large_[35]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0438_),
    .Q(large_[35]),
    .QN(_4608_)
  );
  DFF_X1 \large_[36]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0439_),
    .Q(large_[36]),
    .QN(_4607_)
  );
  DFF_X1 \large_[37]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0440_),
    .Q(large_[37]),
    .QN(_4606_)
  );
  DFF_X1 \large_[38]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0441_),
    .Q(large_[38]),
    .QN(_4605_)
  );
  DFF_X1 \large_[39]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0442_),
    .Q(large_[39]),
    .QN(_4604_)
  );
  DFF_X1 \large_[3]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0598_),
    .Q(large_[3]),
    .QN(_4453_)
  );
  DFF_X1 \large_[40]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0443_),
    .Q(large_[40]),
    .QN(_4603_)
  );
  DFF_X1 \large_[41]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0444_),
    .Q(large_[41]),
    .QN(_4602_)
  );
  DFF_X1 \large_[42]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0445_),
    .Q(large_[42]),
    .QN(_4601_)
  );
  DFF_X1 \large_[43]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0446_),
    .Q(large_[43]),
    .QN(_4600_)
  );
  DFF_X1 \large_[44]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0447_),
    .Q(large_[44]),
    .QN(_4599_)
  );
  DFF_X1 \large_[45]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0448_),
    .Q(large_[45]),
    .QN(_4598_)
  );
  DFF_X1 \large_[46]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0449_),
    .Q(large_[46]),
    .QN(_4597_)
  );
  DFF_X1 \large_[47]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0450_),
    .Q(large_[47]),
    .QN(_4596_)
  );
  DFF_X1 \large_[48]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0451_),
    .Q(large_[48]),
    .QN(_4595_)
  );
  DFF_X1 \large_[49]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0452_),
    .Q(large_[49]),
    .QN(_4594_)
  );
  DFF_X1 \large_[4]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0599_),
    .Q(large_[4]),
    .QN(_4452_)
  );
  DFF_X1 \large_[50]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0453_),
    .Q(large_[50]),
    .QN(_4593_)
  );
  DFF_X1 \large_[51]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0454_),
    .Q(large_[51]),
    .QN(_4592_)
  );
  DFF_X1 \large_[52]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0455_),
    .Q(large_[52]),
    .QN(_4591_)
  );
  DFF_X1 \large_[53]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0456_),
    .Q(large_[53]),
    .QN(_4590_)
  );
  DFF_X1 \large_[54]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0457_),
    .Q(large_[54]),
    .QN(_4589_)
  );
  DFF_X1 \large_[55]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0458_),
    .Q(large_[55]),
    .QN(_4588_)
  );
  DFF_X1 \large_[56]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0459_),
    .Q(large_[56]),
    .QN(_4587_)
  );
  DFF_X1 \large_[57]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0460_),
    .Q(large_[57]),
    .QN(_4586_)
  );
  DFF_X1 \large_[5]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0600_),
    .Q(large_[5]),
    .QN(_4451_)
  );
  DFF_X1 \large_[6]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0601_),
    .Q(large_[6]),
    .QN(_4450_)
  );
  DFF_X1 \large_[7]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0602_),
    .Q(large_[7]),
    .QN(_4449_)
  );
  DFF_X1 \large_[8]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0603_),
    .Q(large_[8]),
    .QN(_4448_)
  );
  DFF_X1 \large_[9]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0604_),
    .Q(large_[9]),
    .QN(_4447_)
  );
  DFF_X1 \reg_bp_0_address[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_0207_),
    .Q(reg_bp_0_address[0]),
    .QN(_4834_)
  );
  DFF_X1 \reg_bp_0_address[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_0217_),
    .Q(reg_bp_0_address[10]),
    .QN(_4824_)
  );
  DFF_X1 \reg_bp_0_address[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_0218_),
    .Q(reg_bp_0_address[11]),
    .QN(_4823_)
  );
  DFF_X1 \reg_bp_0_address[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_0219_),
    .Q(reg_bp_0_address[12]),
    .QN(_4822_)
  );
  DFF_X1 \reg_bp_0_address[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_0220_),
    .Q(reg_bp_0_address[13]),
    .QN(_4821_)
  );
  DFF_X1 \reg_bp_0_address[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_0221_),
    .Q(reg_bp_0_address[14]),
    .QN(_4820_)
  );
  DFF_X1 \reg_bp_0_address[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_0222_),
    .Q(reg_bp_0_address[15]),
    .QN(_4819_)
  );
  DFF_X1 \reg_bp_0_address[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_0223_),
    .Q(reg_bp_0_address[16]),
    .QN(_4818_)
  );
  DFF_X1 \reg_bp_0_address[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_0224_),
    .Q(reg_bp_0_address[17]),
    .QN(_4817_)
  );
  DFF_X1 \reg_bp_0_address[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_0225_),
    .Q(reg_bp_0_address[18]),
    .QN(_4816_)
  );
  DFF_X1 \reg_bp_0_address[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_0226_),
    .Q(reg_bp_0_address[19]),
    .QN(_4815_)
  );
  DFF_X1 \reg_bp_0_address[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_0208_),
    .Q(reg_bp_0_address[1]),
    .QN(_4833_)
  );
  DFF_X1 \reg_bp_0_address[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_0227_),
    .Q(reg_bp_0_address[20]),
    .QN(_4814_)
  );
  DFF_X1 \reg_bp_0_address[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_0228_),
    .Q(reg_bp_0_address[21]),
    .QN(_4813_)
  );
  DFF_X1 \reg_bp_0_address[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_0229_),
    .Q(reg_bp_0_address[22]),
    .QN(_4812_)
  );
  DFF_X1 \reg_bp_0_address[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_0230_),
    .Q(reg_bp_0_address[23]),
    .QN(_4811_)
  );
  DFF_X1 \reg_bp_0_address[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_0231_),
    .Q(reg_bp_0_address[24]),
    .QN(_4810_)
  );
  DFF_X1 \reg_bp_0_address[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_0232_),
    .Q(reg_bp_0_address[25]),
    .QN(_4809_)
  );
  DFF_X1 \reg_bp_0_address[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_0233_),
    .Q(reg_bp_0_address[26]),
    .QN(_4808_)
  );
  DFF_X1 \reg_bp_0_address[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_0234_),
    .Q(reg_bp_0_address[27]),
    .QN(_4807_)
  );
  DFF_X1 \reg_bp_0_address[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_0235_),
    .Q(reg_bp_0_address[28]),
    .QN(_4806_)
  );
  DFF_X1 \reg_bp_0_address[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_0236_),
    .Q(reg_bp_0_address[29]),
    .QN(_4805_)
  );
  DFF_X1 \reg_bp_0_address[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_0209_),
    .Q(reg_bp_0_address[2]),
    .QN(_4832_)
  );
  DFF_X1 \reg_bp_0_address[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_0237_),
    .Q(reg_bp_0_address[30]),
    .QN(_4804_)
  );
  DFF_X1 \reg_bp_0_address[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_0238_),
    .Q(reg_bp_0_address[31]),
    .QN(_4803_)
  );
  DFF_X1 \reg_bp_0_address[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_0210_),
    .Q(reg_bp_0_address[3]),
    .QN(_4831_)
  );
  DFF_X1 \reg_bp_0_address[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_0211_),
    .Q(reg_bp_0_address[4]),
    .QN(_4830_)
  );
  DFF_X1 \reg_bp_0_address[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_0212_),
    .Q(reg_bp_0_address[5]),
    .QN(_4829_)
  );
  DFF_X1 \reg_bp_0_address[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_0213_),
    .Q(reg_bp_0_address[6]),
    .QN(_4828_)
  );
  DFF_X1 \reg_bp_0_address[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_0214_),
    .Q(reg_bp_0_address[7]),
    .QN(_4827_)
  );
  DFF_X1 \reg_bp_0_address[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_0215_),
    .Q(reg_bp_0_address[8]),
    .QN(_4826_)
  );
  DFF_X1 \reg_bp_0_address[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_0216_),
    .Q(reg_bp_0_address[9]),
    .QN(_4825_)
  );
  DFF_X1 \reg_bp_0_control_action$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0248_),
    .Q(reg_bp_0_control_action),
    .QN(_4794_)
  );
  DFF_X1 \reg_bp_0_control_dmode$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0249_),
    .Q(reg_bp_0_control_dmode),
    .QN(_0005_)
  );
  DFF_X1 \reg_bp_0_control_r$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0244_),
    .Q(reg_bp_0_control_r),
    .QN(_4798_)
  );
  DFF_X1 \reg_bp_0_control_tmatch[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_0242_),
    .Q(reg_bp_0_control_tmatch[0]),
    .QN(_4800_)
  );
  DFF_X1 \reg_bp_0_control_tmatch[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_0243_),
    .Q(reg_bp_0_control_tmatch[1]),
    .QN(_4799_)
  );
  DFF_X1 \reg_bp_0_control_w$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0245_),
    .Q(reg_bp_0_control_w),
    .QN(_4797_)
  );
  DFF_X1 \reg_bp_0_control_x$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0246_),
    .Q(reg_bp_0_control_x),
    .QN(_4796_)
  );
  DFF_X1 \reg_custom_0[3]$_SDFFE_PP1P_  (
    .CK(clock),
    .D(_0425_),
    .Q(reg_custom_0[3]),
    .QN(_4620_)
  );
  DFF_X1 \reg_dcsr_cause[0]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0285_),
    .Q(reg_dcsr_cause[0]),
    .QN(_4758_)
  );
  DFF_X1 \reg_dcsr_cause[1]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0286_),
    .Q(reg_dcsr_cause[1]),
    .QN(_4757_)
  );
  DFF_X1 \reg_dcsr_cause[2]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0287_),
    .Q(reg_dcsr_cause[2]),
    .QN(_4756_)
  );
  DFF_X1 \reg_dcsr_ebreakm$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0288_),
    .Q(reg_dcsr_ebreakm),
    .QN(_4755_)
  );
  DFF_X1 \reg_dcsr_step$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0284_),
    .Q(reg_dcsr_step),
    .QN(_4759_)
  );
  DFF_X1 \reg_debug$_SDFF_PP0_  (
    .CK(clock),
    .D(_0282_),
    .Q(reg_debug),
    .QN(_io_decode_0_read_illegal_T_15)
  );
  DFF_X1 \reg_dpc[10]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[10]),
    .Q(reg_dpc[10]),
    .QN(_5019_)
  );
  DFF_X1 \reg_dpc[11]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[11]),
    .Q(reg_dpc[11]),
    .QN(_5020_)
  );
  DFF_X1 \reg_dpc[12]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[12]),
    .Q(reg_dpc[12]),
    .QN(_5021_)
  );
  DFF_X1 \reg_dpc[13]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[13]),
    .Q(reg_dpc[13]),
    .QN(_5022_)
  );
  DFF_X1 \reg_dpc[14]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[14]),
    .Q(reg_dpc[14]),
    .QN(_5023_)
  );
  DFF_X1 \reg_dpc[15]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[15]),
    .Q(reg_dpc[15]),
    .QN(_5024_)
  );
  DFF_X1 \reg_dpc[16]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[16]),
    .Q(reg_dpc[16]),
    .QN(_5025_)
  );
  DFF_X1 \reg_dpc[17]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[17]),
    .Q(reg_dpc[17]),
    .QN(_5026_)
  );
  DFF_X1 \reg_dpc[18]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[18]),
    .Q(reg_dpc[18]),
    .QN(_5027_)
  );
  DFF_X1 \reg_dpc[19]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[19]),
    .Q(reg_dpc[19]),
    .QN(_5028_)
  );
  DFF_X1 \reg_dpc[1]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[1]),
    .Q(reg_dpc[1]),
    .QN(_T_24[1])
  );
  DFF_X1 \reg_dpc[20]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[20]),
    .Q(reg_dpc[20]),
    .QN(_5029_)
  );
  DFF_X1 \reg_dpc[21]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[21]),
    .Q(reg_dpc[21]),
    .QN(_5030_)
  );
  DFF_X1 \reg_dpc[22]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[22]),
    .Q(reg_dpc[22]),
    .QN(_5031_)
  );
  DFF_X1 \reg_dpc[23]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[23]),
    .Q(reg_dpc[23]),
    .QN(_5032_)
  );
  DFF_X1 \reg_dpc[24]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[24]),
    .Q(reg_dpc[24]),
    .QN(_5033_)
  );
  DFF_X1 \reg_dpc[25]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[25]),
    .Q(reg_dpc[25]),
    .QN(_5034_)
  );
  DFF_X1 \reg_dpc[26]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[26]),
    .Q(reg_dpc[26]),
    .QN(_5035_)
  );
  DFF_X1 \reg_dpc[27]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[27]),
    .Q(reg_dpc[27]),
    .QN(_5036_)
  );
  DFF_X1 \reg_dpc[28]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[28]),
    .Q(reg_dpc[28]),
    .QN(_5037_)
  );
  DFF_X1 \reg_dpc[29]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[29]),
    .Q(reg_dpc[29]),
    .QN(_5038_)
  );
  DFF_X1 \reg_dpc[2]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[2]),
    .Q(reg_dpc[2]),
    .QN(_5011_)
  );
  DFF_X1 \reg_dpc[30]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[30]),
    .Q(reg_dpc[30]),
    .QN(_5039_)
  );
  DFF_X1 \reg_dpc[31]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[31]),
    .Q(reg_dpc[31]),
    .QN(_4761_)
  );
  DFF_X1 \reg_dpc[3]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[3]),
    .Q(reg_dpc[3]),
    .QN(_5012_)
  );
  DFF_X1 \reg_dpc[4]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[4]),
    .Q(reg_dpc[4]),
    .QN(_5013_)
  );
  DFF_X1 \reg_dpc[5]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[5]),
    .Q(reg_dpc[5]),
    .QN(_5014_)
  );
  DFF_X1 \reg_dpc[6]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[6]),
    .Q(reg_dpc[6]),
    .QN(_5015_)
  );
  DFF_X1 \reg_dpc[7]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[7]),
    .Q(reg_dpc[7]),
    .QN(_5016_)
  );
  DFF_X1 \reg_dpc[8]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[8]),
    .Q(reg_dpc[8]),
    .QN(_5017_)
  );
  DFF_X1 \reg_dpc[9]$_DFF_P_  (
    .CK(clock),
    .D(_0000_[9]),
    .Q(reg_dpc[9]),
    .QN(_5018_)
  );
  DFF_X1 \reg_dscratch0[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_0250_),
    .Q(reg_dscratch0[0]),
    .QN(_4793_)
  );
  DFF_X1 \reg_dscratch0[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_0260_),
    .Q(reg_dscratch0[10]),
    .QN(_4783_)
  );
  DFF_X1 \reg_dscratch0[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_0261_),
    .Q(reg_dscratch0[11]),
    .QN(_4782_)
  );
  DFF_X1 \reg_dscratch0[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_0262_),
    .Q(reg_dscratch0[12]),
    .QN(_4781_)
  );
  DFF_X1 \reg_dscratch0[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_0263_),
    .Q(reg_dscratch0[13]),
    .QN(_4780_)
  );
  DFF_X1 \reg_dscratch0[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_0264_),
    .Q(reg_dscratch0[14]),
    .QN(_4779_)
  );
  DFF_X1 \reg_dscratch0[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_0265_),
    .Q(reg_dscratch0[15]),
    .QN(_4778_)
  );
  DFF_X1 \reg_dscratch0[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_0266_),
    .Q(reg_dscratch0[16]),
    .QN(_4777_)
  );
  DFF_X1 \reg_dscratch0[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_0267_),
    .Q(reg_dscratch0[17]),
    .QN(_4776_)
  );
  DFF_X1 \reg_dscratch0[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_0268_),
    .Q(reg_dscratch0[18]),
    .QN(_4775_)
  );
  DFF_X1 \reg_dscratch0[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_0269_),
    .Q(reg_dscratch0[19]),
    .QN(_4774_)
  );
  DFF_X1 \reg_dscratch0[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_0251_),
    .Q(reg_dscratch0[1]),
    .QN(_4792_)
  );
  DFF_X1 \reg_dscratch0[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_0270_),
    .Q(reg_dscratch0[20]),
    .QN(_4773_)
  );
  DFF_X1 \reg_dscratch0[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_0271_),
    .Q(reg_dscratch0[21]),
    .QN(_4772_)
  );
  DFF_X1 \reg_dscratch0[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_0272_),
    .Q(reg_dscratch0[22]),
    .QN(_4771_)
  );
  DFF_X1 \reg_dscratch0[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_0273_),
    .Q(reg_dscratch0[23]),
    .QN(_4770_)
  );
  DFF_X1 \reg_dscratch0[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_0274_),
    .Q(reg_dscratch0[24]),
    .QN(_4769_)
  );
  DFF_X1 \reg_dscratch0[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_0275_),
    .Q(reg_dscratch0[25]),
    .QN(_4768_)
  );
  DFF_X1 \reg_dscratch0[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_0276_),
    .Q(reg_dscratch0[26]),
    .QN(_4767_)
  );
  DFF_X1 \reg_dscratch0[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_0277_),
    .Q(reg_dscratch0[27]),
    .QN(_4766_)
  );
  DFF_X1 \reg_dscratch0[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_0278_),
    .Q(reg_dscratch0[28]),
    .QN(_4765_)
  );
  DFF_X1 \reg_dscratch0[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_0279_),
    .Q(reg_dscratch0[29]),
    .QN(_4764_)
  );
  DFF_X1 \reg_dscratch0[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_0252_),
    .Q(reg_dscratch0[2]),
    .QN(_4791_)
  );
  DFF_X1 \reg_dscratch0[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_0280_),
    .Q(reg_dscratch0[30]),
    .QN(_4763_)
  );
  DFF_X1 \reg_dscratch0[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_0281_),
    .Q(reg_dscratch0[31]),
    .QN(_4762_)
  );
  DFF_X1 \reg_dscratch0[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_0253_),
    .Q(reg_dscratch0[3]),
    .QN(_4790_)
  );
  DFF_X1 \reg_dscratch0[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_0254_),
    .Q(reg_dscratch0[4]),
    .QN(_4789_)
  );
  DFF_X1 \reg_dscratch0[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_0255_),
    .Q(reg_dscratch0[5]),
    .QN(_4788_)
  );
  DFF_X1 \reg_dscratch0[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_0256_),
    .Q(reg_dscratch0[6]),
    .QN(_4787_)
  );
  DFF_X1 \reg_dscratch0[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_0257_),
    .Q(reg_dscratch0[7]),
    .QN(_4786_)
  );
  DFF_X1 \reg_dscratch0[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_0258_),
    .Q(reg_dscratch0[8]),
    .QN(_4785_)
  );
  DFF_X1 \reg_dscratch0[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_0259_),
    .Q(reg_dscratch0[9]),
    .QN(_4784_)
  );
  DFF_X1 \reg_mcause[0]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0498_),
    .Q(reg_mcause[0]),
    .QN(_4549_)
  );
  DFF_X1 \reg_mcause[10]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0508_),
    .Q(reg_mcause[10]),
    .QN(_4539_)
  );
  DFF_X1 \reg_mcause[11]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0509_),
    .Q(reg_mcause[11]),
    .QN(_4538_)
  );
  DFF_X1 \reg_mcause[12]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0510_),
    .Q(reg_mcause[12]),
    .QN(_4537_)
  );
  DFF_X1 \reg_mcause[13]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0511_),
    .Q(reg_mcause[13]),
    .QN(_4536_)
  );
  DFF_X1 \reg_mcause[14]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0512_),
    .Q(reg_mcause[14]),
    .QN(_4535_)
  );
  DFF_X1 \reg_mcause[15]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0513_),
    .Q(reg_mcause[15]),
    .QN(_4534_)
  );
  DFF_X1 \reg_mcause[16]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0514_),
    .Q(reg_mcause[16]),
    .QN(_4533_)
  );
  DFF_X1 \reg_mcause[17]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0515_),
    .Q(reg_mcause[17]),
    .QN(_4532_)
  );
  DFF_X1 \reg_mcause[18]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0516_),
    .Q(reg_mcause[18]),
    .QN(_4531_)
  );
  DFF_X1 \reg_mcause[19]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0517_),
    .Q(reg_mcause[19]),
    .QN(_4530_)
  );
  DFF_X1 \reg_mcause[1]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0499_),
    .Q(reg_mcause[1]),
    .QN(_4548_)
  );
  DFF_X1 \reg_mcause[20]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0518_),
    .Q(reg_mcause[20]),
    .QN(_4529_)
  );
  DFF_X1 \reg_mcause[21]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0519_),
    .Q(reg_mcause[21]),
    .QN(_4528_)
  );
  DFF_X1 \reg_mcause[22]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0520_),
    .Q(reg_mcause[22]),
    .QN(_4527_)
  );
  DFF_X1 \reg_mcause[23]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0521_),
    .Q(reg_mcause[23]),
    .QN(_4526_)
  );
  DFF_X1 \reg_mcause[24]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0522_),
    .Q(reg_mcause[24]),
    .QN(_4525_)
  );
  DFF_X1 \reg_mcause[25]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0523_),
    .Q(reg_mcause[25]),
    .QN(_4524_)
  );
  DFF_X1 \reg_mcause[26]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0524_),
    .Q(reg_mcause[26]),
    .QN(_4523_)
  );
  DFF_X1 \reg_mcause[27]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0525_),
    .Q(reg_mcause[27]),
    .QN(_4522_)
  );
  DFF_X1 \reg_mcause[28]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0526_),
    .Q(reg_mcause[28]),
    .QN(_4521_)
  );
  DFF_X1 \reg_mcause[29]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0527_),
    .Q(reg_mcause[29]),
    .QN(_4520_)
  );
  DFF_X1 \reg_mcause[2]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0500_),
    .Q(reg_mcause[2]),
    .QN(_4547_)
  );
  DFF_X1 \reg_mcause[30]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0528_),
    .Q(reg_mcause[30]),
    .QN(_4519_)
  );
  DFF_X1 \reg_mcause[31]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0529_),
    .Q(reg_mcause[31]),
    .QN(_5040_)
  );
  DFF_X1 \reg_mcause[3]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0501_),
    .Q(reg_mcause[3]),
    .QN(_4546_)
  );
  DFF_X1 \reg_mcause[4]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0502_),
    .Q(reg_mcause[4]),
    .QN(_4545_)
  );
  DFF_X1 \reg_mcause[5]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0503_),
    .Q(reg_mcause[5]),
    .QN(_4544_)
  );
  DFF_X1 \reg_mcause[6]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0504_),
    .Q(reg_mcause[6]),
    .QN(_4543_)
  );
  DFF_X1 \reg_mcause[7]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0505_),
    .Q(reg_mcause[7]),
    .QN(_4542_)
  );
  DFF_X1 \reg_mcause[8]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0506_),
    .Q(reg_mcause[8]),
    .QN(_4541_)
  );
  DFF_X1 \reg_mcause[9]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0507_),
    .Q(reg_mcause[9]),
    .QN(_4540_)
  );
  DFF_X1 \reg_mcountinhibit[0]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0290_),
    .Q(reg_mcountinhibit[0]),
    .QN(_T_15)
  );
  DFF_X1 \reg_mcountinhibit[2]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0291_),
    .Q(reg_mcountinhibit[2]),
    .QN(_T_14)
  );
  DFF_X1 \reg_mepc[10]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[10]),
    .Q(reg_mepc[10]),
    .QN(_5081_)
  );
  DFF_X1 \reg_mepc[11]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[11]),
    .Q(reg_mepc[11]),
    .QN(_5082_)
  );
  DFF_X1 \reg_mepc[12]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[12]),
    .Q(reg_mepc[12]),
    .QN(_5083_)
  );
  DFF_X1 \reg_mepc[13]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[13]),
    .Q(reg_mepc[13]),
    .QN(_5084_)
  );
  DFF_X1 \reg_mepc[14]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[14]),
    .Q(reg_mepc[14]),
    .QN(_5085_)
  );
  DFF_X1 \reg_mepc[15]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[15]),
    .Q(reg_mepc[15]),
    .QN(_5086_)
  );
  DFF_X1 \reg_mepc[16]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[16]),
    .Q(reg_mepc[16]),
    .QN(_5087_)
  );
  DFF_X1 \reg_mepc[17]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[17]),
    .Q(reg_mepc[17]),
    .QN(_5088_)
  );
  DFF_X1 \reg_mepc[18]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[18]),
    .Q(reg_mepc[18]),
    .QN(_5089_)
  );
  DFF_X1 \reg_mepc[19]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[19]),
    .Q(reg_mepc[19]),
    .QN(_5090_)
  );
  DFF_X1 \reg_mepc[1]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[1]),
    .Q(reg_mepc[1]),
    .QN(_T_18[1])
  );
  DFF_X1 \reg_mepc[20]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[20]),
    .Q(reg_mepc[20]),
    .QN(_5091_)
  );
  DFF_X1 \reg_mepc[21]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[21]),
    .Q(reg_mepc[21]),
    .QN(_5092_)
  );
  DFF_X1 \reg_mepc[22]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[22]),
    .Q(reg_mepc[22]),
    .QN(_5093_)
  );
  DFF_X1 \reg_mepc[23]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[23]),
    .Q(reg_mepc[23]),
    .QN(_5094_)
  );
  DFF_X1 \reg_mepc[24]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[24]),
    .Q(reg_mepc[24]),
    .QN(_5095_)
  );
  DFF_X1 \reg_mepc[25]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[25]),
    .Q(reg_mepc[25]),
    .QN(_5096_)
  );
  DFF_X1 \reg_mepc[26]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[26]),
    .Q(reg_mepc[26]),
    .QN(_5097_)
  );
  DFF_X1 \reg_mepc[27]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[27]),
    .Q(reg_mepc[27]),
    .QN(_5098_)
  );
  DFF_X1 \reg_mepc[28]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[28]),
    .Q(reg_mepc[28]),
    .QN(_5099_)
  );
  DFF_X1 \reg_mepc[29]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[29]),
    .Q(reg_mepc[29]),
    .QN(_5100_)
  );
  DFF_X1 \reg_mepc[2]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[2]),
    .Q(reg_mepc[2]),
    .QN(_5073_)
  );
  DFF_X1 \reg_mepc[30]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[30]),
    .Q(reg_mepc[30]),
    .QN(_5101_)
  );
  DFF_X1 \reg_mepc[31]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[31]),
    .Q(reg_mepc[31]),
    .QN(_4518_)
  );
  DFF_X1 \reg_mepc[3]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[3]),
    .Q(reg_mepc[3]),
    .QN(_5074_)
  );
  DFF_X1 \reg_mepc[4]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[4]),
    .Q(reg_mepc[4]),
    .QN(_5075_)
  );
  DFF_X1 \reg_mepc[5]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[5]),
    .Q(reg_mepc[5]),
    .QN(_5076_)
  );
  DFF_X1 \reg_mepc[6]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[6]),
    .Q(reg_mepc[6]),
    .QN(_5077_)
  );
  DFF_X1 \reg_mepc[7]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[7]),
    .Q(reg_mepc[7]),
    .QN(_5078_)
  );
  DFF_X1 \reg_mepc[8]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[8]),
    .Q(reg_mepc[8]),
    .QN(_5079_)
  );
  DFF_X1 \reg_mepc[9]$_DFF_P_  (
    .CK(clock),
    .D(_0001_[9]),
    .Q(reg_mepc[9]),
    .QN(_5080_)
  );
  DFF_X1 \reg_mie[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_0532_),
    .Q(reg_mie[11]),
    .QN(_4515_)
  );
  DFF_X1 \reg_mie[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_0530_),
    .Q(reg_mie[3]),
    .QN(_4517_)
  );
  DFF_X1 \reg_mie[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_0531_),
    .Q(reg_mie[7]),
    .QN(_4516_)
  );
  DFF_X1 \reg_misa[0]$_SDFFE_PP1P_  (
    .CK(clock),
    .D(_0426_),
    .Q(reg_misa[0]),
    .QN(_4619_)
  );
  DFF_X1 \reg_misa[12]$_SDFFE_PP1P_  (
    .CK(clock),
    .D(_0428_),
    .Q(reg_misa[12]),
    .QN(_4618_)
  );
  DFF_X1 \reg_misa[2]$_SDFFE_PP1P_  (
    .CK(clock),
    .D(_0427_),
    .Q(reg_misa[2]),
    .QN(_GEN_586[1])
  );
  DFF_X1 \reg_mscratch[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_0332_),
    .Q(reg_mscratch[0]),
    .QN(_4713_)
  );
  DFF_X1 \reg_mscratch[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_0342_),
    .Q(reg_mscratch[10]),
    .QN(_4703_)
  );
  DFF_X1 \reg_mscratch[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_0343_),
    .Q(reg_mscratch[11]),
    .QN(_4702_)
  );
  DFF_X1 \reg_mscratch[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_0344_),
    .Q(reg_mscratch[12]),
    .QN(_4701_)
  );
  DFF_X1 \reg_mscratch[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_0345_),
    .Q(reg_mscratch[13]),
    .QN(_4700_)
  );
  DFF_X1 \reg_mscratch[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_0346_),
    .Q(reg_mscratch[14]),
    .QN(_4699_)
  );
  DFF_X1 \reg_mscratch[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_0347_),
    .Q(reg_mscratch[15]),
    .QN(_4698_)
  );
  DFF_X1 \reg_mscratch[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_0348_),
    .Q(reg_mscratch[16]),
    .QN(_4697_)
  );
  DFF_X1 \reg_mscratch[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_0349_),
    .Q(reg_mscratch[17]),
    .QN(_4696_)
  );
  DFF_X1 \reg_mscratch[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_0350_),
    .Q(reg_mscratch[18]),
    .QN(_4695_)
  );
  DFF_X1 \reg_mscratch[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_0351_),
    .Q(reg_mscratch[19]),
    .QN(_4694_)
  );
  DFF_X1 \reg_mscratch[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_0333_),
    .Q(reg_mscratch[1]),
    .QN(_4712_)
  );
  DFF_X1 \reg_mscratch[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_0352_),
    .Q(reg_mscratch[20]),
    .QN(_4693_)
  );
  DFF_X1 \reg_mscratch[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_0353_),
    .Q(reg_mscratch[21]),
    .QN(_4692_)
  );
  DFF_X1 \reg_mscratch[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_0354_),
    .Q(reg_mscratch[22]),
    .QN(_4691_)
  );
  DFF_X1 \reg_mscratch[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_0355_),
    .Q(reg_mscratch[23]),
    .QN(_4690_)
  );
  DFF_X1 \reg_mscratch[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_0356_),
    .Q(reg_mscratch[24]),
    .QN(_4689_)
  );
  DFF_X1 \reg_mscratch[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_0357_),
    .Q(reg_mscratch[25]),
    .QN(_4688_)
  );
  DFF_X1 \reg_mscratch[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_0358_),
    .Q(reg_mscratch[26]),
    .QN(_4687_)
  );
  DFF_X1 \reg_mscratch[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_0359_),
    .Q(reg_mscratch[27]),
    .QN(_4686_)
  );
  DFF_X1 \reg_mscratch[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_0360_),
    .Q(reg_mscratch[28]),
    .QN(_4685_)
  );
  DFF_X1 \reg_mscratch[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_0361_),
    .Q(reg_mscratch[29]),
    .QN(_4684_)
  );
  DFF_X1 \reg_mscratch[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_0334_),
    .Q(reg_mscratch[2]),
    .QN(_4711_)
  );
  DFF_X1 \reg_mscratch[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_0362_),
    .Q(reg_mscratch[30]),
    .QN(_4683_)
  );
  DFF_X1 \reg_mscratch[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_0363_),
    .Q(reg_mscratch[31]),
    .QN(_4682_)
  );
  DFF_X1 \reg_mscratch[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_0335_),
    .Q(reg_mscratch[3]),
    .QN(_4710_)
  );
  DFF_X1 \reg_mscratch[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_0336_),
    .Q(reg_mscratch[4]),
    .QN(_4709_)
  );
  DFF_X1 \reg_mscratch[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_0337_),
    .Q(reg_mscratch[5]),
    .QN(_4708_)
  );
  DFF_X1 \reg_mscratch[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_0338_),
    .Q(reg_mscratch[6]),
    .QN(_4707_)
  );
  DFF_X1 \reg_mscratch[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_0339_),
    .Q(reg_mscratch[7]),
    .QN(_4706_)
  );
  DFF_X1 \reg_mscratch[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_0340_),
    .Q(reg_mscratch[8]),
    .QN(_4705_)
  );
  DFF_X1 \reg_mscratch[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_0341_),
    .Q(reg_mscratch[9]),
    .QN(_4704_)
  );
  DFF_X1 \reg_mstatus_gva$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0293_),
    .Q(reg_mstatus_gva),
    .QN(_4752_)
  );
  DFF_X1 \reg_mstatus_mie$_SDFF_PP0_  (
    .CK(clock),
    .D(_0283_),
    .Q(reg_mstatus_mie),
    .QN(_4760_)
  );
  DFF_X1 \reg_mstatus_mpie$_SDFF_PP0_  (
    .CK(clock),
    .D(_0289_),
    .Q(reg_mstatus_mpie),
    .QN(_4754_)
  );
  DFF_X1 \reg_mtval[0]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[0]),
    .Q(reg_mtval[0]),
    .QN(_5041_)
  );
  DFF_X1 \reg_mtval[10]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[10]),
    .Q(reg_mtval[10]),
    .QN(_5051_)
  );
  DFF_X1 \reg_mtval[11]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[11]),
    .Q(reg_mtval[11]),
    .QN(_5052_)
  );
  DFF_X1 \reg_mtval[12]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[12]),
    .Q(reg_mtval[12]),
    .QN(_5053_)
  );
  DFF_X1 \reg_mtval[13]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[13]),
    .Q(reg_mtval[13]),
    .QN(_5054_)
  );
  DFF_X1 \reg_mtval[14]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[14]),
    .Q(reg_mtval[14]),
    .QN(_5055_)
  );
  DFF_X1 \reg_mtval[15]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[15]),
    .Q(reg_mtval[15]),
    .QN(_5056_)
  );
  DFF_X1 \reg_mtval[16]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[16]),
    .Q(reg_mtval[16]),
    .QN(_5057_)
  );
  DFF_X1 \reg_mtval[17]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[17]),
    .Q(reg_mtval[17]),
    .QN(_5058_)
  );
  DFF_X1 \reg_mtval[18]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[18]),
    .Q(reg_mtval[18]),
    .QN(_5059_)
  );
  DFF_X1 \reg_mtval[19]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[19]),
    .Q(reg_mtval[19]),
    .QN(_5060_)
  );
  DFF_X1 \reg_mtval[1]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[1]),
    .Q(reg_mtval[1]),
    .QN(_5042_)
  );
  DFF_X1 \reg_mtval[20]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[20]),
    .Q(reg_mtval[20]),
    .QN(_5061_)
  );
  DFF_X1 \reg_mtval[21]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[21]),
    .Q(reg_mtval[21]),
    .QN(_5062_)
  );
  DFF_X1 \reg_mtval[22]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[22]),
    .Q(reg_mtval[22]),
    .QN(_5063_)
  );
  DFF_X1 \reg_mtval[23]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[23]),
    .Q(reg_mtval[23]),
    .QN(_5064_)
  );
  DFF_X1 \reg_mtval[24]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[24]),
    .Q(reg_mtval[24]),
    .QN(_5065_)
  );
  DFF_X1 \reg_mtval[25]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[25]),
    .Q(reg_mtval[25]),
    .QN(_5066_)
  );
  DFF_X1 \reg_mtval[26]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[26]),
    .Q(reg_mtval[26]),
    .QN(_5067_)
  );
  DFF_X1 \reg_mtval[27]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[27]),
    .Q(reg_mtval[27]),
    .QN(_5068_)
  );
  DFF_X1 \reg_mtval[28]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[28]),
    .Q(reg_mtval[28]),
    .QN(_5069_)
  );
  DFF_X1 \reg_mtval[29]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[29]),
    .Q(reg_mtval[29]),
    .QN(_5070_)
  );
  DFF_X1 \reg_mtval[2]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[2]),
    .Q(reg_mtval[2]),
    .QN(_5043_)
  );
  DFF_X1 \reg_mtval[30]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[30]),
    .Q(reg_mtval[30]),
    .QN(_5071_)
  );
  DFF_X1 \reg_mtval[31]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[31]),
    .Q(reg_mtval[31]),
    .QN(_5072_)
  );
  DFF_X1 \reg_mtval[3]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[3]),
    .Q(reg_mtval[3]),
    .QN(_5044_)
  );
  DFF_X1 \reg_mtval[4]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[4]),
    .Q(reg_mtval[4]),
    .QN(_5045_)
  );
  DFF_X1 \reg_mtval[5]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[5]),
    .Q(reg_mtval[5]),
    .QN(_5046_)
  );
  DFF_X1 \reg_mtval[6]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[6]),
    .Q(reg_mtval[6]),
    .QN(_5047_)
  );
  DFF_X1 \reg_mtval[7]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[7]),
    .Q(reg_mtval[7]),
    .QN(_5048_)
  );
  DFF_X1 \reg_mtval[8]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[8]),
    .Q(reg_mtval[8]),
    .QN(_5049_)
  );
  DFF_X1 \reg_mtval[9]$_DFF_P_  (
    .CK(clock),
    .D(_0002_[9]),
    .Q(reg_mtval[9]),
    .QN(_5050_)
  );
  DFF_X1 \reg_mtvec[0]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0467_),
    .Q(reg_mtvec[0]),
    .QN(_read_mtvec_T_4[6])
  );
  DFF_X1 \reg_mtvec[10]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0476_),
    .Q(reg_mtvec[10]),
    .QN(_4571_)
  );
  DFF_X1 \reg_mtvec[11]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0477_),
    .Q(reg_mtvec[11]),
    .QN(_4570_)
  );
  DFF_X1 \reg_mtvec[12]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0478_),
    .Q(reg_mtvec[12]),
    .QN(_4569_)
  );
  DFF_X1 \reg_mtvec[13]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0479_),
    .Q(reg_mtvec[13]),
    .QN(_4568_)
  );
  DFF_X1 \reg_mtvec[14]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0480_),
    .Q(reg_mtvec[14]),
    .QN(_4567_)
  );
  DFF_X1 \reg_mtvec[15]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0481_),
    .Q(reg_mtvec[15]),
    .QN(_4566_)
  );
  DFF_X1 \reg_mtvec[16]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0482_),
    .Q(reg_mtvec[16]),
    .QN(_4565_)
  );
  DFF_X1 \reg_mtvec[17]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0483_),
    .Q(reg_mtvec[17]),
    .QN(_4564_)
  );
  DFF_X1 \reg_mtvec[18]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0484_),
    .Q(reg_mtvec[18]),
    .QN(_4563_)
  );
  DFF_X1 \reg_mtvec[19]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0485_),
    .Q(reg_mtvec[19]),
    .QN(_4562_)
  );
  DFF_X1 \reg_mtvec[20]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0486_),
    .Q(reg_mtvec[20]),
    .QN(_4561_)
  );
  DFF_X1 \reg_mtvec[21]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0487_),
    .Q(reg_mtvec[21]),
    .QN(_4560_)
  );
  DFF_X1 \reg_mtvec[22]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0488_),
    .Q(reg_mtvec[22]),
    .QN(_4559_)
  );
  DFF_X1 \reg_mtvec[23]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0489_),
    .Q(reg_mtvec[23]),
    .QN(_4558_)
  );
  DFF_X1 \reg_mtvec[24]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0490_),
    .Q(reg_mtvec[24]),
    .QN(_4557_)
  );
  DFF_X1 \reg_mtvec[25]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0491_),
    .Q(reg_mtvec[25]),
    .QN(_4556_)
  );
  DFF_X1 \reg_mtvec[26]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0492_),
    .Q(reg_mtvec[26]),
    .QN(_4555_)
  );
  DFF_X1 \reg_mtvec[27]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0493_),
    .Q(reg_mtvec[27]),
    .QN(_4554_)
  );
  DFF_X1 \reg_mtvec[28]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0494_),
    .Q(reg_mtvec[28]),
    .QN(_4553_)
  );
  DFF_X1 \reg_mtvec[29]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0495_),
    .Q(reg_mtvec[29]),
    .QN(_4552_)
  );
  DFF_X1 \reg_mtvec[2]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0468_),
    .Q(reg_mtvec[2]),
    .QN(_4579_)
  );
  DFF_X1 \reg_mtvec[30]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0496_),
    .Q(reg_mtvec[30]),
    .QN(_4551_)
  );
  DFF_X1 \reg_mtvec[31]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0497_),
    .Q(reg_mtvec[31]),
    .QN(_4550_)
  );
  DFF_X1 \reg_mtvec[3]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0469_),
    .Q(reg_mtvec[3]),
    .QN(_4578_)
  );
  DFF_X1 \reg_mtvec[4]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0470_),
    .Q(reg_mtvec[4]),
    .QN(_4577_)
  );
  DFF_X1 \reg_mtvec[5]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0471_),
    .Q(reg_mtvec[5]),
    .QN(_4576_)
  );
  DFF_X1 \reg_mtvec[6]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0472_),
    .Q(reg_mtvec[6]),
    .QN(_4575_)
  );
  DFF_X1 \reg_mtvec[7]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0473_),
    .Q(reg_mtvec[7]),
    .QN(_4574_)
  );
  DFF_X1 \reg_mtvec[8]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0474_),
    .Q(reg_mtvec[8]),
    .QN(_4573_)
  );
  DFF_X1 \reg_mtvec[9]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0475_),
    .Q(reg_mtvec[9]),
    .QN(_4572_)
  );
  DFF_X1 \reg_pmp_0_addr[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_0176_),
    .Q(reg_pmp_0_addr[0]),
    .QN(_4865_)
  );
  DFF_X1 \reg_pmp_0_addr[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_0186_),
    .Q(reg_pmp_0_addr[10]),
    .QN(_4855_)
  );
  DFF_X1 \reg_pmp_0_addr[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_0187_),
    .Q(reg_pmp_0_addr[11]),
    .QN(_4854_)
  );
  DFF_X1 \reg_pmp_0_addr[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_0188_),
    .Q(reg_pmp_0_addr[12]),
    .QN(_4853_)
  );
  DFF_X1 \reg_pmp_0_addr[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_0189_),
    .Q(reg_pmp_0_addr[13]),
    .QN(_4852_)
  );
  DFF_X1 \reg_pmp_0_addr[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_0190_),
    .Q(reg_pmp_0_addr[14]),
    .QN(_4851_)
  );
  DFF_X1 \reg_pmp_0_addr[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_0191_),
    .Q(reg_pmp_0_addr[15]),
    .QN(_4850_)
  );
  DFF_X1 \reg_pmp_0_addr[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_0192_),
    .Q(reg_pmp_0_addr[16]),
    .QN(_4849_)
  );
  DFF_X1 \reg_pmp_0_addr[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_0193_),
    .Q(reg_pmp_0_addr[17]),
    .QN(_4848_)
  );
  DFF_X1 \reg_pmp_0_addr[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_0194_),
    .Q(reg_pmp_0_addr[18]),
    .QN(_4847_)
  );
  DFF_X1 \reg_pmp_0_addr[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_0195_),
    .Q(reg_pmp_0_addr[19]),
    .QN(_4846_)
  );
  DFF_X1 \reg_pmp_0_addr[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_0177_),
    .Q(reg_pmp_0_addr[1]),
    .QN(_4864_)
  );
  DFF_X1 \reg_pmp_0_addr[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_0196_),
    .Q(reg_pmp_0_addr[20]),
    .QN(_4845_)
  );
  DFF_X1 \reg_pmp_0_addr[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_0197_),
    .Q(reg_pmp_0_addr[21]),
    .QN(_4844_)
  );
  DFF_X1 \reg_pmp_0_addr[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_0198_),
    .Q(reg_pmp_0_addr[22]),
    .QN(_4843_)
  );
  DFF_X1 \reg_pmp_0_addr[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_0199_),
    .Q(reg_pmp_0_addr[23]),
    .QN(_4842_)
  );
  DFF_X1 \reg_pmp_0_addr[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_0200_),
    .Q(reg_pmp_0_addr[24]),
    .QN(_4841_)
  );
  DFF_X1 \reg_pmp_0_addr[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_0201_),
    .Q(reg_pmp_0_addr[25]),
    .QN(_4840_)
  );
  DFF_X1 \reg_pmp_0_addr[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_0202_),
    .Q(reg_pmp_0_addr[26]),
    .QN(_4839_)
  );
  DFF_X1 \reg_pmp_0_addr[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_0203_),
    .Q(reg_pmp_0_addr[27]),
    .QN(_4838_)
  );
  DFF_X1 \reg_pmp_0_addr[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_0204_),
    .Q(reg_pmp_0_addr[28]),
    .QN(_4837_)
  );
  DFF_X1 \reg_pmp_0_addr[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_0205_),
    .Q(reg_pmp_0_addr[29]),
    .QN(_4836_)
  );
  DFF_X1 \reg_pmp_0_addr[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_0178_),
    .Q(reg_pmp_0_addr[2]),
    .QN(_4863_)
  );
  DFF_X1 \reg_pmp_0_addr[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_0179_),
    .Q(reg_pmp_0_addr[3]),
    .QN(_4862_)
  );
  DFF_X1 \reg_pmp_0_addr[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_0180_),
    .Q(reg_pmp_0_addr[4]),
    .QN(_4861_)
  );
  DFF_X1 \reg_pmp_0_addr[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_0181_),
    .Q(reg_pmp_0_addr[5]),
    .QN(_4860_)
  );
  DFF_X1 \reg_pmp_0_addr[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_0182_),
    .Q(reg_pmp_0_addr[6]),
    .QN(_4859_)
  );
  DFF_X1 \reg_pmp_0_addr[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_0183_),
    .Q(reg_pmp_0_addr[7]),
    .QN(_4858_)
  );
  DFF_X1 \reg_pmp_0_addr[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_0184_),
    .Q(reg_pmp_0_addr[8]),
    .QN(_4857_)
  );
  DFF_X1 \reg_pmp_0_addr[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_0185_),
    .Q(reg_pmp_0_addr[9]),
    .QN(_4856_)
  );
  DFF_X1 \reg_pmp_0_cfg_a[0]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0239_),
    .Q(reg_pmp_0_cfg_a[0]),
    .QN(_4802_)
  );
  DFF_X1 \reg_pmp_0_cfg_a[1]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0240_),
    .Q(reg_pmp_0_cfg_a[1]),
    .QN(_4801_)
  );
  DFF_X1 \reg_pmp_0_cfg_l$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0241_),
    .Q(reg_pmp_0_cfg_l),
    .QN(_0006_)
  );
  DFF_X1 \reg_pmp_0_cfg_r$_DFFE_PP_  (
    .CK(clock),
    .D(_0175_),
    .Q(reg_pmp_0_cfg_r),
    .QN(_4866_)
  );
  DFF_X1 \reg_pmp_0_cfg_w$_DFFE_PP_  (
    .CK(clock),
    .D(_0057_),
    .Q(reg_pmp_0_cfg_w),
    .QN(_4974_)
  );
  DFF_X1 \reg_pmp_0_cfg_x$_DFFE_PP_  (
    .CK(clock),
    .D(_0206_),
    .Q(reg_pmp_0_cfg_x),
    .QN(_4835_)
  );
  DFF_X1 \reg_pmp_1_addr[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_0365_),
    .Q(reg_pmp_1_addr[0]),
    .QN(_4680_)
  );
  DFF_X1 \reg_pmp_1_addr[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_0375_),
    .Q(reg_pmp_1_addr[10]),
    .QN(_4670_)
  );
  DFF_X1 \reg_pmp_1_addr[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_0376_),
    .Q(reg_pmp_1_addr[11]),
    .QN(_4669_)
  );
  DFF_X1 \reg_pmp_1_addr[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_0377_),
    .Q(reg_pmp_1_addr[12]),
    .QN(_4668_)
  );
  DFF_X1 \reg_pmp_1_addr[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_0378_),
    .Q(reg_pmp_1_addr[13]),
    .QN(_4667_)
  );
  DFF_X1 \reg_pmp_1_addr[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_0379_),
    .Q(reg_pmp_1_addr[14]),
    .QN(_4666_)
  );
  DFF_X1 \reg_pmp_1_addr[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_0380_),
    .Q(reg_pmp_1_addr[15]),
    .QN(_4665_)
  );
  DFF_X1 \reg_pmp_1_addr[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_0381_),
    .Q(reg_pmp_1_addr[16]),
    .QN(_4664_)
  );
  DFF_X1 \reg_pmp_1_addr[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_0382_),
    .Q(reg_pmp_1_addr[17]),
    .QN(_4663_)
  );
  DFF_X1 \reg_pmp_1_addr[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_0383_),
    .Q(reg_pmp_1_addr[18]),
    .QN(_4662_)
  );
  DFF_X1 \reg_pmp_1_addr[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_0384_),
    .Q(reg_pmp_1_addr[19]),
    .QN(_4661_)
  );
  DFF_X1 \reg_pmp_1_addr[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_0366_),
    .Q(reg_pmp_1_addr[1]),
    .QN(_4679_)
  );
  DFF_X1 \reg_pmp_1_addr[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_0385_),
    .Q(reg_pmp_1_addr[20]),
    .QN(_4660_)
  );
  DFF_X1 \reg_pmp_1_addr[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_0386_),
    .Q(reg_pmp_1_addr[21]),
    .QN(_4659_)
  );
  DFF_X1 \reg_pmp_1_addr[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_0387_),
    .Q(reg_pmp_1_addr[22]),
    .QN(_4658_)
  );
  DFF_X1 \reg_pmp_1_addr[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_0388_),
    .Q(reg_pmp_1_addr[23]),
    .QN(_4657_)
  );
  DFF_X1 \reg_pmp_1_addr[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_0389_),
    .Q(reg_pmp_1_addr[24]),
    .QN(_4656_)
  );
  DFF_X1 \reg_pmp_1_addr[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_0390_),
    .Q(reg_pmp_1_addr[25]),
    .QN(_4655_)
  );
  DFF_X1 \reg_pmp_1_addr[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_0391_),
    .Q(reg_pmp_1_addr[26]),
    .QN(_4654_)
  );
  DFF_X1 \reg_pmp_1_addr[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_0392_),
    .Q(reg_pmp_1_addr[27]),
    .QN(_4653_)
  );
  DFF_X1 \reg_pmp_1_addr[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_0393_),
    .Q(reg_pmp_1_addr[28]),
    .QN(_4652_)
  );
  DFF_X1 \reg_pmp_1_addr[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_0394_),
    .Q(reg_pmp_1_addr[29]),
    .QN(_4651_)
  );
  DFF_X1 \reg_pmp_1_addr[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_0367_),
    .Q(reg_pmp_1_addr[2]),
    .QN(_4678_)
  );
  DFF_X1 \reg_pmp_1_addr[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_0368_),
    .Q(reg_pmp_1_addr[3]),
    .QN(_4677_)
  );
  DFF_X1 \reg_pmp_1_addr[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_0369_),
    .Q(reg_pmp_1_addr[4]),
    .QN(_4676_)
  );
  DFF_X1 \reg_pmp_1_addr[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_0370_),
    .Q(reg_pmp_1_addr[5]),
    .QN(_4675_)
  );
  DFF_X1 \reg_pmp_1_addr[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_0371_),
    .Q(reg_pmp_1_addr[6]),
    .QN(_4674_)
  );
  DFF_X1 \reg_pmp_1_addr[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_0372_),
    .Q(reg_pmp_1_addr[7]),
    .QN(_4673_)
  );
  DFF_X1 \reg_pmp_1_addr[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_0373_),
    .Q(reg_pmp_1_addr[8]),
    .QN(_4672_)
  );
  DFF_X1 \reg_pmp_1_addr[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_0374_),
    .Q(reg_pmp_1_addr[9]),
    .QN(_4671_)
  );
  DFF_X1 \reg_pmp_1_cfg_a[0]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0172_),
    .Q(reg_pmp_1_cfg_a[0]),
    .QN(_4867_)
  );
  DFF_X1 \reg_pmp_1_cfg_a[1]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0173_),
    .Q(reg_pmp_1_cfg_a[1]),
    .QN(_0008_)
  );
  DFF_X1 \reg_pmp_1_cfg_l$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0174_),
    .Q(reg_pmp_1_cfg_l),
    .QN(_0007_)
  );
  DFF_X1 \reg_pmp_1_cfg_r$_DFFE_PP_  (
    .CK(clock),
    .D(_0168_),
    .Q(reg_pmp_1_cfg_r),
    .QN(_4871_)
  );
  DFF_X1 \reg_pmp_1_cfg_w$_DFFE_PP_  (
    .CK(clock),
    .D(_0133_),
    .Q(reg_pmp_1_cfg_w),
    .QN(_4904_)
  );
  DFF_X1 \reg_pmp_1_cfg_x$_DFFE_PP_  (
    .CK(clock),
    .D(_0170_),
    .Q(reg_pmp_1_cfg_x),
    .QN(_4869_)
  );
  DFF_X1 \reg_pmp_2_addr[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_0103_),
    .Q(reg_pmp_2_addr[0]),
    .QN(_4934_)
  );
  DFF_X1 \reg_pmp_2_addr[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_0113_),
    .Q(reg_pmp_2_addr[10]),
    .QN(_4924_)
  );
  DFF_X1 \reg_pmp_2_addr[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_0114_),
    .Q(reg_pmp_2_addr[11]),
    .QN(_4923_)
  );
  DFF_X1 \reg_pmp_2_addr[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_0115_),
    .Q(reg_pmp_2_addr[12]),
    .QN(_4922_)
  );
  DFF_X1 \reg_pmp_2_addr[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_0116_),
    .Q(reg_pmp_2_addr[13]),
    .QN(_4921_)
  );
  DFF_X1 \reg_pmp_2_addr[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_0117_),
    .Q(reg_pmp_2_addr[14]),
    .QN(_4920_)
  );
  DFF_X1 \reg_pmp_2_addr[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_0118_),
    .Q(reg_pmp_2_addr[15]),
    .QN(_4919_)
  );
  DFF_X1 \reg_pmp_2_addr[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_0119_),
    .Q(reg_pmp_2_addr[16]),
    .QN(_4918_)
  );
  DFF_X1 \reg_pmp_2_addr[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_0120_),
    .Q(reg_pmp_2_addr[17]),
    .QN(_4917_)
  );
  DFF_X1 \reg_pmp_2_addr[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_0121_),
    .Q(reg_pmp_2_addr[18]),
    .QN(_4916_)
  );
  DFF_X1 \reg_pmp_2_addr[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_0122_),
    .Q(reg_pmp_2_addr[19]),
    .QN(_4915_)
  );
  DFF_X1 \reg_pmp_2_addr[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_0104_),
    .Q(reg_pmp_2_addr[1]),
    .QN(_4933_)
  );
  DFF_X1 \reg_pmp_2_addr[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_0123_),
    .Q(reg_pmp_2_addr[20]),
    .QN(_4914_)
  );
  DFF_X1 \reg_pmp_2_addr[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_0124_),
    .Q(reg_pmp_2_addr[21]),
    .QN(_4913_)
  );
  DFF_X1 \reg_pmp_2_addr[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_0125_),
    .Q(reg_pmp_2_addr[22]),
    .QN(_4912_)
  );
  DFF_X1 \reg_pmp_2_addr[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_0126_),
    .Q(reg_pmp_2_addr[23]),
    .QN(_4911_)
  );
  DFF_X1 \reg_pmp_2_addr[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_0127_),
    .Q(reg_pmp_2_addr[24]),
    .QN(_4910_)
  );
  DFF_X1 \reg_pmp_2_addr[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_0128_),
    .Q(reg_pmp_2_addr[25]),
    .QN(_4909_)
  );
  DFF_X1 \reg_pmp_2_addr[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_0129_),
    .Q(reg_pmp_2_addr[26]),
    .QN(_4908_)
  );
  DFF_X1 \reg_pmp_2_addr[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_0130_),
    .Q(reg_pmp_2_addr[27]),
    .QN(_4907_)
  );
  DFF_X1 \reg_pmp_2_addr[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_0131_),
    .Q(reg_pmp_2_addr[28]),
    .QN(_4906_)
  );
  DFF_X1 \reg_pmp_2_addr[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_0132_),
    .Q(reg_pmp_2_addr[29]),
    .QN(_4905_)
  );
  DFF_X1 \reg_pmp_2_addr[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_0105_),
    .Q(reg_pmp_2_addr[2]),
    .QN(_4932_)
  );
  DFF_X1 \reg_pmp_2_addr[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_0106_),
    .Q(reg_pmp_2_addr[3]),
    .QN(_4931_)
  );
  DFF_X1 \reg_pmp_2_addr[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_0107_),
    .Q(reg_pmp_2_addr[4]),
    .QN(_4930_)
  );
  DFF_X1 \reg_pmp_2_addr[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_0108_),
    .Q(reg_pmp_2_addr[5]),
    .QN(_4929_)
  );
  DFF_X1 \reg_pmp_2_addr[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_0109_),
    .Q(reg_pmp_2_addr[6]),
    .QN(_4928_)
  );
  DFF_X1 \reg_pmp_2_addr[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_0110_),
    .Q(reg_pmp_2_addr[7]),
    .QN(_4927_)
  );
  DFF_X1 \reg_pmp_2_addr[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_0111_),
    .Q(reg_pmp_2_addr[8]),
    .QN(_4926_)
  );
  DFF_X1 \reg_pmp_2_addr[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_0112_),
    .Q(reg_pmp_2_addr[9]),
    .QN(_4925_)
  );
  DFF_X1 \reg_pmp_2_cfg_a[0]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0165_),
    .Q(reg_pmp_2_cfg_a[0]),
    .QN(_4872_)
  );
  DFF_X1 \reg_pmp_2_cfg_a[1]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0166_),
    .Q(reg_pmp_2_cfg_a[1]),
    .QN(_0010_)
  );
  DFF_X1 \reg_pmp_2_cfg_l$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0167_),
    .Q(reg_pmp_2_cfg_l),
    .QN(_0009_)
  );
  DFF_X1 \reg_pmp_2_cfg_r$_DFFE_PP_  (
    .CK(clock),
    .D(_0134_),
    .Q(reg_pmp_2_cfg_r),
    .QN(_4903_)
  );
  DFF_X1 \reg_pmp_2_cfg_w$_DFFE_PP_  (
    .CK(clock),
    .D(_0099_),
    .Q(reg_pmp_2_cfg_w),
    .QN(_4936_)
  );
  DFF_X1 \reg_pmp_2_cfg_x$_DFFE_PP_  (
    .CK(clock),
    .D(_0171_),
    .Q(reg_pmp_2_cfg_x),
    .QN(_4868_)
  );
  DFF_X1 \reg_pmp_3_addr[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_0135_),
    .Q(reg_pmp_3_addr[0]),
    .QN(_4902_)
  );
  DFF_X1 \reg_pmp_3_addr[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_0145_),
    .Q(reg_pmp_3_addr[10]),
    .QN(_4892_)
  );
  DFF_X1 \reg_pmp_3_addr[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_0146_),
    .Q(reg_pmp_3_addr[11]),
    .QN(_4891_)
  );
  DFF_X1 \reg_pmp_3_addr[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_0147_),
    .Q(reg_pmp_3_addr[12]),
    .QN(_4890_)
  );
  DFF_X1 \reg_pmp_3_addr[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_0148_),
    .Q(reg_pmp_3_addr[13]),
    .QN(_4889_)
  );
  DFF_X1 \reg_pmp_3_addr[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_0149_),
    .Q(reg_pmp_3_addr[14]),
    .QN(_4888_)
  );
  DFF_X1 \reg_pmp_3_addr[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_0150_),
    .Q(reg_pmp_3_addr[15]),
    .QN(_4887_)
  );
  DFF_X1 \reg_pmp_3_addr[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_0151_),
    .Q(reg_pmp_3_addr[16]),
    .QN(_4886_)
  );
  DFF_X1 \reg_pmp_3_addr[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_0152_),
    .Q(reg_pmp_3_addr[17]),
    .QN(_4885_)
  );
  DFF_X1 \reg_pmp_3_addr[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_0153_),
    .Q(reg_pmp_3_addr[18]),
    .QN(_4884_)
  );
  DFF_X1 \reg_pmp_3_addr[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_0154_),
    .Q(reg_pmp_3_addr[19]),
    .QN(_4883_)
  );
  DFF_X1 \reg_pmp_3_addr[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_0136_),
    .Q(reg_pmp_3_addr[1]),
    .QN(_4901_)
  );
  DFF_X1 \reg_pmp_3_addr[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_0155_),
    .Q(reg_pmp_3_addr[20]),
    .QN(_4882_)
  );
  DFF_X1 \reg_pmp_3_addr[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_0156_),
    .Q(reg_pmp_3_addr[21]),
    .QN(_4881_)
  );
  DFF_X1 \reg_pmp_3_addr[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_0157_),
    .Q(reg_pmp_3_addr[22]),
    .QN(_4880_)
  );
  DFF_X1 \reg_pmp_3_addr[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_0158_),
    .Q(reg_pmp_3_addr[23]),
    .QN(_4879_)
  );
  DFF_X1 \reg_pmp_3_addr[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_0159_),
    .Q(reg_pmp_3_addr[24]),
    .QN(_4878_)
  );
  DFF_X1 \reg_pmp_3_addr[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_0160_),
    .Q(reg_pmp_3_addr[25]),
    .QN(_4877_)
  );
  DFF_X1 \reg_pmp_3_addr[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_0161_),
    .Q(reg_pmp_3_addr[26]),
    .QN(_4876_)
  );
  DFF_X1 \reg_pmp_3_addr[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_0162_),
    .Q(reg_pmp_3_addr[27]),
    .QN(_4875_)
  );
  DFF_X1 \reg_pmp_3_addr[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_0163_),
    .Q(reg_pmp_3_addr[28]),
    .QN(_4874_)
  );
  DFF_X1 \reg_pmp_3_addr[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_0164_),
    .Q(reg_pmp_3_addr[29]),
    .QN(_4873_)
  );
  DFF_X1 \reg_pmp_3_addr[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_0137_),
    .Q(reg_pmp_3_addr[2]),
    .QN(_4900_)
  );
  DFF_X1 \reg_pmp_3_addr[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_0138_),
    .Q(reg_pmp_3_addr[3]),
    .QN(_4899_)
  );
  DFF_X1 \reg_pmp_3_addr[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_0139_),
    .Q(reg_pmp_3_addr[4]),
    .QN(_4898_)
  );
  DFF_X1 \reg_pmp_3_addr[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_0140_),
    .Q(reg_pmp_3_addr[5]),
    .QN(_4897_)
  );
  DFF_X1 \reg_pmp_3_addr[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_0141_),
    .Q(reg_pmp_3_addr[6]),
    .QN(_4896_)
  );
  DFF_X1 \reg_pmp_3_addr[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_0142_),
    .Q(reg_pmp_3_addr[7]),
    .QN(_4895_)
  );
  DFF_X1 \reg_pmp_3_addr[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_0143_),
    .Q(reg_pmp_3_addr[8]),
    .QN(_4894_)
  );
  DFF_X1 \reg_pmp_3_addr[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_0144_),
    .Q(reg_pmp_3_addr[9]),
    .QN(_4893_)
  );
  DFF_X1 \reg_pmp_3_cfg_a[0]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0100_),
    .Q(reg_pmp_3_cfg_a[0]),
    .QN(_4935_)
  );
  DFF_X1 \reg_pmp_3_cfg_a[1]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0101_),
    .Q(reg_pmp_3_cfg_a[1]),
    .QN(_0012_)
  );
  DFF_X1 \reg_pmp_3_cfg_l$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0102_),
    .Q(reg_pmp_3_cfg_l),
    .QN(_0011_)
  );
  DFF_X1 \reg_pmp_3_cfg_r$_DFFE_PP_  (
    .CK(clock),
    .D(_0098_),
    .Q(reg_pmp_3_cfg_r),
    .QN(_4937_)
  );
  DFF_X1 \reg_pmp_3_cfg_w$_DFFE_PP_  (
    .CK(clock),
    .D(_0096_),
    .Q(reg_pmp_3_cfg_w),
    .QN(_4939_)
  );
  DFF_X1 \reg_pmp_3_cfg_x$_DFFE_PP_  (
    .CK(clock),
    .D(_0097_),
    .Q(reg_pmp_3_cfg_x),
    .QN(_4938_)
  );
  DFF_X1 \reg_pmp_4_addr[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_0061_),
    .Q(reg_pmp_4_addr[0]),
    .QN(_4972_)
  );
  DFF_X1 \reg_pmp_4_addr[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_0071_),
    .Q(reg_pmp_4_addr[10]),
    .QN(_4962_)
  );
  DFF_X1 \reg_pmp_4_addr[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_0072_),
    .Q(reg_pmp_4_addr[11]),
    .QN(_4961_)
  );
  DFF_X1 \reg_pmp_4_addr[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_0073_),
    .Q(reg_pmp_4_addr[12]),
    .QN(_4960_)
  );
  DFF_X1 \reg_pmp_4_addr[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_0074_),
    .Q(reg_pmp_4_addr[13]),
    .QN(_4959_)
  );
  DFF_X1 \reg_pmp_4_addr[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_0075_),
    .Q(reg_pmp_4_addr[14]),
    .QN(_4958_)
  );
  DFF_X1 \reg_pmp_4_addr[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_0076_),
    .Q(reg_pmp_4_addr[15]),
    .QN(_4957_)
  );
  DFF_X1 \reg_pmp_4_addr[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_0077_),
    .Q(reg_pmp_4_addr[16]),
    .QN(_4956_)
  );
  DFF_X1 \reg_pmp_4_addr[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_0078_),
    .Q(reg_pmp_4_addr[17]),
    .QN(_4955_)
  );
  DFF_X1 \reg_pmp_4_addr[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_0079_),
    .Q(reg_pmp_4_addr[18]),
    .QN(_4954_)
  );
  DFF_X1 \reg_pmp_4_addr[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_0080_),
    .Q(reg_pmp_4_addr[19]),
    .QN(_4953_)
  );
  DFF_X1 \reg_pmp_4_addr[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_0062_),
    .Q(reg_pmp_4_addr[1]),
    .QN(_4971_)
  );
  DFF_X1 \reg_pmp_4_addr[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_0081_),
    .Q(reg_pmp_4_addr[20]),
    .QN(_4952_)
  );
  DFF_X1 \reg_pmp_4_addr[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_0082_),
    .Q(reg_pmp_4_addr[21]),
    .QN(_4951_)
  );
  DFF_X1 \reg_pmp_4_addr[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_0083_),
    .Q(reg_pmp_4_addr[22]),
    .QN(_4950_)
  );
  DFF_X1 \reg_pmp_4_addr[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_0084_),
    .Q(reg_pmp_4_addr[23]),
    .QN(_4949_)
  );
  DFF_X1 \reg_pmp_4_addr[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_0085_),
    .Q(reg_pmp_4_addr[24]),
    .QN(_4948_)
  );
  DFF_X1 \reg_pmp_4_addr[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_0086_),
    .Q(reg_pmp_4_addr[25]),
    .QN(_4947_)
  );
  DFF_X1 \reg_pmp_4_addr[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_0087_),
    .Q(reg_pmp_4_addr[26]),
    .QN(_4946_)
  );
  DFF_X1 \reg_pmp_4_addr[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_0088_),
    .Q(reg_pmp_4_addr[27]),
    .QN(_4945_)
  );
  DFF_X1 \reg_pmp_4_addr[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_0089_),
    .Q(reg_pmp_4_addr[28]),
    .QN(_4944_)
  );
  DFF_X1 \reg_pmp_4_addr[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_0090_),
    .Q(reg_pmp_4_addr[29]),
    .QN(_4943_)
  );
  DFF_X1 \reg_pmp_4_addr[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_0063_),
    .Q(reg_pmp_4_addr[2]),
    .QN(_4970_)
  );
  DFF_X1 \reg_pmp_4_addr[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_0064_),
    .Q(reg_pmp_4_addr[3]),
    .QN(_4969_)
  );
  DFF_X1 \reg_pmp_4_addr[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_0065_),
    .Q(reg_pmp_4_addr[4]),
    .QN(_4968_)
  );
  DFF_X1 \reg_pmp_4_addr[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_0066_),
    .Q(reg_pmp_4_addr[5]),
    .QN(_4967_)
  );
  DFF_X1 \reg_pmp_4_addr[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_0067_),
    .Q(reg_pmp_4_addr[6]),
    .QN(_4966_)
  );
  DFF_X1 \reg_pmp_4_addr[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_0068_),
    .Q(reg_pmp_4_addr[7]),
    .QN(_4965_)
  );
  DFF_X1 \reg_pmp_4_addr[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_0069_),
    .Q(reg_pmp_4_addr[8]),
    .QN(_4964_)
  );
  DFF_X1 \reg_pmp_4_addr[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_0070_),
    .Q(reg_pmp_4_addr[9]),
    .QN(_4963_)
  );
  DFF_X1 \reg_pmp_4_cfg_a[0]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0093_),
    .Q(reg_pmp_4_cfg_a[0]),
    .QN(_4940_)
  );
  DFF_X1 \reg_pmp_4_cfg_a[1]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0094_),
    .Q(reg_pmp_4_cfg_a[1]),
    .QN(_0014_)
  );
  DFF_X1 \reg_pmp_4_cfg_l$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0095_),
    .Q(reg_pmp_4_cfg_l),
    .QN(_0013_)
  );
  DFF_X1 \reg_pmp_4_cfg_r$_DFFE_PP_  (
    .CK(clock),
    .D(_0169_),
    .Q(reg_pmp_4_cfg_r),
    .QN(_4870_)
  );
  DFF_X1 \reg_pmp_4_cfg_w$_DFFE_PP_  (
    .CK(clock),
    .D(_0091_),
    .Q(reg_pmp_4_cfg_w),
    .QN(_4942_)
  );
  DFF_X1 \reg_pmp_4_cfg_x$_DFFE_PP_  (
    .CK(clock),
    .D(_0092_),
    .Q(reg_pmp_4_cfg_x),
    .QN(_4941_)
  );
  DFF_X1 \reg_pmp_5_addr[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_0027_),
    .Q(reg_pmp_5_addr[0]),
    .QN(_5004_)
  );
  DFF_X1 \reg_pmp_5_addr[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_0037_),
    .Q(reg_pmp_5_addr[10]),
    .QN(_4994_)
  );
  DFF_X1 \reg_pmp_5_addr[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_0038_),
    .Q(reg_pmp_5_addr[11]),
    .QN(_4993_)
  );
  DFF_X1 \reg_pmp_5_addr[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_0039_),
    .Q(reg_pmp_5_addr[12]),
    .QN(_4992_)
  );
  DFF_X1 \reg_pmp_5_addr[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_0040_),
    .Q(reg_pmp_5_addr[13]),
    .QN(_4991_)
  );
  DFF_X1 \reg_pmp_5_addr[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_0041_),
    .Q(reg_pmp_5_addr[14]),
    .QN(_4990_)
  );
  DFF_X1 \reg_pmp_5_addr[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_0042_),
    .Q(reg_pmp_5_addr[15]),
    .QN(_4989_)
  );
  DFF_X1 \reg_pmp_5_addr[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_0043_),
    .Q(reg_pmp_5_addr[16]),
    .QN(_4988_)
  );
  DFF_X1 \reg_pmp_5_addr[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_0044_),
    .Q(reg_pmp_5_addr[17]),
    .QN(_4987_)
  );
  DFF_X1 \reg_pmp_5_addr[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_0045_),
    .Q(reg_pmp_5_addr[18]),
    .QN(_4986_)
  );
  DFF_X1 \reg_pmp_5_addr[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_0046_),
    .Q(reg_pmp_5_addr[19]),
    .QN(_4985_)
  );
  DFF_X1 \reg_pmp_5_addr[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_0028_),
    .Q(reg_pmp_5_addr[1]),
    .QN(_5003_)
  );
  DFF_X1 \reg_pmp_5_addr[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_0047_),
    .Q(reg_pmp_5_addr[20]),
    .QN(_4984_)
  );
  DFF_X1 \reg_pmp_5_addr[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_0048_),
    .Q(reg_pmp_5_addr[21]),
    .QN(_4983_)
  );
  DFF_X1 \reg_pmp_5_addr[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_0049_),
    .Q(reg_pmp_5_addr[22]),
    .QN(_4982_)
  );
  DFF_X1 \reg_pmp_5_addr[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_0050_),
    .Q(reg_pmp_5_addr[23]),
    .QN(_4981_)
  );
  DFF_X1 \reg_pmp_5_addr[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_0051_),
    .Q(reg_pmp_5_addr[24]),
    .QN(_4980_)
  );
  DFF_X1 \reg_pmp_5_addr[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_0052_),
    .Q(reg_pmp_5_addr[25]),
    .QN(_4979_)
  );
  DFF_X1 \reg_pmp_5_addr[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_0053_),
    .Q(reg_pmp_5_addr[26]),
    .QN(_4978_)
  );
  DFF_X1 \reg_pmp_5_addr[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_0054_),
    .Q(reg_pmp_5_addr[27]),
    .QN(_4977_)
  );
  DFF_X1 \reg_pmp_5_addr[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_0055_),
    .Q(reg_pmp_5_addr[28]),
    .QN(_4976_)
  );
  DFF_X1 \reg_pmp_5_addr[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_0056_),
    .Q(reg_pmp_5_addr[29]),
    .QN(_4975_)
  );
  DFF_X1 \reg_pmp_5_addr[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_0029_),
    .Q(reg_pmp_5_addr[2]),
    .QN(_5002_)
  );
  DFF_X1 \reg_pmp_5_addr[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_0030_),
    .Q(reg_pmp_5_addr[3]),
    .QN(_5001_)
  );
  DFF_X1 \reg_pmp_5_addr[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_0031_),
    .Q(reg_pmp_5_addr[4]),
    .QN(_5000_)
  );
  DFF_X1 \reg_pmp_5_addr[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_0032_),
    .Q(reg_pmp_5_addr[5]),
    .QN(_4999_)
  );
  DFF_X1 \reg_pmp_5_addr[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_0033_),
    .Q(reg_pmp_5_addr[6]),
    .QN(_4998_)
  );
  DFF_X1 \reg_pmp_5_addr[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_0034_),
    .Q(reg_pmp_5_addr[7]),
    .QN(_4997_)
  );
  DFF_X1 \reg_pmp_5_addr[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_0035_),
    .Q(reg_pmp_5_addr[8]),
    .QN(_4996_)
  );
  DFF_X1 \reg_pmp_5_addr[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_0036_),
    .Q(reg_pmp_5_addr[9]),
    .QN(_4995_)
  );
  DFF_X1 \reg_pmp_5_cfg_a[0]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0058_),
    .Q(reg_pmp_5_cfg_a[0]),
    .QN(_4973_)
  );
  DFF_X1 \reg_pmp_5_cfg_a[1]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0059_),
    .Q(reg_pmp_5_cfg_a[1]),
    .QN(_0016_)
  );
  DFF_X1 \reg_pmp_5_cfg_l$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0060_),
    .Q(reg_pmp_5_cfg_l),
    .QN(_0015_)
  );
  DFF_X1 \reg_pmp_5_cfg_r$_DFFE_PP_  (
    .CK(clock),
    .D(_0025_),
    .Q(reg_pmp_5_cfg_r),
    .QN(_5006_)
  );
  DFF_X1 \reg_pmp_5_cfg_w$_DFFE_PP_  (
    .CK(clock),
    .D(_0026_),
    .Q(reg_pmp_5_cfg_w),
    .QN(_5005_)
  );
  DFF_X1 \reg_pmp_5_cfg_x$_DFFE_PP_  (
    .CK(clock),
    .D(_0364_),
    .Q(reg_pmp_5_cfg_x),
    .QN(_4681_)
  );
  DFF_X1 \reg_pmp_6_addr[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_0395_),
    .Q(reg_pmp_6_addr[0]),
    .QN(_4650_)
  );
  DFF_X1 \reg_pmp_6_addr[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_0405_),
    .Q(reg_pmp_6_addr[10]),
    .QN(_4640_)
  );
  DFF_X1 \reg_pmp_6_addr[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_0406_),
    .Q(reg_pmp_6_addr[11]),
    .QN(_4639_)
  );
  DFF_X1 \reg_pmp_6_addr[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_0407_),
    .Q(reg_pmp_6_addr[12]),
    .QN(_4638_)
  );
  DFF_X1 \reg_pmp_6_addr[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_0408_),
    .Q(reg_pmp_6_addr[13]),
    .QN(_4637_)
  );
  DFF_X1 \reg_pmp_6_addr[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_0409_),
    .Q(reg_pmp_6_addr[14]),
    .QN(_4636_)
  );
  DFF_X1 \reg_pmp_6_addr[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_0410_),
    .Q(reg_pmp_6_addr[15]),
    .QN(_4635_)
  );
  DFF_X1 \reg_pmp_6_addr[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_0411_),
    .Q(reg_pmp_6_addr[16]),
    .QN(_4634_)
  );
  DFF_X1 \reg_pmp_6_addr[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_0412_),
    .Q(reg_pmp_6_addr[17]),
    .QN(_4633_)
  );
  DFF_X1 \reg_pmp_6_addr[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_0413_),
    .Q(reg_pmp_6_addr[18]),
    .QN(_4632_)
  );
  DFF_X1 \reg_pmp_6_addr[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_0414_),
    .Q(reg_pmp_6_addr[19]),
    .QN(_4631_)
  );
  DFF_X1 \reg_pmp_6_addr[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_0396_),
    .Q(reg_pmp_6_addr[1]),
    .QN(_4649_)
  );
  DFF_X1 \reg_pmp_6_addr[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_0415_),
    .Q(reg_pmp_6_addr[20]),
    .QN(_4630_)
  );
  DFF_X1 \reg_pmp_6_addr[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_0416_),
    .Q(reg_pmp_6_addr[21]),
    .QN(_4629_)
  );
  DFF_X1 \reg_pmp_6_addr[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_0417_),
    .Q(reg_pmp_6_addr[22]),
    .QN(_4628_)
  );
  DFF_X1 \reg_pmp_6_addr[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_0418_),
    .Q(reg_pmp_6_addr[23]),
    .QN(_4627_)
  );
  DFF_X1 \reg_pmp_6_addr[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_0419_),
    .Q(reg_pmp_6_addr[24]),
    .QN(_4626_)
  );
  DFF_X1 \reg_pmp_6_addr[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_0420_),
    .Q(reg_pmp_6_addr[25]),
    .QN(_4625_)
  );
  DFF_X1 \reg_pmp_6_addr[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_0421_),
    .Q(reg_pmp_6_addr[26]),
    .QN(_4624_)
  );
  DFF_X1 \reg_pmp_6_addr[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_0422_),
    .Q(reg_pmp_6_addr[27]),
    .QN(_4623_)
  );
  DFF_X1 \reg_pmp_6_addr[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_0423_),
    .Q(reg_pmp_6_addr[28]),
    .QN(_4622_)
  );
  DFF_X1 \reg_pmp_6_addr[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_0424_),
    .Q(reg_pmp_6_addr[29]),
    .QN(_4621_)
  );
  DFF_X1 \reg_pmp_6_addr[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_0397_),
    .Q(reg_pmp_6_addr[2]),
    .QN(_4648_)
  );
  DFF_X1 \reg_pmp_6_addr[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_0398_),
    .Q(reg_pmp_6_addr[3]),
    .QN(_4647_)
  );
  DFF_X1 \reg_pmp_6_addr[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_0399_),
    .Q(reg_pmp_6_addr[4]),
    .QN(_4646_)
  );
  DFF_X1 \reg_pmp_6_addr[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_0400_),
    .Q(reg_pmp_6_addr[5]),
    .QN(_4645_)
  );
  DFF_X1 \reg_pmp_6_addr[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_0401_),
    .Q(reg_pmp_6_addr[6]),
    .QN(_4644_)
  );
  DFF_X1 \reg_pmp_6_addr[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_0402_),
    .Q(reg_pmp_6_addr[7]),
    .QN(_4643_)
  );
  DFF_X1 \reg_pmp_6_addr[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_0403_),
    .Q(reg_pmp_6_addr[8]),
    .QN(_4642_)
  );
  DFF_X1 \reg_pmp_6_addr[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_0404_),
    .Q(reg_pmp_6_addr[9]),
    .QN(_4641_)
  );
  DFF_X1 \reg_pmp_6_cfg_a[0]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0022_),
    .Q(reg_pmp_6_cfg_a[0]),
    .QN(_5007_)
  );
  DFF_X1 \reg_pmp_6_cfg_a[1]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0023_),
    .Q(reg_pmp_6_cfg_a[1]),
    .QN(_0018_)
  );
  DFF_X1 \reg_pmp_6_cfg_l$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0024_),
    .Q(reg_pmp_6_cfg_l),
    .QN(_0017_)
  );
  DFF_X1 \reg_pmp_6_cfg_r$_DFFE_PP_  (
    .CK(clock),
    .D(_0019_),
    .Q(reg_pmp_6_cfg_r),
    .QN(_5010_)
  );
  DFF_X1 \reg_pmp_6_cfg_w$_DFFE_PP_  (
    .CK(clock),
    .D(_0621_),
    .Q(reg_pmp_6_cfg_w),
    .QN(_4430_)
  );
  DFF_X1 \reg_pmp_6_cfg_x$_DFFE_PP_  (
    .CK(clock),
    .D(_0020_),
    .Q(reg_pmp_6_cfg_x),
    .QN(_5009_)
  );
  DFF_X1 \reg_pmp_7_addr[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_0536_),
    .Q(reg_pmp_7_addr[0]),
    .QN(_4511_)
  );
  DFF_X1 \reg_pmp_7_addr[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_0546_),
    .Q(reg_pmp_7_addr[10]),
    .QN(_4501_)
  );
  DFF_X1 \reg_pmp_7_addr[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_0547_),
    .Q(reg_pmp_7_addr[11]),
    .QN(_4500_)
  );
  DFF_X1 \reg_pmp_7_addr[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_0548_),
    .Q(reg_pmp_7_addr[12]),
    .QN(_4499_)
  );
  DFF_X1 \reg_pmp_7_addr[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_0549_),
    .Q(reg_pmp_7_addr[13]),
    .QN(_4498_)
  );
  DFF_X1 \reg_pmp_7_addr[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_0550_),
    .Q(reg_pmp_7_addr[14]),
    .QN(_4497_)
  );
  DFF_X1 \reg_pmp_7_addr[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_0551_),
    .Q(reg_pmp_7_addr[15]),
    .QN(_4496_)
  );
  DFF_X1 \reg_pmp_7_addr[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_0552_),
    .Q(reg_pmp_7_addr[16]),
    .QN(_4495_)
  );
  DFF_X1 \reg_pmp_7_addr[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_0553_),
    .Q(reg_pmp_7_addr[17]),
    .QN(_4494_)
  );
  DFF_X1 \reg_pmp_7_addr[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_0554_),
    .Q(reg_pmp_7_addr[18]),
    .QN(_4493_)
  );
  DFF_X1 \reg_pmp_7_addr[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_0555_),
    .Q(reg_pmp_7_addr[19]),
    .QN(_4492_)
  );
  DFF_X1 \reg_pmp_7_addr[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_0537_),
    .Q(reg_pmp_7_addr[1]),
    .QN(_4510_)
  );
  DFF_X1 \reg_pmp_7_addr[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_0556_),
    .Q(reg_pmp_7_addr[20]),
    .QN(_4491_)
  );
  DFF_X1 \reg_pmp_7_addr[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_0557_),
    .Q(reg_pmp_7_addr[21]),
    .QN(_4490_)
  );
  DFF_X1 \reg_pmp_7_addr[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_0558_),
    .Q(reg_pmp_7_addr[22]),
    .QN(_4489_)
  );
  DFF_X1 \reg_pmp_7_addr[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_0559_),
    .Q(reg_pmp_7_addr[23]),
    .QN(_4488_)
  );
  DFF_X1 \reg_pmp_7_addr[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_0560_),
    .Q(reg_pmp_7_addr[24]),
    .QN(_4487_)
  );
  DFF_X1 \reg_pmp_7_addr[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_0561_),
    .Q(reg_pmp_7_addr[25]),
    .QN(_4486_)
  );
  DFF_X1 \reg_pmp_7_addr[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_0562_),
    .Q(reg_pmp_7_addr[26]),
    .QN(_4485_)
  );
  DFF_X1 \reg_pmp_7_addr[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_0563_),
    .Q(reg_pmp_7_addr[27]),
    .QN(_4484_)
  );
  DFF_X1 \reg_pmp_7_addr[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_0564_),
    .Q(reg_pmp_7_addr[28]),
    .QN(_4483_)
  );
  DFF_X1 \reg_pmp_7_addr[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_0565_),
    .Q(reg_pmp_7_addr[29]),
    .QN(_4482_)
  );
  DFF_X1 \reg_pmp_7_addr[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_0538_),
    .Q(reg_pmp_7_addr[2]),
    .QN(_4509_)
  );
  DFF_X1 \reg_pmp_7_addr[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_0539_),
    .Q(reg_pmp_7_addr[3]),
    .QN(_4508_)
  );
  DFF_X1 \reg_pmp_7_addr[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_0540_),
    .Q(reg_pmp_7_addr[4]),
    .QN(_4507_)
  );
  DFF_X1 \reg_pmp_7_addr[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_0541_),
    .Q(reg_pmp_7_addr[5]),
    .QN(_4506_)
  );
  DFF_X1 \reg_pmp_7_addr[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_0542_),
    .Q(reg_pmp_7_addr[6]),
    .QN(_4505_)
  );
  DFF_X1 \reg_pmp_7_addr[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_0543_),
    .Q(reg_pmp_7_addr[7]),
    .QN(_4504_)
  );
  DFF_X1 \reg_pmp_7_addr[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_0544_),
    .Q(reg_pmp_7_addr[8]),
    .QN(_4503_)
  );
  DFF_X1 \reg_pmp_7_addr[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_0545_),
    .Q(reg_pmp_7_addr[9]),
    .QN(_4502_)
  );
  DFF_X1 \reg_pmp_7_cfg_a[0]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0566_),
    .Q(reg_pmp_7_cfg_a[0]),
    .QN(_4481_)
  );
  DFF_X1 \reg_pmp_7_cfg_a[1]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0567_),
    .Q(reg_pmp_7_cfg_a[1]),
    .QN(_0004_)
  );
  DFF_X1 \reg_pmp_7_cfg_l$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0568_),
    .Q(reg_pmp_7_cfg_l),
    .QN(_0003_)
  );
  DFF_X1 \reg_pmp_7_cfg_r$_DFFE_PP_  (
    .CK(clock),
    .D(_0533_),
    .Q(reg_pmp_7_cfg_r),
    .QN(_4514_)
  );
  DFF_X1 \reg_pmp_7_cfg_w$_DFFE_PP_  (
    .CK(clock),
    .D(_0534_),
    .Q(reg_pmp_7_cfg_w),
    .QN(_4513_)
  );
  DFF_X1 \reg_pmp_7_cfg_x$_DFFE_PP_  (
    .CK(clock),
    .D(_0535_),
    .Q(reg_pmp_7_cfg_x),
    .QN(_4512_)
  );
  DFF_X1 \reg_singleStepped$_SDFF_PN0_  (
    .CK(clock),
    .D(_0247_),
    .Q(reg_singleStepped),
    .QN(_4795_)
  );
  DFF_X1 \reg_wfi$_SDFF_PP0_  (
    .CK(io_ungated_clock),
    .D(_0292_),
    .Q(reg_wfi),
    .QN(_4753_)
  );
  DFF_X1 \small_1[0]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0326_),
    .Q(small_1[0]),
    .QN(_4719_)
  );
  DFF_X1 \small_1[1]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0327_),
    .Q(small_1[1]),
    .QN(_4718_)
  );
  DFF_X1 \small_1[2]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0328_),
    .Q(small_1[2]),
    .QN(_4717_)
  );
  DFF_X1 \small_1[3]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0329_),
    .Q(small_1[3]),
    .QN(_4716_)
  );
  DFF_X1 \small_1[4]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0330_),
    .Q(small_1[4]),
    .QN(_4715_)
  );
  DFF_X1 \small_1[5]$_SDFFE_PP0P_  (
    .CK(io_ungated_clock),
    .D(_0331_),
    .Q(small_1[5]),
    .QN(_4714_)
  );
  DFF_X1 \small_[0]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0461_),
    .Q(small_[0]),
    .QN(_4585_)
  );
  DFF_X1 \small_[1]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0462_),
    .Q(small_[1]),
    .QN(_4584_)
  );
  DFF_X1 \small_[2]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0463_),
    .Q(small_[2]),
    .QN(_4583_)
  );
  DFF_X1 \small_[3]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0464_),
    .Q(small_[3]),
    .QN(_4582_)
  );
  DFF_X1 \small_[4]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0465_),
    .Q(small_[4]),
    .QN(_4581_)
  );
  DFF_X1 \small_[5]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0466_),
    .Q(small_[5]),
    .QN(_4580_)
  );
  assign _GEN_170 = 2'h0;
  assign _GEN_207 = 2'h0;
  assign _GEN_239[0] = 1'h0;
  assign _GEN_34 = { 5'h00, io_retire };
  assign _GEN_35[5:1] = 5'h00;
  assign _GEN_40 = { 20'h00000, io_interrupts_meip, 3'h0, io_interrupts_mtip, 3'h0, io_interrupts_msip, 3'h0 };
  assign _GEN_41 = { 28'h0000000, io_interrupt_cause[3:0] };
  assign _GEN_51 = 1'h1;
  assign { _GEN_586[31:2], _GEN_586[0] } = 31'h00000001;
  assign { _GEN_592[31:12], _GEN_592[10:8], _GEN_592[6:4], _GEN_592[2:0] } = 29'h00000000;
  assign _GEN_593[31:1] = 31'h00000000;
  assign { _GEN_594[31:3], _GEN_594[1] } = 30'h00000000;
  assign _GEN_595[63:32] = 32'd0;
  assign _GEN_596[63:32] = 32'd0;
  assign _GEN_597[63:32] = 32'd0;
  assign { _GEN_598[63:32], _GEN_598[30:29], _GEN_598[22:21], _GEN_598[14:13], _GEN_598[6:5] } = 40'h0000000000;
  assign { _GEN_599[63:32], _GEN_599[30:29], _GEN_599[22:21], _GEN_599[14:13], _GEN_599[6:5] } = 40'h0000000000;
  assign _GEN_600[63:30] = 34'h000000000;
  assign _GEN_601[63:30] = 34'h000000000;
  assign _GEN_602[63:30] = 34'h000000000;
  assign _GEN_603[63:30] = 34'h000000000;
  assign _GEN_604[63:30] = 34'h000000000;
  assign _GEN_605[63:30] = 34'h000000000;
  assign _GEN_606[63:30] = 34'h000000000;
  assign _GEN_607[63:30] = 34'h000000000;
  assign { _GEN_608[63:4], _GEN_608[2:0] } = 63'h0000000000000000;
  assign _GEN_609[63:1] = 63'h0000000000000000;
  assign { _GEN_610[63:30], _GEN_610[28:0] } = { 42'h00000000000, _GEN_610[29], _GEN_610[29], 6'h00, _GEN_610[29], 9'h000, _GEN_610[29], 2'h0 };
  assign { _GEN_611[31:4], _GEN_611[2:0] } = 31'h00000000;
  assign _GEN_73 = 2'h0;
  assign _T_16 = { 4'h2, reg_bp_0_control_dmode, 14'h0400, reg_bp_0_control_action, 3'h0, reg_bp_0_control_tmatch, 4'h8, reg_bp_0_control_x, reg_bp_0_control_w, reg_bp_0_control_r };
  assign _T_20 = { _GEN_586[1], 1'h1 };
  assign _T_2000[63:32] = large_1[57:26];
  assign _T_2003 = { _T_2000[31:0], large_1[25:0], small_1 };
  assign _T_2005 = { large_[57:26], _T_2000[31:0] };
  assign _T_2008 = { _T_2000[31:0], large_[25:0], small_ };
  assign { _T_21[31:2], _T_21[0] } = { _T_18[31:2], 1'h1 };
  assign _T_213 = { io_rw_addr, 20'h00000 };
  assign { _T_22[31:2], _T_22[0] } = { reg_mepc[31:2], 1'h0 };
  assign _T_23 = { 16'h4000, reg_dcsr_ebreakm, 6'h00, reg_dcsr_cause, 3'h0, reg_dcsr_step, 2'h3 };
  assign { _T_27[31:2], _T_27[0] } = { _T_24[31:2], 1'h1 };
  assign { _T_28[31:2], _T_28[0] } = { reg_dpc[31:2], 1'h0 };
  assign _T_60 = { reg_pmp_0_cfg_l, 2'h0, reg_pmp_0_cfg_a, reg_pmp_0_cfg_x, reg_pmp_0_cfg_w, reg_pmp_0_cfg_r };
  assign _T_62 = { reg_pmp_2_cfg_l, 2'h0, reg_pmp_2_cfg_a, reg_pmp_2_cfg_x, reg_pmp_2_cfg_w, reg_pmp_2_cfg_r };
  assign _T_64 = { reg_pmp_3_cfg_l, 2'h0, reg_pmp_3_cfg_a, reg_pmp_3_cfg_x, reg_pmp_3_cfg_w, reg_pmp_3_cfg_r, reg_pmp_2_cfg_l, 2'h0, reg_pmp_2_cfg_a, reg_pmp_2_cfg_x, reg_pmp_2_cfg_w, reg_pmp_2_cfg_r, reg_pmp_1_cfg_l, 2'h0, reg_pmp_1_cfg_a, reg_pmp_1_cfg_x, reg_pmp_1_cfg_w, reg_pmp_1_cfg_r, reg_pmp_0_cfg_l, 2'h0, reg_pmp_0_cfg_a, reg_pmp_0_cfg_x, reg_pmp_0_cfg_w, reg_pmp_0_cfg_r };
  assign _T_65 = { reg_pmp_4_cfg_l, 2'h0, reg_pmp_4_cfg_a, reg_pmp_4_cfg_x, reg_pmp_4_cfg_w, reg_pmp_4_cfg_r };
  assign _T_67 = { reg_pmp_6_cfg_l, 2'h0, reg_pmp_6_cfg_a, reg_pmp_6_cfg_x, reg_pmp_6_cfg_w, reg_pmp_6_cfg_r };
  assign _T_69 = { reg_pmp_7_cfg_l, 2'h0, reg_pmp_7_cfg_a, reg_pmp_7_cfg_x, reg_pmp_7_cfg_w, reg_pmp_7_cfg_r, reg_pmp_6_cfg_l, 2'h0, reg_pmp_6_cfg_a, reg_pmp_6_cfg_x, reg_pmp_6_cfg_w, reg_pmp_6_cfg_r, reg_pmp_5_cfg_l, 2'h0, reg_pmp_5_cfg_a, reg_pmp_5_cfg_x, reg_pmp_5_cfg_w, reg_pmp_5_cfg_r, reg_pmp_4_cfg_l, 2'h0, reg_pmp_4_cfg_a, reg_pmp_4_cfg_x, reg_pmp_4_cfg_w, reg_pmp_4_cfg_r };
  assign _any_T_78 = io_interrupts_debug;
  assign _causeIsDebugBreak_T_3 = { reg_dcsr_ebreakm, 3'h0 };
  assign _causeIsDebugBreak_T_4 = { 3'h0, reg_dcsr_ebreakm };
  assign { _debugTVec_T[11:4], _debugTVec_T[2:0] } = 11'h400;
  assign _decoded_T_10[1] = io_rw_addr[10];
  assign _decoded_T_14[11] = io_decode_0_inst[20];
  assign _decoded_T_16[3] = io_decode_0_inst[28];
  assign _decoded_T_18[3:2] = { io_decode_0_inst[28], io_decode_0_inst[29] };
  assign _decoded_T_2[11] = io_rw_addr[0];
  assign { _decoded_T_20[9], _decoded_T_20[3:2] } = { io_decode_0_inst[22], io_decode_0_inst[28], io_decode_0_inst[29] };
  assign _decoded_T_22[1] = io_decode_0_inst[30];
  assign _decoded_T_4[3] = io_rw_addr[8];
  assign _decoded_T_6[3:2] = { io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_T_8[9], _decoded_T_8[3:2] } = { io_rw_addr[2], io_rw_addr[8], io_rw_addr[9] };
  assign _decoded_decoded_T[3:2] = { io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_10[10], _decoded_decoded_T_10[6], _decoded_decoded_T_10[3:2] } = { io_rw_addr[1], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_100[11:9], _decoded_decoded_T_100[7:6], _decoded_decoded_T_100[4:2] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[2], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_102[8:6], _decoded_decoded_T_102[4:2] } = { io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_104[11], _decoded_decoded_T_104[8:6], _decoded_decoded_T_104[4:2] } = { io_rw_addr[0], io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_106[10], _decoded_decoded_T_106[8:6], _decoded_decoded_T_106[4:2] } = { io_rw_addr[1], io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_108[11:10], _decoded_decoded_T_108[8:6], _decoded_decoded_T_108[4:2] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_110[9:6], _decoded_decoded_T_110[4:2] } = { io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_112[11], _decoded_decoded_T_112[9:6], _decoded_decoded_T_112[4:2] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_114[10:6], _decoded_decoded_T_114[4:2] } = { io_rw_addr[1], io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_116[11:6], _decoded_decoded_T_116[4:2] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_118[6], _decoded_decoded_T_118[4:1] } = { io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[10] };
  assign { _decoded_decoded_T_12[9], _decoded_decoded_T_12[6], _decoded_decoded_T_12[3:2] } = { io_rw_addr[2], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_120[11], _decoded_decoded_T_120[6], _decoded_decoded_T_120[4:1] } = { io_rw_addr[0], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[10] };
  assign { _decoded_decoded_T_122[10], _decoded_decoded_T_122[6], _decoded_decoded_T_122[4:1] } = { io_rw_addr[1], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[10] };
  assign { _decoded_decoded_T_124[11:10], _decoded_decoded_T_124[6], _decoded_decoded_T_124[4:1] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[10] };
  assign { _decoded_decoded_T_126[7:6], _decoded_decoded_T_126[4:1] } = { io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[10] };
  assign { _decoded_decoded_T_128[11], _decoded_decoded_T_128[7:6], _decoded_decoded_T_128[4:1] } = { io_rw_addr[0], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[10] };
  assign { _decoded_decoded_T_130[10], _decoded_decoded_T_130[7:6], _decoded_decoded_T_130[4:1] } = { io_rw_addr[1], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[10] };
  assign _decoded_decoded_T_132[5:1] = { io_rw_addr[6], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[10] };
  assign { _decoded_decoded_T_134[3:2], _decoded_decoded_T_134[0] } = { io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_136[10], _decoded_decoded_T_136[3:2], _decoded_decoded_T_136[0] } = { io_rw_addr[1], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_138[11:10], _decoded_decoded_T_138[3:2], _decoded_decoded_T_138[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_14[11], _decoded_decoded_T_14[9], _decoded_decoded_T_14[6], _decoded_decoded_T_14[3:2] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_140[9], _decoded_decoded_T_140[3:2], _decoded_decoded_T_140[0] } = { io_rw_addr[2], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_142[11], _decoded_decoded_T_142[9], _decoded_decoded_T_142[3:2], _decoded_decoded_T_142[0] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_144[10:9], _decoded_decoded_T_144[3:2], _decoded_decoded_T_144[0] } = { io_rw_addr[1], io_rw_addr[2], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_146[11:9], _decoded_decoded_T_146[3:2], _decoded_decoded_T_146[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[2], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_148[8], _decoded_decoded_T_148[3:2], _decoded_decoded_T_148[0] } = { io_rw_addr[3], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_150[11], _decoded_decoded_T_150[8], _decoded_decoded_T_150[3:2], _decoded_decoded_T_150[0] } = { io_rw_addr[0], io_rw_addr[3], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_152[10], _decoded_decoded_T_152[8], _decoded_decoded_T_152[3:2], _decoded_decoded_T_152[0] } = { io_rw_addr[1], io_rw_addr[3], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_154[11:10], _decoded_decoded_T_154[8], _decoded_decoded_T_154[3:2], _decoded_decoded_T_154[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[3], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_156[9:8], _decoded_decoded_T_156[3:2], _decoded_decoded_T_156[0] } = { io_rw_addr[2], io_rw_addr[3], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_158[11], _decoded_decoded_T_158[9:8], _decoded_decoded_T_158[3:2], _decoded_decoded_T_158[0] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[3], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_16[10:9], _decoded_decoded_T_16[6], _decoded_decoded_T_16[3:2] } = { io_rw_addr[1], io_rw_addr[2], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_160[10:8], _decoded_decoded_T_160[3:2], _decoded_decoded_T_160[0] } = { io_rw_addr[1], io_rw_addr[2], io_rw_addr[3], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_162[11:8], _decoded_decoded_T_162[3:2], _decoded_decoded_T_162[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[2], io_rw_addr[3], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_164[7], _decoded_decoded_T_164[3:2], _decoded_decoded_T_164[0] } = { io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_166[11], _decoded_decoded_T_166[7], _decoded_decoded_T_166[3:2], _decoded_decoded_T_166[0] } = { io_rw_addr[0], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_168[10], _decoded_decoded_T_168[7], _decoded_decoded_T_168[3:2], _decoded_decoded_T_168[0] } = { io_rw_addr[1], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_170[11:10], _decoded_decoded_T_170[7], _decoded_decoded_T_170[3:2], _decoded_decoded_T_170[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_172[9], _decoded_decoded_T_172[7], _decoded_decoded_T_172[3:2], _decoded_decoded_T_172[0] } = { io_rw_addr[2], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_174[11], _decoded_decoded_T_174[9], _decoded_decoded_T_174[7], _decoded_decoded_T_174[3:2], _decoded_decoded_T_174[0] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_176[10:9], _decoded_decoded_T_176[7], _decoded_decoded_T_176[3:2], _decoded_decoded_T_176[0] } = { io_rw_addr[1], io_rw_addr[2], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_178[11:9], _decoded_decoded_T_178[7], _decoded_decoded_T_178[3:2], _decoded_decoded_T_178[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[2], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_18[11:9], _decoded_decoded_T_18[6], _decoded_decoded_T_18[3:2] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[2], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_180[8:7], _decoded_decoded_T_180[3:2], _decoded_decoded_T_180[0] } = { io_rw_addr[3], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_182[11], _decoded_decoded_T_182[8:7], _decoded_decoded_T_182[3:2], _decoded_decoded_T_182[0] } = { io_rw_addr[0], io_rw_addr[3], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_184[10], _decoded_decoded_T_184[8:7], _decoded_decoded_T_184[3:2], _decoded_decoded_T_184[0] } = { io_rw_addr[1], io_rw_addr[3], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_186[11:10], _decoded_decoded_T_186[8:7], _decoded_decoded_T_186[3:2], _decoded_decoded_T_186[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[3], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_188[9:7], _decoded_decoded_T_188[3:2], _decoded_decoded_T_188[0] } = { io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_190[11], _decoded_decoded_T_190[9:7], _decoded_decoded_T_190[3:2], _decoded_decoded_T_190[0] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_192[10:7], _decoded_decoded_T_192[3:2], _decoded_decoded_T_192[0] } = { io_rw_addr[1], io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_194[11:7], _decoded_decoded_T_194[3:2], _decoded_decoded_T_194[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_196[4:2], _decoded_decoded_T_196[0] } = { io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_198[10], _decoded_decoded_T_198[4:2], _decoded_decoded_T_198[0] } = { io_rw_addr[1], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_2[11], _decoded_decoded_T_2[3:2] } = { io_rw_addr[0], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_20[8], _decoded_decoded_T_20[6], _decoded_decoded_T_20[3:2] } = { io_rw_addr[3], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_200[11:10], _decoded_decoded_T_200[4:2], _decoded_decoded_T_200[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_202[9], _decoded_decoded_T_202[4:2], _decoded_decoded_T_202[0] } = { io_rw_addr[2], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_204[11], _decoded_decoded_T_204[9], _decoded_decoded_T_204[4:2], _decoded_decoded_T_204[0] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_206[10:9], _decoded_decoded_T_206[4:2], _decoded_decoded_T_206[0] } = { io_rw_addr[1], io_rw_addr[2], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_208[11:9], _decoded_decoded_T_208[4:2], _decoded_decoded_T_208[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[2], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_210[8], _decoded_decoded_T_210[4:2], _decoded_decoded_T_210[0] } = { io_rw_addr[3], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_212[11], _decoded_decoded_T_212[8], _decoded_decoded_T_212[4:2], _decoded_decoded_T_212[0] } = { io_rw_addr[0], io_rw_addr[3], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_214[10], _decoded_decoded_T_214[8], _decoded_decoded_T_214[4:2], _decoded_decoded_T_214[0] } = { io_rw_addr[1], io_rw_addr[3], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_216[11:10], _decoded_decoded_T_216[8], _decoded_decoded_T_216[4:2], _decoded_decoded_T_216[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[3], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_218[9:8], _decoded_decoded_T_218[4:2], _decoded_decoded_T_218[0] } = { io_rw_addr[2], io_rw_addr[3], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_22[11], _decoded_decoded_T_22[8], _decoded_decoded_T_22[6], _decoded_decoded_T_22[3:2] } = { io_rw_addr[0], io_rw_addr[3], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_220[11], _decoded_decoded_T_220[9:8], _decoded_decoded_T_220[4:2], _decoded_decoded_T_220[0] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[3], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_222[10:8], _decoded_decoded_T_222[4:2], _decoded_decoded_T_222[0] } = { io_rw_addr[1], io_rw_addr[2], io_rw_addr[3], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_224[11:8], _decoded_decoded_T_224[4:2], _decoded_decoded_T_224[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[2], io_rw_addr[3], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_226[7], _decoded_decoded_T_226[4:2], _decoded_decoded_T_226[0] } = { io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_228[11], _decoded_decoded_T_228[7], _decoded_decoded_T_228[4:2], _decoded_decoded_T_228[0] } = { io_rw_addr[0], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_230[10], _decoded_decoded_T_230[7], _decoded_decoded_T_230[4:2], _decoded_decoded_T_230[0] } = { io_rw_addr[1], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_232[11:10], _decoded_decoded_T_232[7], _decoded_decoded_T_232[4:2], _decoded_decoded_T_232[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_234[9], _decoded_decoded_T_234[7], _decoded_decoded_T_234[4:2], _decoded_decoded_T_234[0] } = { io_rw_addr[2], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_236[11], _decoded_decoded_T_236[9], _decoded_decoded_T_236[7], _decoded_decoded_T_236[4:2], _decoded_decoded_T_236[0] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_238[10:9], _decoded_decoded_T_238[7], _decoded_decoded_T_238[4:2], _decoded_decoded_T_238[0] } = { io_rw_addr[1], io_rw_addr[2], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_24[10], _decoded_decoded_T_24[8], _decoded_decoded_T_24[6], _decoded_decoded_T_24[3:2] } = { io_rw_addr[1], io_rw_addr[3], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_240[11:9], _decoded_decoded_T_240[7], _decoded_decoded_T_240[4:2], _decoded_decoded_T_240[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[2], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_242[8:7], _decoded_decoded_T_242[4:2], _decoded_decoded_T_242[0] } = { io_rw_addr[3], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_244[11], _decoded_decoded_T_244[8:7], _decoded_decoded_T_244[4:2], _decoded_decoded_T_244[0] } = { io_rw_addr[0], io_rw_addr[3], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_246[10], _decoded_decoded_T_246[8:7], _decoded_decoded_T_246[4:2], _decoded_decoded_T_246[0] } = { io_rw_addr[1], io_rw_addr[3], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_248[11:10], _decoded_decoded_T_248[8:7], _decoded_decoded_T_248[4:2], _decoded_decoded_T_248[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[3], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_250[9:7], _decoded_decoded_T_250[4:2], _decoded_decoded_T_250[0] } = { io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_252[11], _decoded_decoded_T_252[9:7], _decoded_decoded_T_252[4:2], _decoded_decoded_T_252[0] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_254[10:7], _decoded_decoded_T_254[4:2], _decoded_decoded_T_254[0] } = { io_rw_addr[1], io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_256[11:7], _decoded_decoded_T_256[4:2], _decoded_decoded_T_256[0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { _decoded_decoded_T_258[7], _decoded_decoded_T_258[3:0] } = { io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[10], io_rw_addr[11] };
  assign { _decoded_decoded_T_26[11:10], _decoded_decoded_T_26[8], _decoded_decoded_T_26[6], _decoded_decoded_T_26[3:2] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[3], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_260[10], _decoded_decoded_T_260[7], _decoded_decoded_T_260[3:0] } = { io_rw_addr[1], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[10], io_rw_addr[11] };
  assign _decoded_decoded_T_261 = _GEN_609[0];
  assign { _decoded_decoded_T_262[11:10], _decoded_decoded_T_262[7], _decoded_decoded_T_262[3:0] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[10], io_rw_addr[11] };
  assign _decoded_decoded_T_263 = _GEN_610[29];
  assign { _decoded_decoded_T_264[9], _decoded_decoded_T_264[7], _decoded_decoded_T_264[3:0] } = { io_rw_addr[2], io_rw_addr[4], io_rw_addr[8], io_rw_addr[9], io_rw_addr[10], io_rw_addr[11] };
  assign { _decoded_decoded_T_28[9:8], _decoded_decoded_T_28[6], _decoded_decoded_T_28[3:2] } = { io_rw_addr[2], io_rw_addr[3], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_30[11], _decoded_decoded_T_30[9:8], _decoded_decoded_T_30[6], _decoded_decoded_T_30[3:2] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[3], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_32[10:8], _decoded_decoded_T_32[6], _decoded_decoded_T_32[3:2] } = { io_rw_addr[1], io_rw_addr[2], io_rw_addr[3], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_34[11:8], _decoded_decoded_T_34[6], _decoded_decoded_T_34[3:2] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[2], io_rw_addr[3], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_36[7:6], _decoded_decoded_T_36[3:2] } = { io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_38[11], _decoded_decoded_T_38[7:6], _decoded_decoded_T_38[3:2] } = { io_rw_addr[0], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_4[9], _decoded_decoded_T_4[3:2] } = { io_rw_addr[2], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_40[10], _decoded_decoded_T_40[7:6], _decoded_decoded_T_40[3:2] } = { io_rw_addr[1], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_42[11:10], _decoded_decoded_T_42[7:6], _decoded_decoded_T_42[3:2] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_44[9], _decoded_decoded_T_44[7:6], _decoded_decoded_T_44[3:2] } = { io_rw_addr[2], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_46[11], _decoded_decoded_T_46[9], _decoded_decoded_T_46[7:6], _decoded_decoded_T_46[3:2] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_48[10:9], _decoded_decoded_T_48[7:6], _decoded_decoded_T_48[3:2] } = { io_rw_addr[1], io_rw_addr[2], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_50[11:9], _decoded_decoded_T_50[7:6], _decoded_decoded_T_50[3:2] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[2], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_52[8:6], _decoded_decoded_T_52[3:2] } = { io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_54[11], _decoded_decoded_T_54[8:6], _decoded_decoded_T_54[3:2] } = { io_rw_addr[0], io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_56[10], _decoded_decoded_T_56[8:6], _decoded_decoded_T_56[3:2] } = { io_rw_addr[1], io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_58[11:10], _decoded_decoded_T_58[8:6], _decoded_decoded_T_58[3:2] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_6[11], _decoded_decoded_T_6[9], _decoded_decoded_T_6[3:2] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_60[9:6], _decoded_decoded_T_60[3:2] } = { io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_62[11], _decoded_decoded_T_62[9:6], _decoded_decoded_T_62[3:2] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_64[10:6], _decoded_decoded_T_64[3:2] } = { io_rw_addr[1], io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_66[11:6], _decoded_decoded_T_66[3:2] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[2], io_rw_addr[3], io_rw_addr[4], io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_68[5], _decoded_decoded_T_68[3:2] } = { io_rw_addr[6], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_70[11], _decoded_decoded_T_70[5], _decoded_decoded_T_70[3:2] } = { io_rw_addr[0], io_rw_addr[6], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_72[10], _decoded_decoded_T_72[5], _decoded_decoded_T_72[3:2] } = { io_rw_addr[1], io_rw_addr[6], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_74[11:10], _decoded_decoded_T_74[5], _decoded_decoded_T_74[3:2] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[6], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_76[9], _decoded_decoded_T_76[5], _decoded_decoded_T_76[3:2] } = { io_rw_addr[2], io_rw_addr[6], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_78[6], _decoded_decoded_T_78[4:2] } = { io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_8[6], _decoded_decoded_T_8[3:2] } = { io_rw_addr[5], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_80[11], _decoded_decoded_T_80[6], _decoded_decoded_T_80[4:2] } = { io_rw_addr[0], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_82[10], _decoded_decoded_T_82[6], _decoded_decoded_T_82[4:2] } = { io_rw_addr[1], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_84[11:10], _decoded_decoded_T_84[6], _decoded_decoded_T_84[4:2] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_86[7:6], _decoded_decoded_T_86[4:2] } = { io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_88[11], _decoded_decoded_T_88[7:6], _decoded_decoded_T_88[4:2] } = { io_rw_addr[0], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_90[10], _decoded_decoded_T_90[7:6], _decoded_decoded_T_90[4:2] } = { io_rw_addr[1], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_92[11:10], _decoded_decoded_T_92[7:6], _decoded_decoded_T_92[4:2] } = { io_rw_addr[0], io_rw_addr[1], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_94[9], _decoded_decoded_T_94[7:6], _decoded_decoded_T_94[4:2] } = { io_rw_addr[2], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_96[11], _decoded_decoded_T_96[9], _decoded_decoded_T_96[7:6], _decoded_decoded_T_96[4:2] } = { io_rw_addr[0], io_rw_addr[2], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign { _decoded_decoded_T_98[10:9], _decoded_decoded_T_98[7:6], _decoded_decoded_T_98[4:2] } = { io_rw_addr[1], io_rw_addr[2], io_rw_addr[4], io_rw_addr[5], io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign _decoded_decoded_orMatrixOutputs_T = _GEN_610[29];
  assign _decoded_decoded_orMatrixOutputs_T_2 = _GEN_609[0];
  assign _epc_T_1[0] = 1'h1;
  assign { _io_decode_0_read_illegal_T_12[7:6], _io_decode_0_read_illegal_T_12[4:1] } = { io_decode_0_inst[24], io_decode_0_inst[25], io_decode_0_inst[27], io_decode_0_inst[28], io_decode_0_inst[29], io_decode_0_inst[30] };
  assign _io_decode_0_read_illegal_T_17 = io_decode_0_read_illegal;
  assign _io_decode_0_read_illegal_T_21 = 1'h0;
  assign { _io_rw_rdata_T_1[31:30], _io_rw_rdata_T_1[28], _io_rw_rdata_T_1[26:24], _io_rw_rdata_T_1[22:13], _io_rw_rdata_T_1[11:9], _io_rw_rdata_T_1[5:3] } = 22'h000000;
  assign _io_rw_rdata_T_10[0] = 1'h0;
  assign _io_rw_rdata_T_107 = _GEN_596[31:0];
  assign _io_rw_rdata_T_108 = _GEN_597[31:0];
  assign _io_rw_rdata_T_109 = { _GEN_598[31], 2'h0, _GEN_598[28:23], 2'h0, _GEN_598[20:15], 2'h0, _GEN_598[12:7], 2'h0, _GEN_598[4:0] };
  assign _io_rw_rdata_T_110 = { _GEN_599[31], 2'h0, _GEN_599[28:23], 2'h0, _GEN_599[20:15], 2'h0, _GEN_599[12:7], 2'h0, _GEN_599[4:0] };
  assign _io_rw_rdata_T_113 = _GEN_600[29:0];
  assign _io_rw_rdata_T_114 = _GEN_601[29:0];
  assign _io_rw_rdata_T_115 = _GEN_602[29:0];
  assign _io_rw_rdata_T_116 = _GEN_603[29:0];
  assign _io_rw_rdata_T_117 = _GEN_604[29:0];
  assign _io_rw_rdata_T_118 = _GEN_605[29:0];
  assign _io_rw_rdata_T_119 = _GEN_606[29:0];
  assign _io_rw_rdata_T_120 = _GEN_607[29:0];
  assign _io_rw_rdata_T_129 = { 28'h0000000, _GEN_608[3], 3'h0 };
  assign _io_rw_rdata_T_13 = _GEN_593[0];
  assign _io_rw_rdata_T_130 = { 31'h00000000, _GEN_609[0] };
  assign _io_rw_rdata_T_132 = { 2'h0, _GEN_610[29], 8'h00, _GEN_610[29], _GEN_610[29], 6'h00, _GEN_610[29], 9'h000, _GEN_610[29], 2'h0 };
  assign { _io_rw_rdata_T_14[31], _io_rw_rdata_T_14[29:16], _io_rw_rdata_T_14[14:9], _io_rw_rdata_T_14[5:3] } = 24'h000000;
  assign { _io_rw_rdata_T_148[31:3], _io_rw_rdata_T_148[1] } = { _GEN_595[31:3], _GEN_595[1] };
  assign _io_rw_rdata_T_149 = _GEN_595[31:0];
  assign _io_rw_rdata_T_15[0] = 1'h0;
  assign _io_rw_rdata_T_17 = { _GEN_594[2], 1'h0, _GEN_594[0] };
  assign _io_rw_rdata_T_240[30] = io_rw_rdata[30];
  assign { _io_rw_rdata_T_241[30:29], _io_rw_rdata_T_241[22:21], _io_rw_rdata_T_241[14:13], _io_rw_rdata_T_241[6:5] } = { io_rw_rdata[30], _io_rw_rdata_T_240[29], _io_rw_rdata_T_240[22:21], _io_rw_rdata_T_240[14:13], _io_rw_rdata_T_240[6:5] };
  assign { _io_rw_rdata_T_242[31:29], _io_rw_rdata_T_242[22:21], _io_rw_rdata_T_242[14:13], _io_rw_rdata_T_242[6:5] } = { io_rw_rdata[31:30], _io_rw_rdata_T_240[29], _io_rw_rdata_T_240[22:21], _io_rw_rdata_T_240[14:13], _io_rw_rdata_T_240[6:5] };
  assign _io_rw_rdata_T_245[31:30] = io_rw_rdata[31:30];
  assign _io_rw_rdata_T_246[31:30] = io_rw_rdata[31:30];
  assign _io_rw_rdata_T_247[31:30] = io_rw_rdata[31:30];
  assign _io_rw_rdata_T_248[31:30] = io_rw_rdata[31:30];
  assign _io_rw_rdata_T_249[31:30] = io_rw_rdata[31:30];
  assign _io_rw_rdata_T_250[31:30] = io_rw_rdata[31:30];
  assign _io_rw_rdata_T_251[31:30] = io_rw_rdata[31:30];
  assign { _io_rw_rdata_T_252[31:30], _io_rw_rdata_T_252[28:21], _io_rw_rdata_T_252[18:13], _io_rw_rdata_T_252[11:4], _io_rw_rdata_T_252[1] } = { io_rw_rdata[31:30], io_rw_rdata[28:21], io_rw_rdata[18:13], io_rw_rdata[11:4], io_rw_rdata[1] };
  assign _io_rw_rdata_T_261[31:0] = { io_rw_rdata[31:30], _io_rw_rdata_T_252[29], io_rw_rdata[28:21], _io_rw_rdata_T_252[20:19], io_rw_rdata[18:13], _io_rw_rdata_T_252[12], io_rw_rdata[11:3], _io_rw_rdata_T_252[2], io_rw_rdata[1], _io_rw_rdata_T_252[0] };
  assign _io_rw_rdata_T_262[31:0] = { io_rw_rdata[31:30], _io_rw_rdata_T_252[29], io_rw_rdata[28:21], _io_rw_rdata_T_252[20:19], io_rw_rdata[18:13], _io_rw_rdata_T_252[12], io_rw_rdata[11:3], _io_rw_rdata_T_252[2], io_rw_rdata[1:0] };
  assign _io_rw_rdata_T_264[31:0] = io_rw_rdata;
  assign { _io_rw_rdata_T_4[31], _io_rw_rdata_T_4[29:24], _io_rw_rdata_T_4[22:13], _io_rw_rdata_T_4[11:9], _io_rw_rdata_T_4[7:3], _io_rw_rdata_T_4[1] } = 26'h0000000;
  assign { _io_rw_rdata_T_5[31:13], _io_rw_rdata_T_5[10:8], _io_rw_rdata_T_5[6:4], _io_rw_rdata_T_5[2:0] } = 28'h0000000;
  assign _io_rw_rdata_T_6[1] = 1'h0;
  assign _io_rw_rdata_T_7 = { 4'h0, _GEN_592[11], 3'h0, _GEN_592[7], 3'h0, _GEN_592[3], 3'h0 };
  assign { _io_rw_rdata_T_8[31:12], _io_rw_rdata_T_8[10:8], _io_rw_rdata_T_8[6:4], _io_rw_rdata_T_8[2:0] } = 29'h00000000;
  assign { _m_interrupts_T_3[31:12], _m_interrupts_T_3[10:8], _m_interrupts_T_3[6:4], _m_interrupts_T_3[2:0] } = 29'h1fffffff;
  assign { _m_interrupts_T_5[31:12], _m_interrupts_T_5[10:8], _m_interrupts_T_5[6:4], _m_interrupts_T_5[2:0] } = 29'h00000000;
  assign { _newBPC_T_2[31:28], _newBPC_T_2[26:13], _newBPC_T_2[11:9], _newBPC_T_2[6:3] } = { 2'h0, io_rw_cmd[1], 4'h0, io_rw_cmd[1], 13'h0000, io_rw_cmd[1], 3'h0 };
  assign { _newBPC_T_3[31:30], _newBPC_T_3[28], _newBPC_T_3[26:24], _newBPC_T_3[22:13], _newBPC_T_3[11:9], _newBPC_T_3[5:3] } = { io_rw_wdata[31:30], io_rw_wdata[28], io_rw_wdata[26:24], io_rw_wdata[22:13], io_rw_wdata[11:9], io_rw_wdata[5:3] };
  assign _new_mstatus_WIRE = { 73'h0000000000000000000, _T_2000[31:0] };
  assign { _notDebugTVec_T_1[31:7], _notDebugTVec_T_1[1:0] } = { reg_mtvec[31:7], 2'h0 };
  assign _pmp_mask_T_12[0] = reg_pmp_2_cfg_a[0];
  assign _pmp_mask_T_13[29:0] = { io_pmp_2_mask[31:3], reg_pmp_2_cfg_a[0] };
  assign _pmp_mask_T_14 = { _pmp_mask_T_13[30], io_pmp_2_mask[31:3], reg_pmp_2_cfg_a[0], 2'h3 };
  assign _pmp_mask_T_17[0] = reg_pmp_3_cfg_a[0];
  assign _pmp_mask_T_18[29:0] = { io_pmp_3_mask[31:3], reg_pmp_3_cfg_a[0] };
  assign _pmp_mask_T_19 = { _pmp_mask_T_18[30], io_pmp_3_mask[31:3], reg_pmp_3_cfg_a[0], 2'h3 };
  assign _pmp_mask_T_2[0] = reg_pmp_0_cfg_a[0];
  assign _pmp_mask_T_22[0] = reg_pmp_4_cfg_a[0];
  assign _pmp_mask_T_23[29:0] = { io_pmp_4_mask[31:3], reg_pmp_4_cfg_a[0] };
  assign _pmp_mask_T_24 = { _pmp_mask_T_23[30], io_pmp_4_mask[31:3], reg_pmp_4_cfg_a[0], 2'h3 };
  assign _pmp_mask_T_27[0] = reg_pmp_5_cfg_a[0];
  assign _pmp_mask_T_28[29:0] = { io_pmp_5_mask[31:3], reg_pmp_5_cfg_a[0] };
  assign _pmp_mask_T_29 = { _pmp_mask_T_28[30], io_pmp_5_mask[31:3], reg_pmp_5_cfg_a[0], 2'h3 };
  assign _pmp_mask_T_3[29:0] = { io_pmp_0_mask[31:3], reg_pmp_0_cfg_a[0] };
  assign _pmp_mask_T_32[0] = reg_pmp_6_cfg_a[0];
  assign _pmp_mask_T_33[29:0] = { io_pmp_6_mask[31:3], reg_pmp_6_cfg_a[0] };
  assign _pmp_mask_T_34 = { _pmp_mask_T_33[30], io_pmp_6_mask[31:3], reg_pmp_6_cfg_a[0], 2'h3 };
  assign _pmp_mask_T_37[0] = reg_pmp_7_cfg_a[0];
  assign _pmp_mask_T_38[29:0] = { io_pmp_7_mask[31:3], reg_pmp_7_cfg_a[0] };
  assign _pmp_mask_T_39 = { _pmp_mask_T_38[30], io_pmp_7_mask[31:3], reg_pmp_7_cfg_a[0], 2'h3 };
  assign _pmp_mask_T_4 = { _pmp_mask_T_3[30], io_pmp_0_mask[31:3], reg_pmp_0_cfg_a[0], 2'h3 };
  assign _pmp_mask_T_7[0] = reg_pmp_1_cfg_a[0];
  assign _pmp_mask_T_8[29:0] = { io_pmp_1_mask[31:3], reg_pmp_1_cfg_a[0] };
  assign _pmp_mask_T_9 = { _pmp_mask_T_8[30], io_pmp_1_mask[31:3], reg_pmp_1_cfg_a[0], 2'h3 };
  assign _read_mip_T = { 4'h0, io_interrupts_meip, 3'h0, io_interrupts_mtip, 3'h0, io_interrupts_msip, 3'h0 };
  assign _read_mstatus_T = { reg_debug, io_status_cease_r, reg_wfi, 19'h20400, reg_misa[12], 9'h020, reg_misa[2], 1'h0, reg_misa[0], 31'h6c000000, reg_mstatus_gva, 30'h00000018, reg_mstatus_mpie, 3'h0, reg_mstatus_mie, 3'h0 };
  assign _read_mtvec_T_1 = { reg_mtvec[0], reg_mtvec[0], reg_mtvec[0], reg_mtvec[0], reg_mtvec[0], 2'h2 };
  assign _read_mtvec_T_3 = { 25'h0000000, reg_mtvec[0], reg_mtvec[0], reg_mtvec[0], reg_mtvec[0], reg_mtvec[0], 2'h2 };
  assign { _read_mtvec_T_4[31:7], _read_mtvec_T_4[5:0] } = { 25'h1ffffff, _read_mtvec_T_4[6], _read_mtvec_T_4[6], _read_mtvec_T_4[6], _read_mtvec_T_4[6], 2'h1 };
  assign _reg_custom_0_T = { 28'h0000000, _T_2000[3], 3'h0 };
  assign _reg_custom_0_T_2 = 32'd0;
  assign _reg_custom_0_T_3 = { 28'h0000000, _T_2000[3], 3'h0 };
  assign _reg_dcsr_cause_T_2[2] = reg_singleStepped;
  assign _reg_mcause_T = { _T_2000[31], 27'h0000000, _T_2000[3:0] };
  assign _reg_mcountinhibit_T_1 = { _T_2000[31:2], 1'h0, _T_2000[0] };
  assign { _reg_mepc_T_1[5], _reg_mepc_T_1[0] } = { _GEN_611[3], 1'h1 };
  assign _reg_mepc_T_2 = { _T_2000[31:1], 1'h0 };
  assign _reg_mie_T = { 20'h00000, _T_2000[11], 3'h0, _T_2000[7], 3'h0, _T_2000[3], 3'h0 };
  assign _reg_misa_T[31:1] = { _reg_mepc_T_1[31:6], _GEN_611[3], _reg_mepc_T_1[4:1] };
  assign _reg_misa_T_1 = _GEN_611[3];
  assign _reg_misa_T_2 = { _GEN_611[3], 3'h0 };
  assign { _reg_misa_T_3[31:4], _reg_misa_T_3[2:0] } = { _reg_mepc_T_1[31:6], _GEN_611[3], _reg_mepc_T_1[4], _reg_mepc_T_1[2:1], _reg_misa_T[0] };
  assign { _reg_misa_T_4[31:4], _reg_misa_T_4[2:0] } = { _T_2000[31:4], _T_2000[2:0] };
  assign _reg_misa_T_5 = { 19'h00000, _T_2000[12], 9'h000, _T_2000[2], 1'h0, _T_2000[0] };
  assign _reg_misa_T_7 = 32'd1082130688;
  assign _reg_misa_T_8 = { 19'h20400, _T_2000[12], 9'h020, _T_2000[2], 1'h0, _T_2000[0] };
  assign _which_T_100 = 4'h4;
  assign _which_T_101 = 4'h4;
  assign _which_T_102 = 4'h4;
  assign { _which_T_103[3:2], _which_T_103[0] } = { 2'h1, _which_T_103[1] };
  assign { _which_T_104[3], _which_T_104[0] } = { 1'h0, _which_T_104[1] };
  assign _which_T_105[0] = _which_T_105[1];
  assign _which_T_106 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_107 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_108 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_109 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_111 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_112 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_113 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_114 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_115 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_116 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_117 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_118 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_119 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_120 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_121 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_122 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_123 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_124 = { _which_T_105[3:1], _which_T_105[1] };
  assign _which_T_95 = 4'h4;
  assign _which_T_96 = 4'h4;
  assign _which_T_97 = 4'h4;
  assign _which_T_98 = 4'h4;
  assign _which_T_99 = 4'h4;
  assign addr = { 1'h0, io_rw_addr };
  assign addr_1 = io_decode_0_inst[31:20];
  assign d_interrupts = { io_interrupts_debug, 14'h0000 };
  assign { debugTVec[11:4], debugTVec[2:0] } = 11'h400;
  assign decoded_130 = _GEN_609[0];
  assign decoded_132 = _GEN_610[29];
  assign decoded_andMatrixInput_0_1 = io_rw_addr[0];
  assign decoded_andMatrixInput_0_10 = io_decode_0_inst[22];
  assign decoded_andMatrixInput_0_11 = io_decode_0_inst[30];
  assign decoded_andMatrixInput_0_2 = io_rw_addr[8];
  assign decoded_andMatrixInput_0_4 = io_rw_addr[2];
  assign decoded_andMatrixInput_0_5 = io_rw_addr[10];
  assign decoded_andMatrixInput_0_7 = io_decode_0_inst[20];
  assign decoded_andMatrixInput_0_8 = io_decode_0_inst[28];
  assign decoded_andMatrixInput_7_2 = io_rw_addr[9];
  assign decoded_andMatrixInput_7_6 = io_decode_0_inst[29];
  assign decoded_decoded_andMatrixInput_0_1 = io_rw_addr[0];
  assign decoded_decoded_andMatrixInput_0_5 = io_rw_addr[1];
  assign decoded_decoded_andMatrixInput_10_58 = io_rw_addr[10];
  assign decoded_decoded_andMatrixInput_10_65 = io_rw_addr[11];
  assign decoded_decoded_andMatrixInput_2_2 = io_rw_addr[2];
  assign decoded_decoded_andMatrixInput_3_10 = io_rw_addr[3];
  assign decoded_decoded_andMatrixInput_4_18 = io_rw_addr[4];
  assign decoded_decoded_andMatrixInput_4_4 = io_rw_addr[5];
  assign decoded_decoded_andMatrixInput_6_34 = io_rw_addr[6];
  assign decoded_decoded_andMatrixInput_7_39 = io_rw_addr[7];
  assign decoded_decoded_andMatrixInput_8 = io_rw_addr[8];
  assign decoded_decoded_andMatrixInput_9 = io_rw_addr[9];
  assign { decoded_decoded_invMatrixOutputs[2], decoded_decoded_invMatrixOutputs[0] } = { _GEN_609[0], _GEN_610[29] };
  assign { decoded_decoded_invMatrixOutputs_lo_lo[2], decoded_decoded_invMatrixOutputs_lo_lo[0] } = { _GEN_609[0], _GEN_610[29] };
  assign { decoded_decoded_invMatrixOutputs_lo_lo_lo_lo[2], decoded_decoded_invMatrixOutputs_lo_lo_lo_lo[0] } = { _GEN_609[0], _GEN_610[29] };
  assign decoded_decoded_lo[3:2] = { io_rw_addr[8], io_rw_addr[9] };
  assign decoded_decoded_lo_129[3:0] = { io_rw_addr[8], io_rw_addr[9], io_rw_addr[10], io_rw_addr[11] };
  assign decoded_decoded_lo_130[3:0] = { io_rw_addr[8], io_rw_addr[9], io_rw_addr[10], io_rw_addr[11] };
  assign { decoded_decoded_lo_34[5], decoded_decoded_lo_34[3:2] } = { io_rw_addr[6], io_rw_addr[8], io_rw_addr[9] };
  assign decoded_decoded_lo_39[4:2] = { io_rw_addr[7], io_rw_addr[8], io_rw_addr[9] };
  assign decoded_decoded_lo_4[3:2] = { io_rw_addr[8], io_rw_addr[9] };
  assign decoded_decoded_lo_59[4:1] = { io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[10] };
  assign decoded_decoded_lo_65[4:1] = { io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[10] };
  assign { decoded_decoded_lo_67[3:2], decoded_decoded_lo_67[0] } = { io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { decoded_decoded_lo_68[3:2], decoded_decoded_lo_68[0] } = { io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { decoded_decoded_lo_98[4:2], decoded_decoded_lo_98[0] } = { io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { decoded_decoded_lo_99[4:2], decoded_decoded_lo_99[0] } = { io_rw_addr[7], io_rw_addr[8], io_rw_addr[9], io_rw_addr[11] };
  assign { decoded_decoded_orMatrixOutputs[2], decoded_decoded_orMatrixOutputs[0] } = { _GEN_609[0], _GEN_610[29] };
  assign { decoded_decoded_orMatrixOutputs_lo_lo[2], decoded_decoded_orMatrixOutputs_lo_lo[0] } = { _GEN_609[0], _GEN_610[29] };
  assign { decoded_decoded_orMatrixOutputs_lo_lo_lo_lo[2], decoded_decoded_orMatrixOutputs_lo_lo_lo_lo[0] } = { _GEN_609[0], _GEN_610[29] };
  assign decoded_decoded_plaInput = io_rw_addr;
  assign decoded_invInputs[19:0] = 20'hfff8c;
  assign decoded_invMatrixOutputs[3:0] = 4'h0;
  assign decoded_invMatrixOutputs_1[3:0] = 4'h0;
  assign decoded_orMatrixOutputs[3:0] = 4'h0;
  assign decoded_orMatrixOutputs_1[3:0] = 4'h0;
  assign decoded_plaInput = { io_rw_addr, 20'h00073 };
  assign epc = { io_pc[31:1], 1'h0 };
  assign exception = io_trace_0_exception;
  assign f = _T_2000[5];
  assign io_bp_0_address = reg_bp_0_address;
  assign io_bp_0_control_action = reg_bp_0_control_action;
  assign io_bp_0_control_r = reg_bp_0_control_r;
  assign io_bp_0_control_tmatch = reg_bp_0_control_tmatch;
  assign io_bp_0_control_w = reg_bp_0_control_w;
  assign io_bp_0_control_x = reg_bp_0_control_x;
  assign io_customCSRs_0_value = { 28'h0000000, reg_custom_0[3], 3'h0 };
  assign io_decode_0_fp_csr = 1'h0;
  assign io_decode_0_fp_illegal = 1'h1;
  assign io_decode_0_read_illegal_andMatrixInput_0 = io_decode_0_inst[24];
  assign io_decode_0_read_illegal_andMatrixInput_1 = io_decode_0_inst[25];
  assign io_decode_0_read_illegal_andMatrixInput_3 = io_decode_0_inst[27];
  assign io_decode_0_read_illegal_andMatrixInput_4 = io_decode_0_inst[28];
  assign io_decode_0_read_illegal_andMatrixInput_5 = io_decode_0_inst[29];
  assign io_decode_0_read_illegal_andMatrixInput_6 = io_decode_0_inst[30];
  assign io_decode_0_rocc_illegal = 1'h1;
  assign io_decode_0_write_flush_addr_m = { io_decode_0_inst[31:30], 2'h3, io_decode_0_inst[27:20] };
  assign io_evec[0] = 1'h0;
  assign io_inhibit_cycle = reg_mcountinhibit[0];
  assign io_interrupt_cause[31:4] = 28'h8000000;
  assign io_pmp_0_addr = reg_pmp_0_addr;
  assign io_pmp_0_cfg_a = reg_pmp_0_cfg_a;
  assign io_pmp_0_cfg_l = reg_pmp_0_cfg_l;
  assign io_pmp_0_cfg_r = reg_pmp_0_cfg_r;
  assign io_pmp_0_cfg_w = reg_pmp_0_cfg_w;
  assign io_pmp_0_cfg_x = reg_pmp_0_cfg_x;
  assign io_pmp_0_mask[2:0] = { reg_pmp_0_cfg_a[0], 2'h3 };
  assign io_pmp_1_addr = reg_pmp_1_addr;
  assign io_pmp_1_cfg_a = reg_pmp_1_cfg_a;
  assign io_pmp_1_cfg_l = reg_pmp_1_cfg_l;
  assign io_pmp_1_cfg_r = reg_pmp_1_cfg_r;
  assign io_pmp_1_cfg_w = reg_pmp_1_cfg_w;
  assign io_pmp_1_cfg_x = reg_pmp_1_cfg_x;
  assign io_pmp_1_mask[2:0] = { reg_pmp_1_cfg_a[0], 2'h3 };
  assign io_pmp_2_addr = reg_pmp_2_addr;
  assign io_pmp_2_cfg_a = reg_pmp_2_cfg_a;
  assign io_pmp_2_cfg_l = reg_pmp_2_cfg_l;
  assign io_pmp_2_cfg_r = reg_pmp_2_cfg_r;
  assign io_pmp_2_cfg_w = reg_pmp_2_cfg_w;
  assign io_pmp_2_cfg_x = reg_pmp_2_cfg_x;
  assign io_pmp_2_mask[2:0] = { reg_pmp_2_cfg_a[0], 2'h3 };
  assign io_pmp_3_addr = reg_pmp_3_addr;
  assign io_pmp_3_cfg_a = reg_pmp_3_cfg_a;
  assign io_pmp_3_cfg_l = reg_pmp_3_cfg_l;
  assign io_pmp_3_cfg_r = reg_pmp_3_cfg_r;
  assign io_pmp_3_cfg_w = reg_pmp_3_cfg_w;
  assign io_pmp_3_cfg_x = reg_pmp_3_cfg_x;
  assign io_pmp_3_mask[2:0] = { reg_pmp_3_cfg_a[0], 2'h3 };
  assign io_pmp_4_addr = reg_pmp_4_addr;
  assign io_pmp_4_cfg_a = reg_pmp_4_cfg_a;
  assign io_pmp_4_cfg_l = reg_pmp_4_cfg_l;
  assign io_pmp_4_cfg_r = reg_pmp_4_cfg_r;
  assign io_pmp_4_cfg_w = reg_pmp_4_cfg_w;
  assign io_pmp_4_cfg_x = reg_pmp_4_cfg_x;
  assign io_pmp_4_mask[2:0] = { reg_pmp_4_cfg_a[0], 2'h3 };
  assign io_pmp_5_addr = reg_pmp_5_addr;
  assign io_pmp_5_cfg_a = reg_pmp_5_cfg_a;
  assign io_pmp_5_cfg_l = reg_pmp_5_cfg_l;
  assign io_pmp_5_cfg_r = reg_pmp_5_cfg_r;
  assign io_pmp_5_cfg_w = reg_pmp_5_cfg_w;
  assign io_pmp_5_cfg_x = reg_pmp_5_cfg_x;
  assign io_pmp_5_mask[2:0] = { reg_pmp_5_cfg_a[0], 2'h3 };
  assign io_pmp_6_addr = reg_pmp_6_addr;
  assign io_pmp_6_cfg_a = reg_pmp_6_cfg_a;
  assign io_pmp_6_cfg_l = reg_pmp_6_cfg_l;
  assign io_pmp_6_cfg_r = reg_pmp_6_cfg_r;
  assign io_pmp_6_cfg_w = reg_pmp_6_cfg_w;
  assign io_pmp_6_cfg_x = reg_pmp_6_cfg_x;
  assign io_pmp_6_mask[2:0] = { reg_pmp_6_cfg_a[0], 2'h3 };
  assign io_pmp_7_addr = reg_pmp_7_addr;
  assign io_pmp_7_cfg_a = reg_pmp_7_cfg_a;
  assign io_pmp_7_cfg_l = reg_pmp_7_cfg_l;
  assign io_pmp_7_cfg_r = reg_pmp_7_cfg_r;
  assign io_pmp_7_cfg_w = reg_pmp_7_cfg_w;
  assign io_pmp_7_cfg_x = reg_pmp_7_cfg_x;
  assign io_pmp_7_mask[2:0] = { reg_pmp_7_cfg_a[0], 2'h3 };
  assign io_status_cease = io_status_cease_r;
  assign io_status_debug = reg_debug;
  assign io_status_dprv = 2'h3;
  assign io_status_dv = 1'h0;
  assign io_status_fs = 2'h0;
  assign io_status_gva = reg_mstatus_gva;
  assign io_status_hie = 1'h0;
  assign io_status_isa = { 19'h20400, reg_misa[12], 9'h020, reg_misa[2], 1'h0, reg_misa[0] };
  assign io_status_mbe = 1'h0;
  assign io_status_mie = reg_mstatus_mie;
  assign io_status_mpie = reg_mstatus_mpie;
  assign io_status_mpp = 2'h3;
  assign io_status_mprv = 1'h0;
  assign io_status_mpv = 1'h0;
  assign io_status_mxr = 1'h0;
  assign io_status_prv = 2'h3;
  assign io_status_sbe = 1'h0;
  assign io_status_sd = 1'h0;
  assign io_status_sd_rv32 = 1'h0;
  assign io_status_sie = 1'h0;
  assign io_status_spie = 1'h0;
  assign io_status_spp = 1'h0;
  assign io_status_sum = 1'h0;
  assign io_status_sxl = 2'h0;
  assign io_status_tsr = 1'h0;
  assign io_status_tvm = 1'h0;
  assign io_status_tw = 1'h0;
  assign io_status_ube = 1'h0;
  assign io_status_uie = 1'h0;
  assign io_status_upie = 1'h0;
  assign io_status_uxl = 2'h0;
  assign io_status_v = 1'h0;
  assign io_status_vs = 2'h0;
  assign io_status_wfi = reg_wfi;
  assign io_status_xs = 2'h0;
  assign io_status_zero1 = 8'h00;
  assign io_status_zero2 = 23'h000000;
  assign io_time = { large_1[25:0], small_1 };
  assign io_trace_0_iaddr = io_pc;
  assign io_trace_0_insn = io_inst_0;
  assign lo_11 = { reg_pmp_1_cfg_l, 2'h0, reg_pmp_1_cfg_a, reg_pmp_1_cfg_x, reg_pmp_1_cfg_w, reg_pmp_1_cfg_r, reg_pmp_0_cfg_l, 2'h0, reg_pmp_0_cfg_a, reg_pmp_0_cfg_x, reg_pmp_0_cfg_w, reg_pmp_0_cfg_r };
  assign lo_16 = { reg_pmp_5_cfg_l, 2'h0, reg_pmp_5_cfg_a, reg_pmp_5_cfg_x, reg_pmp_5_cfg_w, reg_pmp_5_cfg_r, reg_pmp_4_cfg_l, 2'h0, reg_pmp_4_cfg_a, reg_pmp_4_cfg_x, reg_pmp_4_cfg_w, reg_pmp_4_cfg_r };
  assign lo_4 = { 4'h8, reg_bp_0_control_x, reg_bp_0_control_w, reg_bp_0_control_r };
  assign { m_interrupts[31:4], m_interrupts[2:0] } = { 20'h00000, _which_T_105[3], 3'h0, _which_T_103[1], 6'h00 };
  assign newCfg_1_a = _T_2000[12:11];
  assign newCfg_1_l = _T_2000[15];
  assign newCfg_1_r = _T_2000[8];
  assign newCfg_1_w = _T_2000[9];
  assign newCfg_1_x = _T_2000[10];
  assign newCfg_2_a = _T_2000[20:19];
  assign newCfg_2_l = _T_2000[23];
  assign newCfg_2_r = _T_2000[16];
  assign newCfg_2_w = _T_2000[17];
  assign newCfg_2_x = _T_2000[18];
  assign newCfg_3_a = _T_2000[28:27];
  assign newCfg_3_l = _T_2000[31];
  assign newCfg_3_r = _T_2000[24];
  assign newCfg_3_w = _T_2000[25];
  assign newCfg_3_x = _T_2000[26];
  assign newCfg_a = _T_2000[4:3];
  assign newCfg_l = _T_2000[7];
  assign newCfg_r = _T_2000[0];
  assign newCfg_w = _T_2000[1];
  assign newCfg_x = _T_2000[2];
  assign new_dcsr_ebreakm = _T_2000[15];
  assign new_mstatus_mie = _T_2000[3];
  assign new_mstatus_mpie = _T_2000[7];
  assign { notDebugTVec[31:7], notDebugTVec[1:0] } = { reg_mtvec[31:7], 2'h0 };
  assign notDebugTVec_interruptOffset[1:0] = 2'h0;
  assign { notDebugTVec_interruptVec[31:7], notDebugTVec_interruptVec[1:0] } = { reg_mtvec[31:7], 2'h0 };
  assign pending_interrupts = { 20'h00000, _m_interrupts_T_5[11], 3'h0, _m_interrupts_T_5[7], 3'h0, _m_interrupts_T_5[3], 3'h0 };
  assign pmp_mask_base = { reg_pmp_0_addr, reg_pmp_0_cfg_a[0] };
  assign pmp_mask_base_1 = { reg_pmp_1_addr, reg_pmp_1_cfg_a[0] };
  assign pmp_mask_base_2 = { reg_pmp_2_addr, reg_pmp_2_cfg_a[0] };
  assign pmp_mask_base_3 = { reg_pmp_3_addr, reg_pmp_3_cfg_a[0] };
  assign pmp_mask_base_4 = { reg_pmp_4_addr, reg_pmp_4_cfg_a[0] };
  assign pmp_mask_base_5 = { reg_pmp_5_addr, reg_pmp_5_cfg_a[0] };
  assign pmp_mask_base_6 = { reg_pmp_6_addr, reg_pmp_6_cfg_a[0] };
  assign pmp_mask_base_7 = { reg_pmp_7_addr, reg_pmp_7_cfg_a[0] };
  assign read_mip = { 4'h0, io_interrupts_meip, 3'h0, io_interrupts_mtip, 3'h0, io_interrupts_msip, 3'h0 };
  assign read_mstatus = { 24'h000018, reg_mstatus_mpie, 3'h0, reg_mstatus_mie, 3'h0 };
  assign read_mstatus_hi = { reg_debug, io_status_cease_r, reg_wfi, 19'h20400, reg_misa[12], 9'h020, reg_misa[2], 1'h0, reg_misa[0], 31'h6c000000, reg_mstatus_gva, 16'h0000 };
  assign read_mstatus_hi_hi = { reg_debug, io_status_cease_r, reg_wfi, 19'h20400, reg_misa[12], 9'h020, reg_misa[2], 1'h0, reg_misa[0], 30'h36000000 };
  assign read_mstatus_lo = { 14'h0018, reg_mstatus_mpie, 3'h0, reg_mstatus_mie, 3'h0 };
  assign read_mstatus_lo_lo = { 1'h0, reg_mstatus_mpie, 3'h0, reg_mstatus_mie, 3'h0 };
  assign read_mtvec = { reg_mtvec[31:7], _notDebugTVec_T_1[6:2], 1'h0, reg_mtvec[0] };
  assign { reg_custom_0[31:4], reg_custom_0[2:0] } = 31'h00000000;
  assign reg_mcountinhibit[1] = 1'h0;
  assign { reg_mie[31:12], reg_mie[10:8], reg_mie[6:4], reg_mie[2:0] } = 29'h00000000;
  assign { reg_misa[31:13], reg_misa[11:3], reg_misa[1] } = 29'h08100040;
  assign reg_mstatus_spp = 1'h0;
  assign tvec[1:0] = 2'h0;
  assign value = { large_, small_ };
  assign value_1 = { large_1, small_1 };
  assign wdata = _T_2000[31:0];
  assign whichInterrupt = io_interrupt_cause[3:0];
  assign x79 = reg_mcountinhibit[2];
  assign x86 = _GEN_35[0];
endmodule
module IBuf(clock, reset, io_imem_ready, io_imem_valid, io_imem_bits_pc, io_imem_bits_data, io_imem_bits_xcpt_ae_inst, io_imem_bits_replay, io_kill, io_pc, io_inst_0_ready, io_inst_0_valid, io_inst_0_bits_xcpt0_ae_inst, io_inst_0_bits_xcpt1_pf_inst, io_inst_0_bits_xcpt1_gf_inst, io_inst_0_bits_xcpt1_ae_inst, io_inst_0_bits_replay, io_inst_0_bits_rvc, io_inst_0_bits_inst_bits, io_inst_0_bits_inst_rd, io_inst_0_bits_inst_rs1
, io_inst_0_bits_inst_rs2, io_inst_0_bits_raw);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire [190:0] _GEN_1;
  wire [1:0] _GEN_58;
  wire [1:0] _GEN_59;
  wire [31:0] _GEN_67;
  wire [1:0] _bufMask_T;
  wire [5:0] _buf_data_T;
  wire [31:0] _buf_pc_T_1;
  wire [2:0] _buf_pc_T_2;
  wire [31:0] _buf_pc_T_4;
  wire [31:0] _buf_pc_T_5;
  wire [31:0] _buf_pc_T_6;
  wire [1:0] _full_insn_T_2;
  wire [63:0] _icData_T_2;
  wire [5:0] _icData_T_3;
  wire [190:0] _icData_T_4;
  wire [4:0] _icMask_T_1;
  wire [62:0] _icMask_T_2;
  wire [1:0] _icShiftAmt_T_1;
  wire [1:0] _ic_replay_T;
  wire [1:0] _ic_replay_T_1;
  wire [31:0] _inst_T;
  wire [31:0] _inst_T_1;
  wire [31:0] _inst_T_2;
  wire [2:0] _io_inst_0_bits_xcpt1_T_4;
  wire [2:0] _io_inst_0_bits_xcpt1_T_5;
  wire [1:0] _nReady_T_4;
  wire [1:0] _replay_T_5;
  wire [3:0] _valid_T_2;
  wire [1:0] bufMask;
  wire [31:0] buf__data;
  wire [31:0] buf__pc;
  wire buf__replay;
  wire buf__xcpt_ae_inst;
  wire [63:0] buf_data_data;
  wire [1:0] buf_replay;
  input clock;
  wire clock;
  wire [31:0] exp_io_in;
  wire [31:0] exp_io_out_bits;
  wire [4:0] exp_io_out_rd;
  wire [4:0] exp_io_out_rs1;
  wire [4:0] exp_io_out_rs2;
  wire exp_io_rvc;
  wire [31:0] icData;
  wire [127:0] icData_data;
  wire [31:0] icMask;
  wire [1:0] icShiftAmt;
  input [31:0] io_imem_bits_data;
  wire [31:0] io_imem_bits_data;
  input [31:0] io_imem_bits_pc;
  wire [31:0] io_imem_bits_pc;
  input io_imem_bits_replay;
  wire io_imem_bits_replay;
  input io_imem_bits_xcpt_ae_inst;
  wire io_imem_bits_xcpt_ae_inst;
  output io_imem_ready;
  wire io_imem_ready;
  input io_imem_valid;
  wire io_imem_valid;
  output [31:0] io_inst_0_bits_inst_bits;
  wire [31:0] io_inst_0_bits_inst_bits;
  output [4:0] io_inst_0_bits_inst_rd;
  wire [4:0] io_inst_0_bits_inst_rd;
  output [4:0] io_inst_0_bits_inst_rs1;
  wire [4:0] io_inst_0_bits_inst_rs1;
  output [4:0] io_inst_0_bits_inst_rs2;
  wire [4:0] io_inst_0_bits_inst_rs2;
  output [31:0] io_inst_0_bits_raw;
  wire [31:0] io_inst_0_bits_raw;
  output io_inst_0_bits_replay;
  wire io_inst_0_bits_replay;
  output io_inst_0_bits_rvc;
  wire io_inst_0_bits_rvc;
  output io_inst_0_bits_xcpt0_ae_inst;
  wire io_inst_0_bits_xcpt0_ae_inst;
  output io_inst_0_bits_xcpt1_ae_inst;
  wire io_inst_0_bits_xcpt1_ae_inst;
  output io_inst_0_bits_xcpt1_gf_inst;
  wire io_inst_0_bits_xcpt1_gf_inst;
  output io_inst_0_bits_xcpt1_pf_inst;
  wire io_inst_0_bits_xcpt1_pf_inst;
  input io_inst_0_ready;
  wire io_inst_0_ready;
  output io_inst_0_valid;
  wire io_inst_0_valid;
  input io_kill;
  wire io_kill;
  output [31:0] io_pc;
  wire [31:0] io_pc;
  wire nBufValid;
  wire [1:0] nIC;
  wire [1:0] nICReady;
  wire pcWordBits;
  input reset;
  wire reset;
  wire [1:0] shamt;
  wire [1:0] valid;
  wire xcpt_1_ae_inst;
  INV_X1 _235_ (
    .A(nBufValid),
    .ZN(_051_)
  );
  INV_X1 _236_ (
    .A(io_imem_bits_pc[1]),
    .ZN(_052_)
  );
  INV_X1 _237_ (
    .A(exp_io_rvc),
    .ZN(_053_)
  );
  INV_X1 _238_ (
    .A(_bufMask_T[0]),
    .ZN(_054_)
  );
  AND2_X1 _239_ (
    .A1(_051_),
    .A2(io_imem_bits_pc[1]),
    .ZN(_055_)
  );
  OR2_X1 _240_ (
    .A1(nBufValid),
    .A2(_052_),
    .ZN(_056_)
  );
  AND2_X1 _241_ (
    .A1(io_imem_valid),
    .A2(_056_),
    .ZN(_057_)
  );
  AND2_X1 _242_ (
    .A1(nBufValid),
    .A2(buf__replay),
    .ZN(_058_)
  );
  OR2_X1 _243_ (
    .A1(exp_io_rvc),
    .A2(_058_),
    .ZN(_059_)
  );
  OR2_X1 _244_ (
    .A1(_057_),
    .A2(_059_),
    .ZN(_060_)
  );
  OR2_X1 _245_ (
    .A1(_bufMask_T[0]),
    .A2(_060_),
    .ZN(_061_)
  );
  AND2_X1 _246_ (
    .A1(_053_),
    .A2(_bufMask_T[0]),
    .ZN(_062_)
  );
  OR2_X1 _247_ (
    .A1(exp_io_rvc),
    .A2(_054_),
    .ZN(_063_)
  );
  MUX2_X1 _248_ (
    .A(_bufMask_T[0]),
    .B(_063_),
    .S(_060_),
    .Z(_064_)
  );
  MUX2_X1 _249_ (
    .A(_054_),
    .B(_062_),
    .S(_060_),
    .Z(_065_)
  );
  XOR2_X1 _250_ (
    .A(_053_),
    .B(_bufMask_T[0]),
    .Z(_066_)
  );
  XOR2_X1 _251_ (
    .A(exp_io_rvc),
    .B(_bufMask_T[0]),
    .Z(_067_)
  );
  OR2_X1 _252_ (
    .A1(io_imem_bits_pc[1]),
    .A2(_066_),
    .ZN(_068_)
  );
  OR2_X1 _253_ (
    .A1(_065_),
    .A2(_068_),
    .ZN(_069_)
  );
  AND2_X1 _254_ (
    .A1(io_inst_0_ready),
    .A2(_061_),
    .ZN(_070_)
  );
  INV_X1 _255_ (
    .A(_070_),
    .ZN(_071_)
  );
  AND2_X1 _256_ (
    .A1(_069_),
    .A2(_070_),
    .ZN(io_imem_ready)
  );
  OR2_X1 _257_ (
    .A1(_052_),
    .A2(_067_),
    .ZN(_072_)
  );
  AND2_X1 _258_ (
    .A1(io_imem_valid),
    .A2(_072_),
    .ZN(_073_)
  );
  AND2_X1 _259_ (
    .A1(_064_),
    .A2(_073_),
    .ZN(_074_)
  );
  AND2_X1 _260_ (
    .A1(io_imem_ready),
    .A2(_074_),
    .ZN(_075_)
  );
  MUX2_X1 _261_ (
    .A(buf__replay),
    .B(io_imem_bits_replay),
    .S(_075_),
    .Z(_000_)
  );
  MUX2_X1 _262_ (
    .A(_068_),
    .B(_072_),
    .S(_065_),
    .Z(_076_)
  );
  AND2_X1 _263_ (
    .A1(io_imem_bits_data[16]),
    .A2(_076_),
    .ZN(_077_)
  );
  MUX2_X1 _264_ (
    .A(buf__data[0]),
    .B(_077_),
    .S(_075_),
    .Z(_001_)
  );
  AND2_X1 _265_ (
    .A1(io_imem_bits_data[17]),
    .A2(_076_),
    .ZN(_078_)
  );
  MUX2_X1 _266_ (
    .A(buf__data[1]),
    .B(_078_),
    .S(_075_),
    .Z(_002_)
  );
  AND2_X1 _267_ (
    .A1(io_imem_bits_data[18]),
    .A2(_076_),
    .ZN(_079_)
  );
  MUX2_X1 _268_ (
    .A(buf__data[2]),
    .B(_079_),
    .S(_075_),
    .Z(_003_)
  );
  AND2_X1 _269_ (
    .A1(io_imem_bits_data[19]),
    .A2(_076_),
    .ZN(_080_)
  );
  MUX2_X1 _270_ (
    .A(buf__data[3]),
    .B(_080_),
    .S(_075_),
    .Z(_004_)
  );
  AND2_X1 _271_ (
    .A1(io_imem_bits_data[20]),
    .A2(_076_),
    .ZN(_081_)
  );
  MUX2_X1 _272_ (
    .A(buf__data[4]),
    .B(_081_),
    .S(_075_),
    .Z(_005_)
  );
  AND2_X1 _273_ (
    .A1(io_imem_bits_data[21]),
    .A2(_076_),
    .ZN(_082_)
  );
  MUX2_X1 _274_ (
    .A(buf__data[5]),
    .B(_082_),
    .S(_075_),
    .Z(_006_)
  );
  AND2_X1 _275_ (
    .A1(io_imem_bits_data[22]),
    .A2(_076_),
    .ZN(_083_)
  );
  MUX2_X1 _276_ (
    .A(buf__data[6]),
    .B(_083_),
    .S(_075_),
    .Z(_007_)
  );
  AND2_X1 _277_ (
    .A1(io_imem_bits_data[23]),
    .A2(_076_),
    .ZN(_084_)
  );
  MUX2_X1 _278_ (
    .A(buf__data[7]),
    .B(_084_),
    .S(_075_),
    .Z(_008_)
  );
  AND2_X1 _279_ (
    .A1(io_imem_bits_data[24]),
    .A2(_076_),
    .ZN(_085_)
  );
  MUX2_X1 _280_ (
    .A(buf__data[8]),
    .B(_085_),
    .S(_075_),
    .Z(_009_)
  );
  AND2_X1 _281_ (
    .A1(io_imem_bits_data[25]),
    .A2(_076_),
    .ZN(_086_)
  );
  MUX2_X1 _282_ (
    .A(buf__data[9]),
    .B(_086_),
    .S(_075_),
    .Z(_010_)
  );
  AND2_X1 _283_ (
    .A1(io_imem_bits_data[26]),
    .A2(_076_),
    .ZN(_087_)
  );
  MUX2_X1 _284_ (
    .A(buf__data[10]),
    .B(_087_),
    .S(_075_),
    .Z(_011_)
  );
  AND2_X1 _285_ (
    .A1(io_imem_bits_data[27]),
    .A2(_076_),
    .ZN(_088_)
  );
  MUX2_X1 _286_ (
    .A(buf__data[11]),
    .B(_088_),
    .S(_075_),
    .Z(_012_)
  );
  AND2_X1 _287_ (
    .A1(io_imem_bits_data[28]),
    .A2(_076_),
    .ZN(_089_)
  );
  MUX2_X1 _288_ (
    .A(buf__data[12]),
    .B(_089_),
    .S(_075_),
    .Z(_013_)
  );
  AND2_X1 _289_ (
    .A1(io_imem_bits_data[29]),
    .A2(_076_),
    .ZN(_090_)
  );
  MUX2_X1 _290_ (
    .A(buf__data[13]),
    .B(_090_),
    .S(_075_),
    .Z(_014_)
  );
  AND2_X1 _291_ (
    .A1(io_imem_bits_data[30]),
    .A2(_076_),
    .ZN(_091_)
  );
  MUX2_X1 _292_ (
    .A(buf__data[14]),
    .B(_091_),
    .S(_075_),
    .Z(_015_)
  );
  AND2_X1 _293_ (
    .A1(io_imem_bits_data[31]),
    .A2(_076_),
    .ZN(_092_)
  );
  MUX2_X1 _294_ (
    .A(buf__data[15]),
    .B(_092_),
    .S(_075_),
    .Z(_016_)
  );
  MUX2_X1 _295_ (
    .A(buf__pc[0]),
    .B(io_imem_bits_pc[0]),
    .S(_075_),
    .Z(_017_)
  );
  OR2_X1 _296_ (
    .A1(buf__pc[1]),
    .A2(_075_),
    .ZN(_018_)
  );
  MUX2_X1 _297_ (
    .A(buf__pc[2]),
    .B(io_imem_bits_pc[2]),
    .S(_075_),
    .Z(_019_)
  );
  MUX2_X1 _298_ (
    .A(buf__pc[3]),
    .B(io_imem_bits_pc[3]),
    .S(_075_),
    .Z(_020_)
  );
  MUX2_X1 _299_ (
    .A(buf__pc[4]),
    .B(io_imem_bits_pc[4]),
    .S(_075_),
    .Z(_021_)
  );
  MUX2_X1 _300_ (
    .A(buf__pc[5]),
    .B(io_imem_bits_pc[5]),
    .S(_075_),
    .Z(_022_)
  );
  MUX2_X1 _301_ (
    .A(buf__pc[6]),
    .B(io_imem_bits_pc[6]),
    .S(_075_),
    .Z(_023_)
  );
  MUX2_X1 _302_ (
    .A(buf__pc[7]),
    .B(io_imem_bits_pc[7]),
    .S(_075_),
    .Z(_024_)
  );
  MUX2_X1 _303_ (
    .A(buf__pc[8]),
    .B(io_imem_bits_pc[8]),
    .S(_075_),
    .Z(_025_)
  );
  MUX2_X1 _304_ (
    .A(buf__pc[9]),
    .B(io_imem_bits_pc[9]),
    .S(_075_),
    .Z(_026_)
  );
  MUX2_X1 _305_ (
    .A(buf__pc[10]),
    .B(io_imem_bits_pc[10]),
    .S(_075_),
    .Z(_027_)
  );
  MUX2_X1 _306_ (
    .A(buf__pc[11]),
    .B(io_imem_bits_pc[11]),
    .S(_075_),
    .Z(_028_)
  );
  MUX2_X1 _307_ (
    .A(buf__pc[12]),
    .B(io_imem_bits_pc[12]),
    .S(_075_),
    .Z(_029_)
  );
  MUX2_X1 _308_ (
    .A(buf__pc[13]),
    .B(io_imem_bits_pc[13]),
    .S(_075_),
    .Z(_030_)
  );
  MUX2_X1 _309_ (
    .A(buf__pc[14]),
    .B(io_imem_bits_pc[14]),
    .S(_075_),
    .Z(_031_)
  );
  MUX2_X1 _310_ (
    .A(buf__pc[15]),
    .B(io_imem_bits_pc[15]),
    .S(_075_),
    .Z(_032_)
  );
  MUX2_X1 _311_ (
    .A(buf__pc[16]),
    .B(io_imem_bits_pc[16]),
    .S(_075_),
    .Z(_033_)
  );
  MUX2_X1 _312_ (
    .A(buf__pc[17]),
    .B(io_imem_bits_pc[17]),
    .S(_075_),
    .Z(_034_)
  );
  MUX2_X1 _313_ (
    .A(buf__pc[18]),
    .B(io_imem_bits_pc[18]),
    .S(_075_),
    .Z(_035_)
  );
  MUX2_X1 _314_ (
    .A(buf__pc[19]),
    .B(io_imem_bits_pc[19]),
    .S(_075_),
    .Z(_036_)
  );
  MUX2_X1 _315_ (
    .A(buf__pc[20]),
    .B(io_imem_bits_pc[20]),
    .S(_075_),
    .Z(_037_)
  );
  MUX2_X1 _316_ (
    .A(buf__pc[21]),
    .B(io_imem_bits_pc[21]),
    .S(_075_),
    .Z(_038_)
  );
  MUX2_X1 _317_ (
    .A(buf__pc[22]),
    .B(io_imem_bits_pc[22]),
    .S(_075_),
    .Z(_039_)
  );
  MUX2_X1 _318_ (
    .A(buf__pc[23]),
    .B(io_imem_bits_pc[23]),
    .S(_075_),
    .Z(_040_)
  );
  MUX2_X1 _319_ (
    .A(buf__pc[24]),
    .B(io_imem_bits_pc[24]),
    .S(_075_),
    .Z(_041_)
  );
  MUX2_X1 _320_ (
    .A(buf__pc[25]),
    .B(io_imem_bits_pc[25]),
    .S(_075_),
    .Z(_042_)
  );
  MUX2_X1 _321_ (
    .A(buf__pc[26]),
    .B(io_imem_bits_pc[26]),
    .S(_075_),
    .Z(_043_)
  );
  MUX2_X1 _322_ (
    .A(buf__pc[27]),
    .B(io_imem_bits_pc[27]),
    .S(_075_),
    .Z(_044_)
  );
  MUX2_X1 _323_ (
    .A(buf__pc[28]),
    .B(io_imem_bits_pc[28]),
    .S(_075_),
    .Z(_045_)
  );
  MUX2_X1 _324_ (
    .A(buf__pc[29]),
    .B(io_imem_bits_pc[29]),
    .S(_075_),
    .Z(_046_)
  );
  MUX2_X1 _325_ (
    .A(buf__pc[30]),
    .B(io_imem_bits_pc[30]),
    .S(_075_),
    .Z(_047_)
  );
  MUX2_X1 _326_ (
    .A(buf__pc[31]),
    .B(io_imem_bits_pc[31]),
    .S(_075_),
    .Z(_048_)
  );
  AND2_X1 _327_ (
    .A1(io_inst_0_ready),
    .A2(exp_io_rvc),
    .ZN(_093_)
  );
  XOR2_X1 _328_ (
    .A(nBufValid),
    .B(_093_),
    .Z(_094_)
  );
  AND2_X1 _329_ (
    .A1(_071_),
    .A2(_094_),
    .ZN(_095_)
  );
  OR2_X1 _330_ (
    .A1(_075_),
    .A2(_095_),
    .ZN(_096_)
  );
  OR2_X1 _331_ (
    .A1(reset),
    .A2(io_kill),
    .ZN(_097_)
  );
  INV_X1 _332_ (
    .A(_097_),
    .ZN(_098_)
  );
  AND2_X1 _333_ (
    .A1(_096_),
    .A2(_098_),
    .ZN(_049_)
  );
  MUX2_X1 _334_ (
    .A(buf__xcpt_ae_inst),
    .B(io_imem_bits_xcpt_ae_inst),
    .S(_075_),
    .Z(_050_)
  );
  AND2_X1 _335_ (
    .A1(io_imem_bits_xcpt_ae_inst),
    .A2(_053_),
    .ZN(io_inst_0_bits_xcpt1_ae_inst)
  );
  MUX2_X1 _336_ (
    .A(io_imem_bits_pc[0]),
    .B(buf__pc[0]),
    .S(nBufValid),
    .Z(io_pc[0])
  );
  MUX2_X1 _337_ (
    .A(io_imem_bits_pc[1]),
    .B(buf__pc[1]),
    .S(nBufValid),
    .Z(io_pc[1])
  );
  MUX2_X1 _338_ (
    .A(io_imem_bits_pc[2]),
    .B(buf__pc[2]),
    .S(nBufValid),
    .Z(io_pc[2])
  );
  MUX2_X1 _339_ (
    .A(io_imem_bits_pc[3]),
    .B(buf__pc[3]),
    .S(nBufValid),
    .Z(io_pc[3])
  );
  MUX2_X1 _340_ (
    .A(io_imem_bits_pc[4]),
    .B(buf__pc[4]),
    .S(nBufValid),
    .Z(io_pc[4])
  );
  MUX2_X1 _341_ (
    .A(io_imem_bits_pc[5]),
    .B(buf__pc[5]),
    .S(nBufValid),
    .Z(io_pc[5])
  );
  MUX2_X1 _342_ (
    .A(io_imem_bits_pc[6]),
    .B(buf__pc[6]),
    .S(nBufValid),
    .Z(io_pc[6])
  );
  MUX2_X1 _343_ (
    .A(io_imem_bits_pc[7]),
    .B(buf__pc[7]),
    .S(nBufValid),
    .Z(io_pc[7])
  );
  MUX2_X1 _344_ (
    .A(io_imem_bits_pc[8]),
    .B(buf__pc[8]),
    .S(nBufValid),
    .Z(io_pc[8])
  );
  MUX2_X1 _345_ (
    .A(io_imem_bits_pc[9]),
    .B(buf__pc[9]),
    .S(nBufValid),
    .Z(io_pc[9])
  );
  MUX2_X1 _346_ (
    .A(io_imem_bits_pc[10]),
    .B(buf__pc[10]),
    .S(nBufValid),
    .Z(io_pc[10])
  );
  MUX2_X1 _347_ (
    .A(io_imem_bits_pc[11]),
    .B(buf__pc[11]),
    .S(nBufValid),
    .Z(io_pc[11])
  );
  MUX2_X1 _348_ (
    .A(io_imem_bits_pc[12]),
    .B(buf__pc[12]),
    .S(nBufValid),
    .Z(io_pc[12])
  );
  MUX2_X1 _349_ (
    .A(io_imem_bits_pc[13]),
    .B(buf__pc[13]),
    .S(nBufValid),
    .Z(io_pc[13])
  );
  MUX2_X1 _350_ (
    .A(io_imem_bits_pc[14]),
    .B(buf__pc[14]),
    .S(nBufValid),
    .Z(io_pc[14])
  );
  MUX2_X1 _351_ (
    .A(io_imem_bits_pc[15]),
    .B(buf__pc[15]),
    .S(nBufValid),
    .Z(io_pc[15])
  );
  MUX2_X1 _352_ (
    .A(io_imem_bits_pc[16]),
    .B(buf__pc[16]),
    .S(nBufValid),
    .Z(io_pc[16])
  );
  MUX2_X1 _353_ (
    .A(io_imem_bits_pc[17]),
    .B(buf__pc[17]),
    .S(nBufValid),
    .Z(io_pc[17])
  );
  MUX2_X1 _354_ (
    .A(io_imem_bits_pc[18]),
    .B(buf__pc[18]),
    .S(nBufValid),
    .Z(io_pc[18])
  );
  MUX2_X1 _355_ (
    .A(io_imem_bits_pc[19]),
    .B(buf__pc[19]),
    .S(nBufValid),
    .Z(io_pc[19])
  );
  MUX2_X1 _356_ (
    .A(io_imem_bits_pc[20]),
    .B(buf__pc[20]),
    .S(nBufValid),
    .Z(io_pc[20])
  );
  MUX2_X1 _357_ (
    .A(io_imem_bits_pc[21]),
    .B(buf__pc[21]),
    .S(nBufValid),
    .Z(io_pc[21])
  );
  MUX2_X1 _358_ (
    .A(io_imem_bits_pc[22]),
    .B(buf__pc[22]),
    .S(nBufValid),
    .Z(io_pc[22])
  );
  MUX2_X1 _359_ (
    .A(io_imem_bits_pc[23]),
    .B(buf__pc[23]),
    .S(nBufValid),
    .Z(io_pc[23])
  );
  MUX2_X1 _360_ (
    .A(io_imem_bits_pc[24]),
    .B(buf__pc[24]),
    .S(nBufValid),
    .Z(io_pc[24])
  );
  MUX2_X1 _361_ (
    .A(io_imem_bits_pc[25]),
    .B(buf__pc[25]),
    .S(nBufValid),
    .Z(io_pc[25])
  );
  MUX2_X1 _362_ (
    .A(io_imem_bits_pc[26]),
    .B(buf__pc[26]),
    .S(nBufValid),
    .Z(io_pc[26])
  );
  MUX2_X1 _363_ (
    .A(io_imem_bits_pc[27]),
    .B(buf__pc[27]),
    .S(nBufValid),
    .Z(io_pc[27])
  );
  MUX2_X1 _364_ (
    .A(io_imem_bits_pc[28]),
    .B(buf__pc[28]),
    .S(nBufValid),
    .Z(io_pc[28])
  );
  MUX2_X1 _365_ (
    .A(io_imem_bits_pc[29]),
    .B(buf__pc[29]),
    .S(nBufValid),
    .Z(io_pc[29])
  );
  MUX2_X1 _366_ (
    .A(io_imem_bits_pc[30]),
    .B(buf__pc[30]),
    .S(nBufValid),
    .Z(io_pc[30])
  );
  MUX2_X1 _367_ (
    .A(io_imem_bits_pc[31]),
    .B(buf__pc[31]),
    .S(nBufValid),
    .Z(io_pc[31])
  );
  MUX2_X1 _368_ (
    .A(io_imem_bits_xcpt_ae_inst),
    .B(buf__xcpt_ae_inst),
    .S(nBufValid),
    .Z(io_inst_0_bits_xcpt0_ae_inst)
  );
  OR2_X1 _369_ (
    .A1(nBufValid),
    .A2(io_imem_valid),
    .ZN(_099_)
  );
  AND2_X1 _370_ (
    .A1(_060_),
    .A2(_099_),
    .ZN(io_inst_0_valid)
  );
  AND2_X1 _371_ (
    .A1(_bufMask_T[0]),
    .A2(_099_),
    .ZN(_100_)
  );
  AND2_X1 _372_ (
    .A1(_053_),
    .A2(_057_),
    .ZN(_101_)
  );
  OR2_X1 _373_ (
    .A1(_100_),
    .A2(_101_),
    .ZN(_102_)
  );
  AND2_X1 _374_ (
    .A1(io_imem_bits_replay),
    .A2(_102_),
    .ZN(_103_)
  );
  OR2_X1 _375_ (
    .A1(_058_),
    .A2(_103_),
    .ZN(io_inst_0_bits_replay)
  );
  AND2_X1 _376_ (
    .A1(nBufValid),
    .A2(buf__data[0]),
    .ZN(_104_)
  );
  OR2_X1 _377_ (
    .A1(io_imem_bits_data[0]),
    .A2(_055_),
    .ZN(_105_)
  );
  OR2_X1 _378_ (
    .A1(io_imem_bits_data[16]),
    .A2(_056_),
    .ZN(_106_)
  );
  AND2_X1 _379_ (
    .A1(_bufMask_T[0]),
    .A2(_106_),
    .ZN(_107_)
  );
  AND2_X1 _380_ (
    .A1(_105_),
    .A2(_107_),
    .ZN(_108_)
  );
  OR2_X1 _381_ (
    .A1(_104_),
    .A2(_108_),
    .ZN(exp_io_in[0])
  );
  AND2_X1 _382_ (
    .A1(nBufValid),
    .A2(buf__data[1]),
    .ZN(_109_)
  );
  OR2_X1 _383_ (
    .A1(io_imem_bits_data[1]),
    .A2(_055_),
    .ZN(_110_)
  );
  OR2_X1 _384_ (
    .A1(io_imem_bits_data[17]),
    .A2(_056_),
    .ZN(_111_)
  );
  AND2_X1 _385_ (
    .A1(_bufMask_T[0]),
    .A2(_111_),
    .ZN(_112_)
  );
  AND2_X1 _386_ (
    .A1(_110_),
    .A2(_112_),
    .ZN(_113_)
  );
  OR2_X1 _387_ (
    .A1(_109_),
    .A2(_113_),
    .ZN(exp_io_in[1])
  );
  AND2_X1 _388_ (
    .A1(nBufValid),
    .A2(buf__data[2]),
    .ZN(_114_)
  );
  OR2_X1 _389_ (
    .A1(io_imem_bits_data[2]),
    .A2(_055_),
    .ZN(_115_)
  );
  OR2_X1 _390_ (
    .A1(io_imem_bits_data[18]),
    .A2(_056_),
    .ZN(_116_)
  );
  AND2_X1 _391_ (
    .A1(_bufMask_T[0]),
    .A2(_116_),
    .ZN(_117_)
  );
  AND2_X1 _392_ (
    .A1(_115_),
    .A2(_117_),
    .ZN(_118_)
  );
  OR2_X1 _393_ (
    .A1(_114_),
    .A2(_118_),
    .ZN(exp_io_in[2])
  );
  AND2_X1 _394_ (
    .A1(nBufValid),
    .A2(buf__data[3]),
    .ZN(_119_)
  );
  OR2_X1 _395_ (
    .A1(io_imem_bits_data[19]),
    .A2(_056_),
    .ZN(_120_)
  );
  OR2_X1 _396_ (
    .A1(io_imem_bits_data[3]),
    .A2(_055_),
    .ZN(_121_)
  );
  AND2_X1 _397_ (
    .A1(_bufMask_T[0]),
    .A2(_121_),
    .ZN(_122_)
  );
  AND2_X1 _398_ (
    .A1(_120_),
    .A2(_122_),
    .ZN(_123_)
  );
  OR2_X1 _399_ (
    .A1(_119_),
    .A2(_123_),
    .ZN(exp_io_in[3])
  );
  AND2_X1 _400_ (
    .A1(nBufValid),
    .A2(buf__data[4]),
    .ZN(_124_)
  );
  OR2_X1 _401_ (
    .A1(io_imem_bits_data[4]),
    .A2(_055_),
    .ZN(_125_)
  );
  OR2_X1 _402_ (
    .A1(io_imem_bits_data[20]),
    .A2(_056_),
    .ZN(_126_)
  );
  AND2_X1 _403_ (
    .A1(_bufMask_T[0]),
    .A2(_126_),
    .ZN(_127_)
  );
  AND2_X1 _404_ (
    .A1(_125_),
    .A2(_127_),
    .ZN(_128_)
  );
  OR2_X1 _405_ (
    .A1(_124_),
    .A2(_128_),
    .ZN(exp_io_in[4])
  );
  AND2_X1 _406_ (
    .A1(nBufValid),
    .A2(buf__data[5]),
    .ZN(_129_)
  );
  OR2_X1 _407_ (
    .A1(io_imem_bits_data[21]),
    .A2(_056_),
    .ZN(_130_)
  );
  OR2_X1 _408_ (
    .A1(io_imem_bits_data[5]),
    .A2(_055_),
    .ZN(_131_)
  );
  AND2_X1 _409_ (
    .A1(_bufMask_T[0]),
    .A2(_131_),
    .ZN(_132_)
  );
  AND2_X1 _410_ (
    .A1(_130_),
    .A2(_132_),
    .ZN(_133_)
  );
  OR2_X1 _411_ (
    .A1(_129_),
    .A2(_133_),
    .ZN(exp_io_in[5])
  );
  AND2_X1 _412_ (
    .A1(nBufValid),
    .A2(buf__data[6]),
    .ZN(_134_)
  );
  OR2_X1 _413_ (
    .A1(io_imem_bits_data[6]),
    .A2(_055_),
    .ZN(_135_)
  );
  OR2_X1 _414_ (
    .A1(io_imem_bits_data[22]),
    .A2(_056_),
    .ZN(_136_)
  );
  AND2_X1 _415_ (
    .A1(_bufMask_T[0]),
    .A2(_136_),
    .ZN(_137_)
  );
  AND2_X1 _416_ (
    .A1(_135_),
    .A2(_137_),
    .ZN(_138_)
  );
  OR2_X1 _417_ (
    .A1(_134_),
    .A2(_138_),
    .ZN(exp_io_in[6])
  );
  AND2_X1 _418_ (
    .A1(nBufValid),
    .A2(buf__data[7]),
    .ZN(_139_)
  );
  OR2_X1 _419_ (
    .A1(io_imem_bits_data[7]),
    .A2(_055_),
    .ZN(_140_)
  );
  OR2_X1 _420_ (
    .A1(io_imem_bits_data[23]),
    .A2(_056_),
    .ZN(_141_)
  );
  AND2_X1 _421_ (
    .A1(_bufMask_T[0]),
    .A2(_141_),
    .ZN(_142_)
  );
  AND2_X1 _422_ (
    .A1(_140_),
    .A2(_142_),
    .ZN(_143_)
  );
  OR2_X1 _423_ (
    .A1(_139_),
    .A2(_143_),
    .ZN(exp_io_in[7])
  );
  AND2_X1 _424_ (
    .A1(nBufValid),
    .A2(buf__data[8]),
    .ZN(_144_)
  );
  OR2_X1 _425_ (
    .A1(io_imem_bits_data[8]),
    .A2(_055_),
    .ZN(_145_)
  );
  OR2_X1 _426_ (
    .A1(io_imem_bits_data[24]),
    .A2(_056_),
    .ZN(_146_)
  );
  AND2_X1 _427_ (
    .A1(_bufMask_T[0]),
    .A2(_146_),
    .ZN(_147_)
  );
  AND2_X1 _428_ (
    .A1(_145_),
    .A2(_147_),
    .ZN(_148_)
  );
  OR2_X1 _429_ (
    .A1(_144_),
    .A2(_148_),
    .ZN(exp_io_in[8])
  );
  AND2_X1 _430_ (
    .A1(nBufValid),
    .A2(buf__data[9]),
    .ZN(_149_)
  );
  OR2_X1 _431_ (
    .A1(io_imem_bits_data[9]),
    .A2(_055_),
    .ZN(_150_)
  );
  OR2_X1 _432_ (
    .A1(io_imem_bits_data[25]),
    .A2(_056_),
    .ZN(_151_)
  );
  AND2_X1 _433_ (
    .A1(_bufMask_T[0]),
    .A2(_151_),
    .ZN(_152_)
  );
  AND2_X1 _434_ (
    .A1(_150_),
    .A2(_152_),
    .ZN(_153_)
  );
  OR2_X1 _435_ (
    .A1(_149_),
    .A2(_153_),
    .ZN(exp_io_in[9])
  );
  AND2_X1 _436_ (
    .A1(nBufValid),
    .A2(buf__data[10]),
    .ZN(_154_)
  );
  OR2_X1 _437_ (
    .A1(io_imem_bits_data[10]),
    .A2(_055_),
    .ZN(_155_)
  );
  OR2_X1 _438_ (
    .A1(io_imem_bits_data[26]),
    .A2(_056_),
    .ZN(_156_)
  );
  AND2_X1 _439_ (
    .A1(_bufMask_T[0]),
    .A2(_156_),
    .ZN(_157_)
  );
  AND2_X1 _440_ (
    .A1(_155_),
    .A2(_157_),
    .ZN(_158_)
  );
  OR2_X1 _441_ (
    .A1(_154_),
    .A2(_158_),
    .ZN(exp_io_in[10])
  );
  AND2_X1 _442_ (
    .A1(nBufValid),
    .A2(buf__data[11]),
    .ZN(_159_)
  );
  OR2_X1 _443_ (
    .A1(io_imem_bits_data[11]),
    .A2(_055_),
    .ZN(_160_)
  );
  OR2_X1 _444_ (
    .A1(io_imem_bits_data[27]),
    .A2(_056_),
    .ZN(_161_)
  );
  AND2_X1 _445_ (
    .A1(_bufMask_T[0]),
    .A2(_161_),
    .ZN(_162_)
  );
  AND2_X1 _446_ (
    .A1(_160_),
    .A2(_162_),
    .ZN(_163_)
  );
  OR2_X1 _447_ (
    .A1(_159_),
    .A2(_163_),
    .ZN(exp_io_in[11])
  );
  AND2_X1 _448_ (
    .A1(nBufValid),
    .A2(buf__data[12]),
    .ZN(_164_)
  );
  OR2_X1 _449_ (
    .A1(io_imem_bits_data[12]),
    .A2(_055_),
    .ZN(_165_)
  );
  OR2_X1 _450_ (
    .A1(io_imem_bits_data[28]),
    .A2(_056_),
    .ZN(_166_)
  );
  AND2_X1 _451_ (
    .A1(_bufMask_T[0]),
    .A2(_166_),
    .ZN(_167_)
  );
  AND2_X1 _452_ (
    .A1(_165_),
    .A2(_167_),
    .ZN(_168_)
  );
  OR2_X1 _453_ (
    .A1(_164_),
    .A2(_168_),
    .ZN(exp_io_in[12])
  );
  AND2_X1 _454_ (
    .A1(nBufValid),
    .A2(buf__data[13]),
    .ZN(_169_)
  );
  OR2_X1 _455_ (
    .A1(io_imem_bits_data[29]),
    .A2(_056_),
    .ZN(_170_)
  );
  OR2_X1 _456_ (
    .A1(io_imem_bits_data[13]),
    .A2(_055_),
    .ZN(_171_)
  );
  AND2_X1 _457_ (
    .A1(_bufMask_T[0]),
    .A2(_171_),
    .ZN(_172_)
  );
  AND2_X1 _458_ (
    .A1(_170_),
    .A2(_172_),
    .ZN(_173_)
  );
  OR2_X1 _459_ (
    .A1(_169_),
    .A2(_173_),
    .ZN(exp_io_in[13])
  );
  AND2_X1 _460_ (
    .A1(nBufValid),
    .A2(buf__data[14]),
    .ZN(_174_)
  );
  OR2_X1 _461_ (
    .A1(io_imem_bits_data[14]),
    .A2(_055_),
    .ZN(_175_)
  );
  OR2_X1 _462_ (
    .A1(io_imem_bits_data[30]),
    .A2(_056_),
    .ZN(_176_)
  );
  AND2_X1 _463_ (
    .A1(_bufMask_T[0]),
    .A2(_176_),
    .ZN(_177_)
  );
  AND2_X1 _464_ (
    .A1(_175_),
    .A2(_177_),
    .ZN(_178_)
  );
  OR2_X1 _465_ (
    .A1(_174_),
    .A2(_178_),
    .ZN(exp_io_in[14])
  );
  AND2_X1 _466_ (
    .A1(nBufValid),
    .A2(buf__data[15]),
    .ZN(_179_)
  );
  OR2_X1 _467_ (
    .A1(io_imem_bits_data[15]),
    .A2(_055_),
    .ZN(_180_)
  );
  OR2_X1 _468_ (
    .A1(io_imem_bits_data[31]),
    .A2(_056_),
    .ZN(_181_)
  );
  AND2_X1 _469_ (
    .A1(_bufMask_T[0]),
    .A2(_181_),
    .ZN(_182_)
  );
  AND2_X1 _470_ (
    .A1(_180_),
    .A2(_182_),
    .ZN(_183_)
  );
  OR2_X1 _471_ (
    .A1(_179_),
    .A2(_183_),
    .ZN(exp_io_in[15])
  );
  OR2_X1 _472_ (
    .A1(_051_),
    .A2(io_imem_bits_pc[1]),
    .ZN(_184_)
  );
  MUX2_X1 _473_ (
    .A(io_imem_bits_data[0]),
    .B(io_imem_bits_data[16]),
    .S(_184_),
    .Z(_icData_T_4[80])
  );
  MUX2_X1 _474_ (
    .A(io_imem_bits_data[1]),
    .B(io_imem_bits_data[17]),
    .S(_184_),
    .Z(_icData_T_4[81])
  );
  MUX2_X1 _475_ (
    .A(io_imem_bits_data[2]),
    .B(io_imem_bits_data[18]),
    .S(_184_),
    .Z(_icData_T_4[82])
  );
  MUX2_X1 _476_ (
    .A(io_imem_bits_data[3]),
    .B(io_imem_bits_data[19]),
    .S(_184_),
    .Z(_icData_T_4[83])
  );
  MUX2_X1 _477_ (
    .A(io_imem_bits_data[4]),
    .B(io_imem_bits_data[20]),
    .S(_184_),
    .Z(_icData_T_4[84])
  );
  MUX2_X1 _478_ (
    .A(io_imem_bits_data[5]),
    .B(io_imem_bits_data[21]),
    .S(_184_),
    .Z(_icData_T_4[85])
  );
  MUX2_X1 _479_ (
    .A(io_imem_bits_data[6]),
    .B(io_imem_bits_data[22]),
    .S(_184_),
    .Z(_icData_T_4[86])
  );
  MUX2_X1 _480_ (
    .A(io_imem_bits_data[7]),
    .B(io_imem_bits_data[23]),
    .S(_184_),
    .Z(_icData_T_4[87])
  );
  MUX2_X1 _481_ (
    .A(io_imem_bits_data[8]),
    .B(io_imem_bits_data[24]),
    .S(_184_),
    .Z(_icData_T_4[88])
  );
  MUX2_X1 _482_ (
    .A(io_imem_bits_data[9]),
    .B(io_imem_bits_data[25]),
    .S(_184_),
    .Z(_icData_T_4[89])
  );
  MUX2_X1 _483_ (
    .A(io_imem_bits_data[10]),
    .B(io_imem_bits_data[26]),
    .S(_184_),
    .Z(_icData_T_4[90])
  );
  MUX2_X1 _484_ (
    .A(io_imem_bits_data[11]),
    .B(io_imem_bits_data[27]),
    .S(_184_),
    .Z(_icData_T_4[91])
  );
  MUX2_X1 _485_ (
    .A(io_imem_bits_data[12]),
    .B(io_imem_bits_data[28]),
    .S(_184_),
    .Z(_icData_T_4[92])
  );
  MUX2_X1 _486_ (
    .A(io_imem_bits_data[13]),
    .B(io_imem_bits_data[29]),
    .S(_184_),
    .Z(_icData_T_4[93])
  );
  MUX2_X1 _487_ (
    .A(io_imem_bits_data[14]),
    .B(io_imem_bits_data[30]),
    .S(_184_),
    .Z(_icData_T_4[94])
  );
  MUX2_X1 _488_ (
    .A(io_imem_bits_data[15]),
    .B(io_imem_bits_data[31]),
    .S(_184_),
    .Z(_icData_T_4[95])
  );
  DFF_X1 \buf__data[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_001_),
    .Q(buf__data[0]),
    .QN(_233_)
  );
  DFF_X1 \buf__data[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_011_),
    .Q(buf__data[10]),
    .QN(_223_)
  );
  DFF_X1 \buf__data[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_012_),
    .Q(buf__data[11]),
    .QN(_222_)
  );
  DFF_X1 \buf__data[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_013_),
    .Q(buf__data[12]),
    .QN(_221_)
  );
  DFF_X1 \buf__data[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_014_),
    .Q(buf__data[13]),
    .QN(_220_)
  );
  DFF_X1 \buf__data[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_015_),
    .Q(buf__data[14]),
    .QN(_219_)
  );
  DFF_X1 \buf__data[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_016_),
    .Q(buf__data[15]),
    .QN(_218_)
  );
  DFF_X1 \buf__data[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_002_),
    .Q(buf__data[1]),
    .QN(_232_)
  );
  DFF_X1 \buf__data[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_003_),
    .Q(buf__data[2]),
    .QN(_231_)
  );
  DFF_X1 \buf__data[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_004_),
    .Q(buf__data[3]),
    .QN(_230_)
  );
  DFF_X1 \buf__data[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_005_),
    .Q(buf__data[4]),
    .QN(_229_)
  );
  DFF_X1 \buf__data[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_006_),
    .Q(buf__data[5]),
    .QN(_228_)
  );
  DFF_X1 \buf__data[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_007_),
    .Q(buf__data[6]),
    .QN(_227_)
  );
  DFF_X1 \buf__data[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_008_),
    .Q(buf__data[7]),
    .QN(_226_)
  );
  DFF_X1 \buf__data[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_009_),
    .Q(buf__data[8]),
    .QN(_225_)
  );
  DFF_X1 \buf__data[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_010_),
    .Q(buf__data[9]),
    .QN(_224_)
  );
  DFF_X1 \buf__pc[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_017_),
    .Q(buf__pc[0]),
    .QN(_217_)
  );
  DFF_X1 \buf__pc[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_027_),
    .Q(buf__pc[10]),
    .QN(_207_)
  );
  DFF_X1 \buf__pc[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_028_),
    .Q(buf__pc[11]),
    .QN(_206_)
  );
  DFF_X1 \buf__pc[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_029_),
    .Q(buf__pc[12]),
    .QN(_205_)
  );
  DFF_X1 \buf__pc[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_030_),
    .Q(buf__pc[13]),
    .QN(_204_)
  );
  DFF_X1 \buf__pc[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_031_),
    .Q(buf__pc[14]),
    .QN(_203_)
  );
  DFF_X1 \buf__pc[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_032_),
    .Q(buf__pc[15]),
    .QN(_202_)
  );
  DFF_X1 \buf__pc[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_033_),
    .Q(buf__pc[16]),
    .QN(_201_)
  );
  DFF_X1 \buf__pc[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_034_),
    .Q(buf__pc[17]),
    .QN(_200_)
  );
  DFF_X1 \buf__pc[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_035_),
    .Q(buf__pc[18]),
    .QN(_199_)
  );
  DFF_X1 \buf__pc[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_036_),
    .Q(buf__pc[19]),
    .QN(_198_)
  );
  DFF_X1 \buf__pc[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_018_),
    .Q(buf__pc[1]),
    .QN(_216_)
  );
  DFF_X1 \buf__pc[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_037_),
    .Q(buf__pc[20]),
    .QN(_197_)
  );
  DFF_X1 \buf__pc[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_038_),
    .Q(buf__pc[21]),
    .QN(_196_)
  );
  DFF_X1 \buf__pc[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_039_),
    .Q(buf__pc[22]),
    .QN(_195_)
  );
  DFF_X1 \buf__pc[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_040_),
    .Q(buf__pc[23]),
    .QN(_194_)
  );
  DFF_X1 \buf__pc[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_041_),
    .Q(buf__pc[24]),
    .QN(_193_)
  );
  DFF_X1 \buf__pc[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_042_),
    .Q(buf__pc[25]),
    .QN(_192_)
  );
  DFF_X1 \buf__pc[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_043_),
    .Q(buf__pc[26]),
    .QN(_191_)
  );
  DFF_X1 \buf__pc[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_044_),
    .Q(buf__pc[27]),
    .QN(_190_)
  );
  DFF_X1 \buf__pc[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_045_),
    .Q(buf__pc[28]),
    .QN(_189_)
  );
  DFF_X1 \buf__pc[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_046_),
    .Q(buf__pc[29]),
    .QN(_188_)
  );
  DFF_X1 \buf__pc[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_019_),
    .Q(buf__pc[2]),
    .QN(_215_)
  );
  DFF_X1 \buf__pc[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_047_),
    .Q(buf__pc[30]),
    .QN(_187_)
  );
  DFF_X1 \buf__pc[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_048_),
    .Q(buf__pc[31]),
    .QN(_186_)
  );
  DFF_X1 \buf__pc[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_020_),
    .Q(buf__pc[3]),
    .QN(_214_)
  );
  DFF_X1 \buf__pc[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_021_),
    .Q(buf__pc[4]),
    .QN(_213_)
  );
  DFF_X1 \buf__pc[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_022_),
    .Q(buf__pc[5]),
    .QN(_212_)
  );
  DFF_X1 \buf__pc[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_023_),
    .Q(buf__pc[6]),
    .QN(_211_)
  );
  DFF_X1 \buf__pc[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_024_),
    .Q(buf__pc[7]),
    .QN(_210_)
  );
  DFF_X1 \buf__pc[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_025_),
    .Q(buf__pc[8]),
    .QN(_209_)
  );
  DFF_X1 \buf__pc[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_026_),
    .Q(buf__pc[9]),
    .QN(_208_)
  );
  DFF_X1 \buf__replay$_DFFE_PP_  (
    .CK(clock),
    .D(_000_),
    .Q(buf__replay),
    .QN(_234_)
  );
  DFF_X1 \buf__xcpt_ae_inst$_DFFE_PP_  (
    .CK(clock),
    .D(_050_),
    .Q(buf__xcpt_ae_inst),
    .QN(_185_)
  );
  RVCExpander exp (
    .io_in({ _icData_T_4[95:80], exp_io_in[15:0] }),
    .io_out_bits(exp_io_out_bits),
    .io_out_rd(exp_io_out_rd),
    .io_out_rs1(exp_io_out_rs1),
    .io_out_rs2(exp_io_out_rs2),
    .io_rvc(exp_io_rvc)
  );
  DFF_X1 \nBufValid$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_049_),
    .Q(nBufValid),
    .QN(_bufMask_T[0])
  );
  assign _GEN_1 = { 63'h0000000000000000, io_imem_bits_data[31:16], io_imem_bits_data[31:16], io_imem_bits_data[31:16], io_imem_bits_data[31:16], io_imem_bits_data, io_imem_bits_data[15:0], io_imem_bits_data[15:0] };
  assign _GEN_58 = { 1'h0, io_imem_bits_pc[1] };
  assign _GEN_59 = { 1'h0, nBufValid };
  assign { _GEN_67[31:3], _GEN_67[0] } = 30'h00000000;
  assign _bufMask_T[1] = nBufValid;
  assign _buf_data_T[3:0] = 4'h0;
  assign _buf_pc_T_1 = { io_imem_bits_pc[31:2], 2'h0 };
  assign _buf_pc_T_2 = { _GEN_67[2:1], 1'h0 };
  assign _buf_pc_T_4[1:0] = { _buf_data_T[4], io_imem_bits_pc[0] };
  assign _buf_pc_T_5 = { 30'h00000000, _buf_data_T[4], io_imem_bits_pc[0] };
  assign _buf_pc_T_6 = { io_imem_bits_pc[31:2], _buf_data_T[4], io_imem_bits_pc[0] };
  assign _full_insn_T_2[1] = 1'h0;
  assign _icData_T_2 = { io_imem_bits_data, io_imem_bits_data[15:0], io_imem_bits_data[15:0] };
  assign _icData_T_3[3:0] = 4'h0;
  assign { _icData_T_4[190:176], _icData_T_4[127:96] } = { 15'h0000, io_imem_bits_data[31:16], io_imem_bits_data[31:16] };
  assign _icMask_T_1 = { nBufValid, 4'h0 };
  assign _icMask_T_2 = { 15'h0000, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, 16'hffff, _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0] };
  assign _icShiftAmt_T_1 = { 1'h1, nBufValid };
  assign _ic_replay_T = { 1'h1, _bufMask_T[0] };
  assign _ic_replay_T_1[1] = _full_insn_T_2[0];
  assign _inst_T[31:16] = _icData_T_4[95:80];
  assign _inst_T_1 = { 16'h0000, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid, nBufValid };
  assign _inst_T_2[31:16] = 16'h0000;
  assign _io_inst_0_bits_xcpt1_T_4 = { 2'h0, io_imem_bits_xcpt_ae_inst };
  assign _io_inst_0_bits_xcpt1_T_5 = { 2'h0, io_inst_0_bits_xcpt1_ae_inst };
  assign _nReady_T_4[0] = exp_io_rvc;
  assign _replay_T_5[1] = 1'h0;
  assign _valid_T_2[1] = _full_insn_T_2[0];
  assign bufMask = { 1'h0, nBufValid };
  assign buf__data[31:16] = 16'h0000;
  assign buf_data_data = { io_imem_bits_data[31:16], io_imem_bits_data[31:16], io_imem_bits_data };
  assign buf_replay[1] = 1'h0;
  assign exp_io_in[31:16] = _icData_T_4[95:80];
  assign icData = _icData_T_4[95:64];
  assign icData_data = { io_imem_bits_data[31:16], io_imem_bits_data[31:16], io_imem_bits_data[31:16], io_imem_bits_data[31:16], io_imem_bits_data, io_imem_bits_data[15:0], io_imem_bits_data[15:0] };
  assign icMask = { 16'hffff, _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0], _bufMask_T[0] };
  assign icShiftAmt = _icData_T_3[5:4];
  assign io_inst_0_bits_inst_bits = exp_io_out_bits;
  assign io_inst_0_bits_inst_rd = exp_io_out_rd;
  assign io_inst_0_bits_inst_rs1 = exp_io_out_rs1;
  assign io_inst_0_bits_inst_rs2 = exp_io_out_rs2;
  assign io_inst_0_bits_raw = { _icData_T_4[95:80], exp_io_in[15:0] };
  assign io_inst_0_bits_rvc = exp_io_rvc;
  assign io_inst_0_bits_xcpt1_gf_inst = 1'h0;
  assign io_inst_0_bits_xcpt1_pf_inst = 1'h0;
  assign nIC[0] = io_imem_bits_pc[1];
  assign nICReady = _GEN_67[2:1];
  assign pcWordBits = io_imem_bits_pc[1];
  assign shamt = _buf_data_T[5:4];
  assign valid = { _full_insn_T_2[0], _valid_T_2[0] };
  assign xcpt_1_ae_inst = io_imem_bits_xcpt_ae_inst;
endmodule
module MulDiv(clock, reset, io_req_ready, io_req_valid, io_req_bits_fn, io_req_bits_in1, io_req_bits_in2, io_req_bits_tag, io_kill, io_resp_ready, io_resp_valid, io_resp_bits_data, io_resp_bits_tag);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire _1340_;
  wire _1341_;
  wire _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  wire _1351_;
  wire _1352_;
  wire _1353_;
  wire _1354_;
  wire _1355_;
  wire _1356_;
  wire _1357_;
  wire _1358_;
  wire _1359_;
  wire _1360_;
  wire _1361_;
  wire _1362_;
  wire _1363_;
  wire _1364_;
  wire _1365_;
  wire _1366_;
  wire _1367_;
  wire _1368_;
  wire _1369_;
  wire _1370_;
  wire _1371_;
  wire _1372_;
  wire _1373_;
  wire _1374_;
  wire _1375_;
  wire _1376_;
  wire _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire _1382_;
  wire _1383_;
  wire _1384_;
  wire _1385_;
  wire _1386_;
  wire _1387_;
  wire _1388_;
  wire _1389_;
  wire _1390_;
  wire _1391_;
  wire _1392_;
  wire _1393_;
  wire _1394_;
  wire _1395_;
  wire _1396_;
  wire _1397_;
  wire _1398_;
  wire _1399_;
  wire _1400_;
  wire _1401_;
  wire _1402_;
  wire _1403_;
  wire _1404_;
  wire _1405_;
  wire _1406_;
  wire _1407_;
  wire _1408_;
  wire _1409_;
  wire _1410_;
  wire _1411_;
  wire _1412_;
  wire _1413_;
  wire _1414_;
  wire _1415_;
  wire _1416_;
  wire _1417_;
  wire _1418_;
  wire _1419_;
  wire _1420_;
  wire _1421_;
  wire _1422_;
  wire _1423_;
  wire _1424_;
  wire _1425_;
  wire _1426_;
  wire _1427_;
  wire _1428_;
  wire _1429_;
  wire _1430_;
  wire _1431_;
  wire _1432_;
  wire _1433_;
  wire _1434_;
  wire _1435_;
  wire _1436_;
  wire _1437_;
  wire _1438_;
  wire _1439_;
  wire _1440_;
  wire _1441_;
  wire _1442_;
  wire _1443_;
  wire _1444_;
  wire _1445_;
  wire _1446_;
  wire _1447_;
  wire _1448_;
  wire _1449_;
  wire _1450_;
  wire _1451_;
  wire _1452_;
  wire _1453_;
  wire _1454_;
  wire _1455_;
  wire _1456_;
  wire _1457_;
  wire _1458_;
  wire _1459_;
  wire _1460_;
  wire _1461_;
  wire _1462_;
  wire _1463_;
  wire _1464_;
  wire _1465_;
  wire _1466_;
  wire _1467_;
  wire _1468_;
  wire _1469_;
  wire _1470_;
  wire _1471_;
  wire _1472_;
  wire _1473_;
  wire _1474_;
  wire _1475_;
  wire _1476_;
  wire _1477_;
  wire _1478_;
  wire _1479_;
  wire _1480_;
  wire _1481_;
  wire _1482_;
  wire _1483_;
  wire _1484_;
  wire _1485_;
  wire _1486_;
  wire _1487_;
  wire _1488_;
  wire _1489_;
  wire _1490_;
  wire _1491_;
  wire _1492_;
  wire _1493_;
  wire _1494_;
  wire _1495_;
  wire _1496_;
  wire _1497_;
  wire _1498_;
  wire _1499_;
  wire _1500_;
  wire _1501_;
  wire _1502_;
  wire _1503_;
  wire _1504_;
  wire _1505_;
  wire _1506_;
  wire _1507_;
  wire _1508_;
  wire _1509_;
  wire _1510_;
  wire _1511_;
  wire _1512_;
  wire _1513_;
  wire _1514_;
  wire _1515_;
  wire _1516_;
  wire _1517_;
  wire _1518_;
  wire _1519_;
  wire _1520_;
  wire _1521_;
  wire _1522_;
  wire _1523_;
  wire _1524_;
  wire _1525_;
  wire _1526_;
  wire _1527_;
  wire _1528_;
  wire _1529_;
  wire _1530_;
  wire _1531_;
  wire _1532_;
  wire _1533_;
  wire _1534_;
  wire _1535_;
  wire _1536_;
  wire _1537_;
  wire _1538_;
  wire _1539_;
  wire _1540_;
  wire _1541_;
  wire _1542_;
  wire _1543_;
  wire _1544_;
  wire _1545_;
  wire _1546_;
  wire _1547_;
  wire _1548_;
  wire _1549_;
  wire _1550_;
  wire _1551_;
  wire _1552_;
  wire _1553_;
  wire _1554_;
  wire _1555_;
  wire _1556_;
  wire _1557_;
  wire _1558_;
  wire _1559_;
  wire _1560_;
  wire _1561_;
  wire _1562_;
  wire _1563_;
  wire _1564_;
  wire _1565_;
  wire _1566_;
  wire _1567_;
  wire _1568_;
  wire _1569_;
  wire _1570_;
  wire _1571_;
  wire _1572_;
  wire _1573_;
  wire _1574_;
  wire _1575_;
  wire _1576_;
  wire _1577_;
  wire _1578_;
  wire _1579_;
  wire _1580_;
  wire _1581_;
  wire _1582_;
  wire _1583_;
  wire _1584_;
  wire _1585_;
  wire _1586_;
  wire _1587_;
  wire _1588_;
  wire _1589_;
  wire _1590_;
  wire _1591_;
  wire _1592_;
  wire _1593_;
  wire _1594_;
  wire _1595_;
  wire _1596_;
  wire _1597_;
  wire _1598_;
  wire _1599_;
  wire _1600_;
  wire _1601_;
  wire _1602_;
  wire _1603_;
  wire _1604_;
  wire _1605_;
  wire _1606_;
  wire _1607_;
  wire _1608_;
  wire _1609_;
  wire _1610_;
  wire _1611_;
  wire _1612_;
  wire _1613_;
  wire _1614_;
  wire _1615_;
  wire _1616_;
  wire _1617_;
  wire _1618_;
  wire _1619_;
  wire _1620_;
  wire _1621_;
  wire _1622_;
  wire _1623_;
  wire _1624_;
  wire _1625_;
  wire _1626_;
  wire _1627_;
  wire _1628_;
  wire _1629_;
  wire _1630_;
  wire _1631_;
  wire _1632_;
  wire _1633_;
  wire _1634_;
  wire _1635_;
  wire _1636_;
  wire _1637_;
  wire _1638_;
  wire _1639_;
  wire _1640_;
  wire _1641_;
  wire _1642_;
  wire _1643_;
  wire _1644_;
  wire _1645_;
  wire _1646_;
  wire _1647_;
  wire _1648_;
  wire _1649_;
  wire _1650_;
  wire _1651_;
  wire _1652_;
  wire _1653_;
  wire _1654_;
  wire _1655_;
  wire _1656_;
  wire _1657_;
  wire _1658_;
  wire _1659_;
  wire _1660_;
  wire _1661_;
  wire _1662_;
  wire _1663_;
  wire _1664_;
  wire _1665_;
  wire _1666_;
  wire _1667_;
  wire _1668_;
  wire _1669_;
  wire _1670_;
  wire _1671_;
  wire _1672_;
  wire _1673_;
  wire _1674_;
  wire _1675_;
  wire _1676_;
  wire _1677_;
  wire _1678_;
  wire _1679_;
  wire _1680_;
  wire _1681_;
  wire _1682_;
  wire _1683_;
  wire _1684_;
  wire _1685_;
  wire _1686_;
  wire _1687_;
  wire _1688_;
  wire _1689_;
  wire _1690_;
  wire _1691_;
  wire _1692_;
  wire _1693_;
  wire _1694_;
  wire _1695_;
  wire _1696_;
  wire _1697_;
  wire _1698_;
  wire _1699_;
  wire _1700_;
  wire _1701_;
  wire _1702_;
  wire _1703_;
  wire _1704_;
  wire _1705_;
  wire _1706_;
  wire _1707_;
  wire _1708_;
  wire _1709_;
  wire _1710_;
  wire _1711_;
  wire _1712_;
  wire _1713_;
  wire _1714_;
  wire _1715_;
  wire _1716_;
  wire _1717_;
  wire _1718_;
  wire _1719_;
  wire _1720_;
  wire _1721_;
  wire _1722_;
  wire _1723_;
  wire _1724_;
  wire _1725_;
  wire _1726_;
  wire _1727_;
  wire _1728_;
  wire _1729_;
  wire _1730_;
  wire _1731_;
  wire _1732_;
  wire _1733_;
  wire _1734_;
  wire _1735_;
  wire _1736_;
  wire _1737_;
  wire _1738_;
  wire _1739_;
  wire _1740_;
  wire _1741_;
  wire _1742_;
  wire _1743_;
  wire _1744_;
  wire _1745_;
  wire _1746_;
  wire _1747_;
  wire _1748_;
  wire _1749_;
  wire _1750_;
  wire _1751_;
  wire _1752_;
  wire _1753_;
  wire _1754_;
  wire _1755_;
  wire _1756_;
  wire _1757_;
  wire _1758_;
  wire _1759_;
  wire _1760_;
  wire _1761_;
  wire _1762_;
  wire _1763_;
  wire _1764_;
  wire _1765_;
  wire _1766_;
  wire _1767_;
  wire _1768_;
  wire _1769_;
  wire _1770_;
  wire _1771_;
  wire _1772_;
  wire _1773_;
  wire _1774_;
  wire _1775_;
  wire _1776_;
  wire _1777_;
  wire _1778_;
  wire _1779_;
  wire _1780_;
  wire _1781_;
  wire _1782_;
  wire _1783_;
  wire _1784_;
  wire _1785_;
  wire _1786_;
  wire _1787_;
  wire _1788_;
  wire _1789_;
  wire _1790_;
  wire _1791_;
  wire _1792_;
  wire _1793_;
  wire _1794_;
  wire _1795_;
  wire _1796_;
  wire _1797_;
  wire _1798_;
  wire _1799_;
  wire _1800_;
  wire _1801_;
  wire _1802_;
  wire _1803_;
  wire _1804_;
  wire _1805_;
  wire _1806_;
  wire _1807_;
  wire _1808_;
  wire _1809_;
  wire _1810_;
  wire _1811_;
  wire _1812_;
  wire _1813_;
  wire _1814_;
  wire _1815_;
  wire _1816_;
  wire _1817_;
  wire _1818_;
  wire _1819_;
  wire _1820_;
  wire _1821_;
  wire _1822_;
  wire _1823_;
  wire _1824_;
  wire _1825_;
  wire _1826_;
  wire _1827_;
  wire _1828_;
  wire _1829_;
  wire _1830_;
  wire _1831_;
  wire _1832_;
  wire _1833_;
  wire _1834_;
  wire _1835_;
  wire _1836_;
  wire _1837_;
  wire _1838_;
  wire _1839_;
  wire _1840_;
  wire _1841_;
  wire _1842_;
  wire _1843_;
  wire _1844_;
  wire _1845_;
  wire _1846_;
  wire _1847_;
  wire _1848_;
  wire _1849_;
  wire _1850_;
  wire _1851_;
  wire _1852_;
  wire _1853_;
  wire _1854_;
  wire _1855_;
  wire _1856_;
  wire _1857_;
  wire _1858_;
  wire _1859_;
  wire _1860_;
  wire _1861_;
  wire _1862_;
  wire _1863_;
  wire _1864_;
  wire _1865_;
  wire _1866_;
  wire _1867_;
  wire _1868_;
  wire _1869_;
  wire _1870_;
  wire _1871_;
  wire _1872_;
  wire _1873_;
  wire _1874_;
  wire _1875_;
  wire _1876_;
  wire _1877_;
  wire _1878_;
  wire _1879_;
  wire _1880_;
  wire _1881_;
  wire _1882_;
  wire _1883_;
  wire _1884_;
  wire _1885_;
  wire _1886_;
  wire _1887_;
  wire _1888_;
  wire _1889_;
  wire _1890_;
  wire _1891_;
  wire _1892_;
  wire _1893_;
  wire _1894_;
  wire _1895_;
  wire _1896_;
  wire _1897_;
  wire _1898_;
  wire _1899_;
  wire _1900_;
  wire _1901_;
  wire _1902_;
  wire _1903_;
  wire _1904_;
  wire _1905_;
  wire _1906_;
  wire _1907_;
  wire _1908_;
  wire _1909_;
  wire _1910_;
  wire _1911_;
  wire _1912_;
  wire _1913_;
  wire _1914_;
  wire _1915_;
  wire _1916_;
  wire _1917_;
  wire _1918_;
  wire _1919_;
  wire _1920_;
  wire _1921_;
  wire _1922_;
  wire _1923_;
  wire _1924_;
  wire _1925_;
  wire _1926_;
  wire _1927_;
  wire _1928_;
  wire _1929_;
  wire _1930_;
  wire _1931_;
  wire _1932_;
  wire _1933_;
  wire _1934_;
  wire _1935_;
  wire _1936_;
  wire _1937_;
  wire _1938_;
  wire _1939_;
  wire _1940_;
  wire _1941_;
  wire _1942_;
  wire _1943_;
  wire _1944_;
  wire _1945_;
  wire _1946_;
  wire _1947_;
  wire _1948_;
  wire _1949_;
  wire _1950_;
  wire _1951_;
  wire _1952_;
  wire _1953_;
  wire _1954_;
  wire _1955_;
  wire _1956_;
  wire _1957_;
  wire _1958_;
  wire _1959_;
  wire _1960_;
  wire _1961_;
  wire _1962_;
  wire _1963_;
  wire _1964_;
  wire _1965_;
  wire _1966_;
  wire _1967_;
  wire _1968_;
  wire _1969_;
  wire _1970_;
  wire _1971_;
  wire _1972_;
  wire _1973_;
  wire _1974_;
  wire _1975_;
  wire _1976_;
  wire _1977_;
  wire _1978_;
  wire _1979_;
  wire _1980_;
  wire _1981_;
  wire _1982_;
  wire _1983_;
  wire _1984_;
  wire _1985_;
  wire _1986_;
  wire _1987_;
  wire _1988_;
  wire _1989_;
  wire _1990_;
  wire _1991_;
  wire _1992_;
  wire _1993_;
  wire _1994_;
  wire _1995_;
  wire _1996_;
  wire _1997_;
  wire _1998_;
  wire _1999_;
  wire _2000_;
  wire _2001_;
  wire _2002_;
  wire _2003_;
  wire _2004_;
  wire _2005_;
  wire _2006_;
  wire _2007_;
  wire _2008_;
  wire _2009_;
  wire _2010_;
  wire _2011_;
  wire _2012_;
  wire _2013_;
  wire _2014_;
  wire _2015_;
  wire _2016_;
  wire _2017_;
  wire _2018_;
  wire _2019_;
  wire _2020_;
  wire _2021_;
  wire _2022_;
  wire _2023_;
  wire _2024_;
  wire _2025_;
  wire _2026_;
  wire _2027_;
  wire _2028_;
  wire _2029_;
  wire _2030_;
  wire _2031_;
  wire _2032_;
  wire _2033_;
  wire _2034_;
  wire _2035_;
  wire _2036_;
  wire _2037_;
  wire _2038_;
  wire _2039_;
  wire _2040_;
  wire _2041_;
  wire _2042_;
  wire _2043_;
  wire _2044_;
  wire _2045_;
  wire _2046_;
  wire _2047_;
  wire _2048_;
  wire _2049_;
  wire _2050_;
  wire _2051_;
  wire _2052_;
  wire _2053_;
  wire _2054_;
  wire _2055_;
  wire _2056_;
  wire _2057_;
  wire _2058_;
  wire _2059_;
  wire _2060_;
  wire _2061_;
  wire _2062_;
  wire _2063_;
  wire _2064_;
  wire _2065_;
  wire _2066_;
  wire _2067_;
  wire _2068_;
  wire _2069_;
  wire _2070_;
  wire _2071_;
  wire _2072_;
  wire _2073_;
  wire _2074_;
  wire _2075_;
  wire _2076_;
  wire _2077_;
  wire _2078_;
  wire _2079_;
  wire _2080_;
  wire _2081_;
  wire _2082_;
  wire _2083_;
  wire _2084_;
  wire _2085_;
  wire _2086_;
  wire _2087_;
  wire _2088_;
  wire _2089_;
  wire _2090_;
  wire _2091_;
  wire _2092_;
  wire _2093_;
  wire _2094_;
  wire _2095_;
  wire _2096_;
  wire _2097_;
  wire _2098_;
  wire _2099_;
  wire _2100_;
  wire _2101_;
  wire _2102_;
  wire _2103_;
  wire _2104_;
  wire _2105_;
  wire _2106_;
  wire _2107_;
  wire _2108_;
  wire _2109_;
  wire _2110_;
  wire _2111_;
  wire _2112_;
  wire _2113_;
  wire _2114_;
  wire _2115_;
  wire _2116_;
  wire _2117_;
  wire _2118_;
  wire _2119_;
  wire _2120_;
  wire _2121_;
  wire _2122_;
  wire _2123_;
  wire _2124_;
  wire _2125_;
  wire _2126_;
  wire _2127_;
  wire _2128_;
  wire _2129_;
  wire _2130_;
  wire _2131_;
  wire _2132_;
  wire _2133_;
  wire _2134_;
  wire _2135_;
  wire _2136_;
  wire _2137_;
  wire _2138_;
  wire _2139_;
  wire _2140_;
  wire _2141_;
  wire _2142_;
  wire _2143_;
  wire _2144_;
  wire _2145_;
  wire _2146_;
  wire _2147_;
  wire _2148_;
  wire _2149_;
  wire _2150_;
  wire _2151_;
  wire _2152_;
  wire _2153_;
  wire _2154_;
  wire _2155_;
  wire _2156_;
  wire _2157_;
  wire _2158_;
  wire _2159_;
  wire _2160_;
  wire _2161_;
  wire _2162_;
  wire _2163_;
  wire _2164_;
  wire _2165_;
  wire _2166_;
  wire _2167_;
  wire _2168_;
  wire _2169_;
  wire _2170_;
  wire _2171_;
  wire _2172_;
  wire _2173_;
  wire _2174_;
  wire _2175_;
  wire _2176_;
  wire _2177_;
  wire _2178_;
  wire _2179_;
  wire _2180_;
  wire _2181_;
  wire _2182_;
  wire _2183_;
  wire _2184_;
  wire _2185_;
  wire _2186_;
  wire _2187_;
  wire _2188_;
  wire _2189_;
  wire _2190_;
  wire _2191_;
  wire _2192_;
  wire _2193_;
  wire _2194_;
  wire _2195_;
  wire _2196_;
  wire _2197_;
  wire _2198_;
  wire _2199_;
  wire _2200_;
  wire _2201_;
  wire _2202_;
  wire _2203_;
  wire _2204_;
  wire _2205_;
  wire _2206_;
  wire _2207_;
  wire _2208_;
  wire _2209_;
  wire _2210_;
  wire _2211_;
  wire _2212_;
  wire _2213_;
  wire _2214_;
  wire _2215_;
  wire _2216_;
  wire _2217_;
  wire _2218_;
  wire _2219_;
  wire _2220_;
  wire _2221_;
  wire _2222_;
  wire _2223_;
  wire _2224_;
  wire _2225_;
  wire _2226_;
  wire _2227_;
  wire _2228_;
  wire _2229_;
  wire _2230_;
  wire _2231_;
  wire _2232_;
  wire _2233_;
  wire _2234_;
  wire _2235_;
  wire _2236_;
  wire _2237_;
  wire _2238_;
  wire _2239_;
  wire _2240_;
  wire _2241_;
  wire _2242_;
  wire _2243_;
  wire _2244_;
  wire _2245_;
  wire _2246_;
  wire _2247_;
  wire _2248_;
  wire _2249_;
  wire _2250_;
  wire _2251_;
  wire _2252_;
  wire _2253_;
  wire _2254_;
  wire _2255_;
  wire _2256_;
  wire _2257_;
  wire _2258_;
  wire _2259_;
  wire _2260_;
  wire _2261_;
  wire _2262_;
  wire _2263_;
  wire _2264_;
  wire _2265_;
  wire _2266_;
  wire _2267_;
  wire _2268_;
  wire _2269_;
  wire _2270_;
  wire _2271_;
  wire _2272_;
  wire _2273_;
  wire _2274_;
  wire _2275_;
  wire _2276_;
  wire _2277_;
  wire _2278_;
  wire _2279_;
  wire _2280_;
  wire _2281_;
  wire _2282_;
  wire _2283_;
  wire _2284_;
  wire _2285_;
  wire _2286_;
  wire _2287_;
  wire _2288_;
  wire _2289_;
  wire _2290_;
  wire _2291_;
  wire _2292_;
  wire _2293_;
  wire _2294_;
  wire _2295_;
  wire _2296_;
  wire _2297_;
  wire _2298_;
  wire _2299_;
  wire _2300_;
  wire _2301_;
  wire _2302_;
  wire _2303_;
  wire _2304_;
  wire _2305_;
  wire _2306_;
  wire _2307_;
  wire _2308_;
  wire _2309_;
  wire _2310_;
  wire _2311_;
  wire _2312_;
  wire _2313_;
  wire _2314_;
  wire _2315_;
  wire _2316_;
  wire _2317_;
  wire _2318_;
  wire _2319_;
  wire _2320_;
  wire _2321_;
  wire _2322_;
  wire _2323_;
  wire _2324_;
  wire _2325_;
  wire _2326_;
  wire _2327_;
  wire _2328_;
  wire _2329_;
  wire _2330_;
  wire _2331_;
  wire _2332_;
  wire _2333_;
  wire _2334_;
  wire _2335_;
  wire _2336_;
  wire _2337_;
  wire _2338_;
  wire _2339_;
  wire _2340_;
  wire _2341_;
  wire _2342_;
  wire _2343_;
  wire _2344_;
  wire _2345_;
  wire _2346_;
  wire _2347_;
  wire _2348_;
  wire _2349_;
  wire _2350_;
  wire _2351_;
  wire _2352_;
  wire _2353_;
  wire _2354_;
  wire _2355_;
  wire _2356_;
  wire _2357_;
  wire _2358_;
  wire _2359_;
  wire _2360_;
  wire _2361_;
  wire _2362_;
  wire _2363_;
  wire _2364_;
  wire _2365_;
  wire _2366_;
  wire _2367_;
  wire _2368_;
  wire _2369_;
  wire _2370_;
  wire _2371_;
  wire _2372_;
  wire _2373_;
  wire _2374_;
  wire _2375_;
  wire _2376_;
  wire _2377_;
  wire _2378_;
  wire _2379_;
  wire _2380_;
  wire _2381_;
  wire _2382_;
  wire _2383_;
  wire _2384_;
  wire _2385_;
  wire _2386_;
  wire _2387_;
  wire _2388_;
  wire _2389_;
  wire _2390_;
  wire _2391_;
  wire _2392_;
  wire _2393_;
  wire _2394_;
  wire _2395_;
  wire _2396_;
  wire _2397_;
  wire _2398_;
  wire _2399_;
  wire _2400_;
  wire _2401_;
  wire _2402_;
  wire _2403_;
  wire _2404_;
  wire _2405_;
  wire _2406_;
  wire _2407_;
  wire _2408_;
  wire _2409_;
  wire _2410_;
  wire _2411_;
  wire _2412_;
  wire _2413_;
  wire _2414_;
  wire _2415_;
  wire _2416_;
  wire _2417_;
  wire _2418_;
  wire _2419_;
  wire _2420_;
  wire _2421_;
  wire _2422_;
  wire _2423_;
  wire _2424_;
  wire _2425_;
  wire _2426_;
  wire _2427_;
  wire _2428_;
  wire _2429_;
  wire _2430_;
  wire _2431_;
  wire _2432_;
  wire _2433_;
  wire _2434_;
  wire _2435_;
  wire _2436_;
  wire _2437_;
  wire _2438_;
  wire _2439_;
  wire _2440_;
  wire _2441_;
  wire _2442_;
  wire _2443_;
  wire _2444_;
  wire _2445_;
  wire _2446_;
  wire _2447_;
  wire _2448_;
  wire _2449_;
  wire _2450_;
  wire _2451_;
  wire _2452_;
  wire _2453_;
  wire _2454_;
  wire _2455_;
  wire _2456_;
  wire _2457_;
  wire _2458_;
  wire _2459_;
  wire _2460_;
  wire _2461_;
  wire _2462_;
  wire _2463_;
  wire _2464_;
  wire _2465_;
  wire _2466_;
  wire _2467_;
  wire _2468_;
  wire _2469_;
  wire _2470_;
  wire _2471_;
  wire _2472_;
  wire _2473_;
  wire _2474_;
  wire _2475_;
  wire _2476_;
  wire _2477_;
  wire _2478_;
  wire _2479_;
  wire _2480_;
  wire _2481_;
  wire _2482_;
  wire _2483_;
  wire _2484_;
  wire _2485_;
  wire _2486_;
  wire _2487_;
  wire _2488_;
  wire _2489_;
  wire _2490_;
  wire _2491_;
  wire _2492_;
  wire _2493_;
  wire _2494_;
  wire _2495_;
  wire _2496_;
  wire _2497_;
  wire _2498_;
  wire _2499_;
  wire _2500_;
  wire _2501_;
  wire _2502_;
  wire _2503_;
  wire _2504_;
  wire _2505_;
  wire _2506_;
  wire _2507_;
  wire _2508_;
  wire _2509_;
  wire _2510_;
  wire _2511_;
  wire _2512_;
  wire _2513_;
  wire _2514_;
  wire _2515_;
  wire _2516_;
  wire _2517_;
  wire _2518_;
  wire _2519_;
  wire _2520_;
  wire _2521_;
  wire _2522_;
  wire _2523_;
  wire _2524_;
  wire _2525_;
  wire _2526_;
  wire _2527_;
  wire _2528_;
  wire _2529_;
  wire _2530_;
  wire _2531_;
  wire _2532_;
  wire _2533_;
  wire _2534_;
  wire _2535_;
  wire _2536_;
  wire _2537_;
  wire _2538_;
  wire _2539_;
  wire _2540_;
  wire _2541_;
  wire _2542_;
  wire _2543_;
  wire _2544_;
  wire _2545_;
  wire _2546_;
  wire _2547_;
  wire _2548_;
  wire _2549_;
  wire _2550_;
  wire _2551_;
  wire _2552_;
  wire _2553_;
  wire _2554_;
  wire _2555_;
  wire _2556_;
  wire _2557_;
  wire _2558_;
  wire _2559_;
  wire _2560_;
  wire _2561_;
  wire _2562_;
  wire _2563_;
  wire _2564_;
  wire _2565_;
  wire _2566_;
  wire _2567_;
  wire _2568_;
  wire _2569_;
  wire _2570_;
  wire _2571_;
  wire _2572_;
  wire _2573_;
  wire _2574_;
  wire _2575_;
  wire _2576_;
  wire _2577_;
  wire _2578_;
  wire _2579_;
  wire _2580_;
  wire _2581_;
  wire _2582_;
  wire _2583_;
  wire _2584_;
  wire _2585_;
  wire _2586_;
  wire _2587_;
  wire _2588_;
  wire _2589_;
  wire _2590_;
  wire _2591_;
  wire _2592_;
  wire _2593_;
  wire _2594_;
  wire _2595_;
  wire _2596_;
  wire _2597_;
  wire _2598_;
  wire _2599_;
  wire _2600_;
  wire _2601_;
  wire _2602_;
  wire _2603_;
  wire _2604_;
  wire _2605_;
  wire _2606_;
  wire _2607_;
  wire _2608_;
  wire _2609_;
  wire _2610_;
  wire _2611_;
  wire _2612_;
  wire _2613_;
  wire _2614_;
  wire _2615_;
  wire _2616_;
  wire _2617_;
  wire _2618_;
  wire _2619_;
  wire _2620_;
  wire _2621_;
  wire _2622_;
  wire _2623_;
  wire _2624_;
  wire _2625_;
  wire _2626_;
  wire _2627_;
  wire _2628_;
  wire _2629_;
  wire _2630_;
  wire _2631_;
  wire _2632_;
  wire _2633_;
  wire _2634_;
  wire _2635_;
  wire _2636_;
  wire _2637_;
  wire _2638_;
  wire _2639_;
  wire _2640_;
  wire _2641_;
  wire _2642_;
  wire _2643_;
  wire _2644_;
  wire _2645_;
  wire _2646_;
  wire _2647_;
  wire _2648_;
  wire _2649_;
  wire _2650_;
  wire _2651_;
  wire _2652_;
  wire _2653_;
  wire _2654_;
  wire _2655_;
  wire _2656_;
  wire _2657_;
  wire _2658_;
  wire _2659_;
  wire _2660_;
  wire _2661_;
  wire _2662_;
  wire _2663_;
  wire _2664_;
  wire _2665_;
  wire _2666_;
  wire _2667_;
  wire _2668_;
  wire _2669_;
  wire _2670_;
  wire _2671_;
  wire _2672_;
  wire _2673_;
  wire _2674_;
  wire _2675_;
  wire _2676_;
  wire _2677_;
  wire _2678_;
  wire _2679_;
  wire _2680_;
  wire _2681_;
  wire _2682_;
  wire _2683_;
  wire _2684_;
  wire _2685_;
  wire _2686_;
  wire _2687_;
  wire _2688_;
  wire _2689_;
  wire _2690_;
  wire _2691_;
  wire _2692_;
  wire _2693_;
  wire _2694_;
  wire _2695_;
  wire _2696_;
  wire _2697_;
  wire _2698_;
  wire _2699_;
  wire _2700_;
  wire _2701_;
  wire _2702_;
  wire _2703_;
  wire _2704_;
  wire _2705_;
  wire _2706_;
  wire _2707_;
  wire _2708_;
  wire _2709_;
  wire _2710_;
  wire _2711_;
  wire _2712_;
  wire _2713_;
  wire _2714_;
  wire _2715_;
  wire _2716_;
  wire _2717_;
  wire _2718_;
  wire _2719_;
  wire _2720_;
  wire _2721_;
  wire _2722_;
  wire _2723_;
  wire _2724_;
  wire _2725_;
  wire _2726_;
  wire _2727_;
  wire _2728_;
  wire _2729_;
  wire _2730_;
  wire _2731_;
  wire _2732_;
  wire _2733_;
  wire _2734_;
  wire _2735_;
  wire _2736_;
  wire _2737_;
  wire _2738_;
  wire _2739_;
  wire _2740_;
  wire _2741_;
  wire _2742_;
  wire _2743_;
  wire _2744_;
  wire _2745_;
  wire _2746_;
  wire _2747_;
  wire _2748_;
  wire _2749_;
  wire _2750_;
  wire _2751_;
  wire _2752_;
  wire _2753_;
  wire _2754_;
  wire _2755_;
  wire _2756_;
  wire _2757_;
  wire _2758_;
  wire _2759_;
  wire _2760_;
  wire _2761_;
  wire _2762_;
  wire _2763_;
  wire _2764_;
  wire _2765_;
  wire _2766_;
  wire _2767_;
  wire _2768_;
  wire _2769_;
  wire _2770_;
  wire _2771_;
  wire _2772_;
  wire _2773_;
  wire _2774_;
  wire _2775_;
  wire _2776_;
  wire _2777_;
  wire _2778_;
  wire _2779_;
  wire _2780_;
  wire _2781_;
  wire _2782_;
  wire _2783_;
  wire _2784_;
  wire _2785_;
  wire _2786_;
  wire _2787_;
  wire _2788_;
  wire _2789_;
  wire _2790_;
  wire _2791_;
  wire _2792_;
  wire _2793_;
  wire _2794_;
  wire _2795_;
  wire _2796_;
  wire _2797_;
  wire _2798_;
  wire _2799_;
  wire _2800_;
  wire _2801_;
  wire _2802_;
  wire _2803_;
  wire _2804_;
  wire _2805_;
  wire _2806_;
  wire _2807_;
  wire _2808_;
  wire _2809_;
  wire _2810_;
  wire _2811_;
  wire _2812_;
  wire _2813_;
  wire _2814_;
  wire _2815_;
  wire _2816_;
  wire _2817_;
  wire _2818_;
  wire _2819_;
  wire _2820_;
  wire _2821_;
  wire _2822_;
  wire _2823_;
  wire _2824_;
  wire _2825_;
  wire _2826_;
  wire _2827_;
  wire _2828_;
  wire _2829_;
  wire _2830_;
  wire _2831_;
  wire _2832_;
  wire _2833_;
  wire _2834_;
  wire _2835_;
  wire _2836_;
  wire _2837_;
  wire _2838_;
  wire _2839_;
  wire _2840_;
  wire _2841_;
  wire _2842_;
  wire _2843_;
  wire _2844_;
  wire _2845_;
  wire _2846_;
  wire _2847_;
  wire _2848_;
  wire _2849_;
  wire _2850_;
  wire _2851_;
  wire _2852_;
  wire _2853_;
  wire _2854_;
  wire _2855_;
  wire _2856_;
  wire _2857_;
  wire _2858_;
  wire _2859_;
  wire _2860_;
  wire _2861_;
  wire _2862_;
  wire _2863_;
  wire _2864_;
  wire _2865_;
  wire _2866_;
  wire _2867_;
  wire _2868_;
  wire _2869_;
  wire _2870_;
  wire _2871_;
  wire _2872_;
  wire _2873_;
  wire _2874_;
  wire _2875_;
  wire _2876_;
  wire _2877_;
  wire _2878_;
  wire _2879_;
  wire _2880_;
  wire _2881_;
  wire _2882_;
  wire _2883_;
  wire _2884_;
  wire _2885_;
  wire _2886_;
  wire _2887_;
  wire _2888_;
  wire _2889_;
  wire _2890_;
  wire _2891_;
  wire _2892_;
  wire _2893_;
  wire _2894_;
  wire _2895_;
  wire _2896_;
  wire _2897_;
  wire _2898_;
  wire _2899_;
  wire _2900_;
  wire _2901_;
  wire _2902_;
  wire _2903_;
  wire _2904_;
  wire _2905_;
  wire _2906_;
  wire _2907_;
  wire _2908_;
  wire _2909_;
  wire _2910_;
  wire _2911_;
  wire _2912_;
  wire _2913_;
  wire _2914_;
  wire _2915_;
  wire _2916_;
  wire _2917_;
  wire _2918_;
  wire _2919_;
  wire _2920_;
  wire _2921_;
  wire _2922_;
  wire _2923_;
  wire _2924_;
  wire _2925_;
  wire _2926_;
  wire _2927_;
  wire _2928_;
  wire _2929_;
  wire _2930_;
  wire _2931_;
  wire _2932_;
  wire _2933_;
  wire _2934_;
  wire _2935_;
  wire _2936_;
  wire _2937_;
  wire _2938_;
  wire _2939_;
  wire _2940_;
  wire _2941_;
  wire _2942_;
  wire _2943_;
  wire _2944_;
  wire _2945_;
  wire _2946_;
  wire _2947_;
  wire _2948_;
  wire _2949_;
  wire _2950_;
  wire _2951_;
  wire _2952_;
  wire _2953_;
  wire _2954_;
  wire _2955_;
  wire _2956_;
  wire _2957_;
  wire _2958_;
  wire _2959_;
  wire _2960_;
  wire _2961_;
  wire _2962_;
  wire _2963_;
  wire _2964_;
  wire _2965_;
  wire _2966_;
  wire _2967_;
  wire _2968_;
  wire _2969_;
  wire _2970_;
  wire _2971_;
  wire _2972_;
  wire _2973_;
  wire _2974_;
  wire _2975_;
  wire _2976_;
  wire _2977_;
  wire _2978_;
  wire _2979_;
  wire _2980_;
  wire _2981_;
  wire _2982_;
  wire _2983_;
  wire _2984_;
  wire _2985_;
  wire _2986_;
  wire _2987_;
  wire _2988_;
  wire _2989_;
  wire _2990_;
  wire _2991_;
  wire _2992_;
  wire _2993_;
  wire _2994_;
  wire _2995_;
  wire _2996_;
  wire _2997_;
  wire _2998_;
  wire _2999_;
  wire _3000_;
  wire _3001_;
  wire _3002_;
  wire _3003_;
  wire _3004_;
  wire _3005_;
  wire _3006_;
  wire _3007_;
  wire _3008_;
  wire _3009_;
  wire _3010_;
  wire _3011_;
  wire _3012_;
  wire _3013_;
  wire _3014_;
  wire _3015_;
  wire _3016_;
  wire _3017_;
  wire _3018_;
  wire _3019_;
  wire _3020_;
  wire _3021_;
  wire _3022_;
  wire _3023_;
  wire _3024_;
  wire _3025_;
  wire _3026_;
  wire _3027_;
  wire _3028_;
  wire _3029_;
  wire _3030_;
  wire _3031_;
  wire _3032_;
  wire _3033_;
  wire _3034_;
  wire _3035_;
  wire _3036_;
  wire _3037_;
  wire _3038_;
  wire _3039_;
  wire _3040_;
  wire _3041_;
  wire _3042_;
  wire _3043_;
  wire _3044_;
  wire _3045_;
  wire _3046_;
  wire _3047_;
  wire _3048_;
  wire _3049_;
  wire _3050_;
  wire _3051_;
  wire _3052_;
  wire _3053_;
  wire _3054_;
  wire _3055_;
  wire _3056_;
  wire _3057_;
  wire _3058_;
  wire _3059_;
  wire _3060_;
  wire _3061_;
  wire _3062_;
  wire _3063_;
  wire _3064_;
  wire _3065_;
  wire _3066_;
  wire _3067_;
  wire _3068_;
  wire _3069_;
  wire _3070_;
  wire _3071_;
  wire _3072_;
  wire _3073_;
  wire _3074_;
  wire _3075_;
  wire _3076_;
  wire _3077_;
  wire _3078_;
  wire _3079_;
  wire _3080_;
  wire _3081_;
  wire _3082_;
  wire _3083_;
  wire _3084_;
  wire _3085_;
  wire _3086_;
  wire _3087_;
  wire _3088_;
  wire _3089_;
  wire _3090_;
  wire _3091_;
  wire _3092_;
  wire _3093_;
  wire _3094_;
  wire _3095_;
  wire _3096_;
  wire _3097_;
  wire _3098_;
  wire _3099_;
  wire _3100_;
  wire _3101_;
  wire _3102_;
  wire _3103_;
  wire _3104_;
  wire _3105_;
  wire _3106_;
  wire _3107_;
  wire _3108_;
  wire _3109_;
  wire _3110_;
  wire _3111_;
  wire _3112_;
  wire _3113_;
  wire _3114_;
  wire _3115_;
  wire _3116_;
  wire _3117_;
  wire _3118_;
  wire _3119_;
  wire _3120_;
  wire _3121_;
  wire _3122_;
  wire _3123_;
  wire _3124_;
  wire _3125_;
  wire _3126_;
  wire _3127_;
  wire _3128_;
  wire _3129_;
  wire _3130_;
  wire _3131_;
  wire _3132_;
  wire _3133_;
  wire _3134_;
  wire _3135_;
  wire _3136_;
  wire _3137_;
  wire _3138_;
  wire _3139_;
  wire _3140_;
  wire _3141_;
  wire _3142_;
  wire _3143_;
  wire _3144_;
  wire _3145_;
  wire _3146_;
  wire _3147_;
  wire _3148_;
  wire _3149_;
  wire _3150_;
  wire _3151_;
  wire _3152_;
  wire _3153_;
  wire _3154_;
  wire _3155_;
  wire _3156_;
  wire _3157_;
  wire _3158_;
  wire _3159_;
  wire _3160_;
  wire _3161_;
  wire _3162_;
  wire _3163_;
  wire _3164_;
  wire _3165_;
  wire _3166_;
  wire _3167_;
  wire _3168_;
  wire _3169_;
  wire _3170_;
  wire _3171_;
  wire _3172_;
  wire _3173_;
  wire _3174_;
  wire _3175_;
  wire _3176_;
  wire _3177_;
  wire _3178_;
  wire _3179_;
  wire _3180_;
  wire _3181_;
  wire _3182_;
  wire _3183_;
  wire _3184_;
  wire _3185_;
  wire _3186_;
  wire _3187_;
  wire _3188_;
  wire _3189_;
  wire _3190_;
  wire _3191_;
  wire _3192_;
  wire _3193_;
  wire _3194_;
  wire _3195_;
  wire _3196_;
  wire _3197_;
  wire _3198_;
  wire _3199_;
  wire _3200_;
  wire _3201_;
  wire _3202_;
  wire _3203_;
  wire _3204_;
  wire _3205_;
  wire _3206_;
  wire _3207_;
  wire _3208_;
  wire _3209_;
  wire _3210_;
  wire _3211_;
  wire _3212_;
  wire _3213_;
  wire _3214_;
  wire _3215_;
  wire _3216_;
  wire _3217_;
  wire _3218_;
  wire _3219_;
  wire _3220_;
  wire _3221_;
  wire _3222_;
  wire _3223_;
  wire _3224_;
  wire _3225_;
  wire _3226_;
  wire _3227_;
  wire _3228_;
  wire _3229_;
  wire _3230_;
  wire _3231_;
  wire _3232_;
  wire _3233_;
  wire _3234_;
  wire _3235_;
  wire _3236_;
  wire _3237_;
  wire _3238_;
  wire _3239_;
  wire _3240_;
  wire _3241_;
  wire _3242_;
  wire _3243_;
  wire _3244_;
  wire _3245_;
  wire _3246_;
  wire _3247_;
  wire _3248_;
  wire _3249_;
  wire _3250_;
  wire _3251_;
  wire _3252_;
  wire _3253_;
  wire _3254_;
  wire _3255_;
  wire _3256_;
  wire _3257_;
  wire _3258_;
  wire _3259_;
  wire _3260_;
  wire _3261_;
  wire _3262_;
  wire _3263_;
  wire _3264_;
  wire _3265_;
  wire _3266_;
  wire _3267_;
  wire _3268_;
  wire _3269_;
  wire _3270_;
  wire _3271_;
  wire _3272_;
  wire _3273_;
  wire _3274_;
  wire _3275_;
  wire _3276_;
  wire _3277_;
  wire _3278_;
  wire _3279_;
  wire _3280_;
  wire _3281_;
  wire _3282_;
  wire _3283_;
  wire _3284_;
  wire _3285_;
  wire _3286_;
  wire _3287_;
  wire _3288_;
  wire _3289_;
  wire _3290_;
  wire _3291_;
  wire _3292_;
  wire _3293_;
  wire _3294_;
  wire _3295_;
  wire _3296_;
  wire _3297_;
  wire _3298_;
  wire _3299_;
  wire _3300_;
  wire _3301_;
  wire _3302_;
  wire _3303_;
  wire _3304_;
  wire _3305_;
  wire _3306_;
  wire _3307_;
  wire _3308_;
  wire _3309_;
  wire _3310_;
  wire _3311_;
  wire _3312_;
  wire _3313_;
  wire _3314_;
  wire _3315_;
  wire _3316_;
  wire _3317_;
  wire _3318_;
  wire _3319_;
  wire _3320_;
  wire _3321_;
  wire _3322_;
  wire _3323_;
  wire _3324_;
  wire _3325_;
  wire _3326_;
  wire _3327_;
  wire _3328_;
  wire _3329_;
  wire _3330_;
  wire _3331_;
  wire _3332_;
  wire _3333_;
  wire _3334_;
  wire _3335_;
  wire _3336_;
  wire _3337_;
  wire _3338_;
  wire _3339_;
  wire _3340_;
  wire _3341_;
  wire _3342_;
  wire _3343_;
  wire _3344_;
  wire _3345_;
  wire _3346_;
  wire _3347_;
  wire _3348_;
  wire _3349_;
  wire _3350_;
  wire _3351_;
  wire _3352_;
  wire _3353_;
  wire _3354_;
  wire _3355_;
  wire _3356_;
  wire _3357_;
  wire _3358_;
  wire _3359_;
  wire _3360_;
  wire _3361_;
  wire _3362_;
  wire _3363_;
  wire _3364_;
  wire _3365_;
  wire _3366_;
  wire _3367_;
  wire _3368_;
  wire _3369_;
  wire _3370_;
  wire _3371_;
  wire _3372_;
  wire _3373_;
  wire _3374_;
  wire _3375_;
  wire _3376_;
  wire _3377_;
  wire _3378_;
  wire _3379_;
  wire _3380_;
  wire _3381_;
  wire _3382_;
  wire _3383_;
  wire _3384_;
  wire _3385_;
  wire _3386_;
  wire _3387_;
  wire _3388_;
  wire _3389_;
  wire _3390_;
  wire _3391_;
  wire _3392_;
  wire _3393_;
  wire _3394_;
  wire _3395_;
  wire _3396_;
  wire _3397_;
  wire _3398_;
  wire _3399_;
  wire _3400_;
  wire _3401_;
  wire _3402_;
  wire _3403_;
  wire _3404_;
  wire _3405_;
  wire _3406_;
  wire _3407_;
  wire _3408_;
  wire _3409_;
  wire _3410_;
  wire _3411_;
  wire _3412_;
  wire _3413_;
  wire _3414_;
  wire _3415_;
  wire _3416_;
  wire _3417_;
  wire _3418_;
  wire _3419_;
  wire _3420_;
  wire _3421_;
  wire _3422_;
  wire _3423_;
  wire _3424_;
  wire _3425_;
  wire _3426_;
  wire _3427_;
  wire _3428_;
  wire _3429_;
  wire _3430_;
  wire _3431_;
  wire _3432_;
  wire _3433_;
  wire _3434_;
  wire _3435_;
  wire _3436_;
  wire _3437_;
  wire _3438_;
  wire _3439_;
  wire _3440_;
  wire _3441_;
  wire _3442_;
  wire _3443_;
  wire _3444_;
  wire _3445_;
  wire _3446_;
  wire _3447_;
  wire _3448_;
  wire _3449_;
  wire _3450_;
  wire _3451_;
  wire _3452_;
  wire _3453_;
  wire _3454_;
  wire _3455_;
  wire _3456_;
  wire _3457_;
  wire _3458_;
  wire _3459_;
  wire _3460_;
  wire _3461_;
  wire _3462_;
  wire _3463_;
  wire _3464_;
  wire _3465_;
  wire _3466_;
  wire _3467_;
  wire _3468_;
  wire _3469_;
  wire _3470_;
  wire _3471_;
  wire _3472_;
  wire _3473_;
  wire _3474_;
  wire _3475_;
  wire _3476_;
  wire _3477_;
  wire _3478_;
  wire _3479_;
  wire _3480_;
  wire _3481_;
  wire _3482_;
  wire _3483_;
  wire _3484_;
  wire _3485_;
  wire _3486_;
  wire _3487_;
  wire _3488_;
  wire _3489_;
  wire _3490_;
  wire _3491_;
  wire _3492_;
  wire _3493_;
  wire _3494_;
  wire _3495_;
  wire _3496_;
  wire _3497_;
  wire _3498_;
  wire _3499_;
  wire _3500_;
  wire _3501_;
  wire _3502_;
  wire _3503_;
  wire _3504_;
  wire _3505_;
  wire _3506_;
  wire _3507_;
  wire _3508_;
  wire _3509_;
  wire _3510_;
  wire _3511_;
  wire _3512_;
  wire _3513_;
  wire _3514_;
  wire _3515_;
  wire _3516_;
  wire _3517_;
  wire _3518_;
  wire _3519_;
  wire _3520_;
  wire _3521_;
  wire _3522_;
  wire _3523_;
  wire _3524_;
  wire _3525_;
  wire _3526_;
  wire _3527_;
  wire _3528_;
  wire _3529_;
  wire _3530_;
  wire _3531_;
  wire _3532_;
  wire _3533_;
  wire _3534_;
  wire _3535_;
  wire _3536_;
  wire _3537_;
  wire _3538_;
  wire _3539_;
  wire _3540_;
  wire _3541_;
  wire _3542_;
  wire _3543_;
  wire _3544_;
  wire _3545_;
  wire _3546_;
  wire _3547_;
  wire _3548_;
  wire _3549_;
  wire _3550_;
  wire _3551_;
  wire _3552_;
  wire _3553_;
  wire _3554_;
  wire _3555_;
  wire _3556_;
  wire _3557_;
  wire _3558_;
  wire _3559_;
  wire _3560_;
  wire _3561_;
  wire _3562_;
  wire _3563_;
  wire _3564_;
  wire _3565_;
  wire _3566_;
  wire _3567_;
  wire _3568_;
  wire _3569_;
  wire _3570_;
  wire _3571_;
  wire _3572_;
  wire _3573_;
  wire _3574_;
  wire _3575_;
  wire _3576_;
  wire _3577_;
  wire _3578_;
  wire _3579_;
  wire _3580_;
  wire _3581_;
  wire _3582_;
  wire _3583_;
  wire _3584_;
  wire _3585_;
  wire _3586_;
  wire _3587_;
  wire _3588_;
  wire _3589_;
  wire _3590_;
  wire _3591_;
  wire _3592_;
  wire _3593_;
  wire _3594_;
  wire _3595_;
  wire _3596_;
  wire _3597_;
  wire _3598_;
  wire _3599_;
  wire _3600_;
  wire _3601_;
  wire _3602_;
  wire _3603_;
  wire _3604_;
  wire _3605_;
  wire _3606_;
  wire _3607_;
  wire _3608_;
  wire _3609_;
  wire _3610_;
  wire _3611_;
  wire _3612_;
  wire _3613_;
  wire _3614_;
  wire _3615_;
  wire _3616_;
  wire _3617_;
  wire _3618_;
  wire _3619_;
  wire _3620_;
  wire _3621_;
  wire _3622_;
  wire _3623_;
  wire _3624_;
  wire _3625_;
  wire _3626_;
  wire _3627_;
  wire _3628_;
  wire _3629_;
  wire _3630_;
  wire _3631_;
  wire _3632_;
  wire _3633_;
  wire _3634_;
  wire _3635_;
  wire _3636_;
  wire _3637_;
  wire _3638_;
  wire _3639_;
  wire _3640_;
  wire _3641_;
  wire _3642_;
  wire _3643_;
  wire _3644_;
  wire _3645_;
  wire _3646_;
  wire _3647_;
  wire _3648_;
  wire _3649_;
  wire _3650_;
  wire _3651_;
  wire _3652_;
  wire _3653_;
  wire _3654_;
  wire _3655_;
  wire _3656_;
  wire _3657_;
  wire _3658_;
  wire _3659_;
  wire _3660_;
  wire _3661_;
  wire _3662_;
  wire _3663_;
  wire _3664_;
  wire _3665_;
  wire _3666_;
  wire _3667_;
  wire _3668_;
  wire _3669_;
  wire _3670_;
  wire _3671_;
  wire _3672_;
  wire _3673_;
  wire _3674_;
  wire _3675_;
  wire _3676_;
  wire _3677_;
  wire _3678_;
  wire _3679_;
  wire _3680_;
  wire _3681_;
  wire _3682_;
  wire _3683_;
  wire _3684_;
  wire _3685_;
  wire _3686_;
  wire _3687_;
  wire _3688_;
  wire _3689_;
  wire _3690_;
  wire _3691_;
  wire _3692_;
  wire _3693_;
  wire _3694_;
  wire _3695_;
  wire _3696_;
  wire _3697_;
  wire _3698_;
  wire _3699_;
  wire _3700_;
  wire _3701_;
  wire _3702_;
  wire _3703_;
  wire _3704_;
  wire _3705_;
  wire _3706_;
  wire _3707_;
  wire _3708_;
  wire _3709_;
  wire _3710_;
  wire _3711_;
  wire _3712_;
  wire _3713_;
  wire _3714_;
  wire _3715_;
  wire _3716_;
  wire _3717_;
  wire _3718_;
  wire _3719_;
  wire _3720_;
  wire _3721_;
  wire _3722_;
  wire _3723_;
  wire _3724_;
  wire _3725_;
  wire _3726_;
  wire _3727_;
  wire _3728_;
  wire _3729_;
  wire _3730_;
  wire _3731_;
  wire _3732_;
  wire _3733_;
  wire _3734_;
  wire _3735_;
  wire _3736_;
  wire _3737_;
  wire _3738_;
  wire _3739_;
  wire _3740_;
  wire _3741_;
  wire _3742_;
  wire _3743_;
  wire _3744_;
  wire _3745_;
  wire _3746_;
  wire _3747_;
  wire _3748_;
  wire _3749_;
  wire _3750_;
  wire _3751_;
  wire _3752_;
  wire _3753_;
  wire _3754_;
  wire _3755_;
  wire _3756_;
  wire _3757_;
  wire _3758_;
  wire _3759_;
  wire _3760_;
  wire _3761_;
  wire _3762_;
  wire _3763_;
  wire _3764_;
  wire _3765_;
  wire _3766_;
  wire _3767_;
  wire _3768_;
  wire _3769_;
  wire _3770_;
  wire _3771_;
  wire _3772_;
  wire _3773_;
  wire _3774_;
  wire _3775_;
  wire _3776_;
  wire _3777_;
  wire _3778_;
  wire _3779_;
  wire _3780_;
  wire _3781_;
  wire _3782_;
  wire _3783_;
  wire _3784_;
  wire _3785_;
  wire _3786_;
  wire _3787_;
  wire _3788_;
  wire _3789_;
  wire _3790_;
  wire _3791_;
  wire _3792_;
  wire _3793_;
  wire _3794_;
  wire _3795_;
  wire _3796_;
  wire _3797_;
  wire _3798_;
  wire _3799_;
  wire _3800_;
  wire _3801_;
  wire _3802_;
  wire _3803_;
  wire _3804_;
  wire _3805_;
  wire _3806_;
  wire _3807_;
  wire _3808_;
  wire _3809_;
  wire _3810_;
  wire _3811_;
  wire _3812_;
  wire _3813_;
  wire _3814_;
  wire _3815_;
  wire _3816_;
  wire _3817_;
  wire _3818_;
  wire _3819_;
  wire _3820_;
  wire _3821_;
  wire _3822_;
  wire _3823_;
  wire _3824_;
  wire _3825_;
  wire _3826_;
  wire _3827_;
  wire _3828_;
  wire _3829_;
  wire _3830_;
  wire _3831_;
  wire _3832_;
  wire _3833_;
  wire _3834_;
  wire _3835_;
  wire _3836_;
  wire _3837_;
  wire _3838_;
  wire _3839_;
  wire _3840_;
  wire _3841_;
  wire _3842_;
  wire _3843_;
  wire _3844_;
  wire _3845_;
  wire _3846_;
  wire _3847_;
  wire _3848_;
  wire _3849_;
  wire _3850_;
  wire _3851_;
  wire _3852_;
  wire _3853_;
  wire _3854_;
  wire _3855_;
  wire _3856_;
  wire _3857_;
  wire _3858_;
  wire _3859_;
  wire _3860_;
  wire _3861_;
  wire _3862_;
  wire _3863_;
  wire _3864_;
  wire _3865_;
  wire _3866_;
  wire _3867_;
  wire _3868_;
  wire _3869_;
  wire _3870_;
  wire _3871_;
  wire _3872_;
  wire _3873_;
  wire _3874_;
  wire _3875_;
  wire _3876_;
  wire _3877_;
  wire _3878_;
  wire _3879_;
  wire _3880_;
  wire _3881_;
  wire _3882_;
  wire _3883_;
  wire _3884_;
  wire _3885_;
  wire _3886_;
  wire _3887_;
  wire _3888_;
  wire _3889_;
  wire _3890_;
  wire _3891_;
  wire _3892_;
  wire _3893_;
  wire _3894_;
  wire _3895_;
  wire _3896_;
  wire _3897_;
  wire _3898_;
  wire _3899_;
  wire _3900_;
  wire _3901_;
  wire _3902_;
  wire _3903_;
  wire _3904_;
  wire _3905_;
  wire _3906_;
  wire _3907_;
  wire _3908_;
  wire _3909_;
  wire _3910_;
  wire _3911_;
  wire _3912_;
  wire _3913_;
  wire _3914_;
  wire _3915_;
  wire _3916_;
  wire _3917_;
  wire _3918_;
  wire _3919_;
  wire _3920_;
  wire _3921_;
  wire _3922_;
  wire _3923_;
  wire _3924_;
  wire _3925_;
  wire _3926_;
  wire _3927_;
  wire _3928_;
  wire _3929_;
  wire _3930_;
  wire _3931_;
  wire _3932_;
  wire _3933_;
  wire _3934_;
  wire _3935_;
  wire _3936_;
  wire _3937_;
  wire _3938_;
  wire _3939_;
  wire _3940_;
  wire _3941_;
  wire _3942_;
  wire _3943_;
  wire _3944_;
  wire _3945_;
  wire _3946_;
  wire _3947_;
  wire _3948_;
  wire _3949_;
  wire _3950_;
  wire _3951_;
  wire _3952_;
  wire _3953_;
  wire _3954_;
  wire _3955_;
  wire _3956_;
  wire _3957_;
  wire _3958_;
  wire _3959_;
  wire _3960_;
  wire _3961_;
  wire _3962_;
  wire _3963_;
  wire _3964_;
  wire _3965_;
  wire _3966_;
  wire _3967_;
  wire _3968_;
  wire _3969_;
  wire _3970_;
  wire _3971_;
  wire _3972_;
  wire _3973_;
  wire _3974_;
  wire _3975_;
  wire _3976_;
  wire _3977_;
  wire _3978_;
  wire _3979_;
  wire _3980_;
  wire _3981_;
  wire _3982_;
  wire _3983_;
  wire _3984_;
  wire _3985_;
  wire _3986_;
  wire _3987_;
  wire _3988_;
  wire _3989_;
  wire _3990_;
  wire _3991_;
  wire _3992_;
  wire _3993_;
  wire _3994_;
  wire _3995_;
  wire _3996_;
  wire _3997_;
  wire _3998_;
  wire _3999_;
  wire _4000_;
  wire _4001_;
  wire _4002_;
  wire _4003_;
  wire _4004_;
  wire _4005_;
  wire _4006_;
  wire _4007_;
  wire _4008_;
  wire _4009_;
  wire _4010_;
  wire _4011_;
  wire _4012_;
  wire _4013_;
  wire _4014_;
  wire _4015_;
  wire _4016_;
  wire _4017_;
  wire _4018_;
  wire _4019_;
  wire _4020_;
  wire _4021_;
  wire _4022_;
  wire _4023_;
  wire _4024_;
  wire _4025_;
  wire _4026_;
  wire _4027_;
  wire _4028_;
  wire _4029_;
  wire _4030_;
  wire _4031_;
  wire _4032_;
  wire _4033_;
  wire _4034_;
  wire _4035_;
  wire _4036_;
  wire _4037_;
  wire _4038_;
  wire _4039_;
  wire _4040_;
  wire _4041_;
  wire _4042_;
  wire _4043_;
  wire _4044_;
  wire _4045_;
  wire _4046_;
  wire _4047_;
  wire _4048_;
  wire _4049_;
  wire _4050_;
  wire _4051_;
  wire _4052_;
  wire _4053_;
  wire _4054_;
  wire _4055_;
  wire _4056_;
  wire _4057_;
  wire _4058_;
  wire _4059_;
  wire _4060_;
  wire _4061_;
  wire _4062_;
  wire _4063_;
  wire _4064_;
  wire _4065_;
  wire _4066_;
  wire _4067_;
  wire _4068_;
  wire _4069_;
  wire _4070_;
  wire _4071_;
  wire _4072_;
  wire _4073_;
  wire _4074_;
  wire _4075_;
  wire _4076_;
  wire _4077_;
  wire _4078_;
  wire _4079_;
  wire _4080_;
  wire _4081_;
  wire _4082_;
  wire _4083_;
  wire _4084_;
  wire _4085_;
  wire _4086_;
  wire _4087_;
  wire _4088_;
  wire _4089_;
  wire _4090_;
  wire _4091_;
  wire _4092_;
  wire _4093_;
  wire _4094_;
  wire _4095_;
  wire _4096_;
  wire _4097_;
  wire _4098_;
  wire _4099_;
  wire _4100_;
  wire _4101_;
  wire _4102_;
  wire _4103_;
  wire _4104_;
  wire _4105_;
  wire _4106_;
  wire _4107_;
  wire _4108_;
  wire _4109_;
  wire _4110_;
  wire _4111_;
  wire _4112_;
  wire _4113_;
  wire _4114_;
  wire _4115_;
  wire _4116_;
  wire _4117_;
  wire _4118_;
  wire _4119_;
  wire _4120_;
  wire _4121_;
  wire _4122_;
  wire _4123_;
  wire _4124_;
  wire _4125_;
  wire _4126_;
  wire _4127_;
  wire _4128_;
  wire _4129_;
  wire _4130_;
  wire _4131_;
  wire _4132_;
  wire _4133_;
  wire _4134_;
  wire _4135_;
  wire _4136_;
  wire _4137_;
  wire _4138_;
  wire _4139_;
  wire _4140_;
  wire _4141_;
  wire _4142_;
  wire _4143_;
  wire _4144_;
  wire _4145_;
  wire _4146_;
  wire _4147_;
  wire _4148_;
  wire _4149_;
  wire _4150_;
  wire _4151_;
  wire _4152_;
  wire _4153_;
  wire _4154_;
  wire _4155_;
  wire _4156_;
  wire _4157_;
  wire _4158_;
  wire _4159_;
  wire _4160_;
  wire _4161_;
  wire _4162_;
  wire _4163_;
  wire _4164_;
  wire _4165_;
  wire _4166_;
  wire _4167_;
  wire _4168_;
  wire _4169_;
  wire _4170_;
  wire _4171_;
  wire _4172_;
  wire _4173_;
  wire _4174_;
  wire _4175_;
  wire _4176_;
  wire _4177_;
  wire _4178_;
  wire _4179_;
  wire _4180_;
  wire _4181_;
  wire _4182_;
  wire _4183_;
  wire _4184_;
  wire _4185_;
  wire _4186_;
  wire _4187_;
  wire _4188_;
  wire _4189_;
  wire _4190_;
  wire _4191_;
  wire _4192_;
  wire _4193_;
  wire _4194_;
  wire _4195_;
  wire _4196_;
  wire _4197_;
  wire _4198_;
  wire _4199_;
  wire _4200_;
  wire _4201_;
  wire _4202_;
  wire _4203_;
  wire _4204_;
  wire _4205_;
  wire _4206_;
  wire _4207_;
  wire _4208_;
  wire _4209_;
  wire _4210_;
  wire _4211_;
  wire _4212_;
  wire _4213_;
  wire _4214_;
  wire _4215_;
  wire _4216_;
  wire _4217_;
  wire _4218_;
  wire _4219_;
  wire _4220_;
  wire _4221_;
  wire _4222_;
  wire _4223_;
  wire _4224_;
  wire _4225_;
  wire _4226_;
  wire _4227_;
  wire _4228_;
  wire _4229_;
  wire _4230_;
  wire _4231_;
  wire _4232_;
  wire _4233_;
  wire _4234_;
  wire _4235_;
  wire _4236_;
  wire _4237_;
  wire _4238_;
  wire _4239_;
  wire _4240_;
  wire _4241_;
  wire _4242_;
  wire _4243_;
  wire _4244_;
  wire _4245_;
  wire _4246_;
  wire _4247_;
  wire _4248_;
  wire _4249_;
  wire _4250_;
  wire _4251_;
  wire _4252_;
  wire _4253_;
  wire _4254_;
  wire _4255_;
  wire _4256_;
  wire _4257_;
  wire _4258_;
  wire _4259_;
  wire _4260_;
  wire _4261_;
  wire _4262_;
  wire _4263_;
  wire _4264_;
  wire _4265_;
  wire _4266_;
  wire _4267_;
  wire _4268_;
  wire _4269_;
  wire _4270_;
  wire _4271_;
  wire _4272_;
  wire _4273_;
  wire _4274_;
  wire _4275_;
  wire _4276_;
  wire _4277_;
  wire _4278_;
  wire _4279_;
  wire _4280_;
  wire _4281_;
  wire _4282_;
  wire _4283_;
  wire _4284_;
  wire _4285_;
  wire _4286_;
  wire _4287_;
  wire _4288_;
  wire _4289_;
  wire _4290_;
  wire _4291_;
  wire _4292_;
  wire _4293_;
  wire _4294_;
  wire _4295_;
  wire _4296_;
  wire _4297_;
  wire _4298_;
  wire _4299_;
  wire _4300_;
  wire _4301_;
  wire _4302_;
  wire _4303_;
  wire _4304_;
  wire _4305_;
  wire _4306_;
  wire _4307_;
  wire _4308_;
  wire _4309_;
  wire _4310_;
  wire _4311_;
  wire _4312_;
  wire _4313_;
  wire _4314_;
  wire _4315_;
  wire _4316_;
  wire _4317_;
  wire _4318_;
  wire _4319_;
  wire _4320_;
  wire _4321_;
  wire _4322_;
  wire _4323_;
  wire _4324_;
  wire _4325_;
  wire _4326_;
  wire _4327_;
  wire _4328_;
  wire _4329_;
  wire _4330_;
  wire _4331_;
  wire _4332_;
  wire _4333_;
  wire _4334_;
  wire _4335_;
  wire _4336_;
  wire _4337_;
  wire _4338_;
  wire _4339_;
  wire _4340_;
  wire _4341_;
  wire _4342_;
  wire _4343_;
  wire _4344_;
  wire _4345_;
  wire _4346_;
  wire _4347_;
  wire _4348_;
  wire _4349_;
  wire _4350_;
  wire _4351_;
  wire _4352_;
  wire _4353_;
  wire _4354_;
  wire _4355_;
  wire _4356_;
  wire _4357_;
  wire _4358_;
  wire _4359_;
  wire _4360_;
  wire _4361_;
  wire _4362_;
  wire _4363_;
  wire _4364_;
  wire _4365_;
  wire _4366_;
  wire _4367_;
  wire _4368_;
  wire _4369_;
  wire _4370_;
  wire _4371_;
  wire _4372_;
  wire _4373_;
  wire _4374_;
  wire _4375_;
  wire _4376_;
  wire _4377_;
  wire _4378_;
  wire _4379_;
  wire _4380_;
  wire _4381_;
  wire _4382_;
  wire _4383_;
  wire _4384_;
  wire _4385_;
  wire _4386_;
  wire _4387_;
  wire _4388_;
  wire _4389_;
  wire _4390_;
  wire _4391_;
  wire _4392_;
  wire _4393_;
  wire _4394_;
  wire _4395_;
  wire _4396_;
  wire _4397_;
  wire _4398_;
  wire _4399_;
  wire _4400_;
  wire _4401_;
  wire _4402_;
  wire _4403_;
  wire _4404_;
  wire _4405_;
  wire _4406_;
  wire _4407_;
  wire _4408_;
  wire _4409_;
  wire _4410_;
  wire _4411_;
  wire _4412_;
  wire _4413_;
  wire _4414_;
  wire _4415_;
  wire _4416_;
  wire _4417_;
  wire _4418_;
  wire _4419_;
  wire _4420_;
  wire _4421_;
  wire _4422_;
  wire _4423_;
  wire _4424_;
  wire _4425_;
  wire _4426_;
  wire _4427_;
  wire _4428_;
  wire _4429_;
  wire _4430_;
  wire _4431_;
  wire _4432_;
  wire _4433_;
  wire _4434_;
  wire _4435_;
  wire _4436_;
  wire _4437_;
  wire _4438_;
  wire _4439_;
  wire _4440_;
  wire _4441_;
  wire _4442_;
  wire _4443_;
  wire _4444_;
  wire _4445_;
  wire _4446_;
  wire _4447_;
  wire _4448_;
  wire _4449_;
  wire _4450_;
  wire _4451_;
  wire _4452_;
  wire _4453_;
  wire _4454_;
  wire _4455_;
  wire _4456_;
  wire _4457_;
  wire _4458_;
  wire _4459_;
  wire _4460_;
  wire _4461_;
  wire _4462_;
  wire _4463_;
  wire _4464_;
  wire _4465_;
  wire _4466_;
  wire _4467_;
  wire _4468_;
  wire _4469_;
  wire _4470_;
  wire _4471_;
  wire _4472_;
  wire _4473_;
  wire _4474_;
  wire _4475_;
  wire _4476_;
  wire _4477_;
  wire _4478_;
  wire _4479_;
  wire _4480_;
  wire _4481_;
  wire _4482_;
  wire _4483_;
  wire _4484_;
  wire _4485_;
  wire _4486_;
  wire _4487_;
  wire _4488_;
  wire _4489_;
  wire _4490_;
  wire _4491_;
  wire _4492_;
  wire _4493_;
  wire _4494_;
  wire _4495_;
  wire _4496_;
  wire _4497_;
  wire _4498_;
  wire _4499_;
  wire _4500_;
  wire _4501_;
  wire _4502_;
  wire _4503_;
  wire _4504_;
  wire _4505_;
  wire _4506_;
  wire _4507_;
  wire _4508_;
  wire _4509_;
  wire _4510_;
  wire _4511_;
  wire _4512_;
  wire _4513_;
  wire _4514_;
  wire _4515_;
  wire _4516_;
  wire _4517_;
  wire _4518_;
  wire _4519_;
  wire _4520_;
  wire _4521_;
  wire _4522_;
  wire _4523_;
  wire _4524_;
  wire _4525_;
  wire _4526_;
  wire _4527_;
  wire _4528_;
  wire _4529_;
  wire _4530_;
  wire _4531_;
  wire _4532_;
  wire _4533_;
  wire _4534_;
  wire _4535_;
  wire _4536_;
  wire _4537_;
  wire _4538_;
  wire _4539_;
  wire _4540_;
  wire _4541_;
  wire _4542_;
  wire _4543_;
  wire _4544_;
  wire _4545_;
  wire _4546_;
  wire _4547_;
  wire _4548_;
  wire _4549_;
  wire _4550_;
  wire _4551_;
  wire _4552_;
  wire _4553_;
  wire _4554_;
  wire _4555_;
  wire _4556_;
  wire _4557_;
  wire _4558_;
  wire _4559_;
  wire _4560_;
  wire _4561_;
  wire _4562_;
  wire _4563_;
  wire _4564_;
  wire _4565_;
  wire _4566_;
  wire _4567_;
  wire _4568_;
  wire _4569_;
  wire _4570_;
  wire _4571_;
  wire _4572_;
  wire _4573_;
  wire _4574_;
  wire _4575_;
  wire _4576_;
  wire _4577_;
  wire _4578_;
  wire _4579_;
  wire _4580_;
  wire _4581_;
  wire _4582_;
  wire _4583_;
  wire _4584_;
  wire _4585_;
  wire _4586_;
  wire _4587_;
  wire _4588_;
  wire _4589_;
  wire _4590_;
  wire _4591_;
  wire _4592_;
  wire _4593_;
  wire _4594_;
  wire _4595_;
  wire _4596_;
  wire _4597_;
  wire _4598_;
  wire _4599_;
  wire _4600_;
  wire _4601_;
  wire _4602_;
  wire _4603_;
  wire _4604_;
  wire _4605_;
  wire _4606_;
  wire _4607_;
  wire _4608_;
  wire _4609_;
  wire _4610_;
  wire _4611_;
  wire _4612_;
  wire _4613_;
  wire _4614_;
  wire _4615_;
  wire _4616_;
  wire _4617_;
  wire _4618_;
  wire _4619_;
  wire _4620_;
  wire _4621_;
  wire _4622_;
  wire _4623_;
  wire _4624_;
  wire _4625_;
  wire _4626_;
  wire _4627_;
  wire _4628_;
  wire _4629_;
  wire _4630_;
  wire _4631_;
  wire _4632_;
  wire _4633_;
  wire _4634_;
  wire _4635_;
  wire _4636_;
  wire _4637_;
  wire _4638_;
  wire _4639_;
  wire _4640_;
  wire _4641_;
  wire _4642_;
  wire _4643_;
  wire _4644_;
  wire _4645_;
  wire _4646_;
  wire _4647_;
  wire _4648_;
  wire _4649_;
  wire _4650_;
  wire _4651_;
  wire _4652_;
  wire _4653_;
  wire _4654_;
  wire _4655_;
  wire _4656_;
  wire _4657_;
  wire _4658_;
  wire _4659_;
  wire _4660_;
  wire _4661_;
  wire _4662_;
  wire _4663_;
  wire _4664_;
  wire _4665_;
  wire _4666_;
  wire _4667_;
  wire _4668_;
  wire _4669_;
  wire _4670_;
  wire _4671_;
  wire _4672_;
  wire _4673_;
  wire _4674_;
  wire _4675_;
  wire _4676_;
  wire _4677_;
  wire _4678_;
  wire _4679_;
  wire _4680_;
  wire _4681_;
  wire _4682_;
  wire _4683_;
  wire _4684_;
  wire _4685_;
  wire _4686_;
  wire _4687_;
  wire _4688_;
  wire _4689_;
  wire _4690_;
  wire _4691_;
  wire _4692_;
  wire _4693_;
  wire _4694_;
  wire _4695_;
  wire _4696_;
  wire _4697_;
  wire _4698_;
  wire _4699_;
  wire _4700_;
  wire _4701_;
  wire _4702_;
  wire _4703_;
  wire _4704_;
  wire _4705_;
  wire _4706_;
  wire _4707_;
  wire _4708_;
  wire _4709_;
  wire _4710_;
  wire _4711_;
  wire _4712_;
  wire _4713_;
  wire _4714_;
  wire _4715_;
  wire _4716_;
  wire _4717_;
  wire _4718_;
  wire _4719_;
  wire _4720_;
  wire _4721_;
  wire _4722_;
  wire _4723_;
  wire _4724_;
  wire _4725_;
  wire _4726_;
  wire _4727_;
  wire _4728_;
  wire _4729_;
  wire _4730_;
  wire _4731_;
  wire _4732_;
  wire _4733_;
  wire _4734_;
  wire _4735_;
  wire _4736_;
  wire _4737_;
  wire _4738_;
  wire _4739_;
  wire _4740_;
  wire _4741_;
  wire _4742_;
  wire _4743_;
  wire _4744_;
  wire _4745_;
  wire _4746_;
  wire _4747_;
  wire _4748_;
  wire _4749_;
  wire _4750_;
  wire _4751_;
  wire _4752_;
  wire _4753_;
  wire _4754_;
  wire _4755_;
  wire _4756_;
  wire _4757_;
  wire _4758_;
  wire _4759_;
  wire _4760_;
  wire _4761_;
  wire _4762_;
  wire _4763_;
  wire _4764_;
  wire _4765_;
  wire _4766_;
  wire _4767_;
  wire _4768_;
  wire _4769_;
  wire _4770_;
  wire _4771_;
  wire _4772_;
  wire _4773_;
  wire _4774_;
  wire _4775_;
  wire [32:0] _4776_;
  wire [65:0] _GEN_0;
  wire [65:0] _GEN_2;
  wire [41:0] _GEN_35;
  wire [5:0] _count_T_1;
  wire [1:0] _decoded_T_4;
  wire _decoded_T_6;
  wire [1:0] _decoded_T_7;
  wire [1:0] _decoded_orMatrixOutputs_T_4;
  wire [32:0] _divisor_T;
  wire _eOut_T_4;
  wire [8:0] _prod_T_2;
  wire [65:0] _remainder_T_2;
  wire [2:0] _state_T;
  wire [32:0] accum;
  input clock;
  wire clock;
  wire [5:0] count;
  wire decoded_andMatrixInput_0_3;
  wire decoded_andMatrixInput_0_4;
  wire decoded_andMatrixInput_1_2;
  wire [2:0] decoded_plaInput;
  wire [32:0] divisor;
  wire [15:0] hi;
  wire [15:0] hi_1;
  input io_kill;
  wire io_kill;
  input [3:0] io_req_bits_fn;
  wire [3:0] io_req_bits_fn;
  input [31:0] io_req_bits_in1;
  wire [31:0] io_req_bits_in1;
  input [31:0] io_req_bits_in2;
  wire [31:0] io_req_bits_in2;
  input [4:0] io_req_bits_tag;
  wire [4:0] io_req_bits_tag;
  output io_req_ready;
  wire io_req_ready;
  input io_req_valid;
  wire io_req_valid;
  output [31:0] io_resp_bits_data;
  wire [31:0] io_resp_bits_data;
  output [4:0] io_resp_bits_tag;
  wire [4:0] io_resp_bits_tag;
  input io_resp_ready;
  wire io_resp_ready;
  output io_resp_valid;
  wire io_resp_valid;
  wire isHi;
  wire [31:0] lhs_in;
  wire [15:0] loOut;
  wire [31:0] mplier;
  wire mplierSign;
  wire [64:0] mulReg;
  wire neg_out;
  wire [31:0] negated_remainder;
  wire nextMplierSign;
  wire [65:0] nextMulReg;
  wire [64:0] nextMulReg1;
  wire [41:0] nextMulReg_hi;
  wire [65:0] remainder;
  wire [4:0] req_tag;
  wire resHi;
  input reset;
  wire reset;
  wire [31:0] result;
  wire rhs_sign;
  wire [2:0] state;
  wire [64:0] unrolls_0;
  INV_X1 _4777_ (
    .A(remainder[65]),
    .ZN(_2936_)
  );
  INV_X1 _4778_ (
    .A(remainder[64]),
    .ZN(_2947_)
  );
  INV_X1 _4779_ (
    .A(remainder[62]),
    .ZN(_2958_)
  );
  INV_X1 _4780_ (
    .A(remainder[61]),
    .ZN(_2969_)
  );
  INV_X1 _4781_ (
    .A(remainder[60]),
    .ZN(_2980_)
  );
  INV_X1 _4782_ (
    .A(remainder[59]),
    .ZN(_2991_)
  );
  INV_X1 _4783_ (
    .A(remainder[58]),
    .ZN(_3002_)
  );
  INV_X1 _4784_ (
    .A(remainder[57]),
    .ZN(_3013_)
  );
  INV_X1 _4785_ (
    .A(remainder[55]),
    .ZN(_3023_)
  );
  INV_X1 _4786_ (
    .A(remainder[54]),
    .ZN(_3034_)
  );
  INV_X1 _4787_ (
    .A(remainder[52]),
    .ZN(_3045_)
  );
  INV_X1 _4788_ (
    .A(remainder[50]),
    .ZN(_3056_)
  );
  INV_X1 _4789_ (
    .A(remainder[49]),
    .ZN(_3067_)
  );
  INV_X1 _4790_ (
    .A(remainder[48]),
    .ZN(_3078_)
  );
  INV_X1 _4791_ (
    .A(remainder[47]),
    .ZN(_3089_)
  );
  INV_X1 _4792_ (
    .A(remainder[46]),
    .ZN(_3100_)
  );
  INV_X1 _4793_ (
    .A(remainder[45]),
    .ZN(_3111_)
  );
  INV_X1 _4794_ (
    .A(remainder[44]),
    .ZN(_3122_)
  );
  INV_X1 _4795_ (
    .A(remainder[43]),
    .ZN(_3133_)
  );
  INV_X1 _4796_ (
    .A(remainder[42]),
    .ZN(_3144_)
  );
  INV_X1 _4797_ (
    .A(remainder[41]),
    .ZN(_3155_)
  );
  INV_X1 _4798_ (
    .A(remainder[40]),
    .ZN(_3165_)
  );
  INV_X1 _4799_ (
    .A(remainder[39]),
    .ZN(_3176_)
  );
  INV_X1 _4800_ (
    .A(remainder[37]),
    .ZN(_3187_)
  );
  INV_X1 _4801_ (
    .A(remainder[36]),
    .ZN(_3198_)
  );
  INV_X1 _4802_ (
    .A(remainder[32]),
    .ZN(_3209_)
  );
  INV_X1 _4803_ (
    .A(count[2]),
    .ZN(_3220_)
  );
  INV_X1 _4804_ (
    .A(count[1]),
    .ZN(_3231_)
  );
  INV_X1 _4805_ (
    .A(count[0]),
    .ZN(_3242_)
  );
  INV_X1 _4806_ (
    .A(reset),
    .ZN(_3253_)
  );
  INV_X1 _4807_ (
    .A(divisor[3]),
    .ZN(_3264_)
  );
  INV_X1 _4808_ (
    .A(divisor[5]),
    .ZN(_3274_)
  );
  INV_X1 _4809_ (
    .A(divisor[7]),
    .ZN(_3285_)
  );
  INV_X1 _4810_ (
    .A(divisor[8]),
    .ZN(_3296_)
  );
  INV_X1 _4811_ (
    .A(divisor[10]),
    .ZN(_3307_)
  );
  INV_X1 _4812_ (
    .A(divisor[11]),
    .ZN(_3318_)
  );
  INV_X1 _4813_ (
    .A(divisor[14]),
    .ZN(_3329_)
  );
  INV_X1 _4814_ (
    .A(divisor[16]),
    .ZN(_3340_)
  );
  INV_X1 _4815_ (
    .A(divisor[17]),
    .ZN(_3351_)
  );
  INV_X1 _4816_ (
    .A(divisor[19]),
    .ZN(_3362_)
  );
  INV_X1 _4817_ (
    .A(divisor[20]),
    .ZN(_3373_)
  );
  INV_X1 _4818_ (
    .A(divisor[23]),
    .ZN(_3384_)
  );
  INV_X1 _4819_ (
    .A(divisor[25]),
    .ZN(_3394_)
  );
  INV_X1 _4820_ (
    .A(divisor[26]),
    .ZN(_3405_)
  );
  INV_X1 _4821_ (
    .A(divisor[28]),
    .ZN(_3416_)
  );
  INV_X1 _4822_ (
    .A(divisor[29]),
    .ZN(_3427_)
  );
  INV_X1 _4823_ (
    .A(divisor[31]),
    .ZN(_3438_)
  );
  INV_X1 _4824_ (
    .A(remainder[1]),
    .ZN(_3449_)
  );
  INV_X1 _4825_ (
    .A(remainder[2]),
    .ZN(_3460_)
  );
  INV_X1 _4826_ (
    .A(remainder[4]),
    .ZN(_3471_)
  );
  INV_X1 _4827_ (
    .A(remainder[6]),
    .ZN(_3482_)
  );
  INV_X1 _4828_ (
    .A(remainder[24]),
    .ZN(_3493_)
  );
  INV_X1 _4829_ (
    .A(remainder[31]),
    .ZN(_3504_)
  );
  INV_X1 _4830_ (
    .A(state[2]),
    .ZN(_3514_)
  );
  INV_X1 _4831_ (
    .A(io_req_bits_fn[2]),
    .ZN(_3525_)
  );
  INV_X1 _4832_ (
    .A(_0000_),
    .ZN(_3536_)
  );
  INV_X1 _4833_ (
    .A(io_req_bits_in2[31]),
    .ZN(_3547_)
  );
  INV_X1 _4834_ (
    .A(io_req_bits_in1[31]),
    .ZN(_3558_)
  );
  INV_X1 _4835_ (
    .A(io_resp_ready),
    .ZN(_3569_)
  );
  INV_X1 _4836_ (
    .A(io_req_valid),
    .ZN(_3580_)
  );
  INV_X1 _4837_ (
    .A(io_kill),
    .ZN(_3591_)
  );
  INV_X1 _4838_ (
    .A(_eOut_T_4),
    .ZN(_3602_)
  );
  OR2_X1 _4839_ (
    .A1(count[3]),
    .A2(count[2]),
    .ZN(_3613_)
  );
  OR2_X1 _4840_ (
    .A1(count[1]),
    .A2(count[0]),
    .ZN(_3624_)
  );
  OR2_X1 _4841_ (
    .A1(_3613_),
    .A2(_3624_),
    .ZN(_3634_)
  );
  INV_X1 _4842_ (
    .A(_3634_),
    .ZN(_3645_)
  );
  OR2_X1 _4843_ (
    .A1(_0004_),
    .A2(_0003_),
    .ZN(_3656_)
  );
  INV_X1 _4844_ (
    .A(_3656_),
    .ZN(_3667_)
  );
  AND2_X1 _4845_ (
    .A1(_3514_),
    .A2(_3667_),
    .ZN(_3678_)
  );
  OR2_X1 _4846_ (
    .A1(state[2]),
    .A2(_3656_),
    .ZN(_3689_)
  );
  OR2_X1 _4847_ (
    .A1(count[4]),
    .A2(_0001_),
    .ZN(_3700_)
  );
  OR2_X1 _4848_ (
    .A1(_3689_),
    .A2(_3700_),
    .ZN(_3711_)
  );
  INV_X1 _4849_ (
    .A(_3711_),
    .ZN(_3722_)
  );
  AND2_X1 _4850_ (
    .A1(_3645_),
    .A2(_3722_),
    .ZN(_3733_)
  );
  INV_X1 _4851_ (
    .A(_3733_),
    .ZN(_3744_)
  );
  OR2_X1 _4852_ (
    .A1(count[5]),
    .A2(count[4]),
    .ZN(_3754_)
  );
  OR2_X1 _4853_ (
    .A1(_3613_),
    .A2(_3754_),
    .ZN(_3765_)
  );
  OR2_X1 _4854_ (
    .A1(_0002_),
    .A2(_3765_),
    .ZN(_3776_)
  );
  INV_X1 _4855_ (
    .A(_3776_),
    .ZN(_3787_)
  );
  OR2_X1 _4856_ (
    .A1(state[0]),
    .A2(_0003_),
    .ZN(_3798_)
  );
  INV_X1 _4857_ (
    .A(_3798_),
    .ZN(_3809_)
  );
  AND2_X1 _4858_ (
    .A1(_3514_),
    .A2(_3809_),
    .ZN(_3819_)
  );
  OR2_X1 _4859_ (
    .A1(state[2]),
    .A2(_3798_),
    .ZN(_3829_)
  );
  OR2_X1 _4860_ (
    .A1(_count_T_1[0]),
    .A2(_3829_),
    .ZN(_3838_)
  );
  OR2_X1 _4861_ (
    .A1(_3776_),
    .A2(_3838_),
    .ZN(_3847_)
  );
  INV_X1 _4862_ (
    .A(_3847_),
    .ZN(_3856_)
  );
  OR2_X1 _4863_ (
    .A1(_3733_),
    .A2(_3856_),
    .ZN(_3865_)
  );
  OR2_X1 _4864_ (
    .A1(state[1]),
    .A2(state[2]),
    .ZN(_3875_)
  );
  OR2_X1 _4865_ (
    .A1(state[0]),
    .A2(_3875_),
    .ZN(_3884_)
  );
  INV_X1 _4866_ (
    .A(_3884_),
    .ZN(io_req_ready)
  );
  AND2_X1 _4867_ (
    .A1(io_req_valid),
    .A2(io_req_ready),
    .ZN(_3902_)
  );
  OR2_X1 _4868_ (
    .A1(_3580_),
    .A2(_3884_),
    .ZN(_3911_)
  );
  AND2_X1 _4869_ (
    .A1(isHi),
    .A2(_3911_),
    .ZN(_3921_)
  );
  AND2_X1 _4870_ (
    .A1(resHi),
    .A2(_3911_),
    .ZN(_3931_)
  );
  OR2_X1 _4871_ (
    .A1(state[1]),
    .A2(_0004_),
    .ZN(_3940_)
  );
  INV_X1 _4872_ (
    .A(_3940_),
    .ZN(_3949_)
  );
  AND2_X1 _4873_ (
    .A1(_3536_),
    .A2(_3949_),
    .ZN(_3960_)
  );
  OR2_X1 _4874_ (
    .A1(_0000_),
    .A2(_3940_),
    .ZN(_3969_)
  );
  OR2_X1 _4875_ (
    .A1(_3865_),
    .A2(_3960_),
    .ZN(_3978_)
  );
  AND2_X1 _4876_ (
    .A1(_3931_),
    .A2(_3969_),
    .ZN(_3988_)
  );
  MUX2_X1 _4877_ (
    .A(_3988_),
    .B(_3921_),
    .S(_3865_),
    .Z(_0005_)
  );
  OR2_X1 _4878_ (
    .A1(state[2]),
    .A2(_3940_),
    .ZN(_4006_)
  );
  INV_X1 _4879_ (
    .A(_4006_),
    .ZN(_4015_)
  );
  OR2_X1 _4880_ (
    .A1(_3960_),
    .A2(_4015_),
    .ZN(_4026_)
  );
  OR2_X1 _4881_ (
    .A1(state[0]),
    .A2(_4026_),
    .ZN(_4035_)
  );
  AND2_X1 _4882_ (
    .A1(_3847_),
    .A2(_4035_),
    .ZN(_4044_)
  );
  OR2_X1 _4883_ (
    .A1(_3733_),
    .A2(_4044_),
    .ZN(_4054_)
  );
  AND2_X1 _4884_ (
    .A1(_3656_),
    .A2(_3798_),
    .ZN(_4064_)
  );
  OR2_X1 _4885_ (
    .A1(_0000_),
    .A2(_4064_),
    .ZN(_4073_)
  );
  INV_X1 _4886_ (
    .A(_4073_),
    .ZN(io_resp_valid)
  );
  OR2_X1 _4887_ (
    .A1(_3569_),
    .A2(_4073_),
    .ZN(_4092_)
  );
  AND2_X1 _4888_ (
    .A1(_3591_),
    .A2(_4092_),
    .ZN(_4101_)
  );
  AND2_X1 _4889_ (
    .A1(_3911_),
    .A2(_4101_),
    .ZN(_4110_)
  );
  AND2_X1 _4890_ (
    .A1(_4054_),
    .A2(_4110_),
    .ZN(_4121_)
  );
  AND2_X1 _4891_ (
    .A1(io_req_bits_fn[2]),
    .A2(_3902_),
    .ZN(_4130_)
  );
  INV_X1 _4892_ (
    .A(_4130_),
    .ZN(_4140_)
  );
  OR2_X1 _4893_ (
    .A1(_4121_),
    .A2(_4130_),
    .ZN(_4150_)
  );
  AND2_X1 _4894_ (
    .A1(_3253_),
    .A2(_4150_),
    .ZN(_0006_)
  );
  OR2_X1 _4895_ (
    .A1(state[1]),
    .A2(_4026_),
    .ZN(_4169_)
  );
  OR2_X1 _4896_ (
    .A1(_3865_),
    .A2(_4169_),
    .ZN(_4178_)
  );
  OR2_X1 _4897_ (
    .A1(_state_T[1]),
    .A2(_3744_),
    .ZN(_4189_)
  );
  AND2_X1 _4898_ (
    .A1(_4101_),
    .A2(_4189_),
    .ZN(_4198_)
  );
  AND2_X1 _4899_ (
    .A1(_4178_),
    .A2(_4198_),
    .ZN(_4209_)
  );
  OR2_X1 _4900_ (
    .A1(_3902_),
    .A2(_4209_),
    .ZN(_4218_)
  );
  OR2_X1 _4901_ (
    .A1(io_req_bits_fn[2]),
    .A2(io_req_bits_fn[1]),
    .ZN(_4227_)
  );
  AND2_X1 _4902_ (
    .A1(io_req_bits_fn[0]),
    .A2(_4227_),
    .ZN(_4238_)
  );
  OR2_X1 _4903_ (
    .A1(_3558_),
    .A2(_4238_),
    .ZN(_4247_)
  );
  MUX2_X1 _4904_ (
    .A(io_req_bits_fn[1]),
    .B(io_req_bits_fn[0]),
    .S(io_req_bits_fn[2]),
    .Z(_4257_)
  );
  OR2_X1 _4905_ (
    .A1(_3547_),
    .A2(_4257_),
    .ZN(_4260_)
  );
  INV_X1 _4906_ (
    .A(_4260_),
    .ZN(_4261_)
  );
  AND2_X1 _4907_ (
    .A1(_4247_),
    .A2(_4260_),
    .ZN(_4262_)
  );
  OR2_X1 _4908_ (
    .A1(_4140_),
    .A2(_4262_),
    .ZN(_4263_)
  );
  AND2_X1 _4909_ (
    .A1(_3253_),
    .A2(_4263_),
    .ZN(_4264_)
  );
  AND2_X1 _4910_ (
    .A1(_4218_),
    .A2(_4264_),
    .ZN(_0007_)
  );
  OR2_X1 _4911_ (
    .A1(remainder[63]),
    .A2(_4776_[31]),
    .ZN(_4265_)
  );
  AND2_X1 _4912_ (
    .A1(remainder[63]),
    .A2(_4776_[31]),
    .ZN(_4266_)
  );
  AND2_X1 _4913_ (
    .A1(remainder[62]),
    .A2(_4776_[30]),
    .ZN(_4267_)
  );
  XOR2_X1 _4914_ (
    .A(remainder[62]),
    .B(_4776_[30]),
    .Z(_4268_)
  );
  OR2_X1 _4915_ (
    .A1(remainder[61]),
    .A2(_4776_[29]),
    .ZN(_4269_)
  );
  AND2_X1 _4916_ (
    .A1(remainder[61]),
    .A2(_4776_[29]),
    .ZN(_4270_)
  );
  AND2_X1 _4917_ (
    .A1(remainder[60]),
    .A2(_4776_[28]),
    .ZN(_4271_)
  );
  XOR2_X1 _4918_ (
    .A(remainder[60]),
    .B(_4776_[28]),
    .Z(_4272_)
  );
  AND2_X1 _4919_ (
    .A1(remainder[59]),
    .A2(_4776_[27]),
    .ZN(_4273_)
  );
  OR2_X1 _4920_ (
    .A1(remainder[59]),
    .A2(_4776_[27]),
    .ZN(_4274_)
  );
  AND2_X1 _4921_ (
    .A1(remainder[58]),
    .A2(_4776_[26]),
    .ZN(_4275_)
  );
  XOR2_X1 _4922_ (
    .A(remainder[58]),
    .B(_4776_[26]),
    .Z(_4276_)
  );
  OR2_X1 _4923_ (
    .A1(remainder[57]),
    .A2(_4776_[25]),
    .ZN(_4277_)
  );
  AND2_X1 _4924_ (
    .A1(remainder[57]),
    .A2(_4776_[25]),
    .ZN(_4278_)
  );
  AND2_X1 _4925_ (
    .A1(remainder[56]),
    .A2(_4776_[24]),
    .ZN(_4279_)
  );
  XOR2_X1 _4926_ (
    .A(remainder[56]),
    .B(_4776_[24]),
    .Z(_4280_)
  );
  AND2_X1 _4927_ (
    .A1(remainder[55]),
    .A2(_4776_[23]),
    .ZN(_4281_)
  );
  OR2_X1 _4928_ (
    .A1(remainder[55]),
    .A2(_4776_[23]),
    .ZN(_4282_)
  );
  AND2_X1 _4929_ (
    .A1(remainder[54]),
    .A2(_4776_[22]),
    .ZN(_4283_)
  );
  XOR2_X1 _4930_ (
    .A(remainder[54]),
    .B(_4776_[22]),
    .Z(_4284_)
  );
  AND2_X1 _4931_ (
    .A1(remainder[53]),
    .A2(_4776_[21]),
    .ZN(_4285_)
  );
  OR2_X1 _4932_ (
    .A1(remainder[53]),
    .A2(_4776_[21]),
    .ZN(_4286_)
  );
  AND2_X1 _4933_ (
    .A1(remainder[52]),
    .A2(_4776_[20]),
    .ZN(_4287_)
  );
  XOR2_X1 _4934_ (
    .A(remainder[52]),
    .B(_4776_[20]),
    .Z(_4288_)
  );
  AND2_X1 _4935_ (
    .A1(remainder[51]),
    .A2(_4776_[19]),
    .ZN(_4289_)
  );
  OR2_X1 _4936_ (
    .A1(remainder[51]),
    .A2(_4776_[19]),
    .ZN(_4290_)
  );
  AND2_X1 _4937_ (
    .A1(remainder[50]),
    .A2(_4776_[18]),
    .ZN(_4291_)
  );
  XOR2_X1 _4938_ (
    .A(remainder[50]),
    .B(_4776_[18]),
    .Z(_4292_)
  );
  AND2_X1 _4939_ (
    .A1(remainder[49]),
    .A2(_4776_[17]),
    .ZN(_4293_)
  );
  OR2_X1 _4940_ (
    .A1(remainder[49]),
    .A2(_4776_[17]),
    .ZN(_4294_)
  );
  AND2_X1 _4941_ (
    .A1(remainder[48]),
    .A2(_4776_[16]),
    .ZN(_4295_)
  );
  XOR2_X1 _4942_ (
    .A(remainder[48]),
    .B(_4776_[16]),
    .Z(_4296_)
  );
  AND2_X1 _4943_ (
    .A1(remainder[47]),
    .A2(_4776_[15]),
    .ZN(_4297_)
  );
  OR2_X1 _4944_ (
    .A1(remainder[47]),
    .A2(_4776_[15]),
    .ZN(_4298_)
  );
  AND2_X1 _4945_ (
    .A1(remainder[46]),
    .A2(_4776_[14]),
    .ZN(_4299_)
  );
  XOR2_X1 _4946_ (
    .A(remainder[46]),
    .B(_4776_[14]),
    .Z(_4300_)
  );
  AND2_X1 _4947_ (
    .A1(remainder[45]),
    .A2(_4776_[13]),
    .ZN(_4301_)
  );
  OR2_X1 _4948_ (
    .A1(remainder[45]),
    .A2(_4776_[13]),
    .ZN(_4302_)
  );
  AND2_X1 _4949_ (
    .A1(remainder[44]),
    .A2(_4776_[12]),
    .ZN(_4303_)
  );
  XOR2_X1 _4950_ (
    .A(remainder[44]),
    .B(_4776_[12]),
    .Z(_4304_)
  );
  AND2_X1 _4951_ (
    .A1(remainder[43]),
    .A2(_4776_[11]),
    .ZN(_4305_)
  );
  OR2_X1 _4952_ (
    .A1(remainder[43]),
    .A2(_4776_[11]),
    .ZN(_4306_)
  );
  AND2_X1 _4953_ (
    .A1(remainder[42]),
    .A2(_4776_[10]),
    .ZN(_4307_)
  );
  XOR2_X1 _4954_ (
    .A(remainder[42]),
    .B(_4776_[10]),
    .Z(_4308_)
  );
  AND2_X1 _4955_ (
    .A1(remainder[41]),
    .A2(_4776_[9]),
    .ZN(_4309_)
  );
  OR2_X1 _4956_ (
    .A1(remainder[41]),
    .A2(_4776_[9]),
    .ZN(_4310_)
  );
  AND2_X1 _4957_ (
    .A1(remainder[40]),
    .A2(_4776_[8]),
    .ZN(_4311_)
  );
  XOR2_X1 _4958_ (
    .A(remainder[40]),
    .B(_4776_[8]),
    .Z(_4312_)
  );
  AND2_X1 _4959_ (
    .A1(remainder[39]),
    .A2(_4776_[7]),
    .ZN(_4313_)
  );
  OR2_X1 _4960_ (
    .A1(remainder[39]),
    .A2(_4776_[7]),
    .ZN(_4314_)
  );
  AND2_X1 _4961_ (
    .A1(remainder[38]),
    .A2(_4776_[6]),
    .ZN(_4315_)
  );
  XOR2_X1 _4962_ (
    .A(remainder[38]),
    .B(_4776_[6]),
    .Z(_4316_)
  );
  AND2_X1 _4963_ (
    .A1(remainder[37]),
    .A2(_4776_[5]),
    .ZN(_4317_)
  );
  AND2_X1 _4964_ (
    .A1(remainder[36]),
    .A2(_4776_[4]),
    .ZN(_4318_)
  );
  XOR2_X1 _4965_ (
    .A(remainder[36]),
    .B(_4776_[4]),
    .Z(_4319_)
  );
  AND2_X1 _4966_ (
    .A1(remainder[35]),
    .A2(_4776_[3]),
    .ZN(_4320_)
  );
  OR2_X1 _4967_ (
    .A1(remainder[35]),
    .A2(_4776_[3]),
    .ZN(_4321_)
  );
  AND2_X1 _4968_ (
    .A1(remainder[34]),
    .A2(_4776_[2]),
    .ZN(_4322_)
  );
  AND2_X1 _4969_ (
    .A1(remainder[33]),
    .A2(_4776_[1]),
    .ZN(_4323_)
  );
  OR2_X1 _4970_ (
    .A1(remainder[32]),
    .A2(_4776_[0]),
    .ZN(_4324_)
  );
  XOR2_X1 _4971_ (
    .A(remainder[33]),
    .B(_4776_[1]),
    .Z(_4325_)
  );
  AND2_X1 _4972_ (
    .A1(_4324_),
    .A2(_4325_),
    .ZN(_4326_)
  );
  OR2_X1 _4973_ (
    .A1(_4323_),
    .A2(_4326_),
    .ZN(_4327_)
  );
  XOR2_X1 _4974_ (
    .A(remainder[34]),
    .B(_4776_[2]),
    .Z(_4328_)
  );
  AND2_X1 _4975_ (
    .A1(_4327_),
    .A2(_4328_),
    .ZN(_4329_)
  );
  OR2_X1 _4976_ (
    .A1(_4322_),
    .A2(_4329_),
    .ZN(_4330_)
  );
  AND2_X1 _4977_ (
    .A1(_4321_),
    .A2(_4330_),
    .ZN(_4331_)
  );
  OR2_X1 _4978_ (
    .A1(_4320_),
    .A2(_4331_),
    .ZN(_4332_)
  );
  AND2_X1 _4979_ (
    .A1(_4319_),
    .A2(_4332_),
    .ZN(_4333_)
  );
  OR2_X1 _4980_ (
    .A1(_4318_),
    .A2(_4333_),
    .ZN(_4334_)
  );
  XOR2_X1 _4981_ (
    .A(remainder[37]),
    .B(_4776_[5]),
    .Z(_4335_)
  );
  AND2_X1 _4982_ (
    .A1(_4334_),
    .A2(_4335_),
    .ZN(_4336_)
  );
  OR2_X1 _4983_ (
    .A1(_4317_),
    .A2(_4336_),
    .ZN(_4337_)
  );
  AND2_X1 _4984_ (
    .A1(_4316_),
    .A2(_4337_),
    .ZN(_4338_)
  );
  OR2_X1 _4985_ (
    .A1(_4315_),
    .A2(_4338_),
    .ZN(_4339_)
  );
  AND2_X1 _4986_ (
    .A1(_4314_),
    .A2(_4339_),
    .ZN(_4340_)
  );
  OR2_X1 _4987_ (
    .A1(_4313_),
    .A2(_4340_),
    .ZN(_4341_)
  );
  AND2_X1 _4988_ (
    .A1(_4312_),
    .A2(_4341_),
    .ZN(_4342_)
  );
  OR2_X1 _4989_ (
    .A1(_4311_),
    .A2(_4342_),
    .ZN(_4343_)
  );
  AND2_X1 _4990_ (
    .A1(_4310_),
    .A2(_4343_),
    .ZN(_4344_)
  );
  OR2_X1 _4991_ (
    .A1(_4309_),
    .A2(_4344_),
    .ZN(_4345_)
  );
  AND2_X1 _4992_ (
    .A1(_4308_),
    .A2(_4345_),
    .ZN(_4346_)
  );
  OR2_X1 _4993_ (
    .A1(_4307_),
    .A2(_4346_),
    .ZN(_4347_)
  );
  AND2_X1 _4994_ (
    .A1(_4306_),
    .A2(_4347_),
    .ZN(_4348_)
  );
  OR2_X1 _4995_ (
    .A1(_4305_),
    .A2(_4348_),
    .ZN(_4349_)
  );
  AND2_X1 _4996_ (
    .A1(_4304_),
    .A2(_4349_),
    .ZN(_4350_)
  );
  OR2_X1 _4997_ (
    .A1(_4303_),
    .A2(_4350_),
    .ZN(_4351_)
  );
  AND2_X1 _4998_ (
    .A1(_4302_),
    .A2(_4351_),
    .ZN(_4352_)
  );
  OR2_X1 _4999_ (
    .A1(_4301_),
    .A2(_4352_),
    .ZN(_4353_)
  );
  AND2_X1 _5000_ (
    .A1(_4300_),
    .A2(_4353_),
    .ZN(_4354_)
  );
  OR2_X1 _5001_ (
    .A1(_4299_),
    .A2(_4354_),
    .ZN(_4355_)
  );
  AND2_X1 _5002_ (
    .A1(_4298_),
    .A2(_4355_),
    .ZN(_4356_)
  );
  OR2_X1 _5003_ (
    .A1(_4297_),
    .A2(_4356_),
    .ZN(_4357_)
  );
  AND2_X1 _5004_ (
    .A1(_4296_),
    .A2(_4357_),
    .ZN(_4358_)
  );
  OR2_X1 _5005_ (
    .A1(_4295_),
    .A2(_4358_),
    .ZN(_4359_)
  );
  AND2_X1 _5006_ (
    .A1(_4294_),
    .A2(_4359_),
    .ZN(_4360_)
  );
  OR2_X1 _5007_ (
    .A1(_4293_),
    .A2(_4360_),
    .ZN(_4361_)
  );
  AND2_X1 _5008_ (
    .A1(_4292_),
    .A2(_4361_),
    .ZN(_4362_)
  );
  OR2_X1 _5009_ (
    .A1(_4291_),
    .A2(_4362_),
    .ZN(_4363_)
  );
  AND2_X1 _5010_ (
    .A1(_4290_),
    .A2(_4363_),
    .ZN(_4364_)
  );
  OR2_X1 _5011_ (
    .A1(_4289_),
    .A2(_4364_),
    .ZN(_4365_)
  );
  AND2_X1 _5012_ (
    .A1(_4288_),
    .A2(_4365_),
    .ZN(_4366_)
  );
  OR2_X1 _5013_ (
    .A1(_4287_),
    .A2(_4366_),
    .ZN(_4367_)
  );
  AND2_X1 _5014_ (
    .A1(_4286_),
    .A2(_4367_),
    .ZN(_4368_)
  );
  OR2_X1 _5015_ (
    .A1(_4285_),
    .A2(_4368_),
    .ZN(_4369_)
  );
  AND2_X1 _5016_ (
    .A1(_4284_),
    .A2(_4369_),
    .ZN(_4370_)
  );
  OR2_X1 _5017_ (
    .A1(_4283_),
    .A2(_4370_),
    .ZN(_4371_)
  );
  AND2_X1 _5018_ (
    .A1(_4282_),
    .A2(_4371_),
    .ZN(_4372_)
  );
  OR2_X1 _5019_ (
    .A1(_4281_),
    .A2(_4372_),
    .ZN(_4373_)
  );
  AND2_X1 _5020_ (
    .A1(_4280_),
    .A2(_4373_),
    .ZN(_4374_)
  );
  OR2_X1 _5021_ (
    .A1(_4279_),
    .A2(_4374_),
    .ZN(_4375_)
  );
  OR2_X1 _5022_ (
    .A1(_4278_),
    .A2(_4375_),
    .ZN(_4376_)
  );
  AND2_X1 _5023_ (
    .A1(_4277_),
    .A2(_4376_),
    .ZN(_4377_)
  );
  AND2_X1 _5024_ (
    .A1(_4276_),
    .A2(_4377_),
    .ZN(_4378_)
  );
  OR2_X1 _5025_ (
    .A1(_4275_),
    .A2(_4378_),
    .ZN(_4379_)
  );
  AND2_X1 _5026_ (
    .A1(_4274_),
    .A2(_4379_),
    .ZN(_4380_)
  );
  OR2_X1 _5027_ (
    .A1(_4273_),
    .A2(_4380_),
    .ZN(_4381_)
  );
  AND2_X1 _5028_ (
    .A1(_4272_),
    .A2(_4381_),
    .ZN(_4382_)
  );
  OR2_X1 _5029_ (
    .A1(_4271_),
    .A2(_4382_),
    .ZN(_4383_)
  );
  OR2_X1 _5030_ (
    .A1(_4270_),
    .A2(_4383_),
    .ZN(_4384_)
  );
  AND2_X1 _5031_ (
    .A1(_4269_),
    .A2(_4384_),
    .ZN(_4385_)
  );
  AND2_X1 _5032_ (
    .A1(_4268_),
    .A2(_4385_),
    .ZN(_4386_)
  );
  OR2_X1 _5033_ (
    .A1(_4267_),
    .A2(_4386_),
    .ZN(_4387_)
  );
  OR2_X1 _5034_ (
    .A1(_4266_),
    .A2(_4387_),
    .ZN(_4388_)
  );
  AND2_X1 _5035_ (
    .A1(_4265_),
    .A2(_4388_),
    .ZN(_4389_)
  );
  XOR2_X1 _5036_ (
    .A(remainder[64]),
    .B(_4776_[32]),
    .Z(_4390_)
  );
  XOR2_X1 _5037_ (
    .A(_2947_),
    .B(_4776_[32]),
    .Z(_4391_)
  );
  XOR2_X1 _5038_ (
    .A(_4389_),
    .B(_4390_),
    .Z(_4392_)
  );
  XOR2_X1 _5039_ (
    .A(_4389_),
    .B(_4391_),
    .Z(_4393_)
  );
  OR2_X1 _5040_ (
    .A1(_3689_),
    .A2(_4392_),
    .ZN(_4394_)
  );
  OR2_X1 _5041_ (
    .A1(_3602_),
    .A2(_3754_),
    .ZN(_4395_)
  );
  OR2_X1 _5042_ (
    .A1(_3634_),
    .A2(_4395_),
    .ZN(_4396_)
  );
  OR2_X1 _5043_ (
    .A1(_4394_),
    .A2(_4396_),
    .ZN(_4397_)
  );
  AND2_X1 _5044_ (
    .A1(neg_out),
    .A2(_3911_),
    .ZN(_4398_)
  );
  AND2_X1 _5045_ (
    .A1(_4397_),
    .A2(_4398_),
    .ZN(_4399_)
  );
  AND2_X1 _5046_ (
    .A1(io_req_bits_fn[0]),
    .A2(_3525_),
    .ZN(_4400_)
  );
  OR2_X1 _5047_ (
    .A1(io_req_bits_fn[1]),
    .A2(_4400_),
    .ZN(_4401_)
  );
  OR2_X1 _5048_ (
    .A1(_4260_),
    .A2(_4401_),
    .ZN(_4402_)
  );
  XOR2_X1 _5049_ (
    .A(_4247_),
    .B(_4402_),
    .Z(_4403_)
  );
  AND2_X1 _5050_ (
    .A1(_3902_),
    .A2(_4403_),
    .ZN(_4404_)
  );
  OR2_X1 _5051_ (
    .A1(_4399_),
    .A2(_4404_),
    .ZN(_0008_)
  );
  MUX2_X1 _5052_ (
    .A(io_req_bits_tag[0]),
    .B(req_tag[0]),
    .S(_3911_),
    .Z(_0009_)
  );
  MUX2_X1 _5053_ (
    .A(io_req_bits_tag[1]),
    .B(req_tag[1]),
    .S(_3911_),
    .Z(_0010_)
  );
  MUX2_X1 _5054_ (
    .A(io_req_bits_tag[2]),
    .B(req_tag[2]),
    .S(_3911_),
    .Z(_0011_)
  );
  MUX2_X1 _5055_ (
    .A(io_req_bits_tag[3]),
    .B(req_tag[3]),
    .S(_3911_),
    .Z(_0012_)
  );
  MUX2_X1 _5056_ (
    .A(io_req_bits_tag[4]),
    .B(req_tag[4]),
    .S(_3911_),
    .Z(_0013_)
  );
  OR2_X1 _5057_ (
    .A1(_3678_),
    .A2(_3819_),
    .ZN(_4405_)
  );
  INV_X1 _5058_ (
    .A(_4405_),
    .ZN(_4406_)
  );
  MUX2_X1 _5059_ (
    .A(count[0]),
    .B(_count_T_1[0]),
    .S(_4405_),
    .Z(_4407_)
  );
  AND2_X1 _5060_ (
    .A1(_3911_),
    .A2(_4407_),
    .ZN(_0014_)
  );
  AND2_X1 _5061_ (
    .A1(count[0]),
    .A2(_4405_),
    .ZN(_4408_)
  );
  INV_X1 _5062_ (
    .A(_4408_),
    .ZN(_4409_)
  );
  AND2_X1 _5063_ (
    .A1(count[1]),
    .A2(_4408_),
    .ZN(_4410_)
  );
  OR2_X1 _5064_ (
    .A1(_3231_),
    .A2(_4409_),
    .ZN(_4411_)
  );
  OR2_X1 _5065_ (
    .A1(count[1]),
    .A2(_4408_),
    .ZN(_4412_)
  );
  AND2_X1 _5066_ (
    .A1(_3911_),
    .A2(_4412_),
    .ZN(_4413_)
  );
  AND2_X1 _5067_ (
    .A1(_4411_),
    .A2(_4413_),
    .ZN(_0015_)
  );
  AND2_X1 _5068_ (
    .A1(count[2]),
    .A2(_4410_),
    .ZN(_4414_)
  );
  OR2_X1 _5069_ (
    .A1(_3220_),
    .A2(_4411_),
    .ZN(_4415_)
  );
  OR2_X1 _5070_ (
    .A1(count[2]),
    .A2(_4410_),
    .ZN(_4416_)
  );
  AND2_X1 _5071_ (
    .A1(_3911_),
    .A2(_4416_),
    .ZN(_4417_)
  );
  AND2_X1 _5072_ (
    .A1(_4415_),
    .A2(_4417_),
    .ZN(_0016_)
  );
  AND2_X1 _5073_ (
    .A1(count[3]),
    .A2(_4414_),
    .ZN(_4418_)
  );
  INV_X1 _5074_ (
    .A(_4418_),
    .ZN(_4419_)
  );
  OR2_X1 _5075_ (
    .A1(count[3]),
    .A2(_4414_),
    .ZN(_4420_)
  );
  AND2_X1 _5076_ (
    .A1(_3911_),
    .A2(_4420_),
    .ZN(_4421_)
  );
  AND2_X1 _5077_ (
    .A1(_4419_),
    .A2(_4421_),
    .ZN(_0017_)
  );
  AND2_X1 _5078_ (
    .A1(count[4]),
    .A2(_4418_),
    .ZN(_4422_)
  );
  INV_X1 _5079_ (
    .A(_4422_),
    .ZN(_4423_)
  );
  OR2_X1 _5080_ (
    .A1(count[4]),
    .A2(_4418_),
    .ZN(_4424_)
  );
  AND2_X1 _5081_ (
    .A1(_3911_),
    .A2(_4424_),
    .ZN(_4425_)
  );
  AND2_X1 _5082_ (
    .A1(_4423_),
    .A2(_4425_),
    .ZN(_0018_)
  );
  XOR2_X1 _5083_ (
    .A(count[5]),
    .B(_4422_),
    .Z(_4426_)
  );
  AND2_X1 _5084_ (
    .A1(_3911_),
    .A2(_4426_),
    .ZN(_0019_)
  );
  AND2_X1 _5085_ (
    .A1(divisor[31]),
    .A2(_4015_),
    .ZN(_4427_)
  );
  OR2_X1 _5086_ (
    .A1(_3438_),
    .A2(_4006_),
    .ZN(_4428_)
  );
  AND2_X1 _5087_ (
    .A1(_3911_),
    .A2(_4428_),
    .ZN(_4429_)
  );
  AND2_X1 _5088_ (
    .A1(divisor[0]),
    .A2(_4429_),
    .ZN(_4430_)
  );
  AND2_X1 _5089_ (
    .A1(io_req_bits_in2[0]),
    .A2(_3902_),
    .ZN(_4431_)
  );
  XOR2_X1 _5090_ (
    .A(_3209_),
    .B(_4776_[0]),
    .Z(_4432_)
  );
  AND2_X1 _5091_ (
    .A1(_3911_),
    .A2(_4427_),
    .ZN(_4433_)
  );
  AND2_X1 _5092_ (
    .A1(_4432_),
    .A2(_4433_),
    .ZN(_4434_)
  );
  OR2_X1 _5093_ (
    .A1(_4430_),
    .A2(_4434_),
    .ZN(_4435_)
  );
  OR2_X1 _5094_ (
    .A1(_4431_),
    .A2(_4435_),
    .ZN(_0020_)
  );
  AND2_X1 _5095_ (
    .A1(divisor[1]),
    .A2(_4429_),
    .ZN(_4436_)
  );
  AND2_X1 _5096_ (
    .A1(io_req_bits_in2[1]),
    .A2(_3902_),
    .ZN(_4437_)
  );
  XOR2_X1 _5097_ (
    .A(_4324_),
    .B(_4325_),
    .Z(_4438_)
  );
  AND2_X1 _5098_ (
    .A1(_4433_),
    .A2(_4438_),
    .ZN(_4439_)
  );
  OR2_X1 _5099_ (
    .A1(_4436_),
    .A2(_4439_),
    .ZN(_4440_)
  );
  OR2_X1 _5100_ (
    .A1(_4437_),
    .A2(_4440_),
    .ZN(_0021_)
  );
  XOR2_X1 _5101_ (
    .A(_4327_),
    .B(_4328_),
    .Z(_4441_)
  );
  AND2_X1 _5102_ (
    .A1(_4433_),
    .A2(_4441_),
    .ZN(_4442_)
  );
  AND2_X1 _5103_ (
    .A1(io_req_bits_in2[2]),
    .A2(_3902_),
    .ZN(_4443_)
  );
  AND2_X1 _5104_ (
    .A1(divisor[2]),
    .A2(_4429_),
    .ZN(_4444_)
  );
  OR2_X1 _5105_ (
    .A1(_4443_),
    .A2(_4444_),
    .ZN(_4445_)
  );
  OR2_X1 _5106_ (
    .A1(_4442_),
    .A2(_4445_),
    .ZN(_0022_)
  );
  XOR2_X1 _5107_ (
    .A(remainder[35]),
    .B(_4776_[3]),
    .Z(_4446_)
  );
  XOR2_X1 _5108_ (
    .A(_4330_),
    .B(_4446_),
    .Z(_4447_)
  );
  AND2_X1 _5109_ (
    .A1(_4433_),
    .A2(_4447_),
    .ZN(_4448_)
  );
  AND2_X1 _5110_ (
    .A1(io_req_bits_in2[3]),
    .A2(_3902_),
    .ZN(_4449_)
  );
  AND2_X1 _5111_ (
    .A1(divisor[3]),
    .A2(_4429_),
    .ZN(_4450_)
  );
  OR2_X1 _5112_ (
    .A1(_4449_),
    .A2(_4450_),
    .ZN(_4451_)
  );
  OR2_X1 _5113_ (
    .A1(_4448_),
    .A2(_4451_),
    .ZN(_0023_)
  );
  XOR2_X1 _5114_ (
    .A(_4319_),
    .B(_4332_),
    .Z(_4452_)
  );
  AND2_X1 _5115_ (
    .A1(_4433_),
    .A2(_4452_),
    .ZN(_4453_)
  );
  AND2_X1 _5116_ (
    .A1(divisor[4]),
    .A2(_4429_),
    .ZN(_4454_)
  );
  AND2_X1 _5117_ (
    .A1(io_req_bits_in2[4]),
    .A2(_3902_),
    .ZN(_4455_)
  );
  OR2_X1 _5118_ (
    .A1(_4454_),
    .A2(_4455_),
    .ZN(_4456_)
  );
  OR2_X1 _5119_ (
    .A1(_4453_),
    .A2(_4456_),
    .ZN(_0024_)
  );
  XOR2_X1 _5120_ (
    .A(_4334_),
    .B(_4335_),
    .Z(_4457_)
  );
  AND2_X1 _5121_ (
    .A1(_4433_),
    .A2(_4457_),
    .ZN(_4458_)
  );
  AND2_X1 _5122_ (
    .A1(io_req_bits_in2[5]),
    .A2(_3902_),
    .ZN(_4459_)
  );
  AND2_X1 _5123_ (
    .A1(divisor[5]),
    .A2(_4429_),
    .ZN(_4460_)
  );
  OR2_X1 _5124_ (
    .A1(_4459_),
    .A2(_4460_),
    .ZN(_4461_)
  );
  OR2_X1 _5125_ (
    .A1(_4458_),
    .A2(_4461_),
    .ZN(_0025_)
  );
  XOR2_X1 _5126_ (
    .A(_4316_),
    .B(_4337_),
    .Z(_4462_)
  );
  AND2_X1 _5127_ (
    .A1(_4433_),
    .A2(_4462_),
    .ZN(_4463_)
  );
  AND2_X1 _5128_ (
    .A1(io_req_bits_in2[6]),
    .A2(_3902_),
    .ZN(_4464_)
  );
  AND2_X1 _5129_ (
    .A1(divisor[6]),
    .A2(_4429_),
    .ZN(_4465_)
  );
  OR2_X1 _5130_ (
    .A1(_4464_),
    .A2(_4465_),
    .ZN(_4466_)
  );
  OR2_X1 _5131_ (
    .A1(_4463_),
    .A2(_4466_),
    .ZN(_0026_)
  );
  XOR2_X1 _5132_ (
    .A(remainder[39]),
    .B(_4776_[7]),
    .Z(_4467_)
  );
  XOR2_X1 _5133_ (
    .A(_4339_),
    .B(_4467_),
    .Z(_4468_)
  );
  AND2_X1 _5134_ (
    .A1(_4433_),
    .A2(_4468_),
    .ZN(_4469_)
  );
  AND2_X1 _5135_ (
    .A1(io_req_bits_in2[7]),
    .A2(_3902_),
    .ZN(_4470_)
  );
  AND2_X1 _5136_ (
    .A1(divisor[7]),
    .A2(_4429_),
    .ZN(_4471_)
  );
  OR2_X1 _5137_ (
    .A1(_4470_),
    .A2(_4471_),
    .ZN(_4472_)
  );
  OR2_X1 _5138_ (
    .A1(_4469_),
    .A2(_4472_),
    .ZN(_0027_)
  );
  XOR2_X1 _5139_ (
    .A(_4312_),
    .B(_4341_),
    .Z(_4473_)
  );
  AND2_X1 _5140_ (
    .A1(_4433_),
    .A2(_4473_),
    .ZN(_4474_)
  );
  AND2_X1 _5141_ (
    .A1(divisor[8]),
    .A2(_4429_),
    .ZN(_4475_)
  );
  AND2_X1 _5142_ (
    .A1(io_req_bits_in2[8]),
    .A2(_3902_),
    .ZN(_4476_)
  );
  OR2_X1 _5143_ (
    .A1(_4475_),
    .A2(_4476_),
    .ZN(_4477_)
  );
  OR2_X1 _5144_ (
    .A1(_4474_),
    .A2(_4477_),
    .ZN(_0028_)
  );
  XOR2_X1 _5145_ (
    .A(remainder[41]),
    .B(_4776_[9]),
    .Z(_4478_)
  );
  XOR2_X1 _5146_ (
    .A(_4343_),
    .B(_4478_),
    .Z(_4479_)
  );
  AND2_X1 _5147_ (
    .A1(_4433_),
    .A2(_4479_),
    .ZN(_4480_)
  );
  AND2_X1 _5148_ (
    .A1(io_req_bits_in2[9]),
    .A2(_3902_),
    .ZN(_4481_)
  );
  AND2_X1 _5149_ (
    .A1(divisor[9]),
    .A2(_4429_),
    .ZN(_4482_)
  );
  OR2_X1 _5150_ (
    .A1(_4481_),
    .A2(_4482_),
    .ZN(_4483_)
  );
  OR2_X1 _5151_ (
    .A1(_4480_),
    .A2(_4483_),
    .ZN(_0029_)
  );
  XOR2_X1 _5152_ (
    .A(_4308_),
    .B(_4345_),
    .Z(_4484_)
  );
  AND2_X1 _5153_ (
    .A1(_4433_),
    .A2(_4484_),
    .ZN(_4485_)
  );
  AND2_X1 _5154_ (
    .A1(io_req_bits_in2[10]),
    .A2(_3902_),
    .ZN(_4486_)
  );
  AND2_X1 _5155_ (
    .A1(divisor[10]),
    .A2(_4429_),
    .ZN(_4487_)
  );
  OR2_X1 _5156_ (
    .A1(_4486_),
    .A2(_4487_),
    .ZN(_4488_)
  );
  OR2_X1 _5157_ (
    .A1(_4485_),
    .A2(_4488_),
    .ZN(_0030_)
  );
  XOR2_X1 _5158_ (
    .A(remainder[43]),
    .B(_4776_[11]),
    .Z(_4489_)
  );
  XOR2_X1 _5159_ (
    .A(_4347_),
    .B(_4489_),
    .Z(_4490_)
  );
  AND2_X1 _5160_ (
    .A1(_4433_),
    .A2(_4490_),
    .ZN(_4491_)
  );
  AND2_X1 _5161_ (
    .A1(io_req_bits_in2[11]),
    .A2(_3902_),
    .ZN(_4492_)
  );
  AND2_X1 _5162_ (
    .A1(divisor[11]),
    .A2(_4429_),
    .ZN(_4493_)
  );
  OR2_X1 _5163_ (
    .A1(_4492_),
    .A2(_4493_),
    .ZN(_4494_)
  );
  OR2_X1 _5164_ (
    .A1(_4491_),
    .A2(_4494_),
    .ZN(_0031_)
  );
  XOR2_X1 _5165_ (
    .A(_4304_),
    .B(_4349_),
    .Z(_4495_)
  );
  AND2_X1 _5166_ (
    .A1(_4433_),
    .A2(_4495_),
    .ZN(_4496_)
  );
  AND2_X1 _5167_ (
    .A1(divisor[12]),
    .A2(_4429_),
    .ZN(_4497_)
  );
  AND2_X1 _5168_ (
    .A1(io_req_bits_in2[12]),
    .A2(_3902_),
    .ZN(_4498_)
  );
  OR2_X1 _5169_ (
    .A1(_4497_),
    .A2(_4498_),
    .ZN(_4499_)
  );
  OR2_X1 _5170_ (
    .A1(_4496_),
    .A2(_4499_),
    .ZN(_0032_)
  );
  XOR2_X1 _5171_ (
    .A(remainder[45]),
    .B(_4776_[13]),
    .Z(_4500_)
  );
  XOR2_X1 _5172_ (
    .A(_4351_),
    .B(_4500_),
    .Z(_4501_)
  );
  AND2_X1 _5173_ (
    .A1(_4433_),
    .A2(_4501_),
    .ZN(_4502_)
  );
  AND2_X1 _5174_ (
    .A1(divisor[13]),
    .A2(_4429_),
    .ZN(_4503_)
  );
  AND2_X1 _5175_ (
    .A1(io_req_bits_in2[13]),
    .A2(_3902_),
    .ZN(_4504_)
  );
  OR2_X1 _5176_ (
    .A1(_4503_),
    .A2(_4504_),
    .ZN(_4505_)
  );
  OR2_X1 _5177_ (
    .A1(_4502_),
    .A2(_4505_),
    .ZN(_0033_)
  );
  XOR2_X1 _5178_ (
    .A(_4300_),
    .B(_4353_),
    .Z(_4506_)
  );
  AND2_X1 _5179_ (
    .A1(_4433_),
    .A2(_4506_),
    .ZN(_4507_)
  );
  AND2_X1 _5180_ (
    .A1(io_req_bits_in2[14]),
    .A2(_3902_),
    .ZN(_4508_)
  );
  AND2_X1 _5181_ (
    .A1(divisor[14]),
    .A2(_4429_),
    .ZN(_4509_)
  );
  OR2_X1 _5182_ (
    .A1(_4508_),
    .A2(_4509_),
    .ZN(_4510_)
  );
  OR2_X1 _5183_ (
    .A1(_4507_),
    .A2(_4510_),
    .ZN(_0034_)
  );
  XOR2_X1 _5184_ (
    .A(remainder[47]),
    .B(_4776_[15]),
    .Z(_4511_)
  );
  XOR2_X1 _5185_ (
    .A(_4355_),
    .B(_4511_),
    .Z(_4512_)
  );
  AND2_X1 _5186_ (
    .A1(_4433_),
    .A2(_4512_),
    .ZN(_4513_)
  );
  AND2_X1 _5187_ (
    .A1(divisor[15]),
    .A2(_4429_),
    .ZN(_4514_)
  );
  AND2_X1 _5188_ (
    .A1(io_req_bits_in2[15]),
    .A2(_3902_),
    .ZN(_4515_)
  );
  OR2_X1 _5189_ (
    .A1(_4514_),
    .A2(_4515_),
    .ZN(_4516_)
  );
  OR2_X1 _5190_ (
    .A1(_4513_),
    .A2(_4516_),
    .ZN(_0035_)
  );
  XOR2_X1 _5191_ (
    .A(_4296_),
    .B(_4357_),
    .Z(_4517_)
  );
  AND2_X1 _5192_ (
    .A1(_4433_),
    .A2(_4517_),
    .ZN(_4518_)
  );
  AND2_X1 _5193_ (
    .A1(io_req_bits_in2[16]),
    .A2(_3902_),
    .ZN(_4519_)
  );
  AND2_X1 _5194_ (
    .A1(divisor[16]),
    .A2(_4429_),
    .ZN(_4520_)
  );
  OR2_X1 _5195_ (
    .A1(_4519_),
    .A2(_4520_),
    .ZN(_4521_)
  );
  OR2_X1 _5196_ (
    .A1(_4518_),
    .A2(_4521_),
    .ZN(_0036_)
  );
  XOR2_X1 _5197_ (
    .A(remainder[49]),
    .B(_4776_[17]),
    .Z(_4522_)
  );
  XOR2_X1 _5198_ (
    .A(_4359_),
    .B(_4522_),
    .Z(_4523_)
  );
  AND2_X1 _5199_ (
    .A1(_4433_),
    .A2(_4523_),
    .ZN(_4524_)
  );
  AND2_X1 _5200_ (
    .A1(io_req_bits_in2[17]),
    .A2(_3902_),
    .ZN(_4525_)
  );
  AND2_X1 _5201_ (
    .A1(divisor[17]),
    .A2(_4429_),
    .ZN(_4526_)
  );
  OR2_X1 _5202_ (
    .A1(_4525_),
    .A2(_4526_),
    .ZN(_4527_)
  );
  OR2_X1 _5203_ (
    .A1(_4524_),
    .A2(_4527_),
    .ZN(_0037_)
  );
  XOR2_X1 _5204_ (
    .A(_4292_),
    .B(_4361_),
    .Z(_4528_)
  );
  AND2_X1 _5205_ (
    .A1(_4433_),
    .A2(_4528_),
    .ZN(_4529_)
  );
  AND2_X1 _5206_ (
    .A1(io_req_bits_in2[18]),
    .A2(_3902_),
    .ZN(_4530_)
  );
  AND2_X1 _5207_ (
    .A1(divisor[18]),
    .A2(_4429_),
    .ZN(_4531_)
  );
  OR2_X1 _5208_ (
    .A1(_4530_),
    .A2(_4531_),
    .ZN(_4532_)
  );
  OR2_X1 _5209_ (
    .A1(_4529_),
    .A2(_4532_),
    .ZN(_0038_)
  );
  XOR2_X1 _5210_ (
    .A(remainder[51]),
    .B(_4776_[19]),
    .Z(_4533_)
  );
  XOR2_X1 _5211_ (
    .A(_4363_),
    .B(_4533_),
    .Z(_4534_)
  );
  AND2_X1 _5212_ (
    .A1(_4433_),
    .A2(_4534_),
    .ZN(_4535_)
  );
  AND2_X1 _5213_ (
    .A1(io_req_bits_in2[19]),
    .A2(_3902_),
    .ZN(_4536_)
  );
  AND2_X1 _5214_ (
    .A1(divisor[19]),
    .A2(_4429_),
    .ZN(_4537_)
  );
  OR2_X1 _5215_ (
    .A1(_4536_),
    .A2(_4537_),
    .ZN(_4538_)
  );
  OR2_X1 _5216_ (
    .A1(_4535_),
    .A2(_4538_),
    .ZN(_0039_)
  );
  XOR2_X1 _5217_ (
    .A(_4288_),
    .B(_4365_),
    .Z(_4539_)
  );
  AND2_X1 _5218_ (
    .A1(_4433_),
    .A2(_4539_),
    .ZN(_4540_)
  );
  AND2_X1 _5219_ (
    .A1(divisor[20]),
    .A2(_4429_),
    .ZN(_4541_)
  );
  AND2_X1 _5220_ (
    .A1(io_req_bits_in2[20]),
    .A2(_3902_),
    .ZN(_4542_)
  );
  OR2_X1 _5221_ (
    .A1(_4541_),
    .A2(_4542_),
    .ZN(_4543_)
  );
  OR2_X1 _5222_ (
    .A1(_4540_),
    .A2(_4543_),
    .ZN(_0040_)
  );
  XOR2_X1 _5223_ (
    .A(remainder[53]),
    .B(_4776_[21]),
    .Z(_4544_)
  );
  XOR2_X1 _5224_ (
    .A(_4367_),
    .B(_4544_),
    .Z(_4545_)
  );
  AND2_X1 _5225_ (
    .A1(_4433_),
    .A2(_4545_),
    .ZN(_4546_)
  );
  AND2_X1 _5226_ (
    .A1(io_req_bits_in2[21]),
    .A2(_3902_),
    .ZN(_4547_)
  );
  AND2_X1 _5227_ (
    .A1(divisor[21]),
    .A2(_4429_),
    .ZN(_4548_)
  );
  OR2_X1 _5228_ (
    .A1(_4547_),
    .A2(_4548_),
    .ZN(_4549_)
  );
  OR2_X1 _5229_ (
    .A1(_4546_),
    .A2(_4549_),
    .ZN(_0041_)
  );
  XOR2_X1 _5230_ (
    .A(_4284_),
    .B(_4369_),
    .Z(_4550_)
  );
  AND2_X1 _5231_ (
    .A1(_4433_),
    .A2(_4550_),
    .ZN(_4551_)
  );
  AND2_X1 _5232_ (
    .A1(divisor[22]),
    .A2(_4429_),
    .ZN(_4552_)
  );
  AND2_X1 _5233_ (
    .A1(io_req_bits_in2[22]),
    .A2(_3902_),
    .ZN(_4553_)
  );
  OR2_X1 _5234_ (
    .A1(_4552_),
    .A2(_4553_),
    .ZN(_4554_)
  );
  OR2_X1 _5235_ (
    .A1(_4551_),
    .A2(_4554_),
    .ZN(_0042_)
  );
  XOR2_X1 _5236_ (
    .A(remainder[55]),
    .B(_4776_[23]),
    .Z(_4555_)
  );
  XOR2_X1 _5237_ (
    .A(_4371_),
    .B(_4555_),
    .Z(_4556_)
  );
  AND2_X1 _5238_ (
    .A1(_4433_),
    .A2(_4556_),
    .ZN(_4557_)
  );
  AND2_X1 _5239_ (
    .A1(io_req_bits_in2[23]),
    .A2(_3902_),
    .ZN(_4558_)
  );
  AND2_X1 _5240_ (
    .A1(divisor[23]),
    .A2(_4429_),
    .ZN(_4559_)
  );
  OR2_X1 _5241_ (
    .A1(_4558_),
    .A2(_4559_),
    .ZN(_4560_)
  );
  OR2_X1 _5242_ (
    .A1(_4557_),
    .A2(_4560_),
    .ZN(_0043_)
  );
  XOR2_X1 _5243_ (
    .A(_4280_),
    .B(_4373_),
    .Z(_4561_)
  );
  AND2_X1 _5244_ (
    .A1(_4433_),
    .A2(_4561_),
    .ZN(_4562_)
  );
  AND2_X1 _5245_ (
    .A1(io_req_bits_in2[24]),
    .A2(_3902_),
    .ZN(_4563_)
  );
  AND2_X1 _5246_ (
    .A1(divisor[24]),
    .A2(_4429_),
    .ZN(_4564_)
  );
  OR2_X1 _5247_ (
    .A1(_4563_),
    .A2(_4564_),
    .ZN(_4565_)
  );
  OR2_X1 _5248_ (
    .A1(_4562_),
    .A2(_4565_),
    .ZN(_0044_)
  );
  XOR2_X1 _5249_ (
    .A(remainder[57]),
    .B(_4776_[25]),
    .Z(_4566_)
  );
  XOR2_X1 _5250_ (
    .A(_4375_),
    .B(_4566_),
    .Z(_4567_)
  );
  AND2_X1 _5251_ (
    .A1(_4433_),
    .A2(_4567_),
    .ZN(_4568_)
  );
  AND2_X1 _5252_ (
    .A1(divisor[25]),
    .A2(_4429_),
    .ZN(_4569_)
  );
  AND2_X1 _5253_ (
    .A1(io_req_bits_in2[25]),
    .A2(_3902_),
    .ZN(_4570_)
  );
  OR2_X1 _5254_ (
    .A1(_4569_),
    .A2(_4570_),
    .ZN(_4571_)
  );
  OR2_X1 _5255_ (
    .A1(_4568_),
    .A2(_4571_),
    .ZN(_0045_)
  );
  XOR2_X1 _5256_ (
    .A(_4276_),
    .B(_4377_),
    .Z(_4572_)
  );
  AND2_X1 _5257_ (
    .A1(_4433_),
    .A2(_4572_),
    .ZN(_4573_)
  );
  AND2_X1 _5258_ (
    .A1(divisor[26]),
    .A2(_4429_),
    .ZN(_4574_)
  );
  AND2_X1 _5259_ (
    .A1(io_req_bits_in2[26]),
    .A2(_3902_),
    .ZN(_4575_)
  );
  OR2_X1 _5260_ (
    .A1(_4574_),
    .A2(_4575_),
    .ZN(_4576_)
  );
  OR2_X1 _5261_ (
    .A1(_4573_),
    .A2(_4576_),
    .ZN(_0046_)
  );
  XOR2_X1 _5262_ (
    .A(remainder[59]),
    .B(_4776_[27]),
    .Z(_4577_)
  );
  XOR2_X1 _5263_ (
    .A(_4379_),
    .B(_4577_),
    .Z(_4578_)
  );
  AND2_X1 _5264_ (
    .A1(_4433_),
    .A2(_4578_),
    .ZN(_4579_)
  );
  AND2_X1 _5265_ (
    .A1(io_req_bits_in2[27]),
    .A2(_3902_),
    .ZN(_4580_)
  );
  AND2_X1 _5266_ (
    .A1(divisor[27]),
    .A2(_4429_),
    .ZN(_4581_)
  );
  OR2_X1 _5267_ (
    .A1(_4580_),
    .A2(_4581_),
    .ZN(_4582_)
  );
  OR2_X1 _5268_ (
    .A1(_4579_),
    .A2(_4582_),
    .ZN(_0047_)
  );
  XOR2_X1 _5269_ (
    .A(_4272_),
    .B(_4381_),
    .Z(_4583_)
  );
  AND2_X1 _5270_ (
    .A1(_4433_),
    .A2(_4583_),
    .ZN(_4584_)
  );
  AND2_X1 _5271_ (
    .A1(io_req_bits_in2[28]),
    .A2(_3902_),
    .ZN(_4585_)
  );
  AND2_X1 _5272_ (
    .A1(divisor[28]),
    .A2(_4429_),
    .ZN(_4586_)
  );
  OR2_X1 _5273_ (
    .A1(_4585_),
    .A2(_4586_),
    .ZN(_4587_)
  );
  OR2_X1 _5274_ (
    .A1(_4584_),
    .A2(_4587_),
    .ZN(_0048_)
  );
  XOR2_X1 _5275_ (
    .A(remainder[61]),
    .B(_4776_[29]),
    .Z(_4588_)
  );
  XOR2_X1 _5276_ (
    .A(_4383_),
    .B(_4588_),
    .Z(_4589_)
  );
  AND2_X1 _5277_ (
    .A1(_4433_),
    .A2(_4589_),
    .ZN(_4590_)
  );
  AND2_X1 _5278_ (
    .A1(divisor[29]),
    .A2(_4429_),
    .ZN(_4591_)
  );
  AND2_X1 _5279_ (
    .A1(io_req_bits_in2[29]),
    .A2(_3902_),
    .ZN(_4592_)
  );
  OR2_X1 _5280_ (
    .A1(_4591_),
    .A2(_4592_),
    .ZN(_4593_)
  );
  OR2_X1 _5281_ (
    .A1(_4590_),
    .A2(_4593_),
    .ZN(_0049_)
  );
  XOR2_X1 _5282_ (
    .A(_4268_),
    .B(_4385_),
    .Z(_4594_)
  );
  AND2_X1 _5283_ (
    .A1(_4433_),
    .A2(_4594_),
    .ZN(_4595_)
  );
  AND2_X1 _5284_ (
    .A1(divisor[30]),
    .A2(_4429_),
    .ZN(_4596_)
  );
  AND2_X1 _5285_ (
    .A1(io_req_bits_in2[30]),
    .A2(_3902_),
    .ZN(_4597_)
  );
  OR2_X1 _5286_ (
    .A1(_4596_),
    .A2(_4597_),
    .ZN(_4598_)
  );
  OR2_X1 _5287_ (
    .A1(_4595_),
    .A2(_4598_),
    .ZN(_0050_)
  );
  XOR2_X1 _5288_ (
    .A(remainder[63]),
    .B(_4776_[31]),
    .Z(_4599_)
  );
  XOR2_X1 _5289_ (
    .A(_4387_),
    .B(_4599_),
    .Z(_4600_)
  );
  OR2_X1 _5290_ (
    .A1(_4006_),
    .A2(_4600_),
    .ZN(_4601_)
  );
  AND2_X1 _5291_ (
    .A1(divisor[31]),
    .A2(_4601_),
    .ZN(_4602_)
  );
  MUX2_X1 _5292_ (
    .A(io_req_bits_in2[31]),
    .B(_4602_),
    .S(_3911_),
    .Z(_0051_)
  );
  AND2_X1 _5293_ (
    .A1(_4392_),
    .A2(_4433_),
    .ZN(_4603_)
  );
  AND2_X1 _5294_ (
    .A1(_3902_),
    .A2(_4261_),
    .ZN(_4604_)
  );
  AND2_X1 _5295_ (
    .A1(divisor[32]),
    .A2(_4429_),
    .ZN(_4605_)
  );
  OR2_X1 _5296_ (
    .A1(_4604_),
    .A2(_4605_),
    .ZN(_4606_)
  );
  OR2_X1 _5297_ (
    .A1(_4603_),
    .A2(_4606_),
    .ZN(_0052_)
  );
  OR2_X1 _5298_ (
    .A1(_3504_),
    .A2(_4006_),
    .ZN(_4607_)
  );
  AND2_X1 _5299_ (
    .A1(_3969_),
    .A2(_4607_),
    .ZN(_4608_)
  );
  INV_X1 _5300_ (
    .A(_4608_),
    .ZN(_4609_)
  );
  AND2_X1 _5301_ (
    .A1(_4406_),
    .A2(_4608_),
    .ZN(_4610_)
  );
  AND2_X1 _5302_ (
    .A1(remainder[32]),
    .A2(_4610_),
    .ZN(_4611_)
  );
  AND2_X1 _5303_ (
    .A1(remainder[31]),
    .A2(_3678_),
    .ZN(_4612_)
  );
  AND2_X1 _5304_ (
    .A1(_0004_),
    .A2(_3819_),
    .ZN(_4613_)
  );
  AND2_X1 _5305_ (
    .A1(_3242_),
    .A2(neg_out),
    .ZN(_4614_)
  );
  AND2_X1 _5306_ (
    .A1(_3787_),
    .A2(_4614_),
    .ZN(_4615_)
  );
  AND2_X1 _5307_ (
    .A1(_4613_),
    .A2(_4615_),
    .ZN(_4616_)
  );
  OR2_X1 _5308_ (
    .A1(_4612_),
    .A2(_4616_),
    .ZN(_4617_)
  );
  OR2_X1 _5309_ (
    .A1(_4611_),
    .A2(_4617_),
    .ZN(_4618_)
  );
  AND2_X1 _5310_ (
    .A1(_3911_),
    .A2(_4618_),
    .ZN(_0053_)
  );
  MUX2_X1 _5311_ (
    .A(remainder[32]),
    .B(_4432_),
    .S(_4393_),
    .Z(_4619_)
  );
  AND2_X1 _5312_ (
    .A1(_3678_),
    .A2(_4619_),
    .ZN(_4620_)
  );
  AND2_X1 _5313_ (
    .A1(remainder[33]),
    .A2(_4610_),
    .ZN(_4621_)
  );
  AND2_X1 _5314_ (
    .A1(divisor[3]),
    .A2(remainder[3]),
    .ZN(_4622_)
  );
  INV_X1 _5315_ (
    .A(_4622_),
    .ZN(_4623_)
  );
  AND2_X1 _5316_ (
    .A1(divisor[0]),
    .A2(remainder[4]),
    .ZN(_4624_)
  );
  AND2_X1 _5317_ (
    .A1(divisor[1]),
    .A2(remainder[3]),
    .ZN(_4625_)
  );
  AND2_X1 _5318_ (
    .A1(divisor[1]),
    .A2(remainder[4]),
    .ZN(_4626_)
  );
  AND2_X1 _5319_ (
    .A1(divisor[0]),
    .A2(remainder[3]),
    .ZN(_4627_)
  );
  AND2_X1 _5320_ (
    .A1(_4624_),
    .A2(_4625_),
    .ZN(_4628_)
  );
  AND2_X1 _5321_ (
    .A1(divisor[2]),
    .A2(remainder[2]),
    .ZN(_4629_)
  );
  XOR2_X1 _5322_ (
    .A(_4624_),
    .B(_4625_),
    .Z(_4630_)
  );
  AND2_X1 _5323_ (
    .A1(_4629_),
    .A2(_4630_),
    .ZN(_4631_)
  );
  OR2_X1 _5324_ (
    .A1(_4628_),
    .A2(_4631_),
    .ZN(_4632_)
  );
  AND2_X1 _5325_ (
    .A1(divisor[4]),
    .A2(remainder[0]),
    .ZN(_4633_)
  );
  XOR2_X1 _5326_ (
    .A(_4629_),
    .B(_4630_),
    .Z(_4634_)
  );
  AND2_X1 _5327_ (
    .A1(_4633_),
    .A2(_4634_),
    .ZN(_4635_)
  );
  AND2_X1 _5328_ (
    .A1(divisor[2]),
    .A2(remainder[3]),
    .ZN(_4636_)
  );
  AND2_X1 _5329_ (
    .A1(divisor[0]),
    .A2(remainder[5]),
    .ZN(_4637_)
  );
  AND2_X1 _5330_ (
    .A1(divisor[1]),
    .A2(remainder[5]),
    .ZN(_4638_)
  );
  AND2_X1 _5331_ (
    .A1(_4626_),
    .A2(_4637_),
    .ZN(_4639_)
  );
  XOR2_X1 _5332_ (
    .A(_4626_),
    .B(_4637_),
    .Z(_4640_)
  );
  AND2_X1 _5333_ (
    .A1(_4636_),
    .A2(_4640_),
    .ZN(_4641_)
  );
  XOR2_X1 _5334_ (
    .A(_4636_),
    .B(_4640_),
    .Z(_4642_)
  );
  AND2_X1 _5335_ (
    .A1(divisor[4]),
    .A2(remainder[1]),
    .ZN(_4643_)
  );
  AND2_X1 _5336_ (
    .A1(divisor[5]),
    .A2(remainder[0]),
    .ZN(_4644_)
  );
  AND2_X1 _5337_ (
    .A1(divisor[5]),
    .A2(remainder[1]),
    .ZN(_4645_)
  );
  AND2_X1 _5338_ (
    .A1(_4633_),
    .A2(_4645_),
    .ZN(_4646_)
  );
  XOR2_X1 _5339_ (
    .A(_4643_),
    .B(_4644_),
    .Z(_4647_)
  );
  AND2_X1 _5340_ (
    .A1(_4642_),
    .A2(_4647_),
    .ZN(_4648_)
  );
  XOR2_X1 _5341_ (
    .A(_4642_),
    .B(_4647_),
    .Z(_4649_)
  );
  AND2_X1 _5342_ (
    .A1(_4635_),
    .A2(_4649_),
    .ZN(_4650_)
  );
  XOR2_X1 _5343_ (
    .A(_4635_),
    .B(_4649_),
    .Z(_4651_)
  );
  AND2_X1 _5344_ (
    .A1(_4632_),
    .A2(_4651_),
    .ZN(_4652_)
  );
  OR2_X1 _5345_ (
    .A1(_4639_),
    .A2(_4641_),
    .ZN(_4653_)
  );
  AND2_X1 _5346_ (
    .A1(divisor[2]),
    .A2(remainder[4]),
    .ZN(_4654_)
  );
  AND2_X1 _5347_ (
    .A1(divisor[0]),
    .A2(remainder[6]),
    .ZN(_4655_)
  );
  AND2_X1 _5348_ (
    .A1(divisor[1]),
    .A2(remainder[6]),
    .ZN(_4656_)
  );
  AND2_X1 _5349_ (
    .A1(_4638_),
    .A2(_4655_),
    .ZN(_4657_)
  );
  XOR2_X1 _5350_ (
    .A(_4638_),
    .B(_4655_),
    .Z(_4658_)
  );
  AND2_X1 _5351_ (
    .A1(_4654_),
    .A2(_4658_),
    .ZN(_4659_)
  );
  XOR2_X1 _5352_ (
    .A(_4654_),
    .B(_4658_),
    .Z(_4660_)
  );
  AND2_X1 _5353_ (
    .A1(divisor[4]),
    .A2(remainder[2]),
    .ZN(_4661_)
  );
  AND2_X1 _5354_ (
    .A1(divisor[6]),
    .A2(remainder[0]),
    .ZN(_4662_)
  );
  AND2_X1 _5355_ (
    .A1(divisor[6]),
    .A2(remainder[1]),
    .ZN(_4663_)
  );
  AND2_X1 _5356_ (
    .A1(_4644_),
    .A2(_4663_),
    .ZN(_4664_)
  );
  XOR2_X1 _5357_ (
    .A(_4645_),
    .B(_4662_),
    .Z(_4665_)
  );
  AND2_X1 _5358_ (
    .A1(_4661_),
    .A2(_4665_),
    .ZN(_4666_)
  );
  XOR2_X1 _5359_ (
    .A(_4661_),
    .B(_4665_),
    .Z(_4667_)
  );
  AND2_X1 _5360_ (
    .A1(_4646_),
    .A2(_4667_),
    .ZN(_4668_)
  );
  XOR2_X1 _5361_ (
    .A(_4646_),
    .B(_4667_),
    .Z(_4669_)
  );
  AND2_X1 _5362_ (
    .A1(_4660_),
    .A2(_4669_),
    .ZN(_4670_)
  );
  XOR2_X1 _5363_ (
    .A(_4660_),
    .B(_4669_),
    .Z(_4671_)
  );
  AND2_X1 _5364_ (
    .A1(_4648_),
    .A2(_4671_),
    .ZN(_4672_)
  );
  XOR2_X1 _5365_ (
    .A(_4648_),
    .B(_4671_),
    .Z(_4673_)
  );
  AND2_X1 _5366_ (
    .A1(_4650_),
    .A2(_4673_),
    .ZN(_4674_)
  );
  XOR2_X1 _5367_ (
    .A(_4650_),
    .B(_4673_),
    .Z(_4675_)
  );
  AND2_X1 _5368_ (
    .A1(_4653_),
    .A2(_4675_),
    .ZN(_4676_)
  );
  XOR2_X1 _5369_ (
    .A(_4653_),
    .B(_4675_),
    .Z(_4677_)
  );
  AND2_X1 _5370_ (
    .A1(_4652_),
    .A2(_4677_),
    .ZN(_4678_)
  );
  XOR2_X1 _5371_ (
    .A(_4652_),
    .B(_4677_),
    .Z(_4679_)
  );
  AND2_X1 _5372_ (
    .A1(_4622_),
    .A2(_4679_),
    .ZN(_4680_)
  );
  XOR2_X1 _5373_ (
    .A(_4622_),
    .B(_4679_),
    .Z(_4681_)
  );
  XOR2_X1 _5374_ (
    .A(_4623_),
    .B(_4679_),
    .Z(_4682_)
  );
  AND2_X1 _5375_ (
    .A1(divisor[1]),
    .A2(remainder[2]),
    .ZN(_4683_)
  );
  AND2_X1 _5376_ (
    .A1(divisor[0]),
    .A2(remainder[2]),
    .ZN(_4684_)
  );
  AND2_X1 _5377_ (
    .A1(_4627_),
    .A2(_4683_),
    .ZN(_4685_)
  );
  AND2_X1 _5378_ (
    .A1(divisor[2]),
    .A2(remainder[1]),
    .ZN(_4686_)
  );
  XOR2_X1 _5379_ (
    .A(_4627_),
    .B(_4683_),
    .Z(_4687_)
  );
  AND2_X1 _5380_ (
    .A1(_4686_),
    .A2(_4687_),
    .ZN(_4688_)
  );
  OR2_X1 _5381_ (
    .A1(_4685_),
    .A2(_4688_),
    .ZN(_4689_)
  );
  XOR2_X1 _5382_ (
    .A(_4633_),
    .B(_4634_),
    .Z(_4690_)
  );
  AND2_X1 _5383_ (
    .A1(_4689_),
    .A2(_4690_),
    .ZN(_4691_)
  );
  XOR2_X1 _5384_ (
    .A(_4632_),
    .B(_4651_),
    .Z(_4692_)
  );
  AND2_X1 _5385_ (
    .A1(_4691_),
    .A2(_4692_),
    .ZN(_4693_)
  );
  AND2_X1 _5386_ (
    .A1(divisor[3]),
    .A2(remainder[2]),
    .ZN(_4694_)
  );
  XOR2_X1 _5387_ (
    .A(_4691_),
    .B(_4692_),
    .Z(_4695_)
  );
  AND2_X1 _5388_ (
    .A1(_4694_),
    .A2(_4695_),
    .ZN(_4696_)
  );
  OR2_X1 _5389_ (
    .A1(_4693_),
    .A2(_4696_),
    .ZN(_4697_)
  );
  AND2_X1 _5390_ (
    .A1(_4681_),
    .A2(_4697_),
    .ZN(_4698_)
  );
  OR2_X1 _5391_ (
    .A1(_4657_),
    .A2(_4659_),
    .ZN(_4699_)
  );
  OR2_X1 _5392_ (
    .A1(_4668_),
    .A2(_4670_),
    .ZN(_4700_)
  );
  AND2_X1 _5393_ (
    .A1(divisor[2]),
    .A2(remainder[5]),
    .ZN(_0121_)
  );
  AND2_X1 _5394_ (
    .A1(divisor[0]),
    .A2(remainder[7]),
    .ZN(_0122_)
  );
  AND2_X1 _5395_ (
    .A1(divisor[1]),
    .A2(remainder[7]),
    .ZN(_0123_)
  );
  AND2_X1 _5396_ (
    .A1(_4655_),
    .A2(_0123_),
    .ZN(_0124_)
  );
  XOR2_X1 _5397_ (
    .A(_4656_),
    .B(_0122_),
    .Z(_0125_)
  );
  AND2_X1 _5398_ (
    .A1(_0121_),
    .A2(_0125_),
    .ZN(_0126_)
  );
  XOR2_X1 _5399_ (
    .A(_0121_),
    .B(_0125_),
    .Z(_0127_)
  );
  OR2_X1 _5400_ (
    .A1(_4664_),
    .A2(_4666_),
    .ZN(_0128_)
  );
  AND2_X1 _5401_ (
    .A1(divisor[4]),
    .A2(remainder[3]),
    .ZN(_0129_)
  );
  AND2_X1 _5402_ (
    .A1(divisor[5]),
    .A2(remainder[2]),
    .ZN(_0130_)
  );
  AND2_X1 _5403_ (
    .A1(divisor[6]),
    .A2(remainder[2]),
    .ZN(_0131_)
  );
  AND2_X1 _5404_ (
    .A1(_4645_),
    .A2(_0131_),
    .ZN(_0132_)
  );
  XOR2_X1 _5405_ (
    .A(_4663_),
    .B(_0130_),
    .Z(_0133_)
  );
  AND2_X1 _5406_ (
    .A1(_0129_),
    .A2(_0133_),
    .ZN(_0134_)
  );
  XOR2_X1 _5407_ (
    .A(_0129_),
    .B(_0133_),
    .Z(_0135_)
  );
  AND2_X1 _5408_ (
    .A1(_0128_),
    .A2(_0135_),
    .ZN(_0136_)
  );
  XOR2_X1 _5409_ (
    .A(_0128_),
    .B(_0135_),
    .Z(_0137_)
  );
  AND2_X1 _5410_ (
    .A1(_0127_),
    .A2(_0137_),
    .ZN(_0138_)
  );
  XOR2_X1 _5411_ (
    .A(_0127_),
    .B(_0137_),
    .Z(_0139_)
  );
  AND2_X1 _5412_ (
    .A1(_4700_),
    .A2(_0139_),
    .ZN(_0140_)
  );
  XOR2_X1 _5413_ (
    .A(_4700_),
    .B(_0139_),
    .Z(_0141_)
  );
  OR2_X1 _5414_ (
    .A1(_4672_),
    .A2(_4674_),
    .ZN(_0142_)
  );
  XOR2_X1 _5415_ (
    .A(_0141_),
    .B(_0142_),
    .Z(_0143_)
  );
  AND2_X1 _5416_ (
    .A1(_4699_),
    .A2(_0143_),
    .ZN(_0144_)
  );
  XOR2_X1 _5417_ (
    .A(_4699_),
    .B(_0143_),
    .Z(_0145_)
  );
  AND2_X1 _5418_ (
    .A1(_4676_),
    .A2(_0145_),
    .ZN(_0146_)
  );
  XOR2_X1 _5419_ (
    .A(_4676_),
    .B(_0145_),
    .Z(_0147_)
  );
  AND2_X1 _5420_ (
    .A1(divisor[7]),
    .A2(remainder[0]),
    .ZN(_0148_)
  );
  AND2_X1 _5421_ (
    .A1(divisor[3]),
    .A2(remainder[4]),
    .ZN(_0149_)
  );
  AND2_X1 _5422_ (
    .A1(divisor[3]),
    .A2(remainder[0]),
    .ZN(_0150_)
  );
  INV_X1 _5423_ (
    .A(_0150_),
    .ZN(_0151_)
  );
  AND2_X1 _5424_ (
    .A1(divisor[7]),
    .A2(remainder[4]),
    .ZN(_0152_)
  );
  AND2_X1 _5425_ (
    .A1(_0150_),
    .A2(_0152_),
    .ZN(_0153_)
  );
  XOR2_X1 _5426_ (
    .A(_0148_),
    .B(_0149_),
    .Z(_0154_)
  );
  AND2_X1 _5427_ (
    .A1(_0147_),
    .A2(_0154_),
    .ZN(_0155_)
  );
  XOR2_X1 _5428_ (
    .A(_0147_),
    .B(_0154_),
    .Z(_0156_)
  );
  OR2_X1 _5429_ (
    .A1(_4678_),
    .A2(_4680_),
    .ZN(_0157_)
  );
  AND2_X1 _5430_ (
    .A1(_0156_),
    .A2(_0157_),
    .ZN(_0158_)
  );
  XOR2_X1 _5431_ (
    .A(_0156_),
    .B(_0157_),
    .Z(_0159_)
  );
  AND2_X1 _5432_ (
    .A1(_4698_),
    .A2(_0159_),
    .ZN(_0160_)
  );
  XOR2_X1 _5433_ (
    .A(_4698_),
    .B(_0159_),
    .Z(_0161_)
  );
  XOR2_X1 _5434_ (
    .A(_4682_),
    .B(_4697_),
    .Z(_0162_)
  );
  XOR2_X1 _5435_ (
    .A(_4694_),
    .B(_4695_),
    .Z(_0163_)
  );
  AND2_X1 _5436_ (
    .A1(divisor[1]),
    .A2(remainder[1]),
    .ZN(_0164_)
  );
  AND2_X1 _5437_ (
    .A1(divisor[0]),
    .A2(remainder[1]),
    .ZN(_0165_)
  );
  AND2_X1 _5438_ (
    .A1(_4684_),
    .A2(_0164_),
    .ZN(_0166_)
  );
  AND2_X1 _5439_ (
    .A1(divisor[2]),
    .A2(remainder[0]),
    .ZN(_0167_)
  );
  XOR2_X1 _5440_ (
    .A(_4684_),
    .B(_0164_),
    .Z(_0168_)
  );
  AND2_X1 _5441_ (
    .A1(_0167_),
    .A2(_0168_),
    .ZN(_0169_)
  );
  OR2_X1 _5442_ (
    .A1(_0166_),
    .A2(_0169_),
    .ZN(_0170_)
  );
  XOR2_X1 _5443_ (
    .A(_4686_),
    .B(_4687_),
    .Z(_0171_)
  );
  AND2_X1 _5444_ (
    .A1(_0170_),
    .A2(_0171_),
    .ZN(_0172_)
  );
  XOR2_X1 _5445_ (
    .A(_4689_),
    .B(_4690_),
    .Z(_0173_)
  );
  AND2_X1 _5446_ (
    .A1(_0172_),
    .A2(_0173_),
    .ZN(_0174_)
  );
  AND2_X1 _5447_ (
    .A1(divisor[3]),
    .A2(remainder[1]),
    .ZN(_0175_)
  );
  XOR2_X1 _5448_ (
    .A(_0172_),
    .B(_0173_),
    .Z(_0176_)
  );
  AND2_X1 _5449_ (
    .A1(_0175_),
    .A2(_0176_),
    .ZN(_0177_)
  );
  OR2_X1 _5450_ (
    .A1(_0174_),
    .A2(_0177_),
    .ZN(_0178_)
  );
  AND2_X1 _5451_ (
    .A1(_0163_),
    .A2(_0178_),
    .ZN(_0179_)
  );
  INV_X1 _5452_ (
    .A(_0179_),
    .ZN(_0180_)
  );
  OR2_X1 _5453_ (
    .A1(_0162_),
    .A2(_0180_),
    .ZN(_0181_)
  );
  XOR2_X1 _5454_ (
    .A(_0163_),
    .B(_0178_),
    .Z(_0182_)
  );
  INV_X1 _5455_ (
    .A(_0182_),
    .ZN(_0183_)
  );
  XOR2_X1 _5456_ (
    .A(_0175_),
    .B(_0176_),
    .Z(_0184_)
  );
  AND2_X1 _5457_ (
    .A1(divisor[1]),
    .A2(remainder[0]),
    .ZN(_0185_)
  );
  AND2_X1 _5458_ (
    .A1(divisor[0]),
    .A2(remainder[0]),
    .ZN(_0186_)
  );
  AND2_X1 _5459_ (
    .A1(_0164_),
    .A2(_0186_),
    .ZN(_0187_)
  );
  XOR2_X1 _5460_ (
    .A(_0167_),
    .B(_0168_),
    .Z(_0188_)
  );
  AND2_X1 _5461_ (
    .A1(_0187_),
    .A2(_0188_),
    .ZN(_0189_)
  );
  XOR2_X1 _5462_ (
    .A(_0170_),
    .B(_0171_),
    .Z(_0190_)
  );
  AND2_X1 _5463_ (
    .A1(_0189_),
    .A2(_0190_),
    .ZN(_0191_)
  );
  XOR2_X1 _5464_ (
    .A(_0189_),
    .B(_0190_),
    .Z(_0192_)
  );
  AND2_X1 _5465_ (
    .A1(_0150_),
    .A2(_0192_),
    .ZN(_0193_)
  );
  OR2_X1 _5466_ (
    .A1(_0191_),
    .A2(_0193_),
    .ZN(_0194_)
  );
  AND2_X1 _5467_ (
    .A1(_0184_),
    .A2(_0194_),
    .ZN(_0195_)
  );
  INV_X1 _5468_ (
    .A(_0195_),
    .ZN(_0196_)
  );
  OR2_X1 _5469_ (
    .A1(_0183_),
    .A2(_0196_),
    .ZN(_0197_)
  );
  XOR2_X1 _5470_ (
    .A(_0162_),
    .B(_0179_),
    .Z(_0198_)
  );
  OR2_X1 _5471_ (
    .A1(_0197_),
    .A2(_0198_),
    .ZN(_0199_)
  );
  AND2_X1 _5472_ (
    .A1(_0181_),
    .A2(_0199_),
    .ZN(_0200_)
  );
  INV_X1 _5473_ (
    .A(_0200_),
    .ZN(_0201_)
  );
  AND2_X1 _5474_ (
    .A1(_0161_),
    .A2(_0201_),
    .ZN(_0202_)
  );
  XOR2_X1 _5475_ (
    .A(_0161_),
    .B(_0200_),
    .Z(_0203_)
  );
  INV_X1 _5476_ (
    .A(_0203_),
    .ZN(_0204_)
  );
  AND2_X1 _5477_ (
    .A1(remainder[40]),
    .A2(_0204_),
    .ZN(_0205_)
  );
  OR2_X1 _5478_ (
    .A1(_3165_),
    .A2(_0203_),
    .ZN(_0206_)
  );
  XOR2_X1 _5479_ (
    .A(_0197_),
    .B(_0198_),
    .Z(_0207_)
  );
  AND2_X1 _5480_ (
    .A1(remainder[39]),
    .A2(_0207_),
    .ZN(_0208_)
  );
  INV_X1 _5481_ (
    .A(_0208_),
    .ZN(_0209_)
  );
  XOR2_X1 _5482_ (
    .A(_0182_),
    .B(_0195_),
    .Z(_0210_)
  );
  AND2_X1 _5483_ (
    .A1(remainder[38]),
    .A2(_0210_),
    .ZN(_0211_)
  );
  INV_X1 _5484_ (
    .A(_0211_),
    .ZN(_0212_)
  );
  XOR2_X1 _5485_ (
    .A(remainder[38]),
    .B(_0210_),
    .Z(_0213_)
  );
  INV_X1 _5486_ (
    .A(_0213_),
    .ZN(_0214_)
  );
  XOR2_X1 _5487_ (
    .A(_0184_),
    .B(_0194_),
    .Z(_0215_)
  );
  AND2_X1 _5488_ (
    .A1(remainder[37]),
    .A2(_0215_),
    .ZN(_0216_)
  );
  INV_X1 _5489_ (
    .A(_0216_),
    .ZN(_0217_)
  );
  XOR2_X1 _5490_ (
    .A(remainder[37]),
    .B(_0215_),
    .Z(_0218_)
  );
  XOR2_X1 _5491_ (
    .A(_3187_),
    .B(_0215_),
    .Z(_0219_)
  );
  XOR2_X1 _5492_ (
    .A(_0150_),
    .B(_0192_),
    .Z(_0220_)
  );
  XOR2_X1 _5493_ (
    .A(_0151_),
    .B(_0192_),
    .Z(_0221_)
  );
  AND2_X1 _5494_ (
    .A1(remainder[36]),
    .A2(_0220_),
    .ZN(_0222_)
  );
  INV_X1 _5495_ (
    .A(_0222_),
    .ZN(_0223_)
  );
  AND2_X1 _5496_ (
    .A1(_3198_),
    .A2(_0221_),
    .ZN(_0224_)
  );
  OR2_X1 _5497_ (
    .A1(remainder[36]),
    .A2(_0220_),
    .ZN(_0225_)
  );
  XOR2_X1 _5498_ (
    .A(_0187_),
    .B(_0188_),
    .Z(_0226_)
  );
  AND2_X1 _5499_ (
    .A1(remainder[35]),
    .A2(_0226_),
    .ZN(_0227_)
  );
  INV_X1 _5500_ (
    .A(_0227_),
    .ZN(_0228_)
  );
  XOR2_X1 _5501_ (
    .A(_0165_),
    .B(_0185_),
    .Z(_0229_)
  );
  AND2_X1 _5502_ (
    .A1(remainder[34]),
    .A2(_0229_),
    .ZN(_0230_)
  );
  AND2_X1 _5503_ (
    .A1(remainder[33]),
    .A2(_0186_),
    .ZN(_0231_)
  );
  INV_X1 _5504_ (
    .A(_0231_),
    .ZN(_0232_)
  );
  XOR2_X1 _5505_ (
    .A(remainder[34]),
    .B(_0229_),
    .Z(_0233_)
  );
  AND2_X1 _5506_ (
    .A1(_0231_),
    .A2(_0233_),
    .ZN(_0234_)
  );
  INV_X1 _5507_ (
    .A(_0234_),
    .ZN(_0235_)
  );
  OR2_X1 _5508_ (
    .A1(_0230_),
    .A2(_0234_),
    .ZN(_0236_)
  );
  INV_X1 _5509_ (
    .A(_0236_),
    .ZN(_0237_)
  );
  XOR2_X1 _5510_ (
    .A(remainder[35]),
    .B(_0226_),
    .Z(_0238_)
  );
  INV_X1 _5511_ (
    .A(_0238_),
    .ZN(_0239_)
  );
  AND2_X1 _5512_ (
    .A1(_0236_),
    .A2(_0238_),
    .ZN(_0240_)
  );
  OR2_X1 _5513_ (
    .A1(_0237_),
    .A2(_0239_),
    .ZN(_0241_)
  );
  AND2_X1 _5514_ (
    .A1(_0228_),
    .A2(_0241_),
    .ZN(_0242_)
  );
  OR2_X1 _5515_ (
    .A1(_0227_),
    .A2(_0240_),
    .ZN(_0243_)
  );
  AND2_X1 _5516_ (
    .A1(_0225_),
    .A2(_0243_),
    .ZN(_0244_)
  );
  OR2_X1 _5517_ (
    .A1(_0224_),
    .A2(_0242_),
    .ZN(_0245_)
  );
  AND2_X1 _5518_ (
    .A1(_0223_),
    .A2(_0245_),
    .ZN(_0246_)
  );
  OR2_X1 _5519_ (
    .A1(_0222_),
    .A2(_0244_),
    .ZN(_0247_)
  );
  AND2_X1 _5520_ (
    .A1(_0218_),
    .A2(_0247_),
    .ZN(_0248_)
  );
  OR2_X1 _5521_ (
    .A1(_0219_),
    .A2(_0246_),
    .ZN(_0249_)
  );
  AND2_X1 _5522_ (
    .A1(_0217_),
    .A2(_0249_),
    .ZN(_0250_)
  );
  OR2_X1 _5523_ (
    .A1(_0216_),
    .A2(_0248_),
    .ZN(_0251_)
  );
  AND2_X1 _5524_ (
    .A1(_0213_),
    .A2(_0251_),
    .ZN(_0252_)
  );
  OR2_X1 _5525_ (
    .A1(_0214_),
    .A2(_0250_),
    .ZN(_0253_)
  );
  AND2_X1 _5526_ (
    .A1(_0212_),
    .A2(_0253_),
    .ZN(_0254_)
  );
  OR2_X1 _5527_ (
    .A1(_0211_),
    .A2(_0252_),
    .ZN(_0255_)
  );
  XOR2_X1 _5528_ (
    .A(remainder[39]),
    .B(_0207_),
    .Z(_0256_)
  );
  XOR2_X1 _5529_ (
    .A(_3176_),
    .B(_0207_),
    .Z(_0257_)
  );
  AND2_X1 _5530_ (
    .A1(_0255_),
    .A2(_0256_),
    .ZN(_0258_)
  );
  OR2_X1 _5531_ (
    .A1(_0254_),
    .A2(_0257_),
    .ZN(_0259_)
  );
  AND2_X1 _5532_ (
    .A1(_0209_),
    .A2(_0259_),
    .ZN(_0260_)
  );
  OR2_X1 _5533_ (
    .A1(_0208_),
    .A2(_0258_),
    .ZN(_0261_)
  );
  XOR2_X1 _5534_ (
    .A(_3165_),
    .B(_0203_),
    .Z(_0262_)
  );
  XOR2_X1 _5535_ (
    .A(remainder[40]),
    .B(_0203_),
    .Z(_0263_)
  );
  AND2_X1 _5536_ (
    .A1(_0261_),
    .A2(_0262_),
    .ZN(_0264_)
  );
  OR2_X1 _5537_ (
    .A1(_0260_),
    .A2(_0263_),
    .ZN(_0265_)
  );
  AND2_X1 _5538_ (
    .A1(_0206_),
    .A2(_0265_),
    .ZN(_0266_)
  );
  OR2_X1 _5539_ (
    .A1(_0205_),
    .A2(_0264_),
    .ZN(_0267_)
  );
  AND2_X1 _5540_ (
    .A1(divisor[3]),
    .A2(remainder[5]),
    .ZN(_0268_)
  );
  AND2_X1 _5541_ (
    .A1(divisor[8]),
    .A2(remainder[0]),
    .ZN(_0269_)
  );
  AND2_X1 _5542_ (
    .A1(divisor[7]),
    .A2(remainder[1]),
    .ZN(_0270_)
  );
  AND2_X1 _5543_ (
    .A1(divisor[8]),
    .A2(remainder[1]),
    .ZN(_0271_)
  );
  AND2_X1 _5544_ (
    .A1(_0148_),
    .A2(_0271_),
    .ZN(_0272_)
  );
  XOR2_X1 _5545_ (
    .A(_0269_),
    .B(_0270_),
    .Z(_0273_)
  );
  AND2_X1 _5546_ (
    .A1(_0268_),
    .A2(_0273_),
    .ZN(_0274_)
  );
  XOR2_X1 _5547_ (
    .A(_0268_),
    .B(_0273_),
    .Z(_0275_)
  );
  AND2_X1 _5548_ (
    .A1(_0153_),
    .A2(_0275_),
    .ZN(_0276_)
  );
  XOR2_X1 _5549_ (
    .A(_0153_),
    .B(_0275_),
    .Z(_0277_)
  );
  AND2_X1 _5550_ (
    .A1(_4674_),
    .A2(_0141_),
    .ZN(_0278_)
  );
  OR2_X1 _5551_ (
    .A1(_0144_),
    .A2(_0278_),
    .ZN(_0279_)
  );
  OR2_X1 _5552_ (
    .A1(_0124_),
    .A2(_0126_),
    .ZN(_0280_)
  );
  AND2_X1 _5553_ (
    .A1(_4672_),
    .A2(_0141_),
    .ZN(_0281_)
  );
  OR2_X1 _5554_ (
    .A1(_0136_),
    .A2(_0138_),
    .ZN(_0282_)
  );
  OR2_X1 _5555_ (
    .A1(_0132_),
    .A2(_0134_),
    .ZN(_0283_)
  );
  AND2_X1 _5556_ (
    .A1(divisor[4]),
    .A2(remainder[4]),
    .ZN(_0284_)
  );
  AND2_X1 _5557_ (
    .A1(divisor[5]),
    .A2(remainder[3]),
    .ZN(_0285_)
  );
  AND2_X1 _5558_ (
    .A1(divisor[6]),
    .A2(remainder[3]),
    .ZN(_0286_)
  );
  AND2_X1 _5559_ (
    .A1(_0131_),
    .A2(_0285_),
    .ZN(_0287_)
  );
  XOR2_X1 _5560_ (
    .A(_0131_),
    .B(_0285_),
    .Z(_0288_)
  );
  AND2_X1 _5561_ (
    .A1(_0284_),
    .A2(_0288_),
    .ZN(_0289_)
  );
  XOR2_X1 _5562_ (
    .A(_0284_),
    .B(_0288_),
    .Z(_0290_)
  );
  AND2_X1 _5563_ (
    .A1(_0283_),
    .A2(_0290_),
    .ZN(_0291_)
  );
  XOR2_X1 _5564_ (
    .A(_0283_),
    .B(_0290_),
    .Z(_0292_)
  );
  AND2_X1 _5565_ (
    .A1(divisor[2]),
    .A2(remainder[6]),
    .ZN(_0293_)
  );
  AND2_X1 _5566_ (
    .A1(remainder[32]),
    .A2(divisor[1]),
    .ZN(_0294_)
  );
  AND2_X1 _5567_ (
    .A1(remainder[32]),
    .A2(divisor[0]),
    .ZN(_0295_)
  );
  AND2_X1 _5568_ (
    .A1(divisor[1]),
    .A2(_0295_),
    .ZN(_0296_)
  );
  INV_X1 _5569_ (
    .A(_0296_),
    .ZN(_0297_)
  );
  AND2_X1 _5570_ (
    .A1(_0123_),
    .A2(_0295_),
    .ZN(_0298_)
  );
  XOR2_X1 _5571_ (
    .A(_0123_),
    .B(_0295_),
    .Z(_0299_)
  );
  AND2_X1 _5572_ (
    .A1(_0293_),
    .A2(_0299_),
    .ZN(_0300_)
  );
  XOR2_X1 _5573_ (
    .A(_0293_),
    .B(_0299_),
    .Z(_0301_)
  );
  AND2_X1 _5574_ (
    .A1(_0292_),
    .A2(_0301_),
    .ZN(_0302_)
  );
  XOR2_X1 _5575_ (
    .A(_0292_),
    .B(_0301_),
    .Z(_0303_)
  );
  AND2_X1 _5576_ (
    .A1(_0282_),
    .A2(_0303_),
    .ZN(_0304_)
  );
  XOR2_X1 _5577_ (
    .A(_0282_),
    .B(_0303_),
    .Z(_0305_)
  );
  AND2_X1 _5578_ (
    .A1(_0140_),
    .A2(_0305_),
    .ZN(_0306_)
  );
  XOR2_X1 _5579_ (
    .A(_0140_),
    .B(_0305_),
    .Z(_0307_)
  );
  AND2_X1 _5580_ (
    .A1(_0281_),
    .A2(_0307_),
    .ZN(_0308_)
  );
  XOR2_X1 _5581_ (
    .A(_0281_),
    .B(_0307_),
    .Z(_0309_)
  );
  AND2_X1 _5582_ (
    .A1(_0280_),
    .A2(_0309_),
    .ZN(_0310_)
  );
  XOR2_X1 _5583_ (
    .A(_0280_),
    .B(_0309_),
    .Z(_0311_)
  );
  AND2_X1 _5584_ (
    .A1(_0279_),
    .A2(_0311_),
    .ZN(_0312_)
  );
  XOR2_X1 _5585_ (
    .A(_0279_),
    .B(_0311_),
    .Z(_0313_)
  );
  AND2_X1 _5586_ (
    .A1(_0277_),
    .A2(_0313_),
    .ZN(_0314_)
  );
  XOR2_X1 _5587_ (
    .A(_0277_),
    .B(_0313_),
    .Z(_0315_)
  );
  OR2_X1 _5588_ (
    .A1(_0146_),
    .A2(_0155_),
    .ZN(_0316_)
  );
  AND2_X1 _5589_ (
    .A1(_0315_),
    .A2(_0316_),
    .ZN(_0317_)
  );
  XOR2_X1 _5590_ (
    .A(_0315_),
    .B(_0316_),
    .Z(_0318_)
  );
  AND2_X1 _5591_ (
    .A1(_0160_),
    .A2(_0318_),
    .ZN(_0319_)
  );
  AND2_X1 _5592_ (
    .A1(_0158_),
    .A2(_0318_),
    .ZN(_0320_)
  );
  INV_X1 _5593_ (
    .A(_0320_),
    .ZN(_0321_)
  );
  OR2_X1 _5594_ (
    .A1(_0158_),
    .A2(_0160_),
    .ZN(_0322_)
  );
  XOR2_X1 _5595_ (
    .A(_0318_),
    .B(_0322_),
    .Z(_0323_)
  );
  AND2_X1 _5596_ (
    .A1(_0202_),
    .A2(_0323_),
    .ZN(_0324_)
  );
  XOR2_X1 _5597_ (
    .A(_0202_),
    .B(_0323_),
    .Z(_0325_)
  );
  AND2_X1 _5598_ (
    .A1(remainder[41]),
    .A2(_0325_),
    .ZN(_0326_)
  );
  INV_X1 _5599_ (
    .A(_0326_),
    .ZN(_0327_)
  );
  XOR2_X1 _5600_ (
    .A(remainder[41]),
    .B(_0325_),
    .Z(_0328_)
  );
  XOR2_X1 _5601_ (
    .A(_3155_),
    .B(_0325_),
    .Z(_0329_)
  );
  OR2_X1 _5602_ (
    .A1(_0267_),
    .A2(_0328_),
    .ZN(_0330_)
  );
  AND2_X1 _5603_ (
    .A1(_0267_),
    .A2(_0328_),
    .ZN(_0331_)
  );
  OR2_X1 _5604_ (
    .A1(_0266_),
    .A2(_0329_),
    .ZN(_0332_)
  );
  AND2_X1 _5605_ (
    .A1(_4613_),
    .A2(_0330_),
    .ZN(_0333_)
  );
  AND2_X1 _5606_ (
    .A1(_0332_),
    .A2(_0333_),
    .ZN(_0334_)
  );
  OR2_X1 _5607_ (
    .A1(_4621_),
    .A2(_0334_),
    .ZN(_0335_)
  );
  OR2_X1 _5608_ (
    .A1(_4620_),
    .A2(_0335_),
    .ZN(_0336_)
  );
  AND2_X1 _5609_ (
    .A1(_3911_),
    .A2(_0336_),
    .ZN(_0054_)
  );
  OR2_X1 _5610_ (
    .A1(remainder[33]),
    .A2(_4393_),
    .ZN(_0337_)
  );
  OR2_X1 _5611_ (
    .A1(_4392_),
    .A2(_4438_),
    .ZN(_0338_)
  );
  AND2_X1 _5612_ (
    .A1(_3678_),
    .A2(_0338_),
    .ZN(_0339_)
  );
  AND2_X1 _5613_ (
    .A1(_0337_),
    .A2(_0339_),
    .ZN(_0340_)
  );
  AND2_X1 _5614_ (
    .A1(remainder[34]),
    .A2(_4610_),
    .ZN(_0341_)
  );
  AND2_X1 _5615_ (
    .A1(_0327_),
    .A2(_0332_),
    .ZN(_0342_)
  );
  OR2_X1 _5616_ (
    .A1(_0326_),
    .A2(_0331_),
    .ZN(_0343_)
  );
  OR2_X1 _5617_ (
    .A1(_0319_),
    .A2(_0324_),
    .ZN(_0344_)
  );
  OR2_X1 _5618_ (
    .A1(_0276_),
    .A2(_0314_),
    .ZN(_0345_)
  );
  AND2_X1 _5619_ (
    .A1(divisor[3]),
    .A2(remainder[6]),
    .ZN(_0346_)
  );
  AND2_X1 _5620_ (
    .A1(divisor[7]),
    .A2(remainder[2]),
    .ZN(_0347_)
  );
  AND2_X1 _5621_ (
    .A1(divisor[9]),
    .A2(remainder[0]),
    .ZN(_0348_)
  );
  AND2_X1 _5622_ (
    .A1(divisor[9]),
    .A2(remainder[1]),
    .ZN(_0349_)
  );
  AND2_X1 _5623_ (
    .A1(_0269_),
    .A2(_0349_),
    .ZN(_0350_)
  );
  XOR2_X1 _5624_ (
    .A(_0271_),
    .B(_0348_),
    .Z(_0351_)
  );
  AND2_X1 _5625_ (
    .A1(_0347_),
    .A2(_0351_),
    .ZN(_0352_)
  );
  XOR2_X1 _5626_ (
    .A(_0347_),
    .B(_0351_),
    .Z(_0353_)
  );
  AND2_X1 _5627_ (
    .A1(_0272_),
    .A2(_0353_),
    .ZN(_0354_)
  );
  XOR2_X1 _5628_ (
    .A(_0272_),
    .B(_0353_),
    .Z(_0355_)
  );
  AND2_X1 _5629_ (
    .A1(_0346_),
    .A2(_0355_),
    .ZN(_0356_)
  );
  XOR2_X1 _5630_ (
    .A(_0346_),
    .B(_0355_),
    .Z(_0357_)
  );
  AND2_X1 _5631_ (
    .A1(_0274_),
    .A2(_0357_),
    .ZN(_0358_)
  );
  XOR2_X1 _5632_ (
    .A(_0274_),
    .B(_0357_),
    .Z(_0359_)
  );
  OR2_X1 _5633_ (
    .A1(_0308_),
    .A2(_0310_),
    .ZN(_0360_)
  );
  OR2_X1 _5634_ (
    .A1(_0298_),
    .A2(_0300_),
    .ZN(_0361_)
  );
  OR2_X1 _5635_ (
    .A1(_0291_),
    .A2(_0302_),
    .ZN(_0362_)
  );
  OR2_X1 _5636_ (
    .A1(_0287_),
    .A2(_0289_),
    .ZN(_0363_)
  );
  AND2_X1 _5637_ (
    .A1(divisor[4]),
    .A2(remainder[5]),
    .ZN(_0364_)
  );
  AND2_X1 _5638_ (
    .A1(divisor[5]),
    .A2(remainder[4]),
    .ZN(_0365_)
  );
  AND2_X1 _5639_ (
    .A1(divisor[6]),
    .A2(remainder[4]),
    .ZN(_0366_)
  );
  AND2_X1 _5640_ (
    .A1(_0286_),
    .A2(_0365_),
    .ZN(_0367_)
  );
  XOR2_X1 _5641_ (
    .A(_0286_),
    .B(_0365_),
    .Z(_0368_)
  );
  AND2_X1 _5642_ (
    .A1(_0364_),
    .A2(_0368_),
    .ZN(_0369_)
  );
  XOR2_X1 _5643_ (
    .A(_0364_),
    .B(_0368_),
    .Z(_0370_)
  );
  AND2_X1 _5644_ (
    .A1(_0363_),
    .A2(_0370_),
    .ZN(_0371_)
  );
  XOR2_X1 _5645_ (
    .A(_0363_),
    .B(_0370_),
    .Z(_0372_)
  );
  OR2_X1 _5646_ (
    .A1(_0294_),
    .A2(_0295_),
    .ZN(_0373_)
  );
  AND2_X1 _5647_ (
    .A1(_0297_),
    .A2(_0373_),
    .ZN(_0374_)
  );
  AND2_X1 _5648_ (
    .A1(divisor[2]),
    .A2(remainder[7]),
    .ZN(_0375_)
  );
  AND2_X1 _5649_ (
    .A1(divisor[2]),
    .A2(_0374_),
    .ZN(_0376_)
  );
  INV_X1 _5650_ (
    .A(_0376_),
    .ZN(_0377_)
  );
  AND2_X1 _5651_ (
    .A1(_0374_),
    .A2(_0375_),
    .ZN(_0378_)
  );
  XOR2_X1 _5652_ (
    .A(_0374_),
    .B(_0375_),
    .Z(_0379_)
  );
  AND2_X1 _5653_ (
    .A1(_0372_),
    .A2(_0379_),
    .ZN(_0380_)
  );
  XOR2_X1 _5654_ (
    .A(_0372_),
    .B(_0379_),
    .Z(_0381_)
  );
  AND2_X1 _5655_ (
    .A1(_0362_),
    .A2(_0381_),
    .ZN(_0382_)
  );
  XOR2_X1 _5656_ (
    .A(_0362_),
    .B(_0381_),
    .Z(_0383_)
  );
  AND2_X1 _5657_ (
    .A1(_0304_),
    .A2(_0383_),
    .ZN(_0384_)
  );
  XOR2_X1 _5658_ (
    .A(_0304_),
    .B(_0383_),
    .Z(_0385_)
  );
  AND2_X1 _5659_ (
    .A1(_0306_),
    .A2(_0385_),
    .ZN(_0386_)
  );
  XOR2_X1 _5660_ (
    .A(_0306_),
    .B(_0385_),
    .Z(_0387_)
  );
  AND2_X1 _5661_ (
    .A1(_0361_),
    .A2(_0387_),
    .ZN(_0388_)
  );
  XOR2_X1 _5662_ (
    .A(_0361_),
    .B(_0387_),
    .Z(_0389_)
  );
  AND2_X1 _5663_ (
    .A1(_0360_),
    .A2(_0389_),
    .ZN(_0390_)
  );
  XOR2_X1 _5664_ (
    .A(_0360_),
    .B(_0389_),
    .Z(_0391_)
  );
  AND2_X1 _5665_ (
    .A1(_0359_),
    .A2(_0391_),
    .ZN(_0392_)
  );
  XOR2_X1 _5666_ (
    .A(_0359_),
    .B(_0391_),
    .Z(_0393_)
  );
  AND2_X1 _5667_ (
    .A1(_0345_),
    .A2(_0393_),
    .ZN(_0394_)
  );
  XOR2_X1 _5668_ (
    .A(_0345_),
    .B(_0393_),
    .Z(_0395_)
  );
  AND2_X1 _5669_ (
    .A1(_0312_),
    .A2(_0395_),
    .ZN(_0396_)
  );
  XOR2_X1 _5670_ (
    .A(_0312_),
    .B(_0395_),
    .Z(_0397_)
  );
  AND2_X1 _5671_ (
    .A1(_0317_),
    .A2(_0397_),
    .ZN(_0398_)
  );
  XOR2_X1 _5672_ (
    .A(_0317_),
    .B(_0397_),
    .Z(_0399_)
  );
  AND2_X1 _5673_ (
    .A1(_0320_),
    .A2(_0399_),
    .ZN(_0400_)
  );
  XOR2_X1 _5674_ (
    .A(_0320_),
    .B(_0399_),
    .Z(_0401_)
  );
  XOR2_X1 _5675_ (
    .A(_0321_),
    .B(_0399_),
    .Z(_0402_)
  );
  AND2_X1 _5676_ (
    .A1(_0344_),
    .A2(_0401_),
    .ZN(_0403_)
  );
  XOR2_X1 _5677_ (
    .A(_0344_),
    .B(_0402_),
    .Z(_0404_)
  );
  XOR2_X1 _5678_ (
    .A(_0344_),
    .B(_0401_),
    .Z(_0405_)
  );
  AND2_X1 _5679_ (
    .A1(remainder[42]),
    .A2(_0405_),
    .ZN(_0406_)
  );
  OR2_X1 _5680_ (
    .A1(_3144_),
    .A2(_0404_),
    .ZN(_0407_)
  );
  AND2_X1 _5681_ (
    .A1(_3144_),
    .A2(_0404_),
    .ZN(_0408_)
  );
  INV_X1 _5682_ (
    .A(_0408_),
    .ZN(_0409_)
  );
  AND2_X1 _5683_ (
    .A1(_0407_),
    .A2(_0409_),
    .ZN(_0410_)
  );
  XOR2_X1 _5684_ (
    .A(_0343_),
    .B(_0410_),
    .Z(_0411_)
  );
  AND2_X1 _5685_ (
    .A1(_4613_),
    .A2(_0411_),
    .ZN(_0412_)
  );
  OR2_X1 _5686_ (
    .A1(_0341_),
    .A2(_0412_),
    .ZN(_0413_)
  );
  OR2_X1 _5687_ (
    .A1(_0340_),
    .A2(_0413_),
    .ZN(_0414_)
  );
  AND2_X1 _5688_ (
    .A1(_3911_),
    .A2(_0414_),
    .ZN(_0055_)
  );
  OR2_X1 _5689_ (
    .A1(remainder[34]),
    .A2(_4393_),
    .ZN(_0415_)
  );
  OR2_X1 _5690_ (
    .A1(_4392_),
    .A2(_4441_),
    .ZN(_0416_)
  );
  AND2_X1 _5691_ (
    .A1(_3678_),
    .A2(_0416_),
    .ZN(_0417_)
  );
  AND2_X1 _5692_ (
    .A1(_0415_),
    .A2(_0417_),
    .ZN(_0418_)
  );
  AND2_X1 _5693_ (
    .A1(remainder[35]),
    .A2(_4610_),
    .ZN(_0419_)
  );
  OR2_X1 _5694_ (
    .A1(_0394_),
    .A2(_0396_),
    .ZN(_0420_)
  );
  OR2_X1 _5695_ (
    .A1(_0358_),
    .A2(_0392_),
    .ZN(_0421_)
  );
  AND2_X1 _5696_ (
    .A1(divisor[3]),
    .A2(remainder[7]),
    .ZN(_0422_)
  );
  AND2_X1 _5697_ (
    .A1(divisor[10]),
    .A2(remainder[0]),
    .ZN(_0423_)
  );
  OR2_X1 _5698_ (
    .A1(_0350_),
    .A2(_0352_),
    .ZN(_0424_)
  );
  AND2_X1 _5699_ (
    .A1(divisor[7]),
    .A2(remainder[3]),
    .ZN(_0425_)
  );
  AND2_X1 _5700_ (
    .A1(divisor[8]),
    .A2(remainder[2]),
    .ZN(_0426_)
  );
  AND2_X1 _5701_ (
    .A1(divisor[9]),
    .A2(remainder[2]),
    .ZN(_0427_)
  );
  AND2_X1 _5702_ (
    .A1(_0271_),
    .A2(_0427_),
    .ZN(_0428_)
  );
  XOR2_X1 _5703_ (
    .A(_0349_),
    .B(_0426_),
    .Z(_0429_)
  );
  AND2_X1 _5704_ (
    .A1(_0425_),
    .A2(_0429_),
    .ZN(_0430_)
  );
  XOR2_X1 _5705_ (
    .A(_0425_),
    .B(_0429_),
    .Z(_0431_)
  );
  AND2_X1 _5706_ (
    .A1(_0424_),
    .A2(_0431_),
    .ZN(_0432_)
  );
  XOR2_X1 _5707_ (
    .A(_0424_),
    .B(_0431_),
    .Z(_0433_)
  );
  AND2_X1 _5708_ (
    .A1(_0423_),
    .A2(_0433_),
    .ZN(_0434_)
  );
  XOR2_X1 _5709_ (
    .A(_0423_),
    .B(_0433_),
    .Z(_0435_)
  );
  AND2_X1 _5710_ (
    .A1(_0422_),
    .A2(_0435_),
    .ZN(_0436_)
  );
  XOR2_X1 _5711_ (
    .A(_0422_),
    .B(_0435_),
    .Z(_0437_)
  );
  AND2_X1 _5712_ (
    .A1(_0356_),
    .A2(_0437_),
    .ZN(_0438_)
  );
  XOR2_X1 _5713_ (
    .A(_0356_),
    .B(_0437_),
    .Z(_0439_)
  );
  OR2_X1 _5714_ (
    .A1(_0386_),
    .A2(_0388_),
    .ZN(_0440_)
  );
  OR2_X1 _5715_ (
    .A1(_0296_),
    .A2(_0378_),
    .ZN(_0441_)
  );
  OR2_X1 _5716_ (
    .A1(_0371_),
    .A2(_0380_),
    .ZN(_0442_)
  );
  OR2_X1 _5717_ (
    .A1(_0367_),
    .A2(_0369_),
    .ZN(_0443_)
  );
  AND2_X1 _5718_ (
    .A1(divisor[4]),
    .A2(remainder[6]),
    .ZN(_0444_)
  );
  AND2_X1 _5719_ (
    .A1(divisor[5]),
    .A2(remainder[5]),
    .ZN(_0445_)
  );
  AND2_X1 _5720_ (
    .A1(divisor[6]),
    .A2(remainder[5]),
    .ZN(_0446_)
  );
  AND2_X1 _5721_ (
    .A1(_0366_),
    .A2(_0445_),
    .ZN(_0447_)
  );
  XOR2_X1 _5722_ (
    .A(_0366_),
    .B(_0445_),
    .Z(_0448_)
  );
  AND2_X1 _5723_ (
    .A1(_0444_),
    .A2(_0448_),
    .ZN(_0449_)
  );
  XOR2_X1 _5724_ (
    .A(_0444_),
    .B(_0448_),
    .Z(_0450_)
  );
  AND2_X1 _5725_ (
    .A1(_0443_),
    .A2(_0450_),
    .ZN(_0451_)
  );
  XOR2_X1 _5726_ (
    .A(_0443_),
    .B(_0450_),
    .Z(_0452_)
  );
  AND2_X1 _5727_ (
    .A1(remainder[32]),
    .A2(divisor[2]),
    .ZN(_0453_)
  );
  OR2_X1 _5728_ (
    .A1(_0374_),
    .A2(_0453_),
    .ZN(_0454_)
  );
  AND2_X1 _5729_ (
    .A1(_0377_),
    .A2(_0454_),
    .ZN(_0455_)
  );
  AND2_X1 _5730_ (
    .A1(_0452_),
    .A2(_0455_),
    .ZN(_0456_)
  );
  XOR2_X1 _5731_ (
    .A(_0452_),
    .B(_0455_),
    .Z(_0457_)
  );
  AND2_X1 _5732_ (
    .A1(_0354_),
    .A2(_0457_),
    .ZN(_0458_)
  );
  XOR2_X1 _5733_ (
    .A(_0354_),
    .B(_0457_),
    .Z(_0459_)
  );
  AND2_X1 _5734_ (
    .A1(_0442_),
    .A2(_0459_),
    .ZN(_0460_)
  );
  XOR2_X1 _5735_ (
    .A(_0442_),
    .B(_0459_),
    .Z(_0461_)
  );
  AND2_X1 _5736_ (
    .A1(_0382_),
    .A2(_0461_),
    .ZN(_0462_)
  );
  XOR2_X1 _5737_ (
    .A(_0382_),
    .B(_0461_),
    .Z(_0463_)
  );
  AND2_X1 _5738_ (
    .A1(_0384_),
    .A2(_0463_),
    .ZN(_0464_)
  );
  XOR2_X1 _5739_ (
    .A(_0384_),
    .B(_0463_),
    .Z(_0465_)
  );
  AND2_X1 _5740_ (
    .A1(_0441_),
    .A2(_0465_),
    .ZN(_0466_)
  );
  XOR2_X1 _5741_ (
    .A(_0441_),
    .B(_0465_),
    .Z(_0467_)
  );
  AND2_X1 _5742_ (
    .A1(_0440_),
    .A2(_0467_),
    .ZN(_0468_)
  );
  XOR2_X1 _5743_ (
    .A(_0440_),
    .B(_0467_),
    .Z(_0469_)
  );
  AND2_X1 _5744_ (
    .A1(_0439_),
    .A2(_0469_),
    .ZN(_0470_)
  );
  XOR2_X1 _5745_ (
    .A(_0439_),
    .B(_0469_),
    .Z(_0471_)
  );
  AND2_X1 _5746_ (
    .A1(_0421_),
    .A2(_0471_),
    .ZN(_0472_)
  );
  XOR2_X1 _5747_ (
    .A(_0421_),
    .B(_0471_),
    .Z(_0473_)
  );
  AND2_X1 _5748_ (
    .A1(_0390_),
    .A2(_0473_),
    .ZN(_0474_)
  );
  XOR2_X1 _5749_ (
    .A(_0390_),
    .B(_0473_),
    .Z(_0475_)
  );
  AND2_X1 _5750_ (
    .A1(_0420_),
    .A2(_0475_),
    .ZN(_0476_)
  );
  XOR2_X1 _5751_ (
    .A(_0420_),
    .B(_0475_),
    .Z(_0477_)
  );
  AND2_X1 _5752_ (
    .A1(_0398_),
    .A2(_0477_),
    .ZN(_0478_)
  );
  XOR2_X1 _5753_ (
    .A(_0398_),
    .B(_0477_),
    .Z(_0479_)
  );
  INV_X1 _5754_ (
    .A(_0479_),
    .ZN(_0480_)
  );
  OR2_X1 _5755_ (
    .A1(_0400_),
    .A2(_0403_),
    .ZN(_0481_)
  );
  AND2_X1 _5756_ (
    .A1(_0479_),
    .A2(_0481_),
    .ZN(_0482_)
  );
  XOR2_X1 _5757_ (
    .A(_0480_),
    .B(_0481_),
    .Z(_0483_)
  );
  INV_X1 _5758_ (
    .A(_0483_),
    .ZN(_0484_)
  );
  AND2_X1 _5759_ (
    .A1(remainder[43]),
    .A2(_0484_),
    .ZN(_0485_)
  );
  OR2_X1 _5760_ (
    .A1(_3133_),
    .A2(_0483_),
    .ZN(_0486_)
  );
  XOR2_X1 _5761_ (
    .A(_3133_),
    .B(_0483_),
    .Z(_0487_)
  );
  XOR2_X1 _5762_ (
    .A(remainder[43]),
    .B(_0483_),
    .Z(_0488_)
  );
  AND2_X1 _5763_ (
    .A1(_0342_),
    .A2(_0407_),
    .ZN(_0489_)
  );
  OR2_X1 _5764_ (
    .A1(_0343_),
    .A2(_0406_),
    .ZN(_0490_)
  );
  AND2_X1 _5765_ (
    .A1(_0409_),
    .A2(_0490_),
    .ZN(_0491_)
  );
  OR2_X1 _5766_ (
    .A1(_0408_),
    .A2(_0489_),
    .ZN(_0492_)
  );
  AND2_X1 _5767_ (
    .A1(_0487_),
    .A2(_0491_),
    .ZN(_0493_)
  );
  OR2_X1 _5768_ (
    .A1(_0488_),
    .A2(_0492_),
    .ZN(_0494_)
  );
  OR2_X1 _5769_ (
    .A1(_0487_),
    .A2(_0491_),
    .ZN(_0495_)
  );
  AND2_X1 _5770_ (
    .A1(_4613_),
    .A2(_0495_),
    .ZN(_0496_)
  );
  AND2_X1 _5771_ (
    .A1(_0494_),
    .A2(_0496_),
    .ZN(_0497_)
  );
  OR2_X1 _5772_ (
    .A1(_0419_),
    .A2(_0497_),
    .ZN(_0498_)
  );
  OR2_X1 _5773_ (
    .A1(_0418_),
    .A2(_0498_),
    .ZN(_0499_)
  );
  AND2_X1 _5774_ (
    .A1(_3911_),
    .A2(_0499_),
    .ZN(_0056_)
  );
  OR2_X1 _5775_ (
    .A1(_4392_),
    .A2(_4447_),
    .ZN(_0500_)
  );
  OR2_X1 _5776_ (
    .A1(remainder[35]),
    .A2(_4393_),
    .ZN(_0501_)
  );
  AND2_X1 _5777_ (
    .A1(_3678_),
    .A2(_0500_),
    .ZN(_0502_)
  );
  AND2_X1 _5778_ (
    .A1(_0501_),
    .A2(_0502_),
    .ZN(_0503_)
  );
  AND2_X1 _5779_ (
    .A1(remainder[36]),
    .A2(_4610_),
    .ZN(_0504_)
  );
  AND2_X1 _5780_ (
    .A1(_0486_),
    .A2(_0494_),
    .ZN(_0505_)
  );
  OR2_X1 _5781_ (
    .A1(_0485_),
    .A2(_0493_),
    .ZN(_0506_)
  );
  OR2_X1 _5782_ (
    .A1(_0478_),
    .A2(_0482_),
    .ZN(_0507_)
  );
  OR2_X1 _5783_ (
    .A1(_0472_),
    .A2(_0474_),
    .ZN(_0508_)
  );
  OR2_X1 _5784_ (
    .A1(_0438_),
    .A2(_0470_),
    .ZN(_0509_)
  );
  OR2_X1 _5785_ (
    .A1(_0464_),
    .A2(_0466_),
    .ZN(_0510_)
  );
  AND2_X1 _5786_ (
    .A1(_0297_),
    .A2(_0377_),
    .ZN(_0511_)
  );
  OR2_X1 _5787_ (
    .A1(_0296_),
    .A2(_0376_),
    .ZN(_0512_)
  );
  OR2_X1 _5788_ (
    .A1(_0458_),
    .A2(_0460_),
    .ZN(_0513_)
  );
  OR2_X1 _5789_ (
    .A1(_0451_),
    .A2(_0456_),
    .ZN(_0514_)
  );
  OR2_X1 _5790_ (
    .A1(_0447_),
    .A2(_0449_),
    .ZN(_0515_)
  );
  AND2_X1 _5791_ (
    .A1(divisor[4]),
    .A2(remainder[7]),
    .ZN(_0516_)
  );
  AND2_X1 _5792_ (
    .A1(divisor[5]),
    .A2(remainder[6]),
    .ZN(_0517_)
  );
  AND2_X1 _5793_ (
    .A1(divisor[6]),
    .A2(remainder[6]),
    .ZN(_0518_)
  );
  AND2_X1 _5794_ (
    .A1(_0446_),
    .A2(_0517_),
    .ZN(_0519_)
  );
  XOR2_X1 _5795_ (
    .A(_0446_),
    .B(_0517_),
    .Z(_0520_)
  );
  AND2_X1 _5796_ (
    .A1(_0516_),
    .A2(_0520_),
    .ZN(_0521_)
  );
  XOR2_X1 _5797_ (
    .A(_0516_),
    .B(_0520_),
    .Z(_0522_)
  );
  AND2_X1 _5798_ (
    .A1(_0515_),
    .A2(_0522_),
    .ZN(_0523_)
  );
  XOR2_X1 _5799_ (
    .A(_0515_),
    .B(_0522_),
    .Z(_0524_)
  );
  AND2_X1 _5800_ (
    .A1(_0455_),
    .A2(_0524_),
    .ZN(_0525_)
  );
  XOR2_X1 _5801_ (
    .A(_0455_),
    .B(_0524_),
    .Z(_0526_)
  );
  AND2_X1 _5802_ (
    .A1(_0432_),
    .A2(_0526_),
    .ZN(_0527_)
  );
  XOR2_X1 _5803_ (
    .A(_0432_),
    .B(_0526_),
    .Z(_0528_)
  );
  AND2_X1 _5804_ (
    .A1(_0514_),
    .A2(_0528_),
    .ZN(_0529_)
  );
  XOR2_X1 _5805_ (
    .A(_0514_),
    .B(_0528_),
    .Z(_0530_)
  );
  AND2_X1 _5806_ (
    .A1(_0434_),
    .A2(_0530_),
    .ZN(_0531_)
  );
  XOR2_X1 _5807_ (
    .A(_0434_),
    .B(_0530_),
    .Z(_0532_)
  );
  AND2_X1 _5808_ (
    .A1(_0513_),
    .A2(_0532_),
    .ZN(_0533_)
  );
  XOR2_X1 _5809_ (
    .A(_0513_),
    .B(_0532_),
    .Z(_0534_)
  );
  AND2_X1 _5810_ (
    .A1(_0462_),
    .A2(_0534_),
    .ZN(_0535_)
  );
  XOR2_X1 _5811_ (
    .A(_0462_),
    .B(_0534_),
    .Z(_0536_)
  );
  AND2_X1 _5812_ (
    .A1(_0512_),
    .A2(_0536_),
    .ZN(_0537_)
  );
  XOR2_X1 _5813_ (
    .A(_0512_),
    .B(_0536_),
    .Z(_0538_)
  );
  AND2_X1 _5814_ (
    .A1(_0510_),
    .A2(_0538_),
    .ZN(_0539_)
  );
  XOR2_X1 _5815_ (
    .A(_0510_),
    .B(_0538_),
    .Z(_0540_)
  );
  AND2_X1 _5816_ (
    .A1(remainder[32]),
    .A2(divisor[3]),
    .ZN(_0541_)
  );
  OR2_X1 _5817_ (
    .A1(_3209_),
    .A2(_3264_),
    .ZN(_0542_)
  );
  AND2_X1 _5818_ (
    .A1(divisor[11]),
    .A2(remainder[0]),
    .ZN(_0543_)
  );
  AND2_X1 _5819_ (
    .A1(divisor[10]),
    .A2(remainder[1]),
    .ZN(_0544_)
  );
  AND2_X1 _5820_ (
    .A1(divisor[11]),
    .A2(remainder[1]),
    .ZN(_0545_)
  );
  AND2_X1 _5821_ (
    .A1(_0423_),
    .A2(_0545_),
    .ZN(_0546_)
  );
  XOR2_X1 _5822_ (
    .A(_0543_),
    .B(_0544_),
    .Z(_0547_)
  );
  INV_X1 _5823_ (
    .A(_0547_),
    .ZN(_0548_)
  );
  OR2_X1 _5824_ (
    .A1(_0428_),
    .A2(_0430_),
    .ZN(_0549_)
  );
  AND2_X1 _5825_ (
    .A1(divisor[8]),
    .A2(remainder[3]),
    .ZN(_0550_)
  );
  AND2_X1 _5826_ (
    .A1(divisor[9]),
    .A2(remainder[3]),
    .ZN(_0551_)
  );
  AND2_X1 _5827_ (
    .A1(_0427_),
    .A2(_0550_),
    .ZN(_0552_)
  );
  XOR2_X1 _5828_ (
    .A(_0427_),
    .B(_0550_),
    .Z(_0553_)
  );
  AND2_X1 _5829_ (
    .A1(_0152_),
    .A2(_0553_),
    .ZN(_0554_)
  );
  XOR2_X1 _5830_ (
    .A(_0152_),
    .B(_0553_),
    .Z(_0555_)
  );
  AND2_X1 _5831_ (
    .A1(_0549_),
    .A2(_0555_),
    .ZN(_0556_)
  );
  XOR2_X1 _5832_ (
    .A(_0549_),
    .B(_0555_),
    .Z(_0557_)
  );
  AND2_X1 _5833_ (
    .A1(_0547_),
    .A2(_0557_),
    .ZN(_0558_)
  );
  XOR2_X1 _5834_ (
    .A(_0548_),
    .B(_0557_),
    .Z(_0559_)
  );
  AND2_X1 _5835_ (
    .A1(_0541_),
    .A2(_0559_),
    .ZN(_0560_)
  );
  XOR2_X1 _5836_ (
    .A(_0542_),
    .B(_0559_),
    .Z(_0561_)
  );
  AND2_X1 _5837_ (
    .A1(_0436_),
    .A2(_0561_),
    .ZN(_0562_)
  );
  XOR2_X1 _5838_ (
    .A(_0436_),
    .B(_0561_),
    .Z(_0563_)
  );
  AND2_X1 _5839_ (
    .A1(_0540_),
    .A2(_0563_),
    .ZN(_0564_)
  );
  XOR2_X1 _5840_ (
    .A(_0540_),
    .B(_0563_),
    .Z(_0565_)
  );
  AND2_X1 _5841_ (
    .A1(_0509_),
    .A2(_0565_),
    .ZN(_0566_)
  );
  XOR2_X1 _5842_ (
    .A(_0509_),
    .B(_0565_),
    .Z(_0567_)
  );
  AND2_X1 _5843_ (
    .A1(_0468_),
    .A2(_0567_),
    .ZN(_0568_)
  );
  XOR2_X1 _5844_ (
    .A(_0468_),
    .B(_0567_),
    .Z(_0569_)
  );
  AND2_X1 _5845_ (
    .A1(_0508_),
    .A2(_0569_),
    .ZN(_0570_)
  );
  XOR2_X1 _5846_ (
    .A(_0508_),
    .B(_0569_),
    .Z(_0571_)
  );
  AND2_X1 _5847_ (
    .A1(_0476_),
    .A2(_0571_),
    .ZN(_0572_)
  );
  XOR2_X1 _5848_ (
    .A(_0476_),
    .B(_0571_),
    .Z(_0573_)
  );
  AND2_X1 _5849_ (
    .A1(_0507_),
    .A2(_0573_),
    .ZN(_0574_)
  );
  XOR2_X1 _5850_ (
    .A(_0507_),
    .B(_0573_),
    .Z(_0575_)
  );
  AND2_X1 _5851_ (
    .A1(remainder[44]),
    .A2(_0575_),
    .ZN(_0576_)
  );
  INV_X1 _5852_ (
    .A(_0576_),
    .ZN(_0577_)
  );
  XOR2_X1 _5853_ (
    .A(remainder[44]),
    .B(_0575_),
    .Z(_0578_)
  );
  XOR2_X1 _5854_ (
    .A(_3122_),
    .B(_0575_),
    .Z(_0579_)
  );
  AND2_X1 _5855_ (
    .A1(_0506_),
    .A2(_0578_),
    .ZN(_0580_)
  );
  OR2_X1 _5856_ (
    .A1(_0505_),
    .A2(_0579_),
    .ZN(_0581_)
  );
  OR2_X1 _5857_ (
    .A1(_0506_),
    .A2(_0578_),
    .ZN(_0582_)
  );
  AND2_X1 _5858_ (
    .A1(_4613_),
    .A2(_0582_),
    .ZN(_0583_)
  );
  AND2_X1 _5859_ (
    .A1(_0581_),
    .A2(_0583_),
    .ZN(_0584_)
  );
  OR2_X1 _5860_ (
    .A1(_0504_),
    .A2(_0584_),
    .ZN(_0585_)
  );
  OR2_X1 _5861_ (
    .A1(_0503_),
    .A2(_0585_),
    .ZN(_0586_)
  );
  AND2_X1 _5862_ (
    .A1(_3911_),
    .A2(_0586_),
    .ZN(_0057_)
  );
  OR2_X1 _5863_ (
    .A1(remainder[36]),
    .A2(_4393_),
    .ZN(_0587_)
  );
  OR2_X1 _5864_ (
    .A1(_4392_),
    .A2(_4452_),
    .ZN(_0588_)
  );
  AND2_X1 _5865_ (
    .A1(_3678_),
    .A2(_0588_),
    .ZN(_0589_)
  );
  AND2_X1 _5866_ (
    .A1(_0587_),
    .A2(_0589_),
    .ZN(_0590_)
  );
  AND2_X1 _5867_ (
    .A1(remainder[37]),
    .A2(_4610_),
    .ZN(_0591_)
  );
  AND2_X1 _5868_ (
    .A1(_0577_),
    .A2(_0581_),
    .ZN(_0592_)
  );
  OR2_X1 _5869_ (
    .A1(_0576_),
    .A2(_0580_),
    .ZN(_0593_)
  );
  OR2_X1 _5870_ (
    .A1(_0572_),
    .A2(_0574_),
    .ZN(_0594_)
  );
  OR2_X1 _5871_ (
    .A1(_0566_),
    .A2(_0568_),
    .ZN(_0595_)
  );
  OR2_X1 _5872_ (
    .A1(_0562_),
    .A2(_0564_),
    .ZN(_0596_)
  );
  OR2_X1 _5873_ (
    .A1(_0535_),
    .A2(_0537_),
    .ZN(_0597_)
  );
  OR2_X1 _5874_ (
    .A1(_0531_),
    .A2(_0533_),
    .ZN(_0598_)
  );
  OR2_X1 _5875_ (
    .A1(_0527_),
    .A2(_0529_),
    .ZN(_0599_)
  );
  OR2_X1 _5876_ (
    .A1(_0523_),
    .A2(_0525_),
    .ZN(_0600_)
  );
  OR2_X1 _5877_ (
    .A1(_0519_),
    .A2(_0521_),
    .ZN(_0601_)
  );
  AND2_X1 _5878_ (
    .A1(remainder[32]),
    .A2(divisor[4]),
    .ZN(_0602_)
  );
  INV_X1 _5879_ (
    .A(_0602_),
    .ZN(_0603_)
  );
  AND2_X1 _5880_ (
    .A1(divisor[5]),
    .A2(remainder[7]),
    .ZN(_0604_)
  );
  AND2_X1 _5881_ (
    .A1(divisor[6]),
    .A2(remainder[7]),
    .ZN(_0605_)
  );
  AND2_X1 _5882_ (
    .A1(_0517_),
    .A2(_0605_),
    .ZN(_0606_)
  );
  XOR2_X1 _5883_ (
    .A(_0518_),
    .B(_0604_),
    .Z(_0607_)
  );
  AND2_X1 _5884_ (
    .A1(_0602_),
    .A2(_0607_),
    .ZN(_0608_)
  );
  XOR2_X1 _5885_ (
    .A(_0602_),
    .B(_0607_),
    .Z(_0609_)
  );
  AND2_X1 _5886_ (
    .A1(_0601_),
    .A2(_0609_),
    .ZN(_0610_)
  );
  XOR2_X1 _5887_ (
    .A(_0601_),
    .B(_0609_),
    .Z(_0611_)
  );
  AND2_X1 _5888_ (
    .A1(_0455_),
    .A2(_0611_),
    .ZN(_0612_)
  );
  XOR2_X1 _5889_ (
    .A(_0455_),
    .B(_0611_),
    .Z(_0613_)
  );
  AND2_X1 _5890_ (
    .A1(_0556_),
    .A2(_0613_),
    .ZN(_0614_)
  );
  XOR2_X1 _5891_ (
    .A(_0556_),
    .B(_0613_),
    .Z(_0615_)
  );
  AND2_X1 _5892_ (
    .A1(_0600_),
    .A2(_0615_),
    .ZN(_0616_)
  );
  XOR2_X1 _5893_ (
    .A(_0600_),
    .B(_0615_),
    .Z(_0617_)
  );
  AND2_X1 _5894_ (
    .A1(_0558_),
    .A2(_0617_),
    .ZN(_0618_)
  );
  XOR2_X1 _5895_ (
    .A(_0558_),
    .B(_0617_),
    .Z(_0619_)
  );
  AND2_X1 _5896_ (
    .A1(_0599_),
    .A2(_0619_),
    .ZN(_0620_)
  );
  XOR2_X1 _5897_ (
    .A(_0599_),
    .B(_0619_),
    .Z(_0621_)
  );
  AND2_X1 _5898_ (
    .A1(_0598_),
    .A2(_0621_),
    .ZN(_0622_)
  );
  XOR2_X1 _5899_ (
    .A(_0598_),
    .B(_0621_),
    .Z(_0623_)
  );
  AND2_X1 _5900_ (
    .A1(_0512_),
    .A2(_0623_),
    .ZN(_0624_)
  );
  XOR2_X1 _5901_ (
    .A(_0512_),
    .B(_0623_),
    .Z(_0625_)
  );
  AND2_X1 _5902_ (
    .A1(_0597_),
    .A2(_0625_),
    .ZN(_0626_)
  );
  XOR2_X1 _5903_ (
    .A(_0597_),
    .B(_0625_),
    .Z(_0627_)
  );
  AND2_X1 _5904_ (
    .A1(divisor[10]),
    .A2(remainder[2]),
    .ZN(_0628_)
  );
  AND2_X1 _5905_ (
    .A1(divisor[12]),
    .A2(remainder[0]),
    .ZN(_0629_)
  );
  AND2_X1 _5906_ (
    .A1(divisor[12]),
    .A2(remainder[1]),
    .ZN(_0630_)
  );
  AND2_X1 _5907_ (
    .A1(_0543_),
    .A2(_0630_),
    .ZN(_0631_)
  );
  XOR2_X1 _5908_ (
    .A(_0545_),
    .B(_0629_),
    .Z(_0632_)
  );
  AND2_X1 _5909_ (
    .A1(_0628_),
    .A2(_0632_),
    .ZN(_0633_)
  );
  XOR2_X1 _5910_ (
    .A(_0628_),
    .B(_0632_),
    .Z(_0634_)
  );
  OR2_X1 _5911_ (
    .A1(_0552_),
    .A2(_0554_),
    .ZN(_0635_)
  );
  AND2_X1 _5912_ (
    .A1(divisor[7]),
    .A2(remainder[5]),
    .ZN(_0636_)
  );
  AND2_X1 _5913_ (
    .A1(divisor[8]),
    .A2(remainder[4]),
    .ZN(_0637_)
  );
  AND2_X1 _5914_ (
    .A1(divisor[9]),
    .A2(remainder[4]),
    .ZN(_0638_)
  );
  AND2_X1 _5915_ (
    .A1(_0551_),
    .A2(_0637_),
    .ZN(_0639_)
  );
  XOR2_X1 _5916_ (
    .A(_0551_),
    .B(_0637_),
    .Z(_0640_)
  );
  AND2_X1 _5917_ (
    .A1(_0636_),
    .A2(_0640_),
    .ZN(_0641_)
  );
  XOR2_X1 _5918_ (
    .A(_0636_),
    .B(_0640_),
    .Z(_0642_)
  );
  AND2_X1 _5919_ (
    .A1(_0546_),
    .A2(_0642_),
    .ZN(_0643_)
  );
  XOR2_X1 _5920_ (
    .A(_0546_),
    .B(_0642_),
    .Z(_0644_)
  );
  AND2_X1 _5921_ (
    .A1(_0635_),
    .A2(_0644_),
    .ZN(_0645_)
  );
  XOR2_X1 _5922_ (
    .A(_0635_),
    .B(_0644_),
    .Z(_0646_)
  );
  AND2_X1 _5923_ (
    .A1(_0634_),
    .A2(_0646_),
    .ZN(_0647_)
  );
  XOR2_X1 _5924_ (
    .A(_0634_),
    .B(_0646_),
    .Z(_0648_)
  );
  XOR2_X1 _5925_ (
    .A(_0560_),
    .B(_0648_),
    .Z(_0649_)
  );
  AND2_X1 _5926_ (
    .A1(_0627_),
    .A2(_0649_),
    .ZN(_0650_)
  );
  INV_X1 _5927_ (
    .A(_0650_),
    .ZN(_0651_)
  );
  XOR2_X1 _5928_ (
    .A(_0627_),
    .B(_0649_),
    .Z(_0652_)
  );
  AND2_X1 _5929_ (
    .A1(_0596_),
    .A2(_0652_),
    .ZN(_0653_)
  );
  XOR2_X1 _5930_ (
    .A(_0596_),
    .B(_0652_),
    .Z(_0654_)
  );
  AND2_X1 _5931_ (
    .A1(_0539_),
    .A2(_0654_),
    .ZN(_0655_)
  );
  XOR2_X1 _5932_ (
    .A(_0539_),
    .B(_0654_),
    .Z(_0656_)
  );
  AND2_X1 _5933_ (
    .A1(_0595_),
    .A2(_0656_),
    .ZN(_0657_)
  );
  INV_X1 _5934_ (
    .A(_0657_),
    .ZN(_0658_)
  );
  XOR2_X1 _5935_ (
    .A(_0595_),
    .B(_0656_),
    .Z(_0659_)
  );
  AND2_X1 _5936_ (
    .A1(_0570_),
    .A2(_0659_),
    .ZN(_0660_)
  );
  XOR2_X1 _5937_ (
    .A(_0570_),
    .B(_0659_),
    .Z(_0661_)
  );
  AND2_X1 _5938_ (
    .A1(_0594_),
    .A2(_0661_),
    .ZN(_0662_)
  );
  XOR2_X1 _5939_ (
    .A(_0594_),
    .B(_0661_),
    .Z(_0663_)
  );
  AND2_X1 _5940_ (
    .A1(remainder[45]),
    .A2(_0663_),
    .ZN(_0664_)
  );
  INV_X1 _5941_ (
    .A(_0664_),
    .ZN(_0665_)
  );
  XOR2_X1 _5942_ (
    .A(remainder[45]),
    .B(_0663_),
    .Z(_0666_)
  );
  XOR2_X1 _5943_ (
    .A(_3111_),
    .B(_0663_),
    .Z(_0667_)
  );
  AND2_X1 _5944_ (
    .A1(_0593_),
    .A2(_0666_),
    .ZN(_0668_)
  );
  OR2_X1 _5945_ (
    .A1(_0592_),
    .A2(_0667_),
    .ZN(_0669_)
  );
  OR2_X1 _5946_ (
    .A1(_0593_),
    .A2(_0666_),
    .ZN(_0670_)
  );
  AND2_X1 _5947_ (
    .A1(_4613_),
    .A2(_0670_),
    .ZN(_0671_)
  );
  AND2_X1 _5948_ (
    .A1(_0669_),
    .A2(_0671_),
    .ZN(_0672_)
  );
  OR2_X1 _5949_ (
    .A1(_0591_),
    .A2(_0672_),
    .ZN(_0673_)
  );
  OR2_X1 _5950_ (
    .A1(_0590_),
    .A2(_0673_),
    .ZN(_0674_)
  );
  AND2_X1 _5951_ (
    .A1(_3911_),
    .A2(_0674_),
    .ZN(_0058_)
  );
  OR2_X1 _5952_ (
    .A1(remainder[37]),
    .A2(_4393_),
    .ZN(_0675_)
  );
  OR2_X1 _5953_ (
    .A1(_4392_),
    .A2(_4457_),
    .ZN(_0676_)
  );
  AND2_X1 _5954_ (
    .A1(_3678_),
    .A2(_0676_),
    .ZN(_0677_)
  );
  AND2_X1 _5955_ (
    .A1(_0675_),
    .A2(_0677_),
    .ZN(_0678_)
  );
  AND2_X1 _5956_ (
    .A1(remainder[38]),
    .A2(_4610_),
    .ZN(_0679_)
  );
  AND2_X1 _5957_ (
    .A1(_0665_),
    .A2(_0669_),
    .ZN(_0680_)
  );
  OR2_X1 _5958_ (
    .A1(_0664_),
    .A2(_0668_),
    .ZN(_0681_)
  );
  OR2_X1 _5959_ (
    .A1(_0660_),
    .A2(_0662_),
    .ZN(_0682_)
  );
  OR2_X1 _5960_ (
    .A1(_0653_),
    .A2(_0655_),
    .ZN(_0683_)
  );
  OR2_X1 _5961_ (
    .A1(_0542_),
    .A2(_0648_),
    .ZN(_0684_)
  );
  OR2_X1 _5962_ (
    .A1(_0559_),
    .A2(_0684_),
    .ZN(_0685_)
  );
  AND2_X1 _5963_ (
    .A1(_0651_),
    .A2(_0685_),
    .ZN(_0686_)
  );
  OR2_X1 _5964_ (
    .A1(_0622_),
    .A2(_0624_),
    .ZN(_0687_)
  );
  OR2_X1 _5965_ (
    .A1(_0618_),
    .A2(_0620_),
    .ZN(_0688_)
  );
  OR2_X1 _5966_ (
    .A1(_0614_),
    .A2(_0616_),
    .ZN(_0689_)
  );
  OR2_X1 _5967_ (
    .A1(_0610_),
    .A2(_0612_),
    .ZN(_0690_)
  );
  OR2_X1 _5968_ (
    .A1(_0643_),
    .A2(_0645_),
    .ZN(_0691_)
  );
  OR2_X1 _5969_ (
    .A1(_0606_),
    .A2(_0608_),
    .ZN(_0692_)
  );
  AND2_X1 _5970_ (
    .A1(remainder[32]),
    .A2(divisor[6]),
    .ZN(_0693_)
  );
  AND2_X1 _5971_ (
    .A1(remainder[32]),
    .A2(divisor[5]),
    .ZN(_0694_)
  );
  AND2_X1 _5972_ (
    .A1(_0605_),
    .A2(_0694_),
    .ZN(_0695_)
  );
  XOR2_X1 _5973_ (
    .A(_0605_),
    .B(_0694_),
    .Z(_0696_)
  );
  AND2_X1 _5974_ (
    .A1(_0602_),
    .A2(_0696_),
    .ZN(_0697_)
  );
  XOR2_X1 _5975_ (
    .A(_0602_),
    .B(_0696_),
    .Z(_0698_)
  );
  AND2_X1 _5976_ (
    .A1(_0692_),
    .A2(_0698_),
    .ZN(_0699_)
  );
  XOR2_X1 _5977_ (
    .A(_0692_),
    .B(_0698_),
    .Z(_0700_)
  );
  AND2_X1 _5978_ (
    .A1(_0455_),
    .A2(_0700_),
    .ZN(_0701_)
  );
  XOR2_X1 _5979_ (
    .A(_0455_),
    .B(_0700_),
    .Z(_0702_)
  );
  AND2_X1 _5980_ (
    .A1(_0691_),
    .A2(_0702_),
    .ZN(_0703_)
  );
  XOR2_X1 _5981_ (
    .A(_0691_),
    .B(_0702_),
    .Z(_0704_)
  );
  AND2_X1 _5982_ (
    .A1(_0690_),
    .A2(_0704_),
    .ZN(_0705_)
  );
  XOR2_X1 _5983_ (
    .A(_0690_),
    .B(_0704_),
    .Z(_0706_)
  );
  AND2_X1 _5984_ (
    .A1(_0647_),
    .A2(_0706_),
    .ZN(_0707_)
  );
  XOR2_X1 _5985_ (
    .A(_0647_),
    .B(_0706_),
    .Z(_0708_)
  );
  AND2_X1 _5986_ (
    .A1(_0689_),
    .A2(_0708_),
    .ZN(_0709_)
  );
  XOR2_X1 _5987_ (
    .A(_0689_),
    .B(_0708_),
    .Z(_0710_)
  );
  AND2_X1 _5988_ (
    .A1(_0688_),
    .A2(_0710_),
    .ZN(_0711_)
  );
  XOR2_X1 _5989_ (
    .A(_0688_),
    .B(_0710_),
    .Z(_0712_)
  );
  AND2_X1 _5990_ (
    .A1(_0512_),
    .A2(_0712_),
    .ZN(_0713_)
  );
  XOR2_X1 _5991_ (
    .A(_0512_),
    .B(_0712_),
    .Z(_0714_)
  );
  AND2_X1 _5992_ (
    .A1(_0687_),
    .A2(_0714_),
    .ZN(_0715_)
  );
  XOR2_X1 _5993_ (
    .A(_0687_),
    .B(_0714_),
    .Z(_0716_)
  );
  AND2_X1 _5994_ (
    .A1(divisor[13]),
    .A2(remainder[0]),
    .ZN(_0717_)
  );
  AND2_X1 _5995_ (
    .A1(divisor[10]),
    .A2(remainder[3]),
    .ZN(_0718_)
  );
  AND2_X1 _5996_ (
    .A1(divisor[11]),
    .A2(remainder[2]),
    .ZN(_0719_)
  );
  AND2_X1 _5997_ (
    .A1(divisor[12]),
    .A2(remainder[2]),
    .ZN(_0720_)
  );
  AND2_X1 _5998_ (
    .A1(_0545_),
    .A2(_0720_),
    .ZN(_0721_)
  );
  XOR2_X1 _5999_ (
    .A(_0630_),
    .B(_0719_),
    .Z(_0722_)
  );
  AND2_X1 _6000_ (
    .A1(_0718_),
    .A2(_0722_),
    .ZN(_0723_)
  );
  XOR2_X1 _6001_ (
    .A(_0718_),
    .B(_0722_),
    .Z(_0724_)
  );
  AND2_X1 _6002_ (
    .A1(_0717_),
    .A2(_0724_),
    .ZN(_0725_)
  );
  XOR2_X1 _6003_ (
    .A(_0717_),
    .B(_0724_),
    .Z(_0726_)
  );
  OR2_X1 _6004_ (
    .A1(_0639_),
    .A2(_0641_),
    .ZN(_0727_)
  );
  OR2_X1 _6005_ (
    .A1(_0631_),
    .A2(_0633_),
    .ZN(_0728_)
  );
  AND2_X1 _6006_ (
    .A1(divisor[7]),
    .A2(remainder[6]),
    .ZN(_0729_)
  );
  AND2_X1 _6007_ (
    .A1(divisor[8]),
    .A2(remainder[5]),
    .ZN(_0730_)
  );
  AND2_X1 _6008_ (
    .A1(divisor[9]),
    .A2(remainder[5]),
    .ZN(_0731_)
  );
  AND2_X1 _6009_ (
    .A1(_0638_),
    .A2(_0730_),
    .ZN(_0732_)
  );
  XOR2_X1 _6010_ (
    .A(_0638_),
    .B(_0730_),
    .Z(_0733_)
  );
  AND2_X1 _6011_ (
    .A1(_0729_),
    .A2(_0733_),
    .ZN(_0734_)
  );
  XOR2_X1 _6012_ (
    .A(_0729_),
    .B(_0733_),
    .Z(_0735_)
  );
  AND2_X1 _6013_ (
    .A1(_0728_),
    .A2(_0735_),
    .ZN(_0736_)
  );
  XOR2_X1 _6014_ (
    .A(_0728_),
    .B(_0735_),
    .Z(_0737_)
  );
  AND2_X1 _6015_ (
    .A1(_0727_),
    .A2(_0737_),
    .ZN(_0738_)
  );
  XOR2_X1 _6016_ (
    .A(_0727_),
    .B(_0737_),
    .Z(_0739_)
  );
  AND2_X1 _6017_ (
    .A1(_0726_),
    .A2(_0739_),
    .ZN(_0740_)
  );
  XOR2_X1 _6018_ (
    .A(_0726_),
    .B(_0739_),
    .Z(_0741_)
  );
  INV_X1 _6019_ (
    .A(_0741_),
    .ZN(_0742_)
  );
  XOR2_X1 _6020_ (
    .A(_0684_),
    .B(_0741_),
    .Z(_0743_)
  );
  INV_X1 _6021_ (
    .A(_0743_),
    .ZN(_0744_)
  );
  AND2_X1 _6022_ (
    .A1(_0716_),
    .A2(_0744_),
    .ZN(_0745_)
  );
  XOR2_X1 _6023_ (
    .A(_0716_),
    .B(_0743_),
    .Z(_0746_)
  );
  OR2_X1 _6024_ (
    .A1(_0686_),
    .A2(_0746_),
    .ZN(_0747_)
  );
  INV_X1 _6025_ (
    .A(_0747_),
    .ZN(_0748_)
  );
  XOR2_X1 _6026_ (
    .A(_0686_),
    .B(_0746_),
    .Z(_0749_)
  );
  AND2_X1 _6027_ (
    .A1(_0626_),
    .A2(_0749_),
    .ZN(_0750_)
  );
  XOR2_X1 _6028_ (
    .A(_0626_),
    .B(_0749_),
    .Z(_0751_)
  );
  AND2_X1 _6029_ (
    .A1(_0683_),
    .A2(_0751_),
    .ZN(_0752_)
  );
  INV_X1 _6030_ (
    .A(_0752_),
    .ZN(_0753_)
  );
  XOR2_X1 _6031_ (
    .A(_0683_),
    .B(_0751_),
    .Z(_0754_)
  );
  AND2_X1 _6032_ (
    .A1(_0657_),
    .A2(_0754_),
    .ZN(_0755_)
  );
  XOR2_X1 _6033_ (
    .A(_0657_),
    .B(_0754_),
    .Z(_0756_)
  );
  XOR2_X1 _6034_ (
    .A(_0658_),
    .B(_0754_),
    .Z(_0757_)
  );
  AND2_X1 _6035_ (
    .A1(_0682_),
    .A2(_0756_),
    .ZN(_0758_)
  );
  XOR2_X1 _6036_ (
    .A(_0682_),
    .B(_0757_),
    .Z(_0759_)
  );
  XOR2_X1 _6037_ (
    .A(_0682_),
    .B(_0756_),
    .Z(_0760_)
  );
  AND2_X1 _6038_ (
    .A1(remainder[46]),
    .A2(_0760_),
    .ZN(_0761_)
  );
  OR2_X1 _6039_ (
    .A1(_3100_),
    .A2(_0759_),
    .ZN(_0762_)
  );
  OR2_X1 _6040_ (
    .A1(remainder[46]),
    .A2(_0760_),
    .ZN(_0763_)
  );
  INV_X1 _6041_ (
    .A(_0763_),
    .ZN(_0764_)
  );
  AND2_X1 _6042_ (
    .A1(_0762_),
    .A2(_0763_),
    .ZN(_0765_)
  );
  XOR2_X1 _6043_ (
    .A(_0681_),
    .B(_0765_),
    .Z(_0766_)
  );
  AND2_X1 _6044_ (
    .A1(_4613_),
    .A2(_0766_),
    .ZN(_0767_)
  );
  OR2_X1 _6045_ (
    .A1(_0679_),
    .A2(_0767_),
    .ZN(_0768_)
  );
  OR2_X1 _6046_ (
    .A1(_0678_),
    .A2(_0768_),
    .ZN(_0769_)
  );
  AND2_X1 _6047_ (
    .A1(_3911_),
    .A2(_0769_),
    .ZN(_0059_)
  );
  OR2_X1 _6048_ (
    .A1(remainder[38]),
    .A2(_4393_),
    .ZN(_0770_)
  );
  OR2_X1 _6049_ (
    .A1(_4392_),
    .A2(_4462_),
    .ZN(_0771_)
  );
  AND2_X1 _6050_ (
    .A1(_3678_),
    .A2(_0771_),
    .ZN(_0772_)
  );
  AND2_X1 _6051_ (
    .A1(_0770_),
    .A2(_0772_),
    .ZN(_0773_)
  );
  AND2_X1 _6052_ (
    .A1(remainder[39]),
    .A2(_4610_),
    .ZN(_0774_)
  );
  OR2_X1 _6053_ (
    .A1(_0748_),
    .A2(_0750_),
    .ZN(_0775_)
  );
  AND2_X1 _6054_ (
    .A1(_0541_),
    .A2(_0742_),
    .ZN(_0776_)
  );
  AND2_X1 _6055_ (
    .A1(_0648_),
    .A2(_0776_),
    .ZN(_0777_)
  );
  OR2_X1 _6056_ (
    .A1(_0745_),
    .A2(_0777_),
    .ZN(_0778_)
  );
  OR2_X1 _6057_ (
    .A1(_0711_),
    .A2(_0713_),
    .ZN(_0779_)
  );
  OR2_X1 _6058_ (
    .A1(_0707_),
    .A2(_0709_),
    .ZN(_0780_)
  );
  OR2_X1 _6059_ (
    .A1(_0703_),
    .A2(_0705_),
    .ZN(_0781_)
  );
  OR2_X1 _6060_ (
    .A1(_0699_),
    .A2(_0701_),
    .ZN(_0782_)
  );
  OR2_X1 _6061_ (
    .A1(_0736_),
    .A2(_0738_),
    .ZN(_0783_)
  );
  OR2_X1 _6062_ (
    .A1(_0695_),
    .A2(_0697_),
    .ZN(_0784_)
  );
  OR2_X1 _6063_ (
    .A1(_0693_),
    .A2(_0694_),
    .ZN(_0785_)
  );
  MUX2_X1 _6064_ (
    .A(_0694_),
    .B(_3274_),
    .S(_0693_),
    .Z(_0786_)
  );
  MUX2_X1 _6065_ (
    .A(_0603_),
    .B(divisor[4]),
    .S(_0786_),
    .Z(_0787_)
  );
  INV_X1 _6066_ (
    .A(_0787_),
    .ZN(_0788_)
  );
  AND2_X1 _6067_ (
    .A1(_0784_),
    .A2(_0788_),
    .ZN(_0789_)
  );
  INV_X1 _6068_ (
    .A(_0789_),
    .ZN(_0790_)
  );
  XOR2_X1 _6069_ (
    .A(_0784_),
    .B(_0788_),
    .Z(_0791_)
  );
  AND2_X1 _6070_ (
    .A1(_0455_),
    .A2(_0791_),
    .ZN(_0792_)
  );
  XOR2_X1 _6071_ (
    .A(_0455_),
    .B(_0791_),
    .Z(_0793_)
  );
  AND2_X1 _6072_ (
    .A1(_0783_),
    .A2(_0793_),
    .ZN(_0794_)
  );
  XOR2_X1 _6073_ (
    .A(_0783_),
    .B(_0793_),
    .Z(_0795_)
  );
  AND2_X1 _6074_ (
    .A1(_0782_),
    .A2(_0795_),
    .ZN(_0796_)
  );
  XOR2_X1 _6075_ (
    .A(_0782_),
    .B(_0795_),
    .Z(_0797_)
  );
  AND2_X1 _6076_ (
    .A1(_0740_),
    .A2(_0797_),
    .ZN(_0798_)
  );
  XOR2_X1 _6077_ (
    .A(_0740_),
    .B(_0797_),
    .Z(_0799_)
  );
  AND2_X1 _6078_ (
    .A1(_0781_),
    .A2(_0799_),
    .ZN(_0800_)
  );
  XOR2_X1 _6079_ (
    .A(_0781_),
    .B(_0799_),
    .Z(_0801_)
  );
  AND2_X1 _6080_ (
    .A1(_0780_),
    .A2(_0801_),
    .ZN(_0802_)
  );
  XOR2_X1 _6081_ (
    .A(_0780_),
    .B(_0801_),
    .Z(_0803_)
  );
  AND2_X1 _6082_ (
    .A1(_0512_),
    .A2(_0803_),
    .ZN(_0804_)
  );
  XOR2_X1 _6083_ (
    .A(_0512_),
    .B(_0803_),
    .Z(_0805_)
  );
  AND2_X1 _6084_ (
    .A1(_0779_),
    .A2(_0805_),
    .ZN(_0806_)
  );
  XOR2_X1 _6085_ (
    .A(_0779_),
    .B(_0805_),
    .Z(_0807_)
  );
  AND2_X1 _6086_ (
    .A1(divisor[14]),
    .A2(remainder[0]),
    .ZN(_0808_)
  );
  AND2_X1 _6087_ (
    .A1(divisor[13]),
    .A2(remainder[1]),
    .ZN(_0809_)
  );
  AND2_X1 _6088_ (
    .A1(divisor[14]),
    .A2(remainder[1]),
    .ZN(_0810_)
  );
  AND2_X1 _6089_ (
    .A1(_0717_),
    .A2(_0810_),
    .ZN(_0811_)
  );
  XOR2_X1 _6090_ (
    .A(_0808_),
    .B(_0809_),
    .Z(_0812_)
  );
  AND2_X1 _6091_ (
    .A1(divisor[10]),
    .A2(remainder[4]),
    .ZN(_0813_)
  );
  AND2_X1 _6092_ (
    .A1(divisor[11]),
    .A2(remainder[3]),
    .ZN(_0814_)
  );
  AND2_X1 _6093_ (
    .A1(divisor[12]),
    .A2(remainder[3]),
    .ZN(_0815_)
  );
  AND2_X1 _6094_ (
    .A1(_0720_),
    .A2(_0814_),
    .ZN(_0816_)
  );
  XOR2_X1 _6095_ (
    .A(_0720_),
    .B(_0814_),
    .Z(_0817_)
  );
  AND2_X1 _6096_ (
    .A1(_0813_),
    .A2(_0817_),
    .ZN(_0818_)
  );
  XOR2_X1 _6097_ (
    .A(_0813_),
    .B(_0817_),
    .Z(_0819_)
  );
  AND2_X1 _6098_ (
    .A1(_0812_),
    .A2(_0819_),
    .ZN(_0820_)
  );
  XOR2_X1 _6099_ (
    .A(_0812_),
    .B(_0819_),
    .Z(_0821_)
  );
  AND2_X1 _6100_ (
    .A1(_0725_),
    .A2(_0821_),
    .ZN(_0822_)
  );
  XOR2_X1 _6101_ (
    .A(_0725_),
    .B(_0821_),
    .Z(_0823_)
  );
  OR2_X1 _6102_ (
    .A1(_0732_),
    .A2(_0734_),
    .ZN(_0824_)
  );
  OR2_X1 _6103_ (
    .A1(_0721_),
    .A2(_0723_),
    .ZN(_0825_)
  );
  AND2_X1 _6104_ (
    .A1(divisor[7]),
    .A2(remainder[7]),
    .ZN(_0826_)
  );
  AND2_X1 _6105_ (
    .A1(divisor[8]),
    .A2(remainder[6]),
    .ZN(_0827_)
  );
  AND2_X1 _6106_ (
    .A1(divisor[9]),
    .A2(remainder[6]),
    .ZN(_0828_)
  );
  AND2_X1 _6107_ (
    .A1(_0731_),
    .A2(_0827_),
    .ZN(_0829_)
  );
  XOR2_X1 _6108_ (
    .A(_0731_),
    .B(_0827_),
    .Z(_0830_)
  );
  AND2_X1 _6109_ (
    .A1(_0826_),
    .A2(_0830_),
    .ZN(_0831_)
  );
  XOR2_X1 _6110_ (
    .A(_0826_),
    .B(_0830_),
    .Z(_0832_)
  );
  AND2_X1 _6111_ (
    .A1(_0825_),
    .A2(_0832_),
    .ZN(_0833_)
  );
  XOR2_X1 _6112_ (
    .A(_0825_),
    .B(_0832_),
    .Z(_0834_)
  );
  AND2_X1 _6113_ (
    .A1(_0824_),
    .A2(_0834_),
    .ZN(_0835_)
  );
  XOR2_X1 _6114_ (
    .A(_0824_),
    .B(_0834_),
    .Z(_0836_)
  );
  AND2_X1 _6115_ (
    .A1(_0823_),
    .A2(_0836_),
    .ZN(_0837_)
  );
  XOR2_X1 _6116_ (
    .A(_0823_),
    .B(_0836_),
    .Z(_0838_)
  );
  INV_X1 _6117_ (
    .A(_0838_),
    .ZN(_0839_)
  );
  XOR2_X1 _6118_ (
    .A(_0776_),
    .B(_0839_),
    .Z(_0840_)
  );
  XOR2_X1 _6119_ (
    .A(_0776_),
    .B(_0838_),
    .Z(_0841_)
  );
  AND2_X1 _6120_ (
    .A1(_0807_),
    .A2(_0841_),
    .ZN(_0842_)
  );
  XOR2_X1 _6121_ (
    .A(_0807_),
    .B(_0840_),
    .Z(_0843_)
  );
  INV_X1 _6122_ (
    .A(_0843_),
    .ZN(_0844_)
  );
  AND2_X1 _6123_ (
    .A1(_0778_),
    .A2(_0844_),
    .ZN(_0845_)
  );
  XOR2_X1 _6124_ (
    .A(_0778_),
    .B(_0844_),
    .Z(_0846_)
  );
  AND2_X1 _6125_ (
    .A1(_0715_),
    .A2(_0846_),
    .ZN(_0847_)
  );
  XOR2_X1 _6126_ (
    .A(_0715_),
    .B(_0846_),
    .Z(_0848_)
  );
  AND2_X1 _6127_ (
    .A1(_0775_),
    .A2(_0848_),
    .ZN(_0849_)
  );
  XOR2_X1 _6128_ (
    .A(_0775_),
    .B(_0848_),
    .Z(_0850_)
  );
  AND2_X1 _6129_ (
    .A1(_0752_),
    .A2(_0850_),
    .ZN(_0851_)
  );
  XOR2_X1 _6130_ (
    .A(_0752_),
    .B(_0850_),
    .Z(_0852_)
  );
  XOR2_X1 _6131_ (
    .A(_0753_),
    .B(_0850_),
    .Z(_0853_)
  );
  OR2_X1 _6132_ (
    .A1(_0755_),
    .A2(_0758_),
    .ZN(_0854_)
  );
  AND2_X1 _6133_ (
    .A1(_0852_),
    .A2(_0854_),
    .ZN(_0855_)
  );
  XOR2_X1 _6134_ (
    .A(_0853_),
    .B(_0854_),
    .Z(_0856_)
  );
  INV_X1 _6135_ (
    .A(_0856_),
    .ZN(_0857_)
  );
  AND2_X1 _6136_ (
    .A1(remainder[47]),
    .A2(_0857_),
    .ZN(_0858_)
  );
  OR2_X1 _6137_ (
    .A1(_3089_),
    .A2(_0856_),
    .ZN(_0859_)
  );
  XOR2_X1 _6138_ (
    .A(_3089_),
    .B(_0856_),
    .Z(_0860_)
  );
  XOR2_X1 _6139_ (
    .A(remainder[47]),
    .B(_0856_),
    .Z(_0861_)
  );
  AND2_X1 _6140_ (
    .A1(_0680_),
    .A2(_0762_),
    .ZN(_0862_)
  );
  OR2_X1 _6141_ (
    .A1(_0681_),
    .A2(_0761_),
    .ZN(_0863_)
  );
  AND2_X1 _6142_ (
    .A1(_0763_),
    .A2(_0863_),
    .ZN(_0864_)
  );
  OR2_X1 _6143_ (
    .A1(_0764_),
    .A2(_0862_),
    .ZN(_0865_)
  );
  AND2_X1 _6144_ (
    .A1(_0860_),
    .A2(_0864_),
    .ZN(_0866_)
  );
  OR2_X1 _6145_ (
    .A1(_0861_),
    .A2(_0865_),
    .ZN(_0867_)
  );
  OR2_X1 _6146_ (
    .A1(_0860_),
    .A2(_0864_),
    .ZN(_0868_)
  );
  AND2_X1 _6147_ (
    .A1(_4613_),
    .A2(_0868_),
    .ZN(_0869_)
  );
  AND2_X1 _6148_ (
    .A1(_0867_),
    .A2(_0869_),
    .ZN(_0870_)
  );
  OR2_X1 _6149_ (
    .A1(_0774_),
    .A2(_0870_),
    .ZN(_0871_)
  );
  OR2_X1 _6150_ (
    .A1(_0773_),
    .A2(_0871_),
    .ZN(_0872_)
  );
  AND2_X1 _6151_ (
    .A1(_3911_),
    .A2(_0872_),
    .ZN(_0060_)
  );
  OR2_X1 _6152_ (
    .A1(remainder[39]),
    .A2(_4393_),
    .ZN(_0873_)
  );
  OR2_X1 _6153_ (
    .A1(_4392_),
    .A2(_4468_),
    .ZN(_0874_)
  );
  AND2_X1 _6154_ (
    .A1(_3678_),
    .A2(_0874_),
    .ZN(_0875_)
  );
  AND2_X1 _6155_ (
    .A1(_0873_),
    .A2(_0875_),
    .ZN(_0876_)
  );
  AND2_X1 _6156_ (
    .A1(remainder[40]),
    .A2(_4610_),
    .ZN(_0877_)
  );
  AND2_X1 _6157_ (
    .A1(_0859_),
    .A2(_0867_),
    .ZN(_0878_)
  );
  OR2_X1 _6158_ (
    .A1(_0858_),
    .A2(_0866_),
    .ZN(_0879_)
  );
  OR2_X1 _6159_ (
    .A1(_0851_),
    .A2(_0855_),
    .ZN(_0880_)
  );
  OR2_X1 _6160_ (
    .A1(_0845_),
    .A2(_0847_),
    .ZN(_0881_)
  );
  AND2_X1 _6161_ (
    .A1(_0541_),
    .A2(_0839_),
    .ZN(_0882_)
  );
  AND2_X1 _6162_ (
    .A1(_0741_),
    .A2(_0882_),
    .ZN(_0883_)
  );
  OR2_X1 _6163_ (
    .A1(_0842_),
    .A2(_0883_),
    .ZN(_0884_)
  );
  OR2_X1 _6164_ (
    .A1(_0802_),
    .A2(_0804_),
    .ZN(_0885_)
  );
  OR2_X1 _6165_ (
    .A1(_0798_),
    .A2(_0800_),
    .ZN(_0886_)
  );
  OR2_X1 _6166_ (
    .A1(_0794_),
    .A2(_0796_),
    .ZN(_0887_)
  );
  OR2_X1 _6167_ (
    .A1(_0822_),
    .A2(_0837_),
    .ZN(_0888_)
  );
  OR2_X1 _6168_ (
    .A1(_0789_),
    .A2(_0792_),
    .ZN(_0889_)
  );
  OR2_X1 _6169_ (
    .A1(_0833_),
    .A2(_0835_),
    .ZN(_0890_)
  );
  OR2_X1 _6170_ (
    .A1(_0602_),
    .A2(_0785_),
    .ZN(_0891_)
  );
  AND2_X1 _6171_ (
    .A1(_0790_),
    .A2(_0891_),
    .ZN(_0892_)
  );
  AND2_X1 _6172_ (
    .A1(_0455_),
    .A2(_0892_),
    .ZN(_0893_)
  );
  XOR2_X1 _6173_ (
    .A(_0455_),
    .B(_0892_),
    .Z(_0894_)
  );
  AND2_X1 _6174_ (
    .A1(_0890_),
    .A2(_0894_),
    .ZN(_0895_)
  );
  XOR2_X1 _6175_ (
    .A(_0890_),
    .B(_0894_),
    .Z(_0896_)
  );
  AND2_X1 _6176_ (
    .A1(_0889_),
    .A2(_0896_),
    .ZN(_0897_)
  );
  XOR2_X1 _6177_ (
    .A(_0889_),
    .B(_0896_),
    .Z(_0898_)
  );
  AND2_X1 _6178_ (
    .A1(_0888_),
    .A2(_0898_),
    .ZN(_0899_)
  );
  XOR2_X1 _6179_ (
    .A(_0888_),
    .B(_0898_),
    .Z(_0900_)
  );
  AND2_X1 _6180_ (
    .A1(_0887_),
    .A2(_0900_),
    .ZN(_0901_)
  );
  XOR2_X1 _6181_ (
    .A(_0887_),
    .B(_0900_),
    .Z(_0902_)
  );
  AND2_X1 _6182_ (
    .A1(_0886_),
    .A2(_0902_),
    .ZN(_0903_)
  );
  XOR2_X1 _6183_ (
    .A(_0886_),
    .B(_0902_),
    .Z(_0904_)
  );
  AND2_X1 _6184_ (
    .A1(_0512_),
    .A2(_0904_),
    .ZN(_0905_)
  );
  XOR2_X1 _6185_ (
    .A(_0512_),
    .B(_0904_),
    .Z(_0906_)
  );
  AND2_X1 _6186_ (
    .A1(_0885_),
    .A2(_0906_),
    .ZN(_0907_)
  );
  XOR2_X1 _6187_ (
    .A(_0885_),
    .B(_0906_),
    .Z(_0908_)
  );
  AND2_X1 _6188_ (
    .A1(divisor[13]),
    .A2(remainder[2]),
    .ZN(_0909_)
  );
  AND2_X1 _6189_ (
    .A1(divisor[15]),
    .A2(remainder[0]),
    .ZN(_0910_)
  );
  AND2_X1 _6190_ (
    .A1(divisor[15]),
    .A2(remainder[1]),
    .ZN(_0911_)
  );
  AND2_X1 _6191_ (
    .A1(_0808_),
    .A2(_0911_),
    .ZN(_0912_)
  );
  XOR2_X1 _6192_ (
    .A(_0810_),
    .B(_0910_),
    .Z(_0913_)
  );
  AND2_X1 _6193_ (
    .A1(_0909_),
    .A2(_0913_),
    .ZN(_0914_)
  );
  XOR2_X1 _6194_ (
    .A(_0909_),
    .B(_0913_),
    .Z(_0915_)
  );
  AND2_X1 _6195_ (
    .A1(_0811_),
    .A2(_0915_),
    .ZN(_0916_)
  );
  XOR2_X1 _6196_ (
    .A(_0811_),
    .B(_0915_),
    .Z(_0917_)
  );
  AND2_X1 _6197_ (
    .A1(divisor[10]),
    .A2(remainder[5]),
    .ZN(_0918_)
  );
  AND2_X1 _6198_ (
    .A1(divisor[11]),
    .A2(remainder[4]),
    .ZN(_0919_)
  );
  AND2_X1 _6199_ (
    .A1(divisor[12]),
    .A2(remainder[4]),
    .ZN(_0920_)
  );
  AND2_X1 _6200_ (
    .A1(_0815_),
    .A2(_0919_),
    .ZN(_0921_)
  );
  XOR2_X1 _6201_ (
    .A(_0815_),
    .B(_0919_),
    .Z(_0922_)
  );
  AND2_X1 _6202_ (
    .A1(_0918_),
    .A2(_0922_),
    .ZN(_0923_)
  );
  XOR2_X1 _6203_ (
    .A(_0918_),
    .B(_0922_),
    .Z(_0924_)
  );
  AND2_X1 _6204_ (
    .A1(_0917_),
    .A2(_0924_),
    .ZN(_0925_)
  );
  XOR2_X1 _6205_ (
    .A(_0917_),
    .B(_0924_),
    .Z(_0926_)
  );
  AND2_X1 _6206_ (
    .A1(_0820_),
    .A2(_0926_),
    .ZN(_0927_)
  );
  XOR2_X1 _6207_ (
    .A(_0820_),
    .B(_0926_),
    .Z(_0928_)
  );
  OR2_X1 _6208_ (
    .A1(_0829_),
    .A2(_0831_),
    .ZN(_0929_)
  );
  OR2_X1 _6209_ (
    .A1(_0816_),
    .A2(_0818_),
    .ZN(_0930_)
  );
  AND2_X1 _6210_ (
    .A1(remainder[32]),
    .A2(divisor[7]),
    .ZN(_0931_)
  );
  AND2_X1 _6211_ (
    .A1(divisor[8]),
    .A2(remainder[7]),
    .ZN(_0932_)
  );
  AND2_X1 _6212_ (
    .A1(divisor[9]),
    .A2(remainder[7]),
    .ZN(_0933_)
  );
  AND2_X1 _6213_ (
    .A1(_0827_),
    .A2(_0933_),
    .ZN(_0934_)
  );
  XOR2_X1 _6214_ (
    .A(_0828_),
    .B(_0932_),
    .Z(_0935_)
  );
  AND2_X1 _6215_ (
    .A1(_0931_),
    .A2(_0935_),
    .ZN(_0936_)
  );
  XOR2_X1 _6216_ (
    .A(_0931_),
    .B(_0935_),
    .Z(_0937_)
  );
  AND2_X1 _6217_ (
    .A1(_0930_),
    .A2(_0937_),
    .ZN(_0938_)
  );
  XOR2_X1 _6218_ (
    .A(_0930_),
    .B(_0937_),
    .Z(_0939_)
  );
  AND2_X1 _6219_ (
    .A1(_0929_),
    .A2(_0939_),
    .ZN(_0940_)
  );
  XOR2_X1 _6220_ (
    .A(_0929_),
    .B(_0939_),
    .Z(_0941_)
  );
  AND2_X1 _6221_ (
    .A1(_0928_),
    .A2(_0941_),
    .ZN(_0942_)
  );
  XOR2_X1 _6222_ (
    .A(_0928_),
    .B(_0941_),
    .Z(_0943_)
  );
  INV_X1 _6223_ (
    .A(_0943_),
    .ZN(_0944_)
  );
  XOR2_X1 _6224_ (
    .A(_0882_),
    .B(_0943_),
    .Z(_0945_)
  );
  AND2_X1 _6225_ (
    .A1(_0908_),
    .A2(_0945_),
    .ZN(_0946_)
  );
  XOR2_X1 _6226_ (
    .A(_0908_),
    .B(_0945_),
    .Z(_0947_)
  );
  AND2_X1 _6227_ (
    .A1(_0884_),
    .A2(_0947_),
    .ZN(_0948_)
  );
  XOR2_X1 _6228_ (
    .A(_0884_),
    .B(_0947_),
    .Z(_0949_)
  );
  AND2_X1 _6229_ (
    .A1(_0806_),
    .A2(_0949_),
    .ZN(_0950_)
  );
  XOR2_X1 _6230_ (
    .A(_0806_),
    .B(_0949_),
    .Z(_0951_)
  );
  AND2_X1 _6231_ (
    .A1(_0881_),
    .A2(_0951_),
    .ZN(_0952_)
  );
  XOR2_X1 _6232_ (
    .A(_0881_),
    .B(_0951_),
    .Z(_0953_)
  );
  AND2_X1 _6233_ (
    .A1(_0849_),
    .A2(_0953_),
    .ZN(_0954_)
  );
  XOR2_X1 _6234_ (
    .A(_0849_),
    .B(_0953_),
    .Z(_0955_)
  );
  AND2_X1 _6235_ (
    .A1(_0880_),
    .A2(_0955_),
    .ZN(_0956_)
  );
  XOR2_X1 _6236_ (
    .A(_0880_),
    .B(_0955_),
    .Z(_0957_)
  );
  AND2_X1 _6237_ (
    .A1(remainder[48]),
    .A2(_0957_),
    .ZN(_0958_)
  );
  INV_X1 _6238_ (
    .A(_0958_),
    .ZN(_0959_)
  );
  XOR2_X1 _6239_ (
    .A(remainder[48]),
    .B(_0957_),
    .Z(_0960_)
  );
  XOR2_X1 _6240_ (
    .A(_3078_),
    .B(_0957_),
    .Z(_0961_)
  );
  AND2_X1 _6241_ (
    .A1(_0879_),
    .A2(_0960_),
    .ZN(_0962_)
  );
  OR2_X1 _6242_ (
    .A1(_0878_),
    .A2(_0961_),
    .ZN(_0963_)
  );
  OR2_X1 _6243_ (
    .A1(_0879_),
    .A2(_0960_),
    .ZN(_0964_)
  );
  AND2_X1 _6244_ (
    .A1(_4613_),
    .A2(_0964_),
    .ZN(_0965_)
  );
  AND2_X1 _6245_ (
    .A1(_0963_),
    .A2(_0965_),
    .ZN(_0966_)
  );
  OR2_X1 _6246_ (
    .A1(_0877_),
    .A2(_0966_),
    .ZN(_0967_)
  );
  OR2_X1 _6247_ (
    .A1(_0876_),
    .A2(_0967_),
    .ZN(_0968_)
  );
  AND2_X1 _6248_ (
    .A1(_3911_),
    .A2(_0968_),
    .ZN(_0061_)
  );
  OR2_X1 _6249_ (
    .A1(remainder[40]),
    .A2(_4393_),
    .ZN(_0969_)
  );
  OR2_X1 _6250_ (
    .A1(_4392_),
    .A2(_4473_),
    .ZN(_0970_)
  );
  AND2_X1 _6251_ (
    .A1(_3678_),
    .A2(_0970_),
    .ZN(_0971_)
  );
  AND2_X1 _6252_ (
    .A1(_0969_),
    .A2(_0971_),
    .ZN(_0972_)
  );
  AND2_X1 _6253_ (
    .A1(remainder[41]),
    .A2(_4610_),
    .ZN(_0973_)
  );
  AND2_X1 _6254_ (
    .A1(_0959_),
    .A2(_0963_),
    .ZN(_0974_)
  );
  OR2_X1 _6255_ (
    .A1(_0958_),
    .A2(_0962_),
    .ZN(_0975_)
  );
  OR2_X1 _6256_ (
    .A1(_0954_),
    .A2(_0956_),
    .ZN(_0976_)
  );
  OR2_X1 _6257_ (
    .A1(_0948_),
    .A2(_0950_),
    .ZN(_0977_)
  );
  AND2_X1 _6258_ (
    .A1(_0541_),
    .A2(_0944_),
    .ZN(_0978_)
  );
  AND2_X1 _6259_ (
    .A1(_0838_),
    .A2(_0978_),
    .ZN(_0979_)
  );
  OR2_X1 _6260_ (
    .A1(_0946_),
    .A2(_0979_),
    .ZN(_0980_)
  );
  OR2_X1 _6261_ (
    .A1(_0903_),
    .A2(_0905_),
    .ZN(_0981_)
  );
  OR2_X1 _6262_ (
    .A1(_0899_),
    .A2(_0901_),
    .ZN(_0982_)
  );
  OR2_X1 _6263_ (
    .A1(_0895_),
    .A2(_0897_),
    .ZN(_0983_)
  );
  OR2_X1 _6264_ (
    .A1(_0927_),
    .A2(_0942_),
    .ZN(_0984_)
  );
  OR2_X1 _6265_ (
    .A1(_0789_),
    .A2(_0893_),
    .ZN(_0985_)
  );
  OR2_X1 _6266_ (
    .A1(_0938_),
    .A2(_0940_),
    .ZN(_0986_)
  );
  AND2_X1 _6267_ (
    .A1(_0894_),
    .A2(_0986_),
    .ZN(_0987_)
  );
  XOR2_X1 _6268_ (
    .A(_0894_),
    .B(_0986_),
    .Z(_0988_)
  );
  AND2_X1 _6269_ (
    .A1(_0985_),
    .A2(_0988_),
    .ZN(_0989_)
  );
  XOR2_X1 _6270_ (
    .A(_0985_),
    .B(_0988_),
    .Z(_0990_)
  );
  AND2_X1 _6271_ (
    .A1(_0984_),
    .A2(_0990_),
    .ZN(_0991_)
  );
  XOR2_X1 _6272_ (
    .A(_0984_),
    .B(_0990_),
    .Z(_0992_)
  );
  AND2_X1 _6273_ (
    .A1(_0983_),
    .A2(_0992_),
    .ZN(_0993_)
  );
  XOR2_X1 _6274_ (
    .A(_0983_),
    .B(_0992_),
    .Z(_0994_)
  );
  AND2_X1 _6275_ (
    .A1(_0982_),
    .A2(_0994_),
    .ZN(_0995_)
  );
  XOR2_X1 _6276_ (
    .A(_0982_),
    .B(_0994_),
    .Z(_0996_)
  );
  AND2_X1 _6277_ (
    .A1(_0512_),
    .A2(_0996_),
    .ZN(_0997_)
  );
  XOR2_X1 _6278_ (
    .A(_0512_),
    .B(_0996_),
    .Z(_0998_)
  );
  AND2_X1 _6279_ (
    .A1(_0981_),
    .A2(_0998_),
    .ZN(_0999_)
  );
  XOR2_X1 _6280_ (
    .A(_0981_),
    .B(_0998_),
    .Z(_1000_)
  );
  AND2_X1 _6281_ (
    .A1(divisor[16]),
    .A2(remainder[0]),
    .ZN(_1001_)
  );
  OR2_X1 _6282_ (
    .A1(_0916_),
    .A2(_0925_),
    .ZN(_1002_)
  );
  OR2_X1 _6283_ (
    .A1(_0912_),
    .A2(_0914_),
    .ZN(_1003_)
  );
  AND2_X1 _6284_ (
    .A1(divisor[13]),
    .A2(remainder[3]),
    .ZN(_1004_)
  );
  AND2_X1 _6285_ (
    .A1(divisor[14]),
    .A2(remainder[2]),
    .ZN(_1005_)
  );
  AND2_X1 _6286_ (
    .A1(divisor[15]),
    .A2(remainder[2]),
    .ZN(_1006_)
  );
  AND2_X1 _6287_ (
    .A1(_0810_),
    .A2(_1006_),
    .ZN(_1007_)
  );
  XOR2_X1 _6288_ (
    .A(_0911_),
    .B(_1005_),
    .Z(_1008_)
  );
  AND2_X1 _6289_ (
    .A1(_1004_),
    .A2(_1008_),
    .ZN(_1009_)
  );
  XOR2_X1 _6290_ (
    .A(_1004_),
    .B(_1008_),
    .Z(_1010_)
  );
  AND2_X1 _6291_ (
    .A1(_1003_),
    .A2(_1010_),
    .ZN(_1011_)
  );
  XOR2_X1 _6292_ (
    .A(_1003_),
    .B(_1010_),
    .Z(_1012_)
  );
  AND2_X1 _6293_ (
    .A1(divisor[10]),
    .A2(remainder[6]),
    .ZN(_1013_)
  );
  AND2_X1 _6294_ (
    .A1(divisor[11]),
    .A2(remainder[5]),
    .ZN(_1014_)
  );
  AND2_X1 _6295_ (
    .A1(divisor[12]),
    .A2(remainder[5]),
    .ZN(_1015_)
  );
  AND2_X1 _6296_ (
    .A1(_0920_),
    .A2(_1014_),
    .ZN(_1016_)
  );
  XOR2_X1 _6297_ (
    .A(_0920_),
    .B(_1014_),
    .Z(_1017_)
  );
  AND2_X1 _6298_ (
    .A1(_1013_),
    .A2(_1017_),
    .ZN(_1018_)
  );
  XOR2_X1 _6299_ (
    .A(_1013_),
    .B(_1017_),
    .Z(_1019_)
  );
  AND2_X1 _6300_ (
    .A1(_1012_),
    .A2(_1019_),
    .ZN(_1020_)
  );
  XOR2_X1 _6301_ (
    .A(_1012_),
    .B(_1019_),
    .Z(_1021_)
  );
  AND2_X1 _6302_ (
    .A1(_1002_),
    .A2(_1021_),
    .ZN(_1022_)
  );
  XOR2_X1 _6303_ (
    .A(_1002_),
    .B(_1021_),
    .Z(_1023_)
  );
  OR2_X1 _6304_ (
    .A1(_0934_),
    .A2(_0936_),
    .ZN(_1024_)
  );
  OR2_X1 _6305_ (
    .A1(_0921_),
    .A2(_0923_),
    .ZN(_1025_)
  );
  AND2_X1 _6306_ (
    .A1(remainder[32]),
    .A2(divisor[9]),
    .ZN(_1026_)
  );
  AND2_X1 _6307_ (
    .A1(remainder[32]),
    .A2(divisor[8]),
    .ZN(_1027_)
  );
  AND2_X1 _6308_ (
    .A1(divisor[9]),
    .A2(_1027_),
    .ZN(_1028_)
  );
  AND2_X1 _6309_ (
    .A1(_0933_),
    .A2(_1027_),
    .ZN(_1029_)
  );
  XOR2_X1 _6310_ (
    .A(_0933_),
    .B(_1027_),
    .Z(_1030_)
  );
  AND2_X1 _6311_ (
    .A1(_0931_),
    .A2(_1030_),
    .ZN(_1031_)
  );
  XOR2_X1 _6312_ (
    .A(_0931_),
    .B(_1030_),
    .Z(_1032_)
  );
  AND2_X1 _6313_ (
    .A1(_1025_),
    .A2(_1032_),
    .ZN(_1033_)
  );
  XOR2_X1 _6314_ (
    .A(_1025_),
    .B(_1032_),
    .Z(_1034_)
  );
  AND2_X1 _6315_ (
    .A1(_1024_),
    .A2(_1034_),
    .ZN(_1035_)
  );
  XOR2_X1 _6316_ (
    .A(_1024_),
    .B(_1034_),
    .Z(_1036_)
  );
  AND2_X1 _6317_ (
    .A1(_1023_),
    .A2(_1036_),
    .ZN(_1037_)
  );
  XOR2_X1 _6318_ (
    .A(_1023_),
    .B(_1036_),
    .Z(_1038_)
  );
  AND2_X1 _6319_ (
    .A1(_1001_),
    .A2(_1038_),
    .ZN(_1039_)
  );
  XOR2_X1 _6320_ (
    .A(_1001_),
    .B(_1038_),
    .Z(_1040_)
  );
  XOR2_X1 _6321_ (
    .A(_0978_),
    .B(_1040_),
    .Z(_1041_)
  );
  AND2_X1 _6322_ (
    .A1(_1000_),
    .A2(_1041_),
    .ZN(_1042_)
  );
  INV_X1 _6323_ (
    .A(_1042_),
    .ZN(_1043_)
  );
  XOR2_X1 _6324_ (
    .A(_1000_),
    .B(_1041_),
    .Z(_1044_)
  );
  AND2_X1 _6325_ (
    .A1(_0980_),
    .A2(_1044_),
    .ZN(_1045_)
  );
  XOR2_X1 _6326_ (
    .A(_0980_),
    .B(_1044_),
    .Z(_1046_)
  );
  AND2_X1 _6327_ (
    .A1(_0907_),
    .A2(_1046_),
    .ZN(_1047_)
  );
  XOR2_X1 _6328_ (
    .A(_0907_),
    .B(_1046_),
    .Z(_1048_)
  );
  AND2_X1 _6329_ (
    .A1(_0977_),
    .A2(_1048_),
    .ZN(_1049_)
  );
  XOR2_X1 _6330_ (
    .A(_0977_),
    .B(_1048_),
    .Z(_1050_)
  );
  AND2_X1 _6331_ (
    .A1(_0952_),
    .A2(_1050_),
    .ZN(_1051_)
  );
  XOR2_X1 _6332_ (
    .A(_0952_),
    .B(_1050_),
    .Z(_1052_)
  );
  AND2_X1 _6333_ (
    .A1(_0976_),
    .A2(_1052_),
    .ZN(_1053_)
  );
  XOR2_X1 _6334_ (
    .A(_0976_),
    .B(_1052_),
    .Z(_1054_)
  );
  AND2_X1 _6335_ (
    .A1(remainder[49]),
    .A2(_1054_),
    .ZN(_1055_)
  );
  INV_X1 _6336_ (
    .A(_1055_),
    .ZN(_1056_)
  );
  XOR2_X1 _6337_ (
    .A(remainder[49]),
    .B(_1054_),
    .Z(_1057_)
  );
  XOR2_X1 _6338_ (
    .A(_3067_),
    .B(_1054_),
    .Z(_1058_)
  );
  AND2_X1 _6339_ (
    .A1(_0975_),
    .A2(_1057_),
    .ZN(_1059_)
  );
  OR2_X1 _6340_ (
    .A1(_0974_),
    .A2(_1058_),
    .ZN(_1060_)
  );
  OR2_X1 _6341_ (
    .A1(_0975_),
    .A2(_1057_),
    .ZN(_1061_)
  );
  AND2_X1 _6342_ (
    .A1(_4613_),
    .A2(_1061_),
    .ZN(_1062_)
  );
  AND2_X1 _6343_ (
    .A1(_1060_),
    .A2(_1062_),
    .ZN(_1063_)
  );
  OR2_X1 _6344_ (
    .A1(_0973_),
    .A2(_1063_),
    .ZN(_1064_)
  );
  OR2_X1 _6345_ (
    .A1(_0972_),
    .A2(_1064_),
    .ZN(_1065_)
  );
  AND2_X1 _6346_ (
    .A1(_3911_),
    .A2(_1065_),
    .ZN(_0062_)
  );
  OR2_X1 _6347_ (
    .A1(remainder[41]),
    .A2(_4393_),
    .ZN(_1066_)
  );
  OR2_X1 _6348_ (
    .A1(_4392_),
    .A2(_4479_),
    .ZN(_1067_)
  );
  AND2_X1 _6349_ (
    .A1(_3678_),
    .A2(_1067_),
    .ZN(_1068_)
  );
  AND2_X1 _6350_ (
    .A1(_1066_),
    .A2(_1068_),
    .ZN(_1069_)
  );
  AND2_X1 _6351_ (
    .A1(remainder[42]),
    .A2(_4610_),
    .ZN(_1070_)
  );
  AND2_X1 _6352_ (
    .A1(_1056_),
    .A2(_1060_),
    .ZN(_1071_)
  );
  OR2_X1 _6353_ (
    .A1(_1055_),
    .A2(_1059_),
    .ZN(_1072_)
  );
  OR2_X1 _6354_ (
    .A1(_1051_),
    .A2(_1053_),
    .ZN(_1073_)
  );
  OR2_X1 _6355_ (
    .A1(_1045_),
    .A2(_1047_),
    .ZN(_1074_)
  );
  OR2_X1 _6356_ (
    .A1(_0542_),
    .A2(_1040_),
    .ZN(_1075_)
  );
  OR2_X1 _6357_ (
    .A1(_0944_),
    .A2(_1075_),
    .ZN(_1076_)
  );
  AND2_X1 _6358_ (
    .A1(_1043_),
    .A2(_1076_),
    .ZN(_1077_)
  );
  OR2_X1 _6359_ (
    .A1(_0995_),
    .A2(_0997_),
    .ZN(_1078_)
  );
  OR2_X1 _6360_ (
    .A1(_0991_),
    .A2(_0993_),
    .ZN(_1079_)
  );
  OR2_X1 _6361_ (
    .A1(_0987_),
    .A2(_0989_),
    .ZN(_1080_)
  );
  OR2_X1 _6362_ (
    .A1(_1022_),
    .A2(_1037_),
    .ZN(_1081_)
  );
  OR2_X1 _6363_ (
    .A1(_1033_),
    .A2(_1035_),
    .ZN(_1082_)
  );
  AND2_X1 _6364_ (
    .A1(_0894_),
    .A2(_1082_),
    .ZN(_1083_)
  );
  XOR2_X1 _6365_ (
    .A(_0894_),
    .B(_1082_),
    .Z(_1084_)
  );
  AND2_X1 _6366_ (
    .A1(_0985_),
    .A2(_1084_),
    .ZN(_1085_)
  );
  XOR2_X1 _6367_ (
    .A(_0985_),
    .B(_1084_),
    .Z(_1086_)
  );
  AND2_X1 _6368_ (
    .A1(_1081_),
    .A2(_1086_),
    .ZN(_1087_)
  );
  XOR2_X1 _6369_ (
    .A(_1081_),
    .B(_1086_),
    .Z(_1088_)
  );
  AND2_X1 _6370_ (
    .A1(_1080_),
    .A2(_1088_),
    .ZN(_1089_)
  );
  XOR2_X1 _6371_ (
    .A(_1080_),
    .B(_1088_),
    .Z(_1090_)
  );
  AND2_X1 _6372_ (
    .A1(_1079_),
    .A2(_1090_),
    .ZN(_1091_)
  );
  XOR2_X1 _6373_ (
    .A(_1079_),
    .B(_1090_),
    .Z(_1092_)
  );
  AND2_X1 _6374_ (
    .A1(_0512_),
    .A2(_1092_),
    .ZN(_1093_)
  );
  XOR2_X1 _6375_ (
    .A(_0512_),
    .B(_1092_),
    .Z(_1094_)
  );
  AND2_X1 _6376_ (
    .A1(_1078_),
    .A2(_1094_),
    .ZN(_1095_)
  );
  XOR2_X1 _6377_ (
    .A(_1078_),
    .B(_1094_),
    .Z(_1096_)
  );
  AND2_X1 _6378_ (
    .A1(divisor[17]),
    .A2(remainder[0]),
    .ZN(_1097_)
  );
  AND2_X1 _6379_ (
    .A1(divisor[16]),
    .A2(remainder[1]),
    .ZN(_1098_)
  );
  AND2_X1 _6380_ (
    .A1(divisor[17]),
    .A2(remainder[1]),
    .ZN(_1099_)
  );
  AND2_X1 _6381_ (
    .A1(_1001_),
    .A2(_1099_),
    .ZN(_1100_)
  );
  XOR2_X1 _6382_ (
    .A(_1097_),
    .B(_1098_),
    .Z(_1101_)
  );
  OR2_X1 _6383_ (
    .A1(_1011_),
    .A2(_1020_),
    .ZN(_1102_)
  );
  OR2_X1 _6384_ (
    .A1(_1007_),
    .A2(_1009_),
    .ZN(_1103_)
  );
  AND2_X1 _6385_ (
    .A1(divisor[13]),
    .A2(remainder[4]),
    .ZN(_1104_)
  );
  AND2_X1 _6386_ (
    .A1(divisor[14]),
    .A2(remainder[3]),
    .ZN(_1105_)
  );
  AND2_X1 _6387_ (
    .A1(divisor[15]),
    .A2(remainder[3]),
    .ZN(_1106_)
  );
  AND2_X1 _6388_ (
    .A1(_1006_),
    .A2(_1105_),
    .ZN(_1107_)
  );
  XOR2_X1 _6389_ (
    .A(_1006_),
    .B(_1105_),
    .Z(_1108_)
  );
  AND2_X1 _6390_ (
    .A1(_1104_),
    .A2(_1108_),
    .ZN(_1109_)
  );
  XOR2_X1 _6391_ (
    .A(_1104_),
    .B(_1108_),
    .Z(_1110_)
  );
  AND2_X1 _6392_ (
    .A1(_1103_),
    .A2(_1110_),
    .ZN(_1111_)
  );
  XOR2_X1 _6393_ (
    .A(_1103_),
    .B(_1110_),
    .Z(_1112_)
  );
  AND2_X1 _6394_ (
    .A1(divisor[10]),
    .A2(remainder[7]),
    .ZN(_1113_)
  );
  AND2_X1 _6395_ (
    .A1(divisor[11]),
    .A2(remainder[6]),
    .ZN(_1114_)
  );
  AND2_X1 _6396_ (
    .A1(divisor[12]),
    .A2(remainder[6]),
    .ZN(_1115_)
  );
  AND2_X1 _6397_ (
    .A1(_1015_),
    .A2(_1114_),
    .ZN(_1116_)
  );
  XOR2_X1 _6398_ (
    .A(_1015_),
    .B(_1114_),
    .Z(_1117_)
  );
  AND2_X1 _6399_ (
    .A1(_1113_),
    .A2(_1117_),
    .ZN(_1118_)
  );
  XOR2_X1 _6400_ (
    .A(_1113_),
    .B(_1117_),
    .Z(_1119_)
  );
  AND2_X1 _6401_ (
    .A1(_1112_),
    .A2(_1119_),
    .ZN(_1120_)
  );
  XOR2_X1 _6402_ (
    .A(_1112_),
    .B(_1119_),
    .Z(_1121_)
  );
  AND2_X1 _6403_ (
    .A1(_1102_),
    .A2(_1121_),
    .ZN(_1122_)
  );
  XOR2_X1 _6404_ (
    .A(_1102_),
    .B(_1121_),
    .Z(_1123_)
  );
  OR2_X1 _6405_ (
    .A1(_1029_),
    .A2(_1031_),
    .ZN(_1124_)
  );
  OR2_X1 _6406_ (
    .A1(_1016_),
    .A2(_1018_),
    .ZN(_1125_)
  );
  MUX2_X1 _6407_ (
    .A(_1027_),
    .B(_3296_),
    .S(_1026_),
    .Z(_1126_)
  );
  AND2_X1 _6408_ (
    .A1(divisor[7]),
    .A2(_1126_),
    .ZN(_1127_)
  );
  MUX2_X1 _6409_ (
    .A(_0931_),
    .B(_3285_),
    .S(_1126_),
    .Z(_1128_)
  );
  AND2_X1 _6410_ (
    .A1(_1125_),
    .A2(_1128_),
    .ZN(_1129_)
  );
  XOR2_X1 _6411_ (
    .A(_1125_),
    .B(_1128_),
    .Z(_1130_)
  );
  AND2_X1 _6412_ (
    .A1(_1124_),
    .A2(_1130_),
    .ZN(_1131_)
  );
  XOR2_X1 _6413_ (
    .A(_1124_),
    .B(_1130_),
    .Z(_1132_)
  );
  AND2_X1 _6414_ (
    .A1(_1123_),
    .A2(_1132_),
    .ZN(_1133_)
  );
  XOR2_X1 _6415_ (
    .A(_1123_),
    .B(_1132_),
    .Z(_1134_)
  );
  AND2_X1 _6416_ (
    .A1(_1101_),
    .A2(_1134_),
    .ZN(_1135_)
  );
  XOR2_X1 _6417_ (
    .A(_1101_),
    .B(_1134_),
    .Z(_1136_)
  );
  AND2_X1 _6418_ (
    .A1(_1039_),
    .A2(_1136_),
    .ZN(_1137_)
  );
  XOR2_X1 _6419_ (
    .A(_1039_),
    .B(_1136_),
    .Z(_1138_)
  );
  INV_X1 _6420_ (
    .A(_1138_),
    .ZN(_1139_)
  );
  XOR2_X1 _6421_ (
    .A(_1075_),
    .B(_1138_),
    .Z(_1140_)
  );
  XOR2_X1 _6422_ (
    .A(_1075_),
    .B(_1139_),
    .Z(_1141_)
  );
  AND2_X1 _6423_ (
    .A1(_1096_),
    .A2(_1141_),
    .ZN(_1142_)
  );
  XOR2_X1 _6424_ (
    .A(_1096_),
    .B(_1140_),
    .Z(_1143_)
  );
  OR2_X1 _6425_ (
    .A1(_1077_),
    .A2(_1143_),
    .ZN(_1144_)
  );
  INV_X1 _6426_ (
    .A(_1144_),
    .ZN(_1145_)
  );
  XOR2_X1 _6427_ (
    .A(_1077_),
    .B(_1143_),
    .Z(_1146_)
  );
  AND2_X1 _6428_ (
    .A1(_0999_),
    .A2(_1146_),
    .ZN(_1147_)
  );
  XOR2_X1 _6429_ (
    .A(_0999_),
    .B(_1146_),
    .Z(_1148_)
  );
  AND2_X1 _6430_ (
    .A1(_1074_),
    .A2(_1148_),
    .ZN(_1149_)
  );
  XOR2_X1 _6431_ (
    .A(_1074_),
    .B(_1148_),
    .Z(_1150_)
  );
  AND2_X1 _6432_ (
    .A1(_1049_),
    .A2(_1150_),
    .ZN(_1151_)
  );
  OR2_X1 _6433_ (
    .A1(_1049_),
    .A2(_1150_),
    .ZN(_1152_)
  );
  XOR2_X1 _6434_ (
    .A(_1049_),
    .B(_1150_),
    .Z(_1153_)
  );
  INV_X1 _6435_ (
    .A(_1153_),
    .ZN(_1154_)
  );
  XOR2_X1 _6436_ (
    .A(_1073_),
    .B(_1154_),
    .Z(_1155_)
  );
  XOR2_X1 _6437_ (
    .A(_1073_),
    .B(_1153_),
    .Z(_1156_)
  );
  AND2_X1 _6438_ (
    .A1(remainder[50]),
    .A2(_1156_),
    .ZN(_1157_)
  );
  OR2_X1 _6439_ (
    .A1(_3056_),
    .A2(_1155_),
    .ZN(_1158_)
  );
  OR2_X1 _6440_ (
    .A1(remainder[50]),
    .A2(_1156_),
    .ZN(_1159_)
  );
  INV_X1 _6441_ (
    .A(_1159_),
    .ZN(_1160_)
  );
  AND2_X1 _6442_ (
    .A1(_1158_),
    .A2(_1159_),
    .ZN(_1161_)
  );
  XOR2_X1 _6443_ (
    .A(_1072_),
    .B(_1161_),
    .Z(_1162_)
  );
  AND2_X1 _6444_ (
    .A1(_4613_),
    .A2(_1162_),
    .ZN(_1163_)
  );
  OR2_X1 _6445_ (
    .A1(_1070_),
    .A2(_1163_),
    .ZN(_1164_)
  );
  OR2_X1 _6446_ (
    .A1(_1069_),
    .A2(_1164_),
    .ZN(_1165_)
  );
  AND2_X1 _6447_ (
    .A1(_3911_),
    .A2(_1165_),
    .ZN(_0063_)
  );
  OR2_X1 _6448_ (
    .A1(remainder[42]),
    .A2(_4393_),
    .ZN(_1166_)
  );
  OR2_X1 _6449_ (
    .A1(_4392_),
    .A2(_4484_),
    .ZN(_1167_)
  );
  AND2_X1 _6450_ (
    .A1(_3678_),
    .A2(_1167_),
    .ZN(_1168_)
  );
  AND2_X1 _6451_ (
    .A1(_1166_),
    .A2(_1168_),
    .ZN(_1169_)
  );
  AND2_X1 _6452_ (
    .A1(remainder[43]),
    .A2(_4610_),
    .ZN(_1170_)
  );
  AND2_X1 _6453_ (
    .A1(_1053_),
    .A2(_1153_),
    .ZN(_1171_)
  );
  AND2_X1 _6454_ (
    .A1(_1051_),
    .A2(_1152_),
    .ZN(_1172_)
  );
  OR2_X1 _6455_ (
    .A1(_1151_),
    .A2(_1172_),
    .ZN(_1173_)
  );
  OR2_X1 _6456_ (
    .A1(_1171_),
    .A2(_1173_),
    .ZN(_1174_)
  );
  OR2_X1 _6457_ (
    .A1(_1145_),
    .A2(_1147_),
    .ZN(_1175_)
  );
  AND2_X1 _6458_ (
    .A1(_0541_),
    .A2(_1139_),
    .ZN(_1176_)
  );
  AND2_X1 _6459_ (
    .A1(_1040_),
    .A2(_1176_),
    .ZN(_1177_)
  );
  OR2_X1 _6460_ (
    .A1(_1142_),
    .A2(_1177_),
    .ZN(_1178_)
  );
  OR2_X1 _6461_ (
    .A1(_1091_),
    .A2(_1093_),
    .ZN(_1179_)
  );
  OR2_X1 _6462_ (
    .A1(_1087_),
    .A2(_1089_),
    .ZN(_1180_)
  );
  OR2_X1 _6463_ (
    .A1(_1083_),
    .A2(_1085_),
    .ZN(_1181_)
  );
  INV_X1 _6464_ (
    .A(_1181_),
    .ZN(_1182_)
  );
  OR2_X1 _6465_ (
    .A1(_1122_),
    .A2(_1133_),
    .ZN(_1183_)
  );
  OR2_X1 _6466_ (
    .A1(_1129_),
    .A2(_1131_),
    .ZN(_1184_)
  );
  AND2_X1 _6467_ (
    .A1(_0894_),
    .A2(_1184_),
    .ZN(_1185_)
  );
  XOR2_X1 _6468_ (
    .A(_0894_),
    .B(_1184_),
    .Z(_1186_)
  );
  AND2_X1 _6469_ (
    .A1(_0985_),
    .A2(_1186_),
    .ZN(_1187_)
  );
  XOR2_X1 _6470_ (
    .A(_0985_),
    .B(_1186_),
    .Z(_1188_)
  );
  AND2_X1 _6471_ (
    .A1(_1183_),
    .A2(_1188_),
    .ZN(_1189_)
  );
  XOR2_X1 _6472_ (
    .A(_1183_),
    .B(_1188_),
    .Z(_1190_)
  );
  AND2_X1 _6473_ (
    .A1(_1181_),
    .A2(_1190_),
    .ZN(_1191_)
  );
  XOR2_X1 _6474_ (
    .A(_1181_),
    .B(_1190_),
    .Z(_1192_)
  );
  XOR2_X1 _6475_ (
    .A(_1182_),
    .B(_1190_),
    .Z(_1193_)
  );
  AND2_X1 _6476_ (
    .A1(_1180_),
    .A2(_1192_),
    .ZN(_1194_)
  );
  XOR2_X1 _6477_ (
    .A(_1180_),
    .B(_1193_),
    .Z(_1195_)
  );
  INV_X1 _6478_ (
    .A(_1195_),
    .ZN(_1196_)
  );
  AND2_X1 _6479_ (
    .A1(_0512_),
    .A2(_1196_),
    .ZN(_1197_)
  );
  XOR2_X1 _6480_ (
    .A(_0511_),
    .B(_1195_),
    .Z(_1198_)
  );
  AND2_X1 _6481_ (
    .A1(_1137_),
    .A2(_1198_),
    .ZN(_1199_)
  );
  XOR2_X1 _6482_ (
    .A(_1137_),
    .B(_1198_),
    .Z(_1200_)
  );
  AND2_X1 _6483_ (
    .A1(_1179_),
    .A2(_1200_),
    .ZN(_1201_)
  );
  XOR2_X1 _6484_ (
    .A(_1179_),
    .B(_1200_),
    .Z(_1202_)
  );
  AND2_X1 _6485_ (
    .A1(divisor[16]),
    .A2(remainder[2]),
    .ZN(_1203_)
  );
  AND2_X1 _6486_ (
    .A1(divisor[18]),
    .A2(remainder[0]),
    .ZN(_1204_)
  );
  AND2_X1 _6487_ (
    .A1(divisor[18]),
    .A2(remainder[1]),
    .ZN(_1205_)
  );
  AND2_X1 _6488_ (
    .A1(_1097_),
    .A2(_1205_),
    .ZN(_1206_)
  );
  XOR2_X1 _6489_ (
    .A(_1099_),
    .B(_1204_),
    .Z(_1207_)
  );
  AND2_X1 _6490_ (
    .A1(_1203_),
    .A2(_1207_),
    .ZN(_1208_)
  );
  XOR2_X1 _6491_ (
    .A(_1203_),
    .B(_1207_),
    .Z(_1209_)
  );
  AND2_X1 _6492_ (
    .A1(_1100_),
    .A2(_1209_),
    .ZN(_1210_)
  );
  XOR2_X1 _6493_ (
    .A(_1100_),
    .B(_1209_),
    .Z(_1211_)
  );
  OR2_X1 _6494_ (
    .A1(_1111_),
    .A2(_1120_),
    .ZN(_1212_)
  );
  OR2_X1 _6495_ (
    .A1(_1107_),
    .A2(_1109_),
    .ZN(_1213_)
  );
  AND2_X1 _6496_ (
    .A1(divisor[13]),
    .A2(remainder[5]),
    .ZN(_1214_)
  );
  AND2_X1 _6497_ (
    .A1(divisor[14]),
    .A2(remainder[4]),
    .ZN(_1215_)
  );
  AND2_X1 _6498_ (
    .A1(divisor[15]),
    .A2(remainder[4]),
    .ZN(_1216_)
  );
  AND2_X1 _6499_ (
    .A1(_1106_),
    .A2(_1215_),
    .ZN(_1217_)
  );
  XOR2_X1 _6500_ (
    .A(_1106_),
    .B(_1215_),
    .Z(_1218_)
  );
  AND2_X1 _6501_ (
    .A1(_1214_),
    .A2(_1218_),
    .ZN(_1219_)
  );
  XOR2_X1 _6502_ (
    .A(_1214_),
    .B(_1218_),
    .Z(_1220_)
  );
  AND2_X1 _6503_ (
    .A1(_1213_),
    .A2(_1220_),
    .ZN(_1221_)
  );
  XOR2_X1 _6504_ (
    .A(_1213_),
    .B(_1220_),
    .Z(_1222_)
  );
  AND2_X1 _6505_ (
    .A1(remainder[32]),
    .A2(divisor[10]),
    .ZN(_1223_)
  );
  AND2_X1 _6506_ (
    .A1(divisor[11]),
    .A2(remainder[7]),
    .ZN(_1224_)
  );
  AND2_X1 _6507_ (
    .A1(divisor[12]),
    .A2(remainder[7]),
    .ZN(_1225_)
  );
  AND2_X1 _6508_ (
    .A1(_1114_),
    .A2(_1225_),
    .ZN(_1226_)
  );
  XOR2_X1 _6509_ (
    .A(_1115_),
    .B(_1224_),
    .Z(_1227_)
  );
  AND2_X1 _6510_ (
    .A1(_1223_),
    .A2(_1227_),
    .ZN(_1228_)
  );
  XOR2_X1 _6511_ (
    .A(_1223_),
    .B(_1227_),
    .Z(_1229_)
  );
  AND2_X1 _6512_ (
    .A1(_1222_),
    .A2(_1229_),
    .ZN(_1230_)
  );
  XOR2_X1 _6513_ (
    .A(_1222_),
    .B(_1229_),
    .Z(_1231_)
  );
  AND2_X1 _6514_ (
    .A1(_1212_),
    .A2(_1231_),
    .ZN(_1232_)
  );
  XOR2_X1 _6515_ (
    .A(_1212_),
    .B(_1231_),
    .Z(_1233_)
  );
  OR2_X1 _6516_ (
    .A1(_1028_),
    .A2(_1127_),
    .ZN(_1234_)
  );
  INV_X1 _6517_ (
    .A(_1234_),
    .ZN(_1235_)
  );
  OR2_X1 _6518_ (
    .A1(_1116_),
    .A2(_1118_),
    .ZN(_1236_)
  );
  AND2_X1 _6519_ (
    .A1(_1128_),
    .A2(_1236_),
    .ZN(_1237_)
  );
  XOR2_X1 _6520_ (
    .A(_1128_),
    .B(_1236_),
    .Z(_1238_)
  );
  AND2_X1 _6521_ (
    .A1(_1234_),
    .A2(_1238_),
    .ZN(_1239_)
  );
  XOR2_X1 _6522_ (
    .A(_1234_),
    .B(_1238_),
    .Z(_1240_)
  );
  AND2_X1 _6523_ (
    .A1(_1233_),
    .A2(_1240_),
    .ZN(_1241_)
  );
  XOR2_X1 _6524_ (
    .A(_1233_),
    .B(_1240_),
    .Z(_1242_)
  );
  AND2_X1 _6525_ (
    .A1(_1211_),
    .A2(_1242_),
    .ZN(_1243_)
  );
  XOR2_X1 _6526_ (
    .A(_1211_),
    .B(_1242_),
    .Z(_1244_)
  );
  AND2_X1 _6527_ (
    .A1(_1135_),
    .A2(_1244_),
    .ZN(_1245_)
  );
  XOR2_X1 _6528_ (
    .A(_1135_),
    .B(_1244_),
    .Z(_1246_)
  );
  INV_X1 _6529_ (
    .A(_1246_),
    .ZN(_1247_)
  );
  XOR2_X1 _6530_ (
    .A(_1176_),
    .B(_1246_),
    .Z(_1248_)
  );
  AND2_X1 _6531_ (
    .A1(_1202_),
    .A2(_1248_),
    .ZN(_1249_)
  );
  XOR2_X1 _6532_ (
    .A(_1202_),
    .B(_1248_),
    .Z(_1250_)
  );
  AND2_X1 _6533_ (
    .A1(_1178_),
    .A2(_1250_),
    .ZN(_1251_)
  );
  XOR2_X1 _6534_ (
    .A(_1178_),
    .B(_1250_),
    .Z(_1252_)
  );
  AND2_X1 _6535_ (
    .A1(_1095_),
    .A2(_1252_),
    .ZN(_1253_)
  );
  XOR2_X1 _6536_ (
    .A(_1095_),
    .B(_1252_),
    .Z(_1254_)
  );
  AND2_X1 _6537_ (
    .A1(_1175_),
    .A2(_1254_),
    .ZN(_1255_)
  );
  XOR2_X1 _6538_ (
    .A(_1175_),
    .B(_1254_),
    .Z(_1256_)
  );
  AND2_X1 _6539_ (
    .A1(_1149_),
    .A2(_1256_),
    .ZN(_1257_)
  );
  XOR2_X1 _6540_ (
    .A(_1149_),
    .B(_1256_),
    .Z(_1258_)
  );
  AND2_X1 _6541_ (
    .A1(_1174_),
    .A2(_1258_),
    .ZN(_1259_)
  );
  XOR2_X1 _6542_ (
    .A(_1174_),
    .B(_1258_),
    .Z(_1260_)
  );
  AND2_X1 _6543_ (
    .A1(remainder[51]),
    .A2(_1260_),
    .ZN(_1261_)
  );
  INV_X1 _6544_ (
    .A(_1261_),
    .ZN(_1262_)
  );
  XOR2_X1 _6545_ (
    .A(remainder[51]),
    .B(_1260_),
    .Z(_1263_)
  );
  INV_X1 _6546_ (
    .A(_1263_),
    .ZN(_1264_)
  );
  AND2_X1 _6547_ (
    .A1(_1071_),
    .A2(_1158_),
    .ZN(_1265_)
  );
  OR2_X1 _6548_ (
    .A1(_1072_),
    .A2(_1157_),
    .ZN(_1266_)
  );
  AND2_X1 _6549_ (
    .A1(_1159_),
    .A2(_1266_),
    .ZN(_1267_)
  );
  OR2_X1 _6550_ (
    .A1(_1160_),
    .A2(_1265_),
    .ZN(_1268_)
  );
  AND2_X1 _6551_ (
    .A1(_1263_),
    .A2(_1267_),
    .ZN(_1269_)
  );
  OR2_X1 _6552_ (
    .A1(_1264_),
    .A2(_1268_),
    .ZN(_1270_)
  );
  OR2_X1 _6553_ (
    .A1(_1263_),
    .A2(_1267_),
    .ZN(_1271_)
  );
  AND2_X1 _6554_ (
    .A1(_4613_),
    .A2(_1271_),
    .ZN(_1272_)
  );
  AND2_X1 _6555_ (
    .A1(_1270_),
    .A2(_1272_),
    .ZN(_1273_)
  );
  OR2_X1 _6556_ (
    .A1(_1170_),
    .A2(_1273_),
    .ZN(_1274_)
  );
  OR2_X1 _6557_ (
    .A1(_1169_),
    .A2(_1274_),
    .ZN(_1275_)
  );
  AND2_X1 _6558_ (
    .A1(_3911_),
    .A2(_1275_),
    .ZN(_0064_)
  );
  OR2_X1 _6559_ (
    .A1(_4392_),
    .A2(_4490_),
    .ZN(_1276_)
  );
  OR2_X1 _6560_ (
    .A1(remainder[43]),
    .A2(_4393_),
    .ZN(_1277_)
  );
  AND2_X1 _6561_ (
    .A1(_3678_),
    .A2(_1276_),
    .ZN(_1278_)
  );
  AND2_X1 _6562_ (
    .A1(_1277_),
    .A2(_1278_),
    .ZN(_1279_)
  );
  AND2_X1 _6563_ (
    .A1(remainder[44]),
    .A2(_4610_),
    .ZN(_1280_)
  );
  AND2_X1 _6564_ (
    .A1(_1262_),
    .A2(_1270_),
    .ZN(_1281_)
  );
  OR2_X1 _6565_ (
    .A1(_1261_),
    .A2(_1269_),
    .ZN(_1282_)
  );
  OR2_X1 _6566_ (
    .A1(_1257_),
    .A2(_1259_),
    .ZN(_1283_)
  );
  OR2_X1 _6567_ (
    .A1(_1251_),
    .A2(_1253_),
    .ZN(_1284_)
  );
  OR2_X1 _6568_ (
    .A1(_1199_),
    .A2(_1201_),
    .ZN(_1285_)
  );
  AND2_X1 _6569_ (
    .A1(_0541_),
    .A2(_1138_),
    .ZN(_1286_)
  );
  AND2_X1 _6570_ (
    .A1(_1247_),
    .A2(_1286_),
    .ZN(_1287_)
  );
  OR2_X1 _6571_ (
    .A1(_1249_),
    .A2(_1287_),
    .ZN(_1288_)
  );
  AND2_X1 _6572_ (
    .A1(_0541_),
    .A2(_1246_),
    .ZN(_1289_)
  );
  OR2_X1 _6573_ (
    .A1(_1206_),
    .A2(_1208_),
    .ZN(_1290_)
  );
  AND2_X1 _6574_ (
    .A1(divisor[16]),
    .A2(remainder[3]),
    .ZN(_1291_)
  );
  AND2_X1 _6575_ (
    .A1(divisor[17]),
    .A2(remainder[2]),
    .ZN(_1292_)
  );
  AND2_X1 _6576_ (
    .A1(divisor[18]),
    .A2(remainder[2]),
    .ZN(_1293_)
  );
  AND2_X1 _6577_ (
    .A1(_1099_),
    .A2(_1293_),
    .ZN(_1294_)
  );
  XOR2_X1 _6578_ (
    .A(_1205_),
    .B(_1292_),
    .Z(_1295_)
  );
  AND2_X1 _6579_ (
    .A1(_1291_),
    .A2(_1295_),
    .ZN(_1296_)
  );
  XOR2_X1 _6580_ (
    .A(_1291_),
    .B(_1295_),
    .Z(_1297_)
  );
  AND2_X1 _6581_ (
    .A1(_1290_),
    .A2(_1297_),
    .ZN(_1298_)
  );
  XOR2_X1 _6582_ (
    .A(_1290_),
    .B(_1297_),
    .Z(_1299_)
  );
  AND2_X1 _6583_ (
    .A1(_1210_),
    .A2(_1299_),
    .ZN(_1300_)
  );
  XOR2_X1 _6584_ (
    .A(_1210_),
    .B(_1299_),
    .Z(_1301_)
  );
  OR2_X1 _6585_ (
    .A1(_1221_),
    .A2(_1230_),
    .ZN(_1302_)
  );
  OR2_X1 _6586_ (
    .A1(_1217_),
    .A2(_1219_),
    .ZN(_1303_)
  );
  AND2_X1 _6587_ (
    .A1(divisor[13]),
    .A2(remainder[6]),
    .ZN(_1304_)
  );
  AND2_X1 _6588_ (
    .A1(divisor[14]),
    .A2(remainder[5]),
    .ZN(_1305_)
  );
  AND2_X1 _6589_ (
    .A1(divisor[15]),
    .A2(remainder[5]),
    .ZN(_1306_)
  );
  AND2_X1 _6590_ (
    .A1(_1216_),
    .A2(_1305_),
    .ZN(_1307_)
  );
  XOR2_X1 _6591_ (
    .A(_1216_),
    .B(_1305_),
    .Z(_1308_)
  );
  AND2_X1 _6592_ (
    .A1(_1304_),
    .A2(_1308_),
    .ZN(_1309_)
  );
  XOR2_X1 _6593_ (
    .A(_1304_),
    .B(_1308_),
    .Z(_1310_)
  );
  AND2_X1 _6594_ (
    .A1(_1303_),
    .A2(_1310_),
    .ZN(_1311_)
  );
  XOR2_X1 _6595_ (
    .A(_1303_),
    .B(_1310_),
    .Z(_1312_)
  );
  AND2_X1 _6596_ (
    .A1(remainder[32]),
    .A2(divisor[12]),
    .ZN(_1313_)
  );
  AND2_X1 _6597_ (
    .A1(remainder[32]),
    .A2(divisor[11]),
    .ZN(_1314_)
  );
  AND2_X1 _6598_ (
    .A1(divisor[12]),
    .A2(_1314_),
    .ZN(_1315_)
  );
  AND2_X1 _6599_ (
    .A1(_1225_),
    .A2(_1314_),
    .ZN(_1316_)
  );
  XOR2_X1 _6600_ (
    .A(_1225_),
    .B(_1314_),
    .Z(_1317_)
  );
  AND2_X1 _6601_ (
    .A1(_1223_),
    .A2(_1317_),
    .ZN(_1318_)
  );
  XOR2_X1 _6602_ (
    .A(_1223_),
    .B(_1317_),
    .Z(_1319_)
  );
  AND2_X1 _6603_ (
    .A1(_1312_),
    .A2(_1319_),
    .ZN(_1320_)
  );
  XOR2_X1 _6604_ (
    .A(_1312_),
    .B(_1319_),
    .Z(_1321_)
  );
  AND2_X1 _6605_ (
    .A1(_1302_),
    .A2(_1321_),
    .ZN(_1322_)
  );
  XOR2_X1 _6606_ (
    .A(_1302_),
    .B(_1321_),
    .Z(_1323_)
  );
  OR2_X1 _6607_ (
    .A1(_1226_),
    .A2(_1228_),
    .ZN(_1324_)
  );
  AND2_X1 _6608_ (
    .A1(_1128_),
    .A2(_1324_),
    .ZN(_1325_)
  );
  XOR2_X1 _6609_ (
    .A(_1128_),
    .B(_1324_),
    .Z(_1326_)
  );
  AND2_X1 _6610_ (
    .A1(_1234_),
    .A2(_1326_),
    .ZN(_1327_)
  );
  XOR2_X1 _6611_ (
    .A(_1234_),
    .B(_1326_),
    .Z(_1328_)
  );
  AND2_X1 _6612_ (
    .A1(_1323_),
    .A2(_1328_),
    .ZN(_1329_)
  );
  XOR2_X1 _6613_ (
    .A(_1323_),
    .B(_1328_),
    .Z(_1330_)
  );
  AND2_X1 _6614_ (
    .A1(_1301_),
    .A2(_1330_),
    .ZN(_1331_)
  );
  XOR2_X1 _6615_ (
    .A(_1301_),
    .B(_1330_),
    .Z(_1332_)
  );
  AND2_X1 _6616_ (
    .A1(_1243_),
    .A2(_1332_),
    .ZN(_1333_)
  );
  XOR2_X1 _6617_ (
    .A(_1243_),
    .B(_1332_),
    .Z(_1334_)
  );
  AND2_X1 _6618_ (
    .A1(divisor[19]),
    .A2(remainder[0]),
    .ZN(_1335_)
  );
  OR2_X1 _6619_ (
    .A1(_0542_),
    .A2(_1335_),
    .ZN(_1336_)
  );
  AND2_X1 _6620_ (
    .A1(remainder[32]),
    .A2(divisor[19]),
    .ZN(_1337_)
  );
  XOR2_X1 _6621_ (
    .A(_0542_),
    .B(_1335_),
    .Z(_1338_)
  );
  XOR2_X1 _6622_ (
    .A(_0541_),
    .B(_1335_),
    .Z(_1339_)
  );
  AND2_X1 _6623_ (
    .A1(_1334_),
    .A2(_1339_),
    .ZN(_1340_)
  );
  XOR2_X1 _6624_ (
    .A(_1334_),
    .B(_1338_),
    .Z(_1341_)
  );
  INV_X1 _6625_ (
    .A(_1341_),
    .ZN(_1342_)
  );
  AND2_X1 _6626_ (
    .A1(_1289_),
    .A2(_1342_),
    .ZN(_1343_)
  );
  XOR2_X1 _6627_ (
    .A(_1289_),
    .B(_1342_),
    .Z(_1344_)
  );
  OR2_X1 _6628_ (
    .A1(_1194_),
    .A2(_1197_),
    .ZN(_1345_)
  );
  OR2_X1 _6629_ (
    .A1(_1189_),
    .A2(_1191_),
    .ZN(_1346_)
  );
  OR2_X1 _6630_ (
    .A1(_1185_),
    .A2(_1187_),
    .ZN(_1347_)
  );
  OR2_X1 _6631_ (
    .A1(_1232_),
    .A2(_1241_),
    .ZN(_1348_)
  );
  OR2_X1 _6632_ (
    .A1(_1237_),
    .A2(_1239_),
    .ZN(_1349_)
  );
  AND2_X1 _6633_ (
    .A1(_0894_),
    .A2(_1349_),
    .ZN(_1350_)
  );
  XOR2_X1 _6634_ (
    .A(_0894_),
    .B(_1349_),
    .Z(_1351_)
  );
  AND2_X1 _6635_ (
    .A1(_0985_),
    .A2(_1351_),
    .ZN(_1352_)
  );
  XOR2_X1 _6636_ (
    .A(_0985_),
    .B(_1351_),
    .Z(_1353_)
  );
  AND2_X1 _6637_ (
    .A1(_1348_),
    .A2(_1353_),
    .ZN(_1354_)
  );
  XOR2_X1 _6638_ (
    .A(_1348_),
    .B(_1353_),
    .Z(_1355_)
  );
  AND2_X1 _6639_ (
    .A1(_1347_),
    .A2(_1355_),
    .ZN(_1356_)
  );
  XOR2_X1 _6640_ (
    .A(_1347_),
    .B(_1355_),
    .Z(_1357_)
  );
  AND2_X1 _6641_ (
    .A1(_1346_),
    .A2(_1357_),
    .ZN(_1358_)
  );
  XOR2_X1 _6642_ (
    .A(_1346_),
    .B(_1357_),
    .Z(_1359_)
  );
  AND2_X1 _6643_ (
    .A1(_0512_),
    .A2(_1359_),
    .ZN(_1360_)
  );
  XOR2_X1 _6644_ (
    .A(_0512_),
    .B(_1359_),
    .Z(_1361_)
  );
  AND2_X1 _6645_ (
    .A1(_1245_),
    .A2(_1361_),
    .ZN(_1362_)
  );
  XOR2_X1 _6646_ (
    .A(_1245_),
    .B(_1361_),
    .Z(_1363_)
  );
  AND2_X1 _6647_ (
    .A1(_1345_),
    .A2(_1363_),
    .ZN(_1364_)
  );
  XOR2_X1 _6648_ (
    .A(_1345_),
    .B(_1363_),
    .Z(_1365_)
  );
  AND2_X1 _6649_ (
    .A1(_1344_),
    .A2(_1365_),
    .ZN(_1366_)
  );
  XOR2_X1 _6650_ (
    .A(_1344_),
    .B(_1365_),
    .Z(_1367_)
  );
  AND2_X1 _6651_ (
    .A1(_1288_),
    .A2(_1367_),
    .ZN(_1368_)
  );
  XOR2_X1 _6652_ (
    .A(_1288_),
    .B(_1367_),
    .Z(_1369_)
  );
  AND2_X1 _6653_ (
    .A1(_1285_),
    .A2(_1369_),
    .ZN(_1370_)
  );
  XOR2_X1 _6654_ (
    .A(_1285_),
    .B(_1369_),
    .Z(_1371_)
  );
  AND2_X1 _6655_ (
    .A1(_1284_),
    .A2(_1371_),
    .ZN(_1372_)
  );
  XOR2_X1 _6656_ (
    .A(_1284_),
    .B(_1371_),
    .Z(_1373_)
  );
  AND2_X1 _6657_ (
    .A1(_1255_),
    .A2(_1373_),
    .ZN(_1374_)
  );
  INV_X1 _6658_ (
    .A(_1374_),
    .ZN(_1375_)
  );
  OR2_X1 _6659_ (
    .A1(_1255_),
    .A2(_1373_),
    .ZN(_1376_)
  );
  INV_X1 _6660_ (
    .A(_1376_),
    .ZN(_1377_)
  );
  AND2_X1 _6661_ (
    .A1(_1375_),
    .A2(_1376_),
    .ZN(_1378_)
  );
  OR2_X1 _6662_ (
    .A1(_1374_),
    .A2(_1377_),
    .ZN(_1379_)
  );
  XOR2_X1 _6663_ (
    .A(_1283_),
    .B(_1379_),
    .Z(_1380_)
  );
  XOR2_X1 _6664_ (
    .A(_1283_),
    .B(_1378_),
    .Z(_1381_)
  );
  OR2_X1 _6665_ (
    .A1(_3045_),
    .A2(_1380_),
    .ZN(_1382_)
  );
  INV_X1 _6666_ (
    .A(_1382_),
    .ZN(_1383_)
  );
  OR2_X1 _6667_ (
    .A1(remainder[52]),
    .A2(_1381_),
    .ZN(_1384_)
  );
  INV_X1 _6668_ (
    .A(_1384_),
    .ZN(_1385_)
  );
  AND2_X1 _6669_ (
    .A1(_1382_),
    .A2(_1384_),
    .ZN(_1386_)
  );
  XOR2_X1 _6670_ (
    .A(_1282_),
    .B(_1386_),
    .Z(_1387_)
  );
  AND2_X1 _6671_ (
    .A1(_4613_),
    .A2(_1387_),
    .ZN(_1388_)
  );
  OR2_X1 _6672_ (
    .A1(_1280_),
    .A2(_1388_),
    .ZN(_1389_)
  );
  OR2_X1 _6673_ (
    .A1(_1279_),
    .A2(_1389_),
    .ZN(_1390_)
  );
  AND2_X1 _6674_ (
    .A1(_3911_),
    .A2(_1390_),
    .ZN(_0065_)
  );
  OR2_X1 _6675_ (
    .A1(remainder[44]),
    .A2(_4393_),
    .ZN(_1391_)
  );
  OR2_X1 _6676_ (
    .A1(_4392_),
    .A2(_4495_),
    .ZN(_1392_)
  );
  AND2_X1 _6677_ (
    .A1(_3678_),
    .A2(_1392_),
    .ZN(_1393_)
  );
  AND2_X1 _6678_ (
    .A1(_1391_),
    .A2(_1393_),
    .ZN(_1394_)
  );
  OR2_X1 _6679_ (
    .A1(_1368_),
    .A2(_1370_),
    .ZN(_1395_)
  );
  OR2_X1 _6680_ (
    .A1(_1362_),
    .A2(_1364_),
    .ZN(_1396_)
  );
  OR2_X1 _6681_ (
    .A1(_1343_),
    .A2(_1366_),
    .ZN(_1397_)
  );
  OR2_X1 _6682_ (
    .A1(_1294_),
    .A2(_1296_),
    .ZN(_1398_)
  );
  AND2_X1 _6683_ (
    .A1(divisor[16]),
    .A2(remainder[4]),
    .ZN(_1399_)
  );
  AND2_X1 _6684_ (
    .A1(divisor[17]),
    .A2(remainder[3]),
    .ZN(_1400_)
  );
  AND2_X1 _6685_ (
    .A1(divisor[18]),
    .A2(remainder[3]),
    .ZN(_1401_)
  );
  AND2_X1 _6686_ (
    .A1(_1293_),
    .A2(_1400_),
    .ZN(_1402_)
  );
  XOR2_X1 _6687_ (
    .A(_1293_),
    .B(_1400_),
    .Z(_1403_)
  );
  AND2_X1 _6688_ (
    .A1(_1399_),
    .A2(_1403_),
    .ZN(_1404_)
  );
  XOR2_X1 _6689_ (
    .A(_1399_),
    .B(_1403_),
    .Z(_1405_)
  );
  AND2_X1 _6690_ (
    .A1(_1398_),
    .A2(_1405_),
    .ZN(_1406_)
  );
  XOR2_X1 _6691_ (
    .A(_1398_),
    .B(_1405_),
    .Z(_1407_)
  );
  AND2_X1 _6692_ (
    .A1(_1298_),
    .A2(_1407_),
    .ZN(_1408_)
  );
  XOR2_X1 _6693_ (
    .A(_1298_),
    .B(_1407_),
    .Z(_1409_)
  );
  AND2_X1 _6694_ (
    .A1(_1300_),
    .A2(_1409_),
    .ZN(_1410_)
  );
  INV_X1 _6695_ (
    .A(_1410_),
    .ZN(_1411_)
  );
  XOR2_X1 _6696_ (
    .A(_1300_),
    .B(_1409_),
    .Z(_1412_)
  );
  OR2_X1 _6697_ (
    .A1(_1311_),
    .A2(_1320_),
    .ZN(_1413_)
  );
  OR2_X1 _6698_ (
    .A1(_1307_),
    .A2(_1309_),
    .ZN(_1414_)
  );
  AND2_X1 _6699_ (
    .A1(divisor[13]),
    .A2(remainder[7]),
    .ZN(_1415_)
  );
  AND2_X1 _6700_ (
    .A1(divisor[14]),
    .A2(remainder[6]),
    .ZN(_1416_)
  );
  AND2_X1 _6701_ (
    .A1(divisor[15]),
    .A2(remainder[6]),
    .ZN(_1417_)
  );
  AND2_X1 _6702_ (
    .A1(_1306_),
    .A2(_1416_),
    .ZN(_1418_)
  );
  XOR2_X1 _6703_ (
    .A(_1306_),
    .B(_1416_),
    .Z(_1419_)
  );
  AND2_X1 _6704_ (
    .A1(_1415_),
    .A2(_1419_),
    .ZN(_1420_)
  );
  XOR2_X1 _6705_ (
    .A(_1415_),
    .B(_1419_),
    .Z(_1421_)
  );
  AND2_X1 _6706_ (
    .A1(_1414_),
    .A2(_1421_),
    .ZN(_1422_)
  );
  XOR2_X1 _6707_ (
    .A(_1414_),
    .B(_1421_),
    .Z(_1423_)
  );
  MUX2_X1 _6708_ (
    .A(_1314_),
    .B(_3318_),
    .S(_1313_),
    .Z(_1424_)
  );
  AND2_X1 _6709_ (
    .A1(divisor[10]),
    .A2(_1424_),
    .ZN(_1425_)
  );
  MUX2_X1 _6710_ (
    .A(_1223_),
    .B(_3307_),
    .S(_1424_),
    .Z(_1426_)
  );
  INV_X1 _6711_ (
    .A(_1426_),
    .ZN(_1427_)
  );
  AND2_X1 _6712_ (
    .A1(_1423_),
    .A2(_1426_),
    .ZN(_1428_)
  );
  XOR2_X1 _6713_ (
    .A(_1423_),
    .B(_1426_),
    .Z(_1429_)
  );
  AND2_X1 _6714_ (
    .A1(_1413_),
    .A2(_1429_),
    .ZN(_1430_)
  );
  XOR2_X1 _6715_ (
    .A(_1413_),
    .B(_1429_),
    .Z(_1431_)
  );
  OR2_X1 _6716_ (
    .A1(_1316_),
    .A2(_1318_),
    .ZN(_1432_)
  );
  AND2_X1 _6717_ (
    .A1(_1128_),
    .A2(_1432_),
    .ZN(_1433_)
  );
  XOR2_X1 _6718_ (
    .A(_1128_),
    .B(_1432_),
    .Z(_1434_)
  );
  AND2_X1 _6719_ (
    .A1(_1234_),
    .A2(_1434_),
    .ZN(_1435_)
  );
  XOR2_X1 _6720_ (
    .A(_1234_),
    .B(_1434_),
    .Z(_1436_)
  );
  AND2_X1 _6721_ (
    .A1(_1431_),
    .A2(_1436_),
    .ZN(_1437_)
  );
  XOR2_X1 _6722_ (
    .A(_1431_),
    .B(_1436_),
    .Z(_1438_)
  );
  AND2_X1 _6723_ (
    .A1(_1412_),
    .A2(_1438_),
    .ZN(_1439_)
  );
  INV_X1 _6724_ (
    .A(_1439_),
    .ZN(_1440_)
  );
  XOR2_X1 _6725_ (
    .A(_1412_),
    .B(_1438_),
    .Z(_1441_)
  );
  AND2_X1 _6726_ (
    .A1(_1331_),
    .A2(_1441_),
    .ZN(_1442_)
  );
  XOR2_X1 _6727_ (
    .A(_1331_),
    .B(_1441_),
    .Z(_1443_)
  );
  AND2_X1 _6728_ (
    .A1(divisor[20]),
    .A2(remainder[0]),
    .ZN(_1444_)
  );
  AND2_X1 _6729_ (
    .A1(divisor[19]),
    .A2(remainder[1]),
    .ZN(_1445_)
  );
  AND2_X1 _6730_ (
    .A1(divisor[20]),
    .A2(remainder[1]),
    .ZN(_1446_)
  );
  AND2_X1 _6731_ (
    .A1(_1335_),
    .A2(_1446_),
    .ZN(_1447_)
  );
  XOR2_X1 _6732_ (
    .A(_1444_),
    .B(_1445_),
    .Z(_1448_)
  );
  INV_X1 _6733_ (
    .A(_1448_),
    .ZN(_1449_)
  );
  XOR2_X1 _6734_ (
    .A(_1336_),
    .B(_1449_),
    .Z(_1450_)
  );
  AND2_X1 _6735_ (
    .A1(_1443_),
    .A2(_1450_),
    .ZN(_1451_)
  );
  XOR2_X1 _6736_ (
    .A(_1443_),
    .B(_1450_),
    .Z(_1452_)
  );
  AND2_X1 _6737_ (
    .A1(_1340_),
    .A2(_1452_),
    .ZN(_1453_)
  );
  XOR2_X1 _6738_ (
    .A(_1340_),
    .B(_1452_),
    .Z(_1454_)
  );
  OR2_X1 _6739_ (
    .A1(_1358_),
    .A2(_1360_),
    .ZN(_1455_)
  );
  OR2_X1 _6740_ (
    .A1(_1354_),
    .A2(_1356_),
    .ZN(_1456_)
  );
  OR2_X1 _6741_ (
    .A1(_1350_),
    .A2(_1352_),
    .ZN(_1457_)
  );
  OR2_X1 _6742_ (
    .A1(_1322_),
    .A2(_1329_),
    .ZN(_1458_)
  );
  OR2_X1 _6743_ (
    .A1(_1325_),
    .A2(_1327_),
    .ZN(_1459_)
  );
  AND2_X1 _6744_ (
    .A1(_0894_),
    .A2(_1459_),
    .ZN(_1460_)
  );
  XOR2_X1 _6745_ (
    .A(_0894_),
    .B(_1459_),
    .Z(_1461_)
  );
  AND2_X1 _6746_ (
    .A1(_0985_),
    .A2(_1461_),
    .ZN(_1462_)
  );
  XOR2_X1 _6747_ (
    .A(_0985_),
    .B(_1461_),
    .Z(_1463_)
  );
  AND2_X1 _6748_ (
    .A1(_1458_),
    .A2(_1463_),
    .ZN(_1464_)
  );
  XOR2_X1 _6749_ (
    .A(_1458_),
    .B(_1463_),
    .Z(_1465_)
  );
  AND2_X1 _6750_ (
    .A1(_1457_),
    .A2(_1465_),
    .ZN(_1466_)
  );
  XOR2_X1 _6751_ (
    .A(_1457_),
    .B(_1465_),
    .Z(_1467_)
  );
  AND2_X1 _6752_ (
    .A1(_1456_),
    .A2(_1467_),
    .ZN(_1468_)
  );
  XOR2_X1 _6753_ (
    .A(_1456_),
    .B(_1467_),
    .Z(_1469_)
  );
  AND2_X1 _6754_ (
    .A1(_0512_),
    .A2(_1469_),
    .ZN(_1470_)
  );
  XOR2_X1 _6755_ (
    .A(_0512_),
    .B(_1469_),
    .Z(_1471_)
  );
  AND2_X1 _6756_ (
    .A1(_1333_),
    .A2(_1471_),
    .ZN(_1472_)
  );
  XOR2_X1 _6757_ (
    .A(_1333_),
    .B(_1471_),
    .Z(_1473_)
  );
  AND2_X1 _6758_ (
    .A1(_1455_),
    .A2(_1473_),
    .ZN(_1474_)
  );
  XOR2_X1 _6759_ (
    .A(_1455_),
    .B(_1473_),
    .Z(_1475_)
  );
  AND2_X1 _6760_ (
    .A1(_1454_),
    .A2(_1475_),
    .ZN(_1476_)
  );
  XOR2_X1 _6761_ (
    .A(_1454_),
    .B(_1475_),
    .Z(_1477_)
  );
  AND2_X1 _6762_ (
    .A1(_1397_),
    .A2(_1477_),
    .ZN(_1478_)
  );
  XOR2_X1 _6763_ (
    .A(_1397_),
    .B(_1477_),
    .Z(_1479_)
  );
  AND2_X1 _6764_ (
    .A1(_1396_),
    .A2(_1479_),
    .ZN(_1480_)
  );
  XOR2_X1 _6765_ (
    .A(_1396_),
    .B(_1479_),
    .Z(_1481_)
  );
  AND2_X1 _6766_ (
    .A1(_1395_),
    .A2(_1481_),
    .ZN(_1482_)
  );
  XOR2_X1 _6767_ (
    .A(_1395_),
    .B(_1481_),
    .Z(_1483_)
  );
  AND2_X1 _6768_ (
    .A1(_1372_),
    .A2(_1483_),
    .ZN(_1484_)
  );
  XOR2_X1 _6769_ (
    .A(_1372_),
    .B(_1483_),
    .Z(_1485_)
  );
  OR2_X1 _6770_ (
    .A1(_1257_),
    .A2(_1374_),
    .ZN(_1486_)
  );
  OR2_X1 _6771_ (
    .A1(_1259_),
    .A2(_1486_),
    .ZN(_1487_)
  );
  AND2_X1 _6772_ (
    .A1(_1376_),
    .A2(_1487_),
    .ZN(_1488_)
  );
  AND2_X1 _6773_ (
    .A1(_1485_),
    .A2(_1488_),
    .ZN(_1489_)
  );
  XOR2_X1 _6774_ (
    .A(_1485_),
    .B(_1488_),
    .Z(_1490_)
  );
  AND2_X1 _6775_ (
    .A1(remainder[53]),
    .A2(_1490_),
    .ZN(_1491_)
  );
  INV_X1 _6776_ (
    .A(_1491_),
    .ZN(_1492_)
  );
  XOR2_X1 _6777_ (
    .A(remainder[53]),
    .B(_1490_),
    .Z(_1493_)
  );
  INV_X1 _6778_ (
    .A(_1493_),
    .ZN(_1494_)
  );
  AND2_X1 _6779_ (
    .A1(_1282_),
    .A2(_1384_),
    .ZN(_1495_)
  );
  OR2_X1 _6780_ (
    .A1(_1281_),
    .A2(_1385_),
    .ZN(_1496_)
  );
  AND2_X1 _6781_ (
    .A1(_1382_),
    .A2(_1496_),
    .ZN(_1497_)
  );
  OR2_X1 _6782_ (
    .A1(_1383_),
    .A2(_1495_),
    .ZN(_1498_)
  );
  AND2_X1 _6783_ (
    .A1(_1493_),
    .A2(_1498_),
    .ZN(_1499_)
  );
  OR2_X1 _6784_ (
    .A1(_1494_),
    .A2(_1497_),
    .ZN(_1500_)
  );
  OR2_X1 _6785_ (
    .A1(_1493_),
    .A2(_1498_),
    .ZN(_1501_)
  );
  AND2_X1 _6786_ (
    .A1(_4613_),
    .A2(_1501_),
    .ZN(_1502_)
  );
  AND2_X1 _6787_ (
    .A1(_1500_),
    .A2(_1502_),
    .ZN(_1503_)
  );
  AND2_X1 _6788_ (
    .A1(remainder[45]),
    .A2(_4610_),
    .ZN(_1504_)
  );
  OR2_X1 _6789_ (
    .A1(_1503_),
    .A2(_1504_),
    .ZN(_1505_)
  );
  OR2_X1 _6790_ (
    .A1(_1394_),
    .A2(_1505_),
    .ZN(_1506_)
  );
  AND2_X1 _6791_ (
    .A1(_3911_),
    .A2(_1506_),
    .ZN(_0066_)
  );
  OR2_X1 _6792_ (
    .A1(remainder[45]),
    .A2(_4393_),
    .ZN(_1507_)
  );
  OR2_X1 _6793_ (
    .A1(_4392_),
    .A2(_4501_),
    .ZN(_1508_)
  );
  AND2_X1 _6794_ (
    .A1(_3678_),
    .A2(_1508_),
    .ZN(_1509_)
  );
  AND2_X1 _6795_ (
    .A1(_1507_),
    .A2(_1509_),
    .ZN(_1510_)
  );
  AND2_X1 _6796_ (
    .A1(remainder[46]),
    .A2(_4610_),
    .ZN(_1511_)
  );
  AND2_X1 _6797_ (
    .A1(_1492_),
    .A2(_1500_),
    .ZN(_1512_)
  );
  OR2_X1 _6798_ (
    .A1(_1491_),
    .A2(_1499_),
    .ZN(_1513_)
  );
  OR2_X1 _6799_ (
    .A1(_1484_),
    .A2(_1489_),
    .ZN(_1514_)
  );
  OR2_X1 _6800_ (
    .A1(_1478_),
    .A2(_1480_),
    .ZN(_1515_)
  );
  OR2_X1 _6801_ (
    .A1(_1472_),
    .A2(_1474_),
    .ZN(_1516_)
  );
  OR2_X1 _6802_ (
    .A1(_1453_),
    .A2(_1476_),
    .ZN(_1517_)
  );
  AND2_X1 _6803_ (
    .A1(_0541_),
    .A2(_1449_),
    .ZN(_1518_)
  );
  AND2_X1 _6804_ (
    .A1(_1335_),
    .A2(_1518_),
    .ZN(_1519_)
  );
  OR2_X1 _6805_ (
    .A1(_1451_),
    .A2(_1519_),
    .ZN(_1520_)
  );
  AND2_X1 _6806_ (
    .A1(_1411_),
    .A2(_1440_),
    .ZN(_1521_)
  );
  OR2_X1 _6807_ (
    .A1(_1422_),
    .A2(_1428_),
    .ZN(_1522_)
  );
  OR2_X1 _6808_ (
    .A1(_1418_),
    .A2(_1420_),
    .ZN(_1523_)
  );
  AND2_X1 _6809_ (
    .A1(remainder[32]),
    .A2(divisor[13]),
    .ZN(_1524_)
  );
  INV_X1 _6810_ (
    .A(_1524_),
    .ZN(_1525_)
  );
  AND2_X1 _6811_ (
    .A1(divisor[14]),
    .A2(remainder[7]),
    .ZN(_1526_)
  );
  AND2_X1 _6812_ (
    .A1(divisor[15]),
    .A2(remainder[7]),
    .ZN(_1527_)
  );
  AND2_X1 _6813_ (
    .A1(_1416_),
    .A2(_1527_),
    .ZN(_1528_)
  );
  XOR2_X1 _6814_ (
    .A(_1417_),
    .B(_1526_),
    .Z(_1529_)
  );
  AND2_X1 _6815_ (
    .A1(_1524_),
    .A2(_1529_),
    .ZN(_1530_)
  );
  XOR2_X1 _6816_ (
    .A(_1524_),
    .B(_1529_),
    .Z(_1531_)
  );
  AND2_X1 _6817_ (
    .A1(_1523_),
    .A2(_1531_),
    .ZN(_1532_)
  );
  XOR2_X1 _6818_ (
    .A(_1523_),
    .B(_1531_),
    .Z(_1533_)
  );
  AND2_X1 _6819_ (
    .A1(_1426_),
    .A2(_1533_),
    .ZN(_1534_)
  );
  XOR2_X1 _6820_ (
    .A(_1426_),
    .B(_1533_),
    .Z(_1535_)
  );
  AND2_X1 _6821_ (
    .A1(_1522_),
    .A2(_1535_),
    .ZN(_1536_)
  );
  XOR2_X1 _6822_ (
    .A(_1522_),
    .B(_1535_),
    .Z(_1537_)
  );
  OR2_X1 _6823_ (
    .A1(_1315_),
    .A2(_1425_),
    .ZN(_1538_)
  );
  AND2_X1 _6824_ (
    .A1(_1128_),
    .A2(_1538_),
    .ZN(_1539_)
  );
  XOR2_X1 _6825_ (
    .A(_1128_),
    .B(_1538_),
    .Z(_1540_)
  );
  AND2_X1 _6826_ (
    .A1(_1234_),
    .A2(_1540_),
    .ZN(_1541_)
  );
  XOR2_X1 _6827_ (
    .A(_1234_),
    .B(_1540_),
    .Z(_1542_)
  );
  XOR2_X1 _6828_ (
    .A(_1235_),
    .B(_1540_),
    .Z(_1543_)
  );
  AND2_X1 _6829_ (
    .A1(_1537_),
    .A2(_1542_),
    .ZN(_1544_)
  );
  XOR2_X1 _6830_ (
    .A(_1537_),
    .B(_1542_),
    .Z(_1545_)
  );
  XOR2_X1 _6831_ (
    .A(_1537_),
    .B(_1543_),
    .Z(_1546_)
  );
  OR2_X1 _6832_ (
    .A1(_1402_),
    .A2(_1404_),
    .ZN(_1547_)
  );
  AND2_X1 _6833_ (
    .A1(divisor[16]),
    .A2(remainder[5]),
    .ZN(_1548_)
  );
  AND2_X1 _6834_ (
    .A1(divisor[17]),
    .A2(remainder[4]),
    .ZN(_1549_)
  );
  AND2_X1 _6835_ (
    .A1(divisor[18]),
    .A2(remainder[4]),
    .ZN(_1550_)
  );
  AND2_X1 _6836_ (
    .A1(_1401_),
    .A2(_1549_),
    .ZN(_1551_)
  );
  XOR2_X1 _6837_ (
    .A(_1401_),
    .B(_1549_),
    .Z(_1552_)
  );
  AND2_X1 _6838_ (
    .A1(_1548_),
    .A2(_1552_),
    .ZN(_1553_)
  );
  XOR2_X1 _6839_ (
    .A(_1548_),
    .B(_1552_),
    .Z(_1554_)
  );
  AND2_X1 _6840_ (
    .A1(_1447_),
    .A2(_1554_),
    .ZN(_1555_)
  );
  XOR2_X1 _6841_ (
    .A(_1447_),
    .B(_1554_),
    .Z(_1556_)
  );
  AND2_X1 _6842_ (
    .A1(_1547_),
    .A2(_1556_),
    .ZN(_1557_)
  );
  XOR2_X1 _6843_ (
    .A(_1547_),
    .B(_1556_),
    .Z(_1558_)
  );
  OR2_X1 _6844_ (
    .A1(_1406_),
    .A2(_1408_),
    .ZN(_1559_)
  );
  XOR2_X1 _6845_ (
    .A(_1558_),
    .B(_1559_),
    .Z(_1560_)
  );
  AND2_X1 _6846_ (
    .A1(_1545_),
    .A2(_1560_),
    .ZN(_1561_)
  );
  XOR2_X1 _6847_ (
    .A(_1546_),
    .B(_1560_),
    .Z(_1562_)
  );
  OR2_X1 _6848_ (
    .A1(_1521_),
    .A2(_1562_),
    .ZN(_1563_)
  );
  INV_X1 _6849_ (
    .A(_1563_),
    .ZN(_1564_)
  );
  XOR2_X1 _6850_ (
    .A(_1521_),
    .B(_1562_),
    .Z(_1565_)
  );
  AND2_X1 _6851_ (
    .A1(divisor[19]),
    .A2(remainder[2]),
    .ZN(_1566_)
  );
  AND2_X1 _6852_ (
    .A1(divisor[21]),
    .A2(remainder[0]),
    .ZN(_1567_)
  );
  AND2_X1 _6853_ (
    .A1(divisor[21]),
    .A2(remainder[1]),
    .ZN(_1568_)
  );
  AND2_X1 _6854_ (
    .A1(_1444_),
    .A2(_1568_),
    .ZN(_1569_)
  );
  XOR2_X1 _6855_ (
    .A(_1446_),
    .B(_1567_),
    .Z(_1570_)
  );
  AND2_X1 _6856_ (
    .A1(_1566_),
    .A2(_1570_),
    .ZN(_1571_)
  );
  XOR2_X1 _6857_ (
    .A(_1566_),
    .B(_1570_),
    .Z(_1572_)
  );
  INV_X1 _6858_ (
    .A(_1572_),
    .ZN(_1573_)
  );
  XOR2_X1 _6859_ (
    .A(_1518_),
    .B(_1573_),
    .Z(_1574_)
  );
  INV_X1 _6860_ (
    .A(_1574_),
    .ZN(_1575_)
  );
  AND2_X1 _6861_ (
    .A1(_1565_),
    .A2(_1575_),
    .ZN(_1576_)
  );
  XOR2_X1 _6862_ (
    .A(_1565_),
    .B(_1575_),
    .Z(_1577_)
  );
  AND2_X1 _6863_ (
    .A1(_1520_),
    .A2(_1577_),
    .ZN(_1578_)
  );
  XOR2_X1 _6864_ (
    .A(_1520_),
    .B(_1577_),
    .Z(_1579_)
  );
  OR2_X1 _6865_ (
    .A1(_1468_),
    .A2(_1470_),
    .ZN(_1580_)
  );
  OR2_X1 _6866_ (
    .A1(_1464_),
    .A2(_1466_),
    .ZN(_1581_)
  );
  OR2_X1 _6867_ (
    .A1(_1460_),
    .A2(_1462_),
    .ZN(_1582_)
  );
  OR2_X1 _6868_ (
    .A1(_1430_),
    .A2(_1437_),
    .ZN(_1583_)
  );
  OR2_X1 _6869_ (
    .A1(_1433_),
    .A2(_1435_),
    .ZN(_1584_)
  );
  AND2_X1 _6870_ (
    .A1(_0894_),
    .A2(_1584_),
    .ZN(_1585_)
  );
  XOR2_X1 _6871_ (
    .A(_0894_),
    .B(_1584_),
    .Z(_1586_)
  );
  AND2_X1 _6872_ (
    .A1(_0985_),
    .A2(_1586_),
    .ZN(_1587_)
  );
  XOR2_X1 _6873_ (
    .A(_0985_),
    .B(_1586_),
    .Z(_1588_)
  );
  AND2_X1 _6874_ (
    .A1(_1583_),
    .A2(_1588_),
    .ZN(_1589_)
  );
  XOR2_X1 _6875_ (
    .A(_1583_),
    .B(_1588_),
    .Z(_1590_)
  );
  AND2_X1 _6876_ (
    .A1(_1582_),
    .A2(_1590_),
    .ZN(_1591_)
  );
  XOR2_X1 _6877_ (
    .A(_1582_),
    .B(_1590_),
    .Z(_1592_)
  );
  AND2_X1 _6878_ (
    .A1(_1581_),
    .A2(_1592_),
    .ZN(_1593_)
  );
  XOR2_X1 _6879_ (
    .A(_1581_),
    .B(_1592_),
    .Z(_1594_)
  );
  AND2_X1 _6880_ (
    .A1(_0512_),
    .A2(_1594_),
    .ZN(_1595_)
  );
  XOR2_X1 _6881_ (
    .A(_0512_),
    .B(_1594_),
    .Z(_1596_)
  );
  AND2_X1 _6882_ (
    .A1(_1442_),
    .A2(_1596_),
    .ZN(_1597_)
  );
  XOR2_X1 _6883_ (
    .A(_1442_),
    .B(_1596_),
    .Z(_1598_)
  );
  AND2_X1 _6884_ (
    .A1(_1580_),
    .A2(_1598_),
    .ZN(_1599_)
  );
  XOR2_X1 _6885_ (
    .A(_1580_),
    .B(_1598_),
    .Z(_1600_)
  );
  AND2_X1 _6886_ (
    .A1(_1579_),
    .A2(_1600_),
    .ZN(_1601_)
  );
  XOR2_X1 _6887_ (
    .A(_1579_),
    .B(_1600_),
    .Z(_1602_)
  );
  AND2_X1 _6888_ (
    .A1(_1517_),
    .A2(_1602_),
    .ZN(_1603_)
  );
  XOR2_X1 _6889_ (
    .A(_1517_),
    .B(_1602_),
    .Z(_1604_)
  );
  AND2_X1 _6890_ (
    .A1(_1516_),
    .A2(_1604_),
    .ZN(_1605_)
  );
  XOR2_X1 _6891_ (
    .A(_1516_),
    .B(_1604_),
    .Z(_1606_)
  );
  AND2_X1 _6892_ (
    .A1(_1515_),
    .A2(_1606_),
    .ZN(_1607_)
  );
  XOR2_X1 _6893_ (
    .A(_1515_),
    .B(_1606_),
    .Z(_1608_)
  );
  AND2_X1 _6894_ (
    .A1(_1482_),
    .A2(_1608_),
    .ZN(_1609_)
  );
  INV_X1 _6895_ (
    .A(_1609_),
    .ZN(_1610_)
  );
  OR2_X1 _6896_ (
    .A1(_1482_),
    .A2(_1608_),
    .ZN(_1611_)
  );
  INV_X1 _6897_ (
    .A(_1611_),
    .ZN(_1612_)
  );
  AND2_X1 _6898_ (
    .A1(_1610_),
    .A2(_1611_),
    .ZN(_1613_)
  );
  OR2_X1 _6899_ (
    .A1(_1609_),
    .A2(_1612_),
    .ZN(_1614_)
  );
  AND2_X1 _6900_ (
    .A1(_1514_),
    .A2(_1613_),
    .ZN(_1615_)
  );
  XOR2_X1 _6901_ (
    .A(_1514_),
    .B(_1613_),
    .Z(_1616_)
  );
  XOR2_X1 _6902_ (
    .A(_1514_),
    .B(_1614_),
    .Z(_1617_)
  );
  OR2_X1 _6903_ (
    .A1(_3034_),
    .A2(_1617_),
    .ZN(_1618_)
  );
  INV_X1 _6904_ (
    .A(_1618_),
    .ZN(_1619_)
  );
  OR2_X1 _6905_ (
    .A1(remainder[54]),
    .A2(_1616_),
    .ZN(_1620_)
  );
  INV_X1 _6906_ (
    .A(_1620_),
    .ZN(_1621_)
  );
  AND2_X1 _6907_ (
    .A1(_1618_),
    .A2(_1620_),
    .ZN(_1622_)
  );
  XOR2_X1 _6908_ (
    .A(_1513_),
    .B(_1622_),
    .Z(_1623_)
  );
  AND2_X1 _6909_ (
    .A1(_4613_),
    .A2(_1623_),
    .ZN(_1624_)
  );
  OR2_X1 _6910_ (
    .A1(_1511_),
    .A2(_1624_),
    .ZN(_1625_)
  );
  OR2_X1 _6911_ (
    .A1(_1510_),
    .A2(_1625_),
    .ZN(_1626_)
  );
  AND2_X1 _6912_ (
    .A1(_3911_),
    .A2(_1626_),
    .ZN(_0067_)
  );
  OR2_X1 _6913_ (
    .A1(_4392_),
    .A2(_4506_),
    .ZN(_1627_)
  );
  OR2_X1 _6914_ (
    .A1(remainder[46]),
    .A2(_4393_),
    .ZN(_1628_)
  );
  AND2_X1 _6915_ (
    .A1(_3678_),
    .A2(_1627_),
    .ZN(_1629_)
  );
  AND2_X1 _6916_ (
    .A1(_1628_),
    .A2(_1629_),
    .ZN(_1630_)
  );
  AND2_X1 _6917_ (
    .A1(remainder[47]),
    .A2(_4610_),
    .ZN(_1631_)
  );
  OR2_X1 _6918_ (
    .A1(_1603_),
    .A2(_1605_),
    .ZN(_1632_)
  );
  OR2_X1 _6919_ (
    .A1(_1597_),
    .A2(_1599_),
    .ZN(_1633_)
  );
  OR2_X1 _6920_ (
    .A1(_1578_),
    .A2(_1601_),
    .ZN(_1634_)
  );
  AND2_X1 _6921_ (
    .A1(_0541_),
    .A2(_1573_),
    .ZN(_1635_)
  );
  AND2_X1 _6922_ (
    .A1(_1448_),
    .A2(_1635_),
    .ZN(_1636_)
  );
  OR2_X1 _6923_ (
    .A1(_1576_),
    .A2(_1636_),
    .ZN(_1637_)
  );
  AND2_X1 _6924_ (
    .A1(_1408_),
    .A2(_1558_),
    .ZN(_1638_)
  );
  OR2_X1 _6925_ (
    .A1(_1561_),
    .A2(_1638_),
    .ZN(_1639_)
  );
  AND2_X1 _6926_ (
    .A1(_1406_),
    .A2(_1558_),
    .ZN(_1640_)
  );
  OR2_X1 _6927_ (
    .A1(_1555_),
    .A2(_1557_),
    .ZN(_1641_)
  );
  OR2_X1 _6928_ (
    .A1(_1551_),
    .A2(_1553_),
    .ZN(_1642_)
  );
  OR2_X1 _6929_ (
    .A1(_1569_),
    .A2(_1571_),
    .ZN(_1643_)
  );
  AND2_X1 _6930_ (
    .A1(divisor[16]),
    .A2(remainder[6]),
    .ZN(_1644_)
  );
  AND2_X1 _6931_ (
    .A1(divisor[17]),
    .A2(remainder[5]),
    .ZN(_1645_)
  );
  AND2_X1 _6932_ (
    .A1(divisor[18]),
    .A2(remainder[5]),
    .ZN(_1646_)
  );
  AND2_X1 _6933_ (
    .A1(_1550_),
    .A2(_1645_),
    .ZN(_1647_)
  );
  XOR2_X1 _6934_ (
    .A(_1550_),
    .B(_1645_),
    .Z(_1648_)
  );
  AND2_X1 _6935_ (
    .A1(_1644_),
    .A2(_1648_),
    .ZN(_1649_)
  );
  XOR2_X1 _6936_ (
    .A(_1644_),
    .B(_1648_),
    .Z(_1650_)
  );
  AND2_X1 _6937_ (
    .A1(_1643_),
    .A2(_1650_),
    .ZN(_1651_)
  );
  XOR2_X1 _6938_ (
    .A(_1643_),
    .B(_1650_),
    .Z(_1652_)
  );
  AND2_X1 _6939_ (
    .A1(_1642_),
    .A2(_1652_),
    .ZN(_1653_)
  );
  XOR2_X1 _6940_ (
    .A(_1642_),
    .B(_1652_),
    .Z(_1654_)
  );
  AND2_X1 _6941_ (
    .A1(_1641_),
    .A2(_1654_),
    .ZN(_1655_)
  );
  XOR2_X1 _6942_ (
    .A(_1641_),
    .B(_1654_),
    .Z(_1656_)
  );
  AND2_X1 _6943_ (
    .A1(_1640_),
    .A2(_1656_),
    .ZN(_1657_)
  );
  XOR2_X1 _6944_ (
    .A(_1640_),
    .B(_1656_),
    .Z(_1658_)
  );
  OR2_X1 _6945_ (
    .A1(_1532_),
    .A2(_1534_),
    .ZN(_1659_)
  );
  OR2_X1 _6946_ (
    .A1(_1528_),
    .A2(_1530_),
    .ZN(_1660_)
  );
  AND2_X1 _6947_ (
    .A1(remainder[32]),
    .A2(divisor[15]),
    .ZN(_1661_)
  );
  AND2_X1 _6948_ (
    .A1(remainder[32]),
    .A2(divisor[14]),
    .ZN(_1662_)
  );
  AND2_X1 _6949_ (
    .A1(_1527_),
    .A2(_1662_),
    .ZN(_1663_)
  );
  XOR2_X1 _6950_ (
    .A(_1527_),
    .B(_1662_),
    .Z(_1664_)
  );
  AND2_X1 _6951_ (
    .A1(_1524_),
    .A2(_1664_),
    .ZN(_1665_)
  );
  XOR2_X1 _6952_ (
    .A(_1524_),
    .B(_1664_),
    .Z(_1666_)
  );
  AND2_X1 _6953_ (
    .A1(_1660_),
    .A2(_1666_),
    .ZN(_1667_)
  );
  XOR2_X1 _6954_ (
    .A(_1660_),
    .B(_1666_),
    .Z(_1668_)
  );
  AND2_X1 _6955_ (
    .A1(_1426_),
    .A2(_1668_),
    .ZN(_1669_)
  );
  XOR2_X1 _6956_ (
    .A(_1426_),
    .B(_1668_),
    .Z(_1670_)
  );
  AND2_X1 _6957_ (
    .A1(_1659_),
    .A2(_1670_),
    .ZN(_1671_)
  );
  XOR2_X1 _6958_ (
    .A(_1659_),
    .B(_1670_),
    .Z(_1672_)
  );
  AND2_X1 _6959_ (
    .A1(_1542_),
    .A2(_1672_),
    .ZN(_1673_)
  );
  XOR2_X1 _6960_ (
    .A(_1542_),
    .B(_1672_),
    .Z(_1674_)
  );
  AND2_X1 _6961_ (
    .A1(_1658_),
    .A2(_1674_),
    .ZN(_1675_)
  );
  XOR2_X1 _6962_ (
    .A(_1658_),
    .B(_1674_),
    .Z(_1676_)
  );
  AND2_X1 _6963_ (
    .A1(_1639_),
    .A2(_1676_),
    .ZN(_1677_)
  );
  XOR2_X1 _6964_ (
    .A(_1639_),
    .B(_1676_),
    .Z(_1678_)
  );
  AND2_X1 _6965_ (
    .A1(divisor[22]),
    .A2(remainder[0]),
    .ZN(_1679_)
  );
  AND2_X1 _6966_ (
    .A1(divisor[19]),
    .A2(remainder[3]),
    .ZN(_1680_)
  );
  AND2_X1 _6967_ (
    .A1(divisor[20]),
    .A2(remainder[2]),
    .ZN(_1681_)
  );
  AND2_X1 _6968_ (
    .A1(divisor[21]),
    .A2(remainder[2]),
    .ZN(_1682_)
  );
  AND2_X1 _6969_ (
    .A1(_1446_),
    .A2(_1682_),
    .ZN(_1683_)
  );
  XOR2_X1 _6970_ (
    .A(_1568_),
    .B(_1681_),
    .Z(_1684_)
  );
  AND2_X1 _6971_ (
    .A1(_1680_),
    .A2(_1684_),
    .ZN(_1685_)
  );
  XOR2_X1 _6972_ (
    .A(_1680_),
    .B(_1684_),
    .Z(_1686_)
  );
  AND2_X1 _6973_ (
    .A1(_1679_),
    .A2(_1686_),
    .ZN(_1687_)
  );
  XOR2_X1 _6974_ (
    .A(_1679_),
    .B(_1686_),
    .Z(_1688_)
  );
  INV_X1 _6975_ (
    .A(_1688_),
    .ZN(_1689_)
  );
  XOR2_X1 _6976_ (
    .A(_1635_),
    .B(_1688_),
    .Z(_1690_)
  );
  AND2_X1 _6977_ (
    .A1(_1678_),
    .A2(_1690_),
    .ZN(_1691_)
  );
  XOR2_X1 _6978_ (
    .A(_1678_),
    .B(_1690_),
    .Z(_1692_)
  );
  AND2_X1 _6979_ (
    .A1(_1637_),
    .A2(_1692_),
    .ZN(_1693_)
  );
  XOR2_X1 _6980_ (
    .A(_1637_),
    .B(_1692_),
    .Z(_1694_)
  );
  OR2_X1 _6981_ (
    .A1(_1593_),
    .A2(_1595_),
    .ZN(_1695_)
  );
  OR2_X1 _6982_ (
    .A1(_1589_),
    .A2(_1591_),
    .ZN(_1696_)
  );
  OR2_X1 _6983_ (
    .A1(_1585_),
    .A2(_1587_),
    .ZN(_1697_)
  );
  OR2_X1 _6984_ (
    .A1(_1536_),
    .A2(_1544_),
    .ZN(_1698_)
  );
  OR2_X1 _6985_ (
    .A1(_1539_),
    .A2(_1541_),
    .ZN(_1699_)
  );
  AND2_X1 _6986_ (
    .A1(_0894_),
    .A2(_1699_),
    .ZN(_1700_)
  );
  XOR2_X1 _6987_ (
    .A(_0894_),
    .B(_1699_),
    .Z(_1701_)
  );
  AND2_X1 _6988_ (
    .A1(_0985_),
    .A2(_1701_),
    .ZN(_1702_)
  );
  XOR2_X1 _6989_ (
    .A(_0985_),
    .B(_1701_),
    .Z(_1703_)
  );
  INV_X1 _6990_ (
    .A(_1703_),
    .ZN(_1704_)
  );
  AND2_X1 _6991_ (
    .A1(_1698_),
    .A2(_1703_),
    .ZN(_1705_)
  );
  XOR2_X1 _6992_ (
    .A(_1698_),
    .B(_1703_),
    .Z(_1706_)
  );
  AND2_X1 _6993_ (
    .A1(_1697_),
    .A2(_1706_),
    .ZN(_1707_)
  );
  XOR2_X1 _6994_ (
    .A(_1697_),
    .B(_1706_),
    .Z(_1708_)
  );
  AND2_X1 _6995_ (
    .A1(_1696_),
    .A2(_1708_),
    .ZN(_1709_)
  );
  XOR2_X1 _6996_ (
    .A(_1696_),
    .B(_1708_),
    .Z(_1710_)
  );
  AND2_X1 _6997_ (
    .A1(_0512_),
    .A2(_1710_),
    .ZN(_1711_)
  );
  XOR2_X1 _6998_ (
    .A(_0512_),
    .B(_1710_),
    .Z(_1712_)
  );
  AND2_X1 _6999_ (
    .A1(_1564_),
    .A2(_1712_),
    .ZN(_1713_)
  );
  XOR2_X1 _7000_ (
    .A(_1564_),
    .B(_1712_),
    .Z(_1714_)
  );
  AND2_X1 _7001_ (
    .A1(_1695_),
    .A2(_1714_),
    .ZN(_1715_)
  );
  XOR2_X1 _7002_ (
    .A(_1695_),
    .B(_1714_),
    .Z(_1716_)
  );
  AND2_X1 _7003_ (
    .A1(_1694_),
    .A2(_1716_),
    .ZN(_1717_)
  );
  XOR2_X1 _7004_ (
    .A(_1694_),
    .B(_1716_),
    .Z(_1718_)
  );
  AND2_X1 _7005_ (
    .A1(_1634_),
    .A2(_1718_),
    .ZN(_1719_)
  );
  XOR2_X1 _7006_ (
    .A(_1634_),
    .B(_1718_),
    .Z(_1720_)
  );
  AND2_X1 _7007_ (
    .A1(_1633_),
    .A2(_1720_),
    .ZN(_1721_)
  );
  XOR2_X1 _7008_ (
    .A(_1633_),
    .B(_1720_),
    .Z(_1722_)
  );
  AND2_X1 _7009_ (
    .A1(_1632_),
    .A2(_1722_),
    .ZN(_1723_)
  );
  INV_X1 _7010_ (
    .A(_1723_),
    .ZN(_1724_)
  );
  XOR2_X1 _7011_ (
    .A(_1632_),
    .B(_1722_),
    .Z(_1725_)
  );
  AND2_X1 _7012_ (
    .A1(_1607_),
    .A2(_1725_),
    .ZN(_1726_)
  );
  XOR2_X1 _7013_ (
    .A(_1607_),
    .B(_1725_),
    .Z(_1727_)
  );
  INV_X1 _7014_ (
    .A(_1727_),
    .ZN(_1728_)
  );
  OR2_X1 _7015_ (
    .A1(_1609_),
    .A2(_1615_),
    .ZN(_1729_)
  );
  AND2_X1 _7016_ (
    .A1(_1727_),
    .A2(_1729_),
    .ZN(_1730_)
  );
  XOR2_X1 _7017_ (
    .A(_1727_),
    .B(_1729_),
    .Z(_1731_)
  );
  XOR2_X1 _7018_ (
    .A(_1728_),
    .B(_1729_),
    .Z(_1732_)
  );
  AND2_X1 _7019_ (
    .A1(remainder[55]),
    .A2(_1731_),
    .ZN(_1733_)
  );
  OR2_X1 _7020_ (
    .A1(_3023_),
    .A2(_1732_),
    .ZN(_1734_)
  );
  XOR2_X1 _7021_ (
    .A(remainder[55]),
    .B(_1731_),
    .Z(_1735_)
  );
  INV_X1 _7022_ (
    .A(_1735_),
    .ZN(_1736_)
  );
  AND2_X1 _7023_ (
    .A1(_1512_),
    .A2(_1618_),
    .ZN(_1737_)
  );
  OR2_X1 _7024_ (
    .A1(_1513_),
    .A2(_1619_),
    .ZN(_1738_)
  );
  AND2_X1 _7025_ (
    .A1(_1620_),
    .A2(_1738_),
    .ZN(_1739_)
  );
  OR2_X1 _7026_ (
    .A1(_1621_),
    .A2(_1737_),
    .ZN(_1740_)
  );
  OR2_X1 _7027_ (
    .A1(_1735_),
    .A2(_1739_),
    .ZN(_1741_)
  );
  AND2_X1 _7028_ (
    .A1(_1735_),
    .A2(_1739_),
    .ZN(_1742_)
  );
  OR2_X1 _7029_ (
    .A1(_1736_),
    .A2(_1740_),
    .ZN(_1743_)
  );
  AND2_X1 _7030_ (
    .A1(_4613_),
    .A2(_1741_),
    .ZN(_1744_)
  );
  AND2_X1 _7031_ (
    .A1(_1743_),
    .A2(_1744_),
    .ZN(_1745_)
  );
  OR2_X1 _7032_ (
    .A1(_1631_),
    .A2(_1745_),
    .ZN(_1746_)
  );
  OR2_X1 _7033_ (
    .A1(_1630_),
    .A2(_1746_),
    .ZN(_1747_)
  );
  AND2_X1 _7034_ (
    .A1(_3911_),
    .A2(_1747_),
    .ZN(_0068_)
  );
  OR2_X1 _7035_ (
    .A1(remainder[47]),
    .A2(_4393_),
    .ZN(_1748_)
  );
  OR2_X1 _7036_ (
    .A1(_4392_),
    .A2(_4512_),
    .ZN(_1749_)
  );
  AND2_X1 _7037_ (
    .A1(_3678_),
    .A2(_1749_),
    .ZN(_1750_)
  );
  AND2_X1 _7038_ (
    .A1(_1748_),
    .A2(_1750_),
    .ZN(_1751_)
  );
  AND2_X1 _7039_ (
    .A1(remainder[48]),
    .A2(_4610_),
    .ZN(_1752_)
  );
  AND2_X1 _7040_ (
    .A1(_1734_),
    .A2(_1743_),
    .ZN(_1753_)
  );
  OR2_X1 _7041_ (
    .A1(_1733_),
    .A2(_1742_),
    .ZN(_1754_)
  );
  OR2_X1 _7042_ (
    .A1(_1726_),
    .A2(_1730_),
    .ZN(_1755_)
  );
  OR2_X1 _7043_ (
    .A1(_1719_),
    .A2(_1721_),
    .ZN(_1756_)
  );
  INV_X1 _7044_ (
    .A(_1756_),
    .ZN(_1757_)
  );
  OR2_X1 _7045_ (
    .A1(_1713_),
    .A2(_1715_),
    .ZN(_1758_)
  );
  OR2_X1 _7046_ (
    .A1(_1693_),
    .A2(_1717_),
    .ZN(_1759_)
  );
  AND2_X1 _7047_ (
    .A1(_0541_),
    .A2(_1689_),
    .ZN(_1760_)
  );
  AND2_X1 _7048_ (
    .A1(_1572_),
    .A2(_1760_),
    .ZN(_1761_)
  );
  OR2_X1 _7049_ (
    .A1(_1691_),
    .A2(_1761_),
    .ZN(_1762_)
  );
  OR2_X1 _7050_ (
    .A1(_1657_),
    .A2(_1675_),
    .ZN(_1763_)
  );
  OR2_X1 _7051_ (
    .A1(_1667_),
    .A2(_1669_),
    .ZN(_1764_)
  );
  OR2_X1 _7052_ (
    .A1(_1663_),
    .A2(_1665_),
    .ZN(_1765_)
  );
  INV_X1 _7053_ (
    .A(_1765_),
    .ZN(_1766_)
  );
  OR2_X1 _7054_ (
    .A1(_1661_),
    .A2(_1662_),
    .ZN(_1767_)
  );
  MUX2_X1 _7055_ (
    .A(_1662_),
    .B(_3329_),
    .S(_1661_),
    .Z(_1768_)
  );
  MUX2_X1 _7056_ (
    .A(_1525_),
    .B(divisor[13]),
    .S(_1768_),
    .Z(_1769_)
  );
  OR2_X1 _7057_ (
    .A1(_1766_),
    .A2(_1769_),
    .ZN(_1770_)
  );
  AND2_X1 _7058_ (
    .A1(_1766_),
    .A2(_1769_),
    .ZN(_1771_)
  );
  XOR2_X1 _7059_ (
    .A(_1765_),
    .B(_1769_),
    .Z(_1772_)
  );
  AND2_X1 _7060_ (
    .A1(_1426_),
    .A2(_1772_),
    .ZN(_1773_)
  );
  OR2_X1 _7061_ (
    .A1(_1427_),
    .A2(_1771_),
    .ZN(_1774_)
  );
  XOR2_X1 _7062_ (
    .A(_1426_),
    .B(_1772_),
    .Z(_1775_)
  );
  XOR2_X1 _7063_ (
    .A(_1427_),
    .B(_1772_),
    .Z(_1776_)
  );
  AND2_X1 _7064_ (
    .A1(_1764_),
    .A2(_1776_),
    .ZN(_1777_)
  );
  XOR2_X1 _7065_ (
    .A(_1764_),
    .B(_1775_),
    .Z(_1778_)
  );
  INV_X1 _7066_ (
    .A(_1778_),
    .ZN(_1779_)
  );
  AND2_X1 _7067_ (
    .A1(_1542_),
    .A2(_1779_),
    .ZN(_1780_)
  );
  XOR2_X1 _7068_ (
    .A(_1543_),
    .B(_1778_),
    .Z(_1781_)
  );
  OR2_X1 _7069_ (
    .A1(_1651_),
    .A2(_1653_),
    .ZN(_1782_)
  );
  OR2_X1 _7070_ (
    .A1(_1647_),
    .A2(_1649_),
    .ZN(_1783_)
  );
  OR2_X1 _7071_ (
    .A1(_1683_),
    .A2(_1685_),
    .ZN(_1784_)
  );
  AND2_X1 _7072_ (
    .A1(divisor[16]),
    .A2(remainder[7]),
    .ZN(_1785_)
  );
  AND2_X1 _7073_ (
    .A1(divisor[17]),
    .A2(remainder[6]),
    .ZN(_1786_)
  );
  AND2_X1 _7074_ (
    .A1(divisor[18]),
    .A2(remainder[6]),
    .ZN(_1787_)
  );
  AND2_X1 _7075_ (
    .A1(_1646_),
    .A2(_1786_),
    .ZN(_1788_)
  );
  XOR2_X1 _7076_ (
    .A(_1646_),
    .B(_1786_),
    .Z(_1789_)
  );
  AND2_X1 _7077_ (
    .A1(_1785_),
    .A2(_1789_),
    .ZN(_1790_)
  );
  XOR2_X1 _7078_ (
    .A(_1785_),
    .B(_1789_),
    .Z(_1791_)
  );
  AND2_X1 _7079_ (
    .A1(_1784_),
    .A2(_1791_),
    .ZN(_1792_)
  );
  XOR2_X1 _7080_ (
    .A(_1784_),
    .B(_1791_),
    .Z(_1793_)
  );
  AND2_X1 _7081_ (
    .A1(_1783_),
    .A2(_1793_),
    .ZN(_1794_)
  );
  XOR2_X1 _7082_ (
    .A(_1783_),
    .B(_1793_),
    .Z(_1795_)
  );
  AND2_X1 _7083_ (
    .A1(_1687_),
    .A2(_1795_),
    .ZN(_1796_)
  );
  XOR2_X1 _7084_ (
    .A(_1687_),
    .B(_1795_),
    .Z(_1797_)
  );
  AND2_X1 _7085_ (
    .A1(_1782_),
    .A2(_1797_),
    .ZN(_1798_)
  );
  XOR2_X1 _7086_ (
    .A(_1782_),
    .B(_1797_),
    .Z(_1799_)
  );
  AND2_X1 _7087_ (
    .A1(_1655_),
    .A2(_1799_),
    .ZN(_1800_)
  );
  XOR2_X1 _7088_ (
    .A(_1655_),
    .B(_1799_),
    .Z(_1801_)
  );
  AND2_X1 _7089_ (
    .A1(_1781_),
    .A2(_1801_),
    .ZN(_1802_)
  );
  XOR2_X1 _7090_ (
    .A(_1781_),
    .B(_1801_),
    .Z(_1803_)
  );
  AND2_X1 _7091_ (
    .A1(_1763_),
    .A2(_1803_),
    .ZN(_1804_)
  );
  XOR2_X1 _7092_ (
    .A(_1763_),
    .B(_1803_),
    .Z(_1805_)
  );
  AND2_X1 _7093_ (
    .A1(divisor[23]),
    .A2(remainder[0]),
    .ZN(_1806_)
  );
  AND2_X1 _7094_ (
    .A1(divisor[22]),
    .A2(remainder[1]),
    .ZN(_1807_)
  );
  AND2_X1 _7095_ (
    .A1(divisor[23]),
    .A2(remainder[1]),
    .ZN(_1808_)
  );
  AND2_X1 _7096_ (
    .A1(_1679_),
    .A2(_1808_),
    .ZN(_1809_)
  );
  XOR2_X1 _7097_ (
    .A(_1806_),
    .B(_1807_),
    .Z(_1810_)
  );
  AND2_X1 _7098_ (
    .A1(divisor[19]),
    .A2(remainder[4]),
    .ZN(_1811_)
  );
  AND2_X1 _7099_ (
    .A1(divisor[20]),
    .A2(remainder[3]),
    .ZN(_1812_)
  );
  AND2_X1 _7100_ (
    .A1(divisor[21]),
    .A2(remainder[3]),
    .ZN(_1813_)
  );
  AND2_X1 _7101_ (
    .A1(_1682_),
    .A2(_1812_),
    .ZN(_1814_)
  );
  XOR2_X1 _7102_ (
    .A(_1682_),
    .B(_1812_),
    .Z(_1815_)
  );
  AND2_X1 _7103_ (
    .A1(_1811_),
    .A2(_1815_),
    .ZN(_1816_)
  );
  XOR2_X1 _7104_ (
    .A(_1811_),
    .B(_1815_),
    .Z(_1817_)
  );
  AND2_X1 _7105_ (
    .A1(_1810_),
    .A2(_1817_),
    .ZN(_1818_)
  );
  XOR2_X1 _7106_ (
    .A(_1810_),
    .B(_1817_),
    .Z(_1819_)
  );
  INV_X1 _7107_ (
    .A(_1819_),
    .ZN(_1820_)
  );
  XOR2_X1 _7108_ (
    .A(_1760_),
    .B(_1820_),
    .Z(_1821_)
  );
  INV_X1 _7109_ (
    .A(_1821_),
    .ZN(_1822_)
  );
  AND2_X1 _7110_ (
    .A1(_1805_),
    .A2(_1822_),
    .ZN(_1823_)
  );
  XOR2_X1 _7111_ (
    .A(_1805_),
    .B(_1822_),
    .Z(_1824_)
  );
  AND2_X1 _7112_ (
    .A1(_1762_),
    .A2(_1824_),
    .ZN(_1825_)
  );
  XOR2_X1 _7113_ (
    .A(_1762_),
    .B(_1824_),
    .Z(_1826_)
  );
  OR2_X1 _7114_ (
    .A1(_1709_),
    .A2(_1711_),
    .ZN(_1827_)
  );
  OR2_X1 _7115_ (
    .A1(_1705_),
    .A2(_1707_),
    .ZN(_1828_)
  );
  OR2_X1 _7116_ (
    .A1(_1700_),
    .A2(_1702_),
    .ZN(_1829_)
  );
  INV_X1 _7117_ (
    .A(_1829_),
    .ZN(_1830_)
  );
  OR2_X1 _7118_ (
    .A1(_1671_),
    .A2(_1673_),
    .ZN(_1831_)
  );
  AND2_X1 _7119_ (
    .A1(_1703_),
    .A2(_1831_),
    .ZN(_1832_)
  );
  XOR2_X1 _7120_ (
    .A(_1703_),
    .B(_1831_),
    .Z(_1833_)
  );
  AND2_X1 _7121_ (
    .A1(_1829_),
    .A2(_1833_),
    .ZN(_1834_)
  );
  XOR2_X1 _7122_ (
    .A(_1829_),
    .B(_1833_),
    .Z(_1835_)
  );
  AND2_X1 _7123_ (
    .A1(_1828_),
    .A2(_1835_),
    .ZN(_1836_)
  );
  XOR2_X1 _7124_ (
    .A(_1828_),
    .B(_1835_),
    .Z(_1837_)
  );
  AND2_X1 _7125_ (
    .A1(_0512_),
    .A2(_1837_),
    .ZN(_1838_)
  );
  XOR2_X1 _7126_ (
    .A(_0512_),
    .B(_1837_),
    .Z(_1839_)
  );
  AND2_X1 _7127_ (
    .A1(_1677_),
    .A2(_1839_),
    .ZN(_1840_)
  );
  XOR2_X1 _7128_ (
    .A(_1677_),
    .B(_1839_),
    .Z(_1841_)
  );
  AND2_X1 _7129_ (
    .A1(_1827_),
    .A2(_1841_),
    .ZN(_1842_)
  );
  XOR2_X1 _7130_ (
    .A(_1827_),
    .B(_1841_),
    .Z(_1843_)
  );
  AND2_X1 _7131_ (
    .A1(_1826_),
    .A2(_1843_),
    .ZN(_1844_)
  );
  XOR2_X1 _7132_ (
    .A(_1826_),
    .B(_1843_),
    .Z(_1845_)
  );
  AND2_X1 _7133_ (
    .A1(_1759_),
    .A2(_1845_),
    .ZN(_1846_)
  );
  XOR2_X1 _7134_ (
    .A(_1759_),
    .B(_1845_),
    .Z(_1847_)
  );
  AND2_X1 _7135_ (
    .A1(_1758_),
    .A2(_1847_),
    .ZN(_1848_)
  );
  XOR2_X1 _7136_ (
    .A(_1758_),
    .B(_1847_),
    .Z(_1849_)
  );
  AND2_X1 _7137_ (
    .A1(_1756_),
    .A2(_1849_),
    .ZN(_1850_)
  );
  INV_X1 _7138_ (
    .A(_1850_),
    .ZN(_1851_)
  );
  XOR2_X1 _7139_ (
    .A(_1757_),
    .B(_1849_),
    .Z(_1852_)
  );
  OR2_X1 _7140_ (
    .A1(_1724_),
    .A2(_1852_),
    .ZN(_1853_)
  );
  INV_X1 _7141_ (
    .A(_1853_),
    .ZN(_1854_)
  );
  XOR2_X1 _7142_ (
    .A(_1724_),
    .B(_1852_),
    .Z(_1855_)
  );
  AND2_X1 _7143_ (
    .A1(_1755_),
    .A2(_1855_),
    .ZN(_1856_)
  );
  XOR2_X1 _7144_ (
    .A(_1755_),
    .B(_1855_),
    .Z(_1857_)
  );
  AND2_X1 _7145_ (
    .A1(remainder[56]),
    .A2(_1857_),
    .ZN(_1858_)
  );
  INV_X1 _7146_ (
    .A(_1858_),
    .ZN(_1859_)
  );
  XOR2_X1 _7147_ (
    .A(remainder[56]),
    .B(_1857_),
    .Z(_1860_)
  );
  INV_X1 _7148_ (
    .A(_1860_),
    .ZN(_1861_)
  );
  AND2_X1 _7149_ (
    .A1(_1754_),
    .A2(_1860_),
    .ZN(_1862_)
  );
  OR2_X1 _7150_ (
    .A1(_1753_),
    .A2(_1861_),
    .ZN(_1863_)
  );
  OR2_X1 _7151_ (
    .A1(_1754_),
    .A2(_1860_),
    .ZN(_1864_)
  );
  AND2_X1 _7152_ (
    .A1(_4613_),
    .A2(_1864_),
    .ZN(_1865_)
  );
  AND2_X1 _7153_ (
    .A1(_1863_),
    .A2(_1865_),
    .ZN(_1866_)
  );
  OR2_X1 _7154_ (
    .A1(_1752_),
    .A2(_1866_),
    .ZN(_1867_)
  );
  OR2_X1 _7155_ (
    .A1(_1751_),
    .A2(_1867_),
    .ZN(_1868_)
  );
  AND2_X1 _7156_ (
    .A1(_3911_),
    .A2(_1868_),
    .ZN(_0069_)
  );
  OR2_X1 _7157_ (
    .A1(remainder[48]),
    .A2(_4393_),
    .ZN(_1869_)
  );
  OR2_X1 _7158_ (
    .A1(_4392_),
    .A2(_4517_),
    .ZN(_1870_)
  );
  AND2_X1 _7159_ (
    .A1(_3678_),
    .A2(_1870_),
    .ZN(_1871_)
  );
  AND2_X1 _7160_ (
    .A1(_1869_),
    .A2(_1871_),
    .ZN(_1872_)
  );
  AND2_X1 _7161_ (
    .A1(_1859_),
    .A2(_1863_),
    .ZN(_1873_)
  );
  OR2_X1 _7162_ (
    .A1(_1858_),
    .A2(_1862_),
    .ZN(_1874_)
  );
  OR2_X1 _7163_ (
    .A1(_1846_),
    .A2(_1848_),
    .ZN(_1875_)
  );
  OR2_X1 _7164_ (
    .A1(_1840_),
    .A2(_1842_),
    .ZN(_1876_)
  );
  OR2_X1 _7165_ (
    .A1(_1825_),
    .A2(_1844_),
    .ZN(_1877_)
  );
  AND2_X1 _7166_ (
    .A1(_0541_),
    .A2(_1820_),
    .ZN(_1878_)
  );
  AND2_X1 _7167_ (
    .A1(_1688_),
    .A2(_1878_),
    .ZN(_1879_)
  );
  OR2_X1 _7168_ (
    .A1(_1823_),
    .A2(_1879_),
    .ZN(_1880_)
  );
  OR2_X1 _7169_ (
    .A1(_1800_),
    .A2(_1802_),
    .ZN(_1881_)
  );
  OR2_X1 _7170_ (
    .A1(_1796_),
    .A2(_1798_),
    .ZN(_1882_)
  );
  OR2_X1 _7171_ (
    .A1(_1792_),
    .A2(_1794_),
    .ZN(_1883_)
  );
  OR2_X1 _7172_ (
    .A1(_1788_),
    .A2(_1790_),
    .ZN(_1884_)
  );
  OR2_X1 _7173_ (
    .A1(_1814_),
    .A2(_1816_),
    .ZN(_1885_)
  );
  AND2_X1 _7174_ (
    .A1(remainder[32]),
    .A2(divisor[16]),
    .ZN(_1886_)
  );
  AND2_X1 _7175_ (
    .A1(divisor[17]),
    .A2(remainder[7]),
    .ZN(_1887_)
  );
  AND2_X1 _7176_ (
    .A1(divisor[18]),
    .A2(remainder[7]),
    .ZN(_1888_)
  );
  AND2_X1 _7177_ (
    .A1(_1786_),
    .A2(_1888_),
    .ZN(_1889_)
  );
  XOR2_X1 _7178_ (
    .A(_1787_),
    .B(_1887_),
    .Z(_1890_)
  );
  AND2_X1 _7179_ (
    .A1(_1886_),
    .A2(_1890_),
    .ZN(_1891_)
  );
  XOR2_X1 _7180_ (
    .A(_1886_),
    .B(_1890_),
    .Z(_1892_)
  );
  AND2_X1 _7181_ (
    .A1(_1885_),
    .A2(_1892_),
    .ZN(_1893_)
  );
  XOR2_X1 _7182_ (
    .A(_1885_),
    .B(_1892_),
    .Z(_1894_)
  );
  AND2_X1 _7183_ (
    .A1(_1884_),
    .A2(_1894_),
    .ZN(_1895_)
  );
  XOR2_X1 _7184_ (
    .A(_1884_),
    .B(_1894_),
    .Z(_1896_)
  );
  AND2_X1 _7185_ (
    .A1(_1818_),
    .A2(_1896_),
    .ZN(_1897_)
  );
  XOR2_X1 _7186_ (
    .A(_1818_),
    .B(_1896_),
    .Z(_1898_)
  );
  AND2_X1 _7187_ (
    .A1(_1883_),
    .A2(_1898_),
    .ZN(_1899_)
  );
  XOR2_X1 _7188_ (
    .A(_1883_),
    .B(_1898_),
    .Z(_1900_)
  );
  AND2_X1 _7189_ (
    .A1(_1882_),
    .A2(_1900_),
    .ZN(_1901_)
  );
  XOR2_X1 _7190_ (
    .A(_1882_),
    .B(_1900_),
    .Z(_1902_)
  );
  OR2_X1 _7191_ (
    .A1(_1524_),
    .A2(_1767_),
    .ZN(_1903_)
  );
  OR2_X1 _7192_ (
    .A1(_1426_),
    .A2(_1903_),
    .ZN(_1904_)
  );
  INV_X1 _7193_ (
    .A(_1904_),
    .ZN(_1905_)
  );
  AND2_X1 _7194_ (
    .A1(_1773_),
    .A2(_1903_),
    .ZN(_1906_)
  );
  AND2_X1 _7195_ (
    .A1(_1770_),
    .A2(_1903_),
    .ZN(_1907_)
  );
  OR2_X1 _7196_ (
    .A1(_1774_),
    .A2(_1907_),
    .ZN(_1908_)
  );
  INV_X1 _7197_ (
    .A(_1908_),
    .ZN(_1909_)
  );
  OR2_X1 _7198_ (
    .A1(_1905_),
    .A2(_1906_),
    .ZN(_1910_)
  );
  OR2_X1 _7199_ (
    .A1(_1543_),
    .A2(_1910_),
    .ZN(_1911_)
  );
  XOR2_X1 _7200_ (
    .A(_1543_),
    .B(_1910_),
    .Z(_1912_)
  );
  AND2_X1 _7201_ (
    .A1(_1902_),
    .A2(_1912_),
    .ZN(_1913_)
  );
  XOR2_X1 _7202_ (
    .A(_1902_),
    .B(_1912_),
    .Z(_1914_)
  );
  AND2_X1 _7203_ (
    .A1(_1881_),
    .A2(_1914_),
    .ZN(_1915_)
  );
  XOR2_X1 _7204_ (
    .A(_1881_),
    .B(_1914_),
    .Z(_1916_)
  );
  AND2_X1 _7205_ (
    .A1(divisor[22]),
    .A2(remainder[2]),
    .ZN(_1917_)
  );
  AND2_X1 _7206_ (
    .A1(divisor[24]),
    .A2(remainder[0]),
    .ZN(_1918_)
  );
  AND2_X1 _7207_ (
    .A1(divisor[24]),
    .A2(remainder[1]),
    .ZN(_1919_)
  );
  AND2_X1 _7208_ (
    .A1(_1806_),
    .A2(_1919_),
    .ZN(_1920_)
  );
  XOR2_X1 _7209_ (
    .A(_1808_),
    .B(_1918_),
    .Z(_1921_)
  );
  AND2_X1 _7210_ (
    .A1(_1917_),
    .A2(_1921_),
    .ZN(_1922_)
  );
  XOR2_X1 _7211_ (
    .A(_1917_),
    .B(_1921_),
    .Z(_1923_)
  );
  AND2_X1 _7212_ (
    .A1(_1809_),
    .A2(_1923_),
    .ZN(_1924_)
  );
  XOR2_X1 _7213_ (
    .A(_1809_),
    .B(_1923_),
    .Z(_1925_)
  );
  AND2_X1 _7214_ (
    .A1(divisor[19]),
    .A2(remainder[5]),
    .ZN(_1926_)
  );
  AND2_X1 _7215_ (
    .A1(divisor[20]),
    .A2(remainder[4]),
    .ZN(_1927_)
  );
  AND2_X1 _7216_ (
    .A1(divisor[21]),
    .A2(remainder[4]),
    .ZN(_1928_)
  );
  AND2_X1 _7217_ (
    .A1(_1813_),
    .A2(_1927_),
    .ZN(_1929_)
  );
  XOR2_X1 _7218_ (
    .A(_1813_),
    .B(_1927_),
    .Z(_1930_)
  );
  AND2_X1 _7219_ (
    .A1(_1926_),
    .A2(_1930_),
    .ZN(_1931_)
  );
  XOR2_X1 _7220_ (
    .A(_1926_),
    .B(_1930_),
    .Z(_1932_)
  );
  AND2_X1 _7221_ (
    .A1(_1925_),
    .A2(_1932_),
    .ZN(_1933_)
  );
  XOR2_X1 _7222_ (
    .A(_1925_),
    .B(_1932_),
    .Z(_1934_)
  );
  INV_X1 _7223_ (
    .A(_1934_),
    .ZN(_1935_)
  );
  XOR2_X1 _7224_ (
    .A(_1878_),
    .B(_1935_),
    .Z(_1936_)
  );
  XOR2_X1 _7225_ (
    .A(_1878_),
    .B(_1934_),
    .Z(_1937_)
  );
  AND2_X1 _7226_ (
    .A1(_1916_),
    .A2(_1937_),
    .ZN(_1938_)
  );
  XOR2_X1 _7227_ (
    .A(_1916_),
    .B(_1936_),
    .Z(_1939_)
  );
  INV_X1 _7228_ (
    .A(_1939_),
    .ZN(_1940_)
  );
  AND2_X1 _7229_ (
    .A1(_1880_),
    .A2(_1940_),
    .ZN(_1941_)
  );
  XOR2_X1 _7230_ (
    .A(_1880_),
    .B(_1940_),
    .Z(_1942_)
  );
  OR2_X1 _7231_ (
    .A1(_1836_),
    .A2(_1838_),
    .ZN(_1943_)
  );
  OR2_X1 _7232_ (
    .A1(_1832_),
    .A2(_1834_),
    .ZN(_1944_)
  );
  OR2_X1 _7233_ (
    .A1(_1777_),
    .A2(_1780_),
    .ZN(_1945_)
  );
  AND2_X1 _7234_ (
    .A1(_1703_),
    .A2(_1945_),
    .ZN(_1946_)
  );
  XOR2_X1 _7235_ (
    .A(_1703_),
    .B(_1945_),
    .Z(_1947_)
  );
  AND2_X1 _7236_ (
    .A1(_1829_),
    .A2(_1947_),
    .ZN(_1948_)
  );
  XOR2_X1 _7237_ (
    .A(_1829_),
    .B(_1947_),
    .Z(_1949_)
  );
  AND2_X1 _7238_ (
    .A1(_1944_),
    .A2(_1949_),
    .ZN(_1950_)
  );
  XOR2_X1 _7239_ (
    .A(_1944_),
    .B(_1949_),
    .Z(_1951_)
  );
  AND2_X1 _7240_ (
    .A1(_0512_),
    .A2(_1951_),
    .ZN(_1952_)
  );
  XOR2_X1 _7241_ (
    .A(_0512_),
    .B(_1951_),
    .Z(_1953_)
  );
  AND2_X1 _7242_ (
    .A1(_1804_),
    .A2(_1953_),
    .ZN(_1954_)
  );
  XOR2_X1 _7243_ (
    .A(_1804_),
    .B(_1953_),
    .Z(_1955_)
  );
  AND2_X1 _7244_ (
    .A1(_1943_),
    .A2(_1955_),
    .ZN(_1956_)
  );
  XOR2_X1 _7245_ (
    .A(_1943_),
    .B(_1955_),
    .Z(_1957_)
  );
  AND2_X1 _7246_ (
    .A1(_1942_),
    .A2(_1957_),
    .ZN(_1958_)
  );
  XOR2_X1 _7247_ (
    .A(_1942_),
    .B(_1957_),
    .Z(_1959_)
  );
  AND2_X1 _7248_ (
    .A1(_1877_),
    .A2(_1959_),
    .ZN(_1960_)
  );
  XOR2_X1 _7249_ (
    .A(_1877_),
    .B(_1959_),
    .Z(_1961_)
  );
  AND2_X1 _7250_ (
    .A1(_1876_),
    .A2(_1961_),
    .ZN(_1962_)
  );
  XOR2_X1 _7251_ (
    .A(_1876_),
    .B(_1961_),
    .Z(_1963_)
  );
  AND2_X1 _7252_ (
    .A1(_1875_),
    .A2(_1963_),
    .ZN(_1964_)
  );
  INV_X1 _7253_ (
    .A(_1964_),
    .ZN(_1965_)
  );
  XOR2_X1 _7254_ (
    .A(_1875_),
    .B(_1963_),
    .Z(_1966_)
  );
  AND2_X1 _7255_ (
    .A1(_1850_),
    .A2(_1966_),
    .ZN(_1967_)
  );
  XOR2_X1 _7256_ (
    .A(_1850_),
    .B(_1966_),
    .Z(_1968_)
  );
  XOR2_X1 _7257_ (
    .A(_1851_),
    .B(_1966_),
    .Z(_1969_)
  );
  OR2_X1 _7258_ (
    .A1(_1854_),
    .A2(_1856_),
    .ZN(_1970_)
  );
  AND2_X1 _7259_ (
    .A1(_1968_),
    .A2(_1970_),
    .ZN(_1971_)
  );
  XOR2_X1 _7260_ (
    .A(_1968_),
    .B(_1970_),
    .Z(_1972_)
  );
  XOR2_X1 _7261_ (
    .A(_1969_),
    .B(_1970_),
    .Z(_1973_)
  );
  AND2_X1 _7262_ (
    .A1(remainder[57]),
    .A2(_1972_),
    .ZN(_1974_)
  );
  OR2_X1 _7263_ (
    .A1(_3013_),
    .A2(_1973_),
    .ZN(_1975_)
  );
  XOR2_X1 _7264_ (
    .A(remainder[57]),
    .B(_1972_),
    .Z(_1976_)
  );
  INV_X1 _7265_ (
    .A(_1976_),
    .ZN(_1977_)
  );
  AND2_X1 _7266_ (
    .A1(_1874_),
    .A2(_1976_),
    .ZN(_1978_)
  );
  OR2_X1 _7267_ (
    .A1(_1873_),
    .A2(_1977_),
    .ZN(_1979_)
  );
  OR2_X1 _7268_ (
    .A1(_1874_),
    .A2(_1976_),
    .ZN(_1980_)
  );
  AND2_X1 _7269_ (
    .A1(_4613_),
    .A2(_1980_),
    .ZN(_1981_)
  );
  AND2_X1 _7270_ (
    .A1(_1979_),
    .A2(_1981_),
    .ZN(_1982_)
  );
  AND2_X1 _7271_ (
    .A1(remainder[49]),
    .A2(_4610_),
    .ZN(_1983_)
  );
  OR2_X1 _7272_ (
    .A1(_1982_),
    .A2(_1983_),
    .ZN(_1984_)
  );
  OR2_X1 _7273_ (
    .A1(_1872_),
    .A2(_1984_),
    .ZN(_1985_)
  );
  AND2_X1 _7274_ (
    .A1(_3911_),
    .A2(_1985_),
    .ZN(_0070_)
  );
  MUX2_X1 _7275_ (
    .A(remainder[49]),
    .B(_4523_),
    .S(_4393_),
    .Z(_1986_)
  );
  AND2_X1 _7276_ (
    .A1(_3678_),
    .A2(_1986_),
    .ZN(_1987_)
  );
  AND2_X1 _7277_ (
    .A1(remainder[50]),
    .A2(_4610_),
    .ZN(_1988_)
  );
  AND2_X1 _7278_ (
    .A1(_1975_),
    .A2(_1979_),
    .ZN(_1989_)
  );
  OR2_X1 _7279_ (
    .A1(_1974_),
    .A2(_1978_),
    .ZN(_1990_)
  );
  OR2_X1 _7280_ (
    .A1(_1967_),
    .A2(_1971_),
    .ZN(_1991_)
  );
  INV_X1 _7281_ (
    .A(_1991_),
    .ZN(_1992_)
  );
  OR2_X1 _7282_ (
    .A1(_1960_),
    .A2(_1962_),
    .ZN(_1993_)
  );
  INV_X1 _7283_ (
    .A(_1993_),
    .ZN(_1994_)
  );
  OR2_X1 _7284_ (
    .A1(_1954_),
    .A2(_1956_),
    .ZN(_1995_)
  );
  OR2_X1 _7285_ (
    .A1(_1941_),
    .A2(_1958_),
    .ZN(_1996_)
  );
  AND2_X1 _7286_ (
    .A1(_0541_),
    .A2(_1935_),
    .ZN(_1997_)
  );
  AND2_X1 _7287_ (
    .A1(_1819_),
    .A2(_1997_),
    .ZN(_1998_)
  );
  OR2_X1 _7288_ (
    .A1(_1938_),
    .A2(_1998_),
    .ZN(_1999_)
  );
  OR2_X1 _7289_ (
    .A1(_1901_),
    .A2(_1913_),
    .ZN(_2000_)
  );
  OR2_X1 _7290_ (
    .A1(_1897_),
    .A2(_1899_),
    .ZN(_2001_)
  );
  OR2_X1 _7291_ (
    .A1(_1893_),
    .A2(_1895_),
    .ZN(_2002_)
  );
  OR2_X1 _7292_ (
    .A1(_1924_),
    .A2(_1933_),
    .ZN(_2003_)
  );
  OR2_X1 _7293_ (
    .A1(_1889_),
    .A2(_1891_),
    .ZN(_2004_)
  );
  OR2_X1 _7294_ (
    .A1(_1929_),
    .A2(_1931_),
    .ZN(_2005_)
  );
  AND2_X1 _7295_ (
    .A1(remainder[32]),
    .A2(divisor[18]),
    .ZN(_2006_)
  );
  AND2_X1 _7296_ (
    .A1(remainder[32]),
    .A2(divisor[17]),
    .ZN(_2007_)
  );
  AND2_X1 _7297_ (
    .A1(divisor[18]),
    .A2(_2007_),
    .ZN(_2008_)
  );
  AND2_X1 _7298_ (
    .A1(_1888_),
    .A2(_2007_),
    .ZN(_2009_)
  );
  XOR2_X1 _7299_ (
    .A(_1888_),
    .B(_2007_),
    .Z(_2010_)
  );
  AND2_X1 _7300_ (
    .A1(_1886_),
    .A2(_2010_),
    .ZN(_2011_)
  );
  XOR2_X1 _7301_ (
    .A(_1886_),
    .B(_2010_),
    .Z(_2012_)
  );
  AND2_X1 _7302_ (
    .A1(_2005_),
    .A2(_2012_),
    .ZN(_2013_)
  );
  XOR2_X1 _7303_ (
    .A(_2005_),
    .B(_2012_),
    .Z(_2014_)
  );
  AND2_X1 _7304_ (
    .A1(_2004_),
    .A2(_2014_),
    .ZN(_2015_)
  );
  XOR2_X1 _7305_ (
    .A(_2004_),
    .B(_2014_),
    .Z(_2016_)
  );
  AND2_X1 _7306_ (
    .A1(_2003_),
    .A2(_2016_),
    .ZN(_2017_)
  );
  XOR2_X1 _7307_ (
    .A(_2003_),
    .B(_2016_),
    .Z(_2018_)
  );
  AND2_X1 _7308_ (
    .A1(_2002_),
    .A2(_2018_),
    .ZN(_2019_)
  );
  XOR2_X1 _7309_ (
    .A(_2002_),
    .B(_2018_),
    .Z(_2020_)
  );
  AND2_X1 _7310_ (
    .A1(_2001_),
    .A2(_2020_),
    .ZN(_2021_)
  );
  XOR2_X1 _7311_ (
    .A(_2001_),
    .B(_2020_),
    .Z(_2022_)
  );
  OR2_X1 _7312_ (
    .A1(_1905_),
    .A2(_1909_),
    .ZN(_2023_)
  );
  OR2_X1 _7313_ (
    .A1(_1543_),
    .A2(_2023_),
    .ZN(_2024_)
  );
  XOR2_X1 _7314_ (
    .A(_1543_),
    .B(_2023_),
    .Z(_2025_)
  );
  AND2_X1 _7315_ (
    .A1(_2022_),
    .A2(_2025_),
    .ZN(_2026_)
  );
  XOR2_X1 _7316_ (
    .A(_2022_),
    .B(_2025_),
    .Z(_2027_)
  );
  AND2_X1 _7317_ (
    .A1(_2000_),
    .A2(_2027_),
    .ZN(_2028_)
  );
  XOR2_X1 _7318_ (
    .A(_2000_),
    .B(_2027_),
    .Z(_2029_)
  );
  AND2_X1 _7319_ (
    .A1(divisor[25]),
    .A2(remainder[0]),
    .ZN(_2030_)
  );
  OR2_X1 _7320_ (
    .A1(_1920_),
    .A2(_1922_),
    .ZN(_2031_)
  );
  AND2_X1 _7321_ (
    .A1(divisor[22]),
    .A2(remainder[3]),
    .ZN(_2032_)
  );
  AND2_X1 _7322_ (
    .A1(divisor[23]),
    .A2(remainder[2]),
    .ZN(_2033_)
  );
  AND2_X1 _7323_ (
    .A1(divisor[24]),
    .A2(remainder[2]),
    .ZN(_2034_)
  );
  AND2_X1 _7324_ (
    .A1(_1808_),
    .A2(_2034_),
    .ZN(_2035_)
  );
  XOR2_X1 _7325_ (
    .A(_1919_),
    .B(_2033_),
    .Z(_2036_)
  );
  AND2_X1 _7326_ (
    .A1(_2032_),
    .A2(_2036_),
    .ZN(_2037_)
  );
  XOR2_X1 _7327_ (
    .A(_2032_),
    .B(_2036_),
    .Z(_2038_)
  );
  AND2_X1 _7328_ (
    .A1(_2031_),
    .A2(_2038_),
    .ZN(_2039_)
  );
  XOR2_X1 _7329_ (
    .A(_2031_),
    .B(_2038_),
    .Z(_2040_)
  );
  AND2_X1 _7330_ (
    .A1(divisor[19]),
    .A2(remainder[6]),
    .ZN(_2041_)
  );
  AND2_X1 _7331_ (
    .A1(divisor[20]),
    .A2(remainder[5]),
    .ZN(_2042_)
  );
  AND2_X1 _7332_ (
    .A1(divisor[21]),
    .A2(remainder[5]),
    .ZN(_2043_)
  );
  AND2_X1 _7333_ (
    .A1(_1928_),
    .A2(_2042_),
    .ZN(_2044_)
  );
  XOR2_X1 _7334_ (
    .A(_1928_),
    .B(_2042_),
    .Z(_2045_)
  );
  AND2_X1 _7335_ (
    .A1(_2041_),
    .A2(_2045_),
    .ZN(_2046_)
  );
  XOR2_X1 _7336_ (
    .A(_2041_),
    .B(_2045_),
    .Z(_2047_)
  );
  AND2_X1 _7337_ (
    .A1(_2040_),
    .A2(_2047_),
    .ZN(_2048_)
  );
  XOR2_X1 _7338_ (
    .A(_2040_),
    .B(_2047_),
    .Z(_2049_)
  );
  AND2_X1 _7339_ (
    .A1(_2030_),
    .A2(_2049_),
    .ZN(_2050_)
  );
  XOR2_X1 _7340_ (
    .A(_2030_),
    .B(_2049_),
    .Z(_2051_)
  );
  XOR2_X1 _7341_ (
    .A(_1997_),
    .B(_2051_),
    .Z(_2052_)
  );
  AND2_X1 _7342_ (
    .A1(_2029_),
    .A2(_2052_),
    .ZN(_2053_)
  );
  INV_X1 _7343_ (
    .A(_2053_),
    .ZN(_2054_)
  );
  XOR2_X1 _7344_ (
    .A(_2029_),
    .B(_2052_),
    .Z(_2055_)
  );
  AND2_X1 _7345_ (
    .A1(_1999_),
    .A2(_2055_),
    .ZN(_2056_)
  );
  XOR2_X1 _7346_ (
    .A(_1999_),
    .B(_2055_),
    .Z(_2057_)
  );
  OR2_X1 _7347_ (
    .A1(_1950_),
    .A2(_1952_),
    .ZN(_2058_)
  );
  OR2_X1 _7348_ (
    .A1(_1946_),
    .A2(_1948_),
    .ZN(_2059_)
  );
  AND2_X1 _7349_ (
    .A1(_1908_),
    .A2(_1911_),
    .ZN(_2060_)
  );
  OR2_X1 _7350_ (
    .A1(_1704_),
    .A2(_2060_),
    .ZN(_2061_)
  );
  XOR2_X1 _7351_ (
    .A(_1703_),
    .B(_2060_),
    .Z(_2062_)
  );
  OR2_X1 _7352_ (
    .A1(_1830_),
    .A2(_2062_),
    .ZN(_2063_)
  );
  XOR2_X1 _7353_ (
    .A(_1830_),
    .B(_2062_),
    .Z(_2064_)
  );
  AND2_X1 _7354_ (
    .A1(_2059_),
    .A2(_2064_),
    .ZN(_2065_)
  );
  XOR2_X1 _7355_ (
    .A(_2059_),
    .B(_2064_),
    .Z(_2066_)
  );
  AND2_X1 _7356_ (
    .A1(_0512_),
    .A2(_2066_),
    .ZN(_2067_)
  );
  XOR2_X1 _7357_ (
    .A(_0512_),
    .B(_2066_),
    .Z(_2068_)
  );
  AND2_X1 _7358_ (
    .A1(_1915_),
    .A2(_2068_),
    .ZN(_2069_)
  );
  XOR2_X1 _7359_ (
    .A(_1915_),
    .B(_2068_),
    .Z(_2070_)
  );
  AND2_X1 _7360_ (
    .A1(_2058_),
    .A2(_2070_),
    .ZN(_2071_)
  );
  XOR2_X1 _7361_ (
    .A(_2058_),
    .B(_2070_),
    .Z(_2072_)
  );
  AND2_X1 _7362_ (
    .A1(_2057_),
    .A2(_2072_),
    .ZN(_2073_)
  );
  XOR2_X1 _7363_ (
    .A(_2057_),
    .B(_2072_),
    .Z(_2074_)
  );
  AND2_X1 _7364_ (
    .A1(_1996_),
    .A2(_2074_),
    .ZN(_2075_)
  );
  XOR2_X1 _7365_ (
    .A(_1996_),
    .B(_2074_),
    .Z(_2076_)
  );
  AND2_X1 _7366_ (
    .A1(_1995_),
    .A2(_2076_),
    .ZN(_2077_)
  );
  XOR2_X1 _7367_ (
    .A(_1995_),
    .B(_2076_),
    .Z(_2078_)
  );
  AND2_X1 _7368_ (
    .A1(_1993_),
    .A2(_2078_),
    .ZN(_2079_)
  );
  INV_X1 _7369_ (
    .A(_2079_),
    .ZN(_2080_)
  );
  XOR2_X1 _7370_ (
    .A(_1994_),
    .B(_2078_),
    .Z(_2081_)
  );
  OR2_X1 _7371_ (
    .A1(_1965_),
    .A2(_2081_),
    .ZN(_2082_)
  );
  INV_X1 _7372_ (
    .A(_2082_),
    .ZN(_2083_)
  );
  XOR2_X1 _7373_ (
    .A(_1965_),
    .B(_2081_),
    .Z(_2084_)
  );
  AND2_X1 _7374_ (
    .A1(_1991_),
    .A2(_2084_),
    .ZN(_2085_)
  );
  XOR2_X1 _7375_ (
    .A(_1991_),
    .B(_2084_),
    .Z(_2086_)
  );
  XOR2_X1 _7376_ (
    .A(_1992_),
    .B(_2084_),
    .Z(_2087_)
  );
  OR2_X1 _7377_ (
    .A1(_3002_),
    .A2(_2087_),
    .ZN(_2088_)
  );
  INV_X1 _7378_ (
    .A(_2088_),
    .ZN(_2089_)
  );
  OR2_X1 _7379_ (
    .A1(remainder[58]),
    .A2(_2086_),
    .ZN(_2090_)
  );
  INV_X1 _7380_ (
    .A(_2090_),
    .ZN(_2091_)
  );
  AND2_X1 _7381_ (
    .A1(_2088_),
    .A2(_2090_),
    .ZN(_2092_)
  );
  XOR2_X1 _7382_ (
    .A(_1990_),
    .B(_2092_),
    .Z(_2093_)
  );
  AND2_X1 _7383_ (
    .A1(_4613_),
    .A2(_2093_),
    .ZN(_2094_)
  );
  OR2_X1 _7384_ (
    .A1(_1988_),
    .A2(_2094_),
    .ZN(_2095_)
  );
  OR2_X1 _7385_ (
    .A1(_1987_),
    .A2(_2095_),
    .ZN(_2096_)
  );
  AND2_X1 _7386_ (
    .A1(_3911_),
    .A2(_2096_),
    .ZN(_0071_)
  );
  OR2_X1 _7387_ (
    .A1(_2075_),
    .A2(_2077_),
    .ZN(_2097_)
  );
  OR2_X1 _7388_ (
    .A1(_2069_),
    .A2(_2071_),
    .ZN(_2098_)
  );
  OR2_X1 _7389_ (
    .A1(_2056_),
    .A2(_2073_),
    .ZN(_2099_)
  );
  OR2_X1 _7390_ (
    .A1(_0542_),
    .A2(_2051_),
    .ZN(_2100_)
  );
  OR2_X1 _7391_ (
    .A1(_1935_),
    .A2(_2100_),
    .ZN(_2101_)
  );
  AND2_X1 _7392_ (
    .A1(_2054_),
    .A2(_2101_),
    .ZN(_2102_)
  );
  OR2_X1 _7393_ (
    .A1(_2021_),
    .A2(_2026_),
    .ZN(_2103_)
  );
  OR2_X1 _7394_ (
    .A1(_2017_),
    .A2(_2019_),
    .ZN(_2104_)
  );
  OR2_X1 _7395_ (
    .A1(_2013_),
    .A2(_2015_),
    .ZN(_2105_)
  );
  OR2_X1 _7396_ (
    .A1(_2039_),
    .A2(_2048_),
    .ZN(_2106_)
  );
  OR2_X1 _7397_ (
    .A1(_2009_),
    .A2(_2011_),
    .ZN(_2107_)
  );
  OR2_X1 _7398_ (
    .A1(_2044_),
    .A2(_2046_),
    .ZN(_2108_)
  );
  MUX2_X1 _7399_ (
    .A(_2007_),
    .B(_3351_),
    .S(_2006_),
    .Z(_2109_)
  );
  AND2_X1 _7400_ (
    .A1(divisor[16]),
    .A2(_2109_),
    .ZN(_2110_)
  );
  MUX2_X1 _7401_ (
    .A(_1886_),
    .B(_3340_),
    .S(_2109_),
    .Z(_2111_)
  );
  AND2_X1 _7402_ (
    .A1(_2108_),
    .A2(_2111_),
    .ZN(_2112_)
  );
  XOR2_X1 _7403_ (
    .A(_2108_),
    .B(_2111_),
    .Z(_2113_)
  );
  AND2_X1 _7404_ (
    .A1(_2107_),
    .A2(_2113_),
    .ZN(_2114_)
  );
  XOR2_X1 _7405_ (
    .A(_2107_),
    .B(_2113_),
    .Z(_2115_)
  );
  AND2_X1 _7406_ (
    .A1(_2106_),
    .A2(_2115_),
    .ZN(_2116_)
  );
  XOR2_X1 _7407_ (
    .A(_2106_),
    .B(_2115_),
    .Z(_2117_)
  );
  AND2_X1 _7408_ (
    .A1(_2105_),
    .A2(_2117_),
    .ZN(_2118_)
  );
  XOR2_X1 _7409_ (
    .A(_2105_),
    .B(_2117_),
    .Z(_2119_)
  );
  AND2_X1 _7410_ (
    .A1(_2104_),
    .A2(_2119_),
    .ZN(_2120_)
  );
  XOR2_X1 _7411_ (
    .A(_2104_),
    .B(_2119_),
    .Z(_2121_)
  );
  AND2_X1 _7412_ (
    .A1(_2025_),
    .A2(_2121_),
    .ZN(_2122_)
  );
  XOR2_X1 _7413_ (
    .A(_2025_),
    .B(_2121_),
    .Z(_2123_)
  );
  AND2_X1 _7414_ (
    .A1(_2103_),
    .A2(_2123_),
    .ZN(_2124_)
  );
  XOR2_X1 _7415_ (
    .A(_2103_),
    .B(_2123_),
    .Z(_2125_)
  );
  AND2_X1 _7416_ (
    .A1(divisor[26]),
    .A2(remainder[0]),
    .ZN(_2126_)
  );
  AND2_X1 _7417_ (
    .A1(divisor[25]),
    .A2(remainder[1]),
    .ZN(_2127_)
  );
  AND2_X1 _7418_ (
    .A1(divisor[26]),
    .A2(remainder[1]),
    .ZN(_2128_)
  );
  AND2_X1 _7419_ (
    .A1(_2030_),
    .A2(_2128_),
    .ZN(_2129_)
  );
  XOR2_X1 _7420_ (
    .A(_2126_),
    .B(_2127_),
    .Z(_2130_)
  );
  OR2_X1 _7421_ (
    .A1(_2035_),
    .A2(_2037_),
    .ZN(_2131_)
  );
  AND2_X1 _7422_ (
    .A1(divisor[22]),
    .A2(remainder[4]),
    .ZN(_2132_)
  );
  AND2_X1 _7423_ (
    .A1(divisor[23]),
    .A2(remainder[3]),
    .ZN(_2133_)
  );
  AND2_X1 _7424_ (
    .A1(divisor[24]),
    .A2(remainder[3]),
    .ZN(_2134_)
  );
  AND2_X1 _7425_ (
    .A1(_2034_),
    .A2(_2133_),
    .ZN(_2135_)
  );
  XOR2_X1 _7426_ (
    .A(_2034_),
    .B(_2133_),
    .Z(_2136_)
  );
  AND2_X1 _7427_ (
    .A1(_2132_),
    .A2(_2136_),
    .ZN(_2137_)
  );
  XOR2_X1 _7428_ (
    .A(_2132_),
    .B(_2136_),
    .Z(_2138_)
  );
  AND2_X1 _7429_ (
    .A1(_2131_),
    .A2(_2138_),
    .ZN(_2139_)
  );
  XOR2_X1 _7430_ (
    .A(_2131_),
    .B(_2138_),
    .Z(_2140_)
  );
  AND2_X1 _7431_ (
    .A1(divisor[19]),
    .A2(remainder[7]),
    .ZN(_2141_)
  );
  AND2_X1 _7432_ (
    .A1(divisor[20]),
    .A2(remainder[6]),
    .ZN(_2142_)
  );
  AND2_X1 _7433_ (
    .A1(divisor[21]),
    .A2(remainder[6]),
    .ZN(_2143_)
  );
  AND2_X1 _7434_ (
    .A1(_2043_),
    .A2(_2142_),
    .ZN(_2144_)
  );
  XOR2_X1 _7435_ (
    .A(_2043_),
    .B(_2142_),
    .Z(_2145_)
  );
  AND2_X1 _7436_ (
    .A1(_2141_),
    .A2(_2145_),
    .ZN(_2146_)
  );
  XOR2_X1 _7437_ (
    .A(_2141_),
    .B(_2145_),
    .Z(_2147_)
  );
  AND2_X1 _7438_ (
    .A1(_2140_),
    .A2(_2147_),
    .ZN(_2148_)
  );
  XOR2_X1 _7439_ (
    .A(_2140_),
    .B(_2147_),
    .Z(_2149_)
  );
  AND2_X1 _7440_ (
    .A1(_2130_),
    .A2(_2149_),
    .ZN(_2150_)
  );
  XOR2_X1 _7441_ (
    .A(_2130_),
    .B(_2149_),
    .Z(_2151_)
  );
  AND2_X1 _7442_ (
    .A1(_2050_),
    .A2(_2151_),
    .ZN(_2152_)
  );
  XOR2_X1 _7443_ (
    .A(_2050_),
    .B(_2151_),
    .Z(_2153_)
  );
  INV_X1 _7444_ (
    .A(_2153_),
    .ZN(_2154_)
  );
  XOR2_X1 _7445_ (
    .A(_2100_),
    .B(_2153_),
    .Z(_2155_)
  );
  XOR2_X1 _7446_ (
    .A(_2100_),
    .B(_2154_),
    .Z(_2156_)
  );
  AND2_X1 _7447_ (
    .A1(_2125_),
    .A2(_2156_),
    .ZN(_2157_)
  );
  XOR2_X1 _7448_ (
    .A(_2125_),
    .B(_2155_),
    .Z(_2158_)
  );
  OR2_X1 _7449_ (
    .A1(_2102_),
    .A2(_2158_),
    .ZN(_2159_)
  );
  INV_X1 _7450_ (
    .A(_2159_),
    .ZN(_2160_)
  );
  XOR2_X1 _7451_ (
    .A(_2102_),
    .B(_2158_),
    .Z(_2161_)
  );
  OR2_X1 _7452_ (
    .A1(_2065_),
    .A2(_2067_),
    .ZN(_2162_)
  );
  AND2_X1 _7453_ (
    .A1(_2061_),
    .A2(_2063_),
    .ZN(_2163_)
  );
  INV_X1 _7454_ (
    .A(_2163_),
    .ZN(_2164_)
  );
  AND2_X1 _7455_ (
    .A1(_1908_),
    .A2(_2024_),
    .ZN(_2165_)
  );
  AND2_X1 _7456_ (
    .A1(_1704_),
    .A2(_2165_),
    .ZN(_2166_)
  );
  XOR2_X1 _7457_ (
    .A(_1704_),
    .B(_2165_),
    .Z(_2167_)
  );
  XOR2_X1 _7458_ (
    .A(_1829_),
    .B(_2167_),
    .Z(_2168_)
  );
  AND2_X1 _7459_ (
    .A1(_2164_),
    .A2(_2168_),
    .ZN(_2169_)
  );
  INV_X1 _7460_ (
    .A(_2169_),
    .ZN(_2170_)
  );
  XOR2_X1 _7461_ (
    .A(_2163_),
    .B(_2168_),
    .Z(_2171_)
  );
  INV_X1 _7462_ (
    .A(_2171_),
    .ZN(_2172_)
  );
  AND2_X1 _7463_ (
    .A1(_0512_),
    .A2(_2172_),
    .ZN(_2173_)
  );
  XOR2_X1 _7464_ (
    .A(_0511_),
    .B(_2171_),
    .Z(_2174_)
  );
  AND2_X1 _7465_ (
    .A1(_2028_),
    .A2(_2174_),
    .ZN(_2175_)
  );
  XOR2_X1 _7466_ (
    .A(_2028_),
    .B(_2174_),
    .Z(_2176_)
  );
  AND2_X1 _7467_ (
    .A1(_2162_),
    .A2(_2176_),
    .ZN(_2177_)
  );
  XOR2_X1 _7468_ (
    .A(_2162_),
    .B(_2176_),
    .Z(_2178_)
  );
  AND2_X1 _7469_ (
    .A1(_2161_),
    .A2(_2178_),
    .ZN(_2179_)
  );
  XOR2_X1 _7470_ (
    .A(_2161_),
    .B(_2178_),
    .Z(_2180_)
  );
  AND2_X1 _7471_ (
    .A1(_2099_),
    .A2(_2180_),
    .ZN(_2181_)
  );
  XOR2_X1 _7472_ (
    .A(_2099_),
    .B(_2180_),
    .Z(_2182_)
  );
  AND2_X1 _7473_ (
    .A1(_2098_),
    .A2(_2182_),
    .ZN(_2183_)
  );
  XOR2_X1 _7474_ (
    .A(_2098_),
    .B(_2182_),
    .Z(_2184_)
  );
  AND2_X1 _7475_ (
    .A1(_2097_),
    .A2(_2184_),
    .ZN(_2185_)
  );
  XOR2_X1 _7476_ (
    .A(_2097_),
    .B(_2184_),
    .Z(_2186_)
  );
  AND2_X1 _7477_ (
    .A1(_2079_),
    .A2(_2186_),
    .ZN(_2187_)
  );
  XOR2_X1 _7478_ (
    .A(_2079_),
    .B(_2186_),
    .Z(_2188_)
  );
  XOR2_X1 _7479_ (
    .A(_2080_),
    .B(_2186_),
    .Z(_2189_)
  );
  OR2_X1 _7480_ (
    .A1(_2083_),
    .A2(_2085_),
    .ZN(_2190_)
  );
  AND2_X1 _7481_ (
    .A1(_2188_),
    .A2(_2190_),
    .ZN(_2191_)
  );
  XOR2_X1 _7482_ (
    .A(_2188_),
    .B(_2190_),
    .Z(_2192_)
  );
  XOR2_X1 _7483_ (
    .A(_2189_),
    .B(_2190_),
    .Z(_2193_)
  );
  AND2_X1 _7484_ (
    .A1(remainder[59]),
    .A2(_2192_),
    .ZN(_2194_)
  );
  OR2_X1 _7485_ (
    .A1(_2991_),
    .A2(_2193_),
    .ZN(_2195_)
  );
  XOR2_X1 _7486_ (
    .A(remainder[59]),
    .B(_2192_),
    .Z(_2196_)
  );
  INV_X1 _7487_ (
    .A(_2196_),
    .ZN(_2197_)
  );
  AND2_X1 _7488_ (
    .A1(_1989_),
    .A2(_2088_),
    .ZN(_2198_)
  );
  OR2_X1 _7489_ (
    .A1(_1990_),
    .A2(_2089_),
    .ZN(_2199_)
  );
  AND2_X1 _7490_ (
    .A1(_2090_),
    .A2(_2199_),
    .ZN(_2200_)
  );
  OR2_X1 _7491_ (
    .A1(_2091_),
    .A2(_2198_),
    .ZN(_2201_)
  );
  AND2_X1 _7492_ (
    .A1(_2196_),
    .A2(_2200_),
    .ZN(_2202_)
  );
  OR2_X1 _7493_ (
    .A1(_2197_),
    .A2(_2201_),
    .ZN(_2203_)
  );
  OR2_X1 _7494_ (
    .A1(_2196_),
    .A2(_2200_),
    .ZN(_2204_)
  );
  AND2_X1 _7495_ (
    .A1(_4613_),
    .A2(_2204_),
    .ZN(_2205_)
  );
  AND2_X1 _7496_ (
    .A1(_2203_),
    .A2(_2205_),
    .ZN(_2206_)
  );
  AND2_X1 _7497_ (
    .A1(remainder[51]),
    .A2(_4610_),
    .ZN(_2207_)
  );
  MUX2_X1 _7498_ (
    .A(remainder[50]),
    .B(_4528_),
    .S(_4393_),
    .Z(_2208_)
  );
  AND2_X1 _7499_ (
    .A1(_3678_),
    .A2(_2208_),
    .ZN(_2209_)
  );
  OR2_X1 _7500_ (
    .A1(_2206_),
    .A2(_2209_),
    .ZN(_2210_)
  );
  OR2_X1 _7501_ (
    .A1(_2207_),
    .A2(_2210_),
    .ZN(_2211_)
  );
  AND2_X1 _7502_ (
    .A1(_3911_),
    .A2(_2211_),
    .ZN(_0072_)
  );
  AND2_X1 _7503_ (
    .A1(_2195_),
    .A2(_2203_),
    .ZN(_2212_)
  );
  OR2_X1 _7504_ (
    .A1(_2194_),
    .A2(_2202_),
    .ZN(_2213_)
  );
  OR2_X1 _7505_ (
    .A1(_2187_),
    .A2(_2191_),
    .ZN(_2214_)
  );
  OR2_X1 _7506_ (
    .A1(_2181_),
    .A2(_2183_),
    .ZN(_2215_)
  );
  OR2_X1 _7507_ (
    .A1(_2175_),
    .A2(_2177_),
    .ZN(_2216_)
  );
  OR2_X1 _7508_ (
    .A1(_2160_),
    .A2(_2179_),
    .ZN(_2217_)
  );
  AND2_X1 _7509_ (
    .A1(_0541_),
    .A2(_2154_),
    .ZN(_2218_)
  );
  AND2_X1 _7510_ (
    .A1(_2051_),
    .A2(_2218_),
    .ZN(_2219_)
  );
  OR2_X1 _7511_ (
    .A1(_2157_),
    .A2(_2219_),
    .ZN(_2220_)
  );
  OR2_X1 _7512_ (
    .A1(_2120_),
    .A2(_2122_),
    .ZN(_2221_)
  );
  OR2_X1 _7513_ (
    .A1(_2116_),
    .A2(_2118_),
    .ZN(_2222_)
  );
  OR2_X1 _7514_ (
    .A1(_2112_),
    .A2(_2114_),
    .ZN(_2223_)
  );
  OR2_X1 _7515_ (
    .A1(_2139_),
    .A2(_2148_),
    .ZN(_2224_)
  );
  OR2_X1 _7516_ (
    .A1(_2008_),
    .A2(_2110_),
    .ZN(_2225_)
  );
  OR2_X1 _7517_ (
    .A1(_2144_),
    .A2(_2146_),
    .ZN(_2226_)
  );
  AND2_X1 _7518_ (
    .A1(_2111_),
    .A2(_2226_),
    .ZN(_2227_)
  );
  XOR2_X1 _7519_ (
    .A(_2111_),
    .B(_2226_),
    .Z(_2228_)
  );
  AND2_X1 _7520_ (
    .A1(_2225_),
    .A2(_2228_),
    .ZN(_2229_)
  );
  XOR2_X1 _7521_ (
    .A(_2225_),
    .B(_2228_),
    .Z(_2230_)
  );
  AND2_X1 _7522_ (
    .A1(_2224_),
    .A2(_2230_),
    .ZN(_2231_)
  );
  XOR2_X1 _7523_ (
    .A(_2224_),
    .B(_2230_),
    .Z(_2232_)
  );
  AND2_X1 _7524_ (
    .A1(_2223_),
    .A2(_2232_),
    .ZN(_2233_)
  );
  XOR2_X1 _7525_ (
    .A(_2223_),
    .B(_2232_),
    .Z(_2234_)
  );
  AND2_X1 _7526_ (
    .A1(_2222_),
    .A2(_2234_),
    .ZN(_2235_)
  );
  XOR2_X1 _7527_ (
    .A(_2222_),
    .B(_2234_),
    .Z(_2236_)
  );
  AND2_X1 _7528_ (
    .A1(_2025_),
    .A2(_2236_),
    .ZN(_2237_)
  );
  XOR2_X1 _7529_ (
    .A(_2025_),
    .B(_2236_),
    .Z(_2238_)
  );
  AND2_X1 _7530_ (
    .A1(_2152_),
    .A2(_2238_),
    .ZN(_2239_)
  );
  XOR2_X1 _7531_ (
    .A(_2152_),
    .B(_2238_),
    .Z(_2240_)
  );
  AND2_X1 _7532_ (
    .A1(_2221_),
    .A2(_2240_),
    .ZN(_2241_)
  );
  XOR2_X1 _7533_ (
    .A(_2221_),
    .B(_2240_),
    .Z(_2242_)
  );
  AND2_X1 _7534_ (
    .A1(divisor[25]),
    .A2(remainder[2]),
    .ZN(_2243_)
  );
  AND2_X1 _7535_ (
    .A1(divisor[27]),
    .A2(remainder[0]),
    .ZN(_2244_)
  );
  AND2_X1 _7536_ (
    .A1(divisor[27]),
    .A2(remainder[1]),
    .ZN(_2245_)
  );
  AND2_X1 _7537_ (
    .A1(_2126_),
    .A2(_2245_),
    .ZN(_2246_)
  );
  XOR2_X1 _7538_ (
    .A(_2128_),
    .B(_2244_),
    .Z(_2247_)
  );
  AND2_X1 _7539_ (
    .A1(_2243_),
    .A2(_2247_),
    .ZN(_2248_)
  );
  XOR2_X1 _7540_ (
    .A(_2243_),
    .B(_2247_),
    .Z(_2249_)
  );
  AND2_X1 _7541_ (
    .A1(_2129_),
    .A2(_2249_),
    .ZN(_2250_)
  );
  XOR2_X1 _7542_ (
    .A(_2129_),
    .B(_2249_),
    .Z(_2251_)
  );
  OR2_X1 _7543_ (
    .A1(_2135_),
    .A2(_2137_),
    .ZN(_2252_)
  );
  AND2_X1 _7544_ (
    .A1(divisor[22]),
    .A2(remainder[5]),
    .ZN(_2253_)
  );
  AND2_X1 _7545_ (
    .A1(divisor[23]),
    .A2(remainder[4]),
    .ZN(_2254_)
  );
  AND2_X1 _7546_ (
    .A1(divisor[24]),
    .A2(remainder[4]),
    .ZN(_2255_)
  );
  AND2_X1 _7547_ (
    .A1(_2134_),
    .A2(_2254_),
    .ZN(_2256_)
  );
  XOR2_X1 _7548_ (
    .A(_2134_),
    .B(_2254_),
    .Z(_2257_)
  );
  AND2_X1 _7549_ (
    .A1(_2253_),
    .A2(_2257_),
    .ZN(_2258_)
  );
  XOR2_X1 _7550_ (
    .A(_2253_),
    .B(_2257_),
    .Z(_2259_)
  );
  AND2_X1 _7551_ (
    .A1(_2252_),
    .A2(_2259_),
    .ZN(_2260_)
  );
  XOR2_X1 _7552_ (
    .A(_2252_),
    .B(_2259_),
    .Z(_2261_)
  );
  AND2_X1 _7553_ (
    .A1(divisor[20]),
    .A2(remainder[7]),
    .ZN(_2262_)
  );
  AND2_X1 _7554_ (
    .A1(divisor[21]),
    .A2(remainder[7]),
    .ZN(_2263_)
  );
  AND2_X1 _7555_ (
    .A1(_2142_),
    .A2(_2263_),
    .ZN(_2264_)
  );
  XOR2_X1 _7556_ (
    .A(_2143_),
    .B(_2262_),
    .Z(_2265_)
  );
  AND2_X1 _7557_ (
    .A1(_1337_),
    .A2(_2265_),
    .ZN(_2266_)
  );
  XOR2_X1 _7558_ (
    .A(_1337_),
    .B(_2265_),
    .Z(_2267_)
  );
  AND2_X1 _7559_ (
    .A1(_2261_),
    .A2(_2267_),
    .ZN(_2268_)
  );
  XOR2_X1 _7560_ (
    .A(_2261_),
    .B(_2267_),
    .Z(_2269_)
  );
  AND2_X1 _7561_ (
    .A1(_2251_),
    .A2(_2269_),
    .ZN(_2270_)
  );
  XOR2_X1 _7562_ (
    .A(_2251_),
    .B(_2269_),
    .Z(_2271_)
  );
  AND2_X1 _7563_ (
    .A1(_2150_),
    .A2(_2271_),
    .ZN(_2272_)
  );
  XOR2_X1 _7564_ (
    .A(_2150_),
    .B(_2271_),
    .Z(_2273_)
  );
  INV_X1 _7565_ (
    .A(_2273_),
    .ZN(_2274_)
  );
  XOR2_X1 _7566_ (
    .A(_2218_),
    .B(_2273_),
    .Z(_2275_)
  );
  AND2_X1 _7567_ (
    .A1(_2242_),
    .A2(_2275_),
    .ZN(_2276_)
  );
  XOR2_X1 _7568_ (
    .A(_2242_),
    .B(_2275_),
    .Z(_2277_)
  );
  AND2_X1 _7569_ (
    .A1(_2220_),
    .A2(_2277_),
    .ZN(_2278_)
  );
  XOR2_X1 _7570_ (
    .A(_2220_),
    .B(_2277_),
    .Z(_2279_)
  );
  OR2_X1 _7571_ (
    .A1(_2169_),
    .A2(_2173_),
    .ZN(_2280_)
  );
  AND2_X1 _7572_ (
    .A1(_1830_),
    .A2(_2166_),
    .ZN(_2281_)
  );
  OR2_X1 _7573_ (
    .A1(_2169_),
    .A2(_2281_),
    .ZN(_2282_)
  );
  INV_X1 _7574_ (
    .A(_2282_),
    .ZN(_2283_)
  );
  AND2_X1 _7575_ (
    .A1(_0512_),
    .A2(_2283_),
    .ZN(_2284_)
  );
  INV_X1 _7576_ (
    .A(_2284_),
    .ZN(_2285_)
  );
  AND2_X1 _7577_ (
    .A1(_0511_),
    .A2(_2282_),
    .ZN(_2286_)
  );
  XOR2_X1 _7578_ (
    .A(_0511_),
    .B(_2282_),
    .Z(_2287_)
  );
  OR2_X1 _7579_ (
    .A1(_2284_),
    .A2(_2286_),
    .ZN(_2288_)
  );
  AND2_X1 _7580_ (
    .A1(_2124_),
    .A2(_2287_),
    .ZN(_2289_)
  );
  XOR2_X1 _7581_ (
    .A(_2124_),
    .B(_2287_),
    .Z(_2290_)
  );
  AND2_X1 _7582_ (
    .A1(_2280_),
    .A2(_2290_),
    .ZN(_2291_)
  );
  XOR2_X1 _7583_ (
    .A(_2280_),
    .B(_2290_),
    .Z(_2292_)
  );
  AND2_X1 _7584_ (
    .A1(_2279_),
    .A2(_2292_),
    .ZN(_2293_)
  );
  XOR2_X1 _7585_ (
    .A(_2279_),
    .B(_2292_),
    .Z(_2294_)
  );
  AND2_X1 _7586_ (
    .A1(_2217_),
    .A2(_2294_),
    .ZN(_2295_)
  );
  XOR2_X1 _7587_ (
    .A(_2217_),
    .B(_2294_),
    .Z(_2296_)
  );
  AND2_X1 _7588_ (
    .A1(_2216_),
    .A2(_2296_),
    .ZN(_2297_)
  );
  XOR2_X1 _7589_ (
    .A(_2216_),
    .B(_2296_),
    .Z(_2298_)
  );
  AND2_X1 _7590_ (
    .A1(_2215_),
    .A2(_2298_),
    .ZN(_2299_)
  );
  XOR2_X1 _7591_ (
    .A(_2215_),
    .B(_2298_),
    .Z(_2300_)
  );
  AND2_X1 _7592_ (
    .A1(_2185_),
    .A2(_2300_),
    .ZN(_2301_)
  );
  INV_X1 _7593_ (
    .A(_2301_),
    .ZN(_2302_)
  );
  OR2_X1 _7594_ (
    .A1(_2185_),
    .A2(_2300_),
    .ZN(_2303_)
  );
  INV_X1 _7595_ (
    .A(_2303_),
    .ZN(_2304_)
  );
  AND2_X1 _7596_ (
    .A1(_2302_),
    .A2(_2303_),
    .ZN(_2305_)
  );
  OR2_X1 _7597_ (
    .A1(_2301_),
    .A2(_2304_),
    .ZN(_2306_)
  );
  AND2_X1 _7598_ (
    .A1(_2214_),
    .A2(_2305_),
    .ZN(_2307_)
  );
  XOR2_X1 _7599_ (
    .A(_2214_),
    .B(_2305_),
    .Z(_2308_)
  );
  XOR2_X1 _7600_ (
    .A(_2214_),
    .B(_2306_),
    .Z(_2309_)
  );
  OR2_X1 _7601_ (
    .A1(_2980_),
    .A2(_2309_),
    .ZN(_2310_)
  );
  INV_X1 _7602_ (
    .A(_2310_),
    .ZN(_2311_)
  );
  OR2_X1 _7603_ (
    .A1(remainder[60]),
    .A2(_2308_),
    .ZN(_2312_)
  );
  INV_X1 _7604_ (
    .A(_2312_),
    .ZN(_2313_)
  );
  AND2_X1 _7605_ (
    .A1(_2310_),
    .A2(_2312_),
    .ZN(_2314_)
  );
  XOR2_X1 _7606_ (
    .A(_2213_),
    .B(_2314_),
    .Z(_2315_)
  );
  AND2_X1 _7607_ (
    .A1(_4613_),
    .A2(_2315_),
    .ZN(_2316_)
  );
  AND2_X1 _7608_ (
    .A1(remainder[52]),
    .A2(_4610_),
    .ZN(_2317_)
  );
  OR2_X1 _7609_ (
    .A1(remainder[51]),
    .A2(_4393_),
    .ZN(_2318_)
  );
  OR2_X1 _7610_ (
    .A1(_4392_),
    .A2(_4534_),
    .ZN(_2319_)
  );
  AND2_X1 _7611_ (
    .A1(_3678_),
    .A2(_2319_),
    .ZN(_2320_)
  );
  AND2_X1 _7612_ (
    .A1(_2318_),
    .A2(_2320_),
    .ZN(_2321_)
  );
  OR2_X1 _7613_ (
    .A1(_2316_),
    .A2(_2321_),
    .ZN(_2322_)
  );
  OR2_X1 _7614_ (
    .A1(_2317_),
    .A2(_2322_),
    .ZN(_2323_)
  );
  AND2_X1 _7615_ (
    .A1(_3911_),
    .A2(_2323_),
    .ZN(_0073_)
  );
  OR2_X1 _7616_ (
    .A1(_2295_),
    .A2(_2297_),
    .ZN(_2324_)
  );
  OR2_X1 _7617_ (
    .A1(_2289_),
    .A2(_2291_),
    .ZN(_2325_)
  );
  OR2_X1 _7618_ (
    .A1(_2278_),
    .A2(_2293_),
    .ZN(_2326_)
  );
  AND2_X1 _7619_ (
    .A1(_0541_),
    .A2(_2153_),
    .ZN(_2327_)
  );
  AND2_X1 _7620_ (
    .A1(_2274_),
    .A2(_2327_),
    .ZN(_2328_)
  );
  OR2_X1 _7621_ (
    .A1(_2276_),
    .A2(_2328_),
    .ZN(_2329_)
  );
  AND2_X1 _7622_ (
    .A1(_0541_),
    .A2(_2273_),
    .ZN(_2330_)
  );
  OR2_X1 _7623_ (
    .A1(_2246_),
    .A2(_2248_),
    .ZN(_2331_)
  );
  AND2_X1 _7624_ (
    .A1(divisor[25]),
    .A2(remainder[3]),
    .ZN(_2332_)
  );
  AND2_X1 _7625_ (
    .A1(divisor[26]),
    .A2(remainder[2]),
    .ZN(_2333_)
  );
  AND2_X1 _7626_ (
    .A1(divisor[27]),
    .A2(remainder[2]),
    .ZN(_2334_)
  );
  AND2_X1 _7627_ (
    .A1(_2128_),
    .A2(_2334_),
    .ZN(_2335_)
  );
  XOR2_X1 _7628_ (
    .A(_2245_),
    .B(_2333_),
    .Z(_2336_)
  );
  AND2_X1 _7629_ (
    .A1(_2332_),
    .A2(_2336_),
    .ZN(_2337_)
  );
  XOR2_X1 _7630_ (
    .A(_2332_),
    .B(_2336_),
    .Z(_2338_)
  );
  AND2_X1 _7631_ (
    .A1(_2331_),
    .A2(_2338_),
    .ZN(_2339_)
  );
  XOR2_X1 _7632_ (
    .A(_2331_),
    .B(_2338_),
    .Z(_2340_)
  );
  AND2_X1 _7633_ (
    .A1(_2250_),
    .A2(_2340_),
    .ZN(_2341_)
  );
  XOR2_X1 _7634_ (
    .A(_2250_),
    .B(_2340_),
    .Z(_2342_)
  );
  OR2_X1 _7635_ (
    .A1(_2256_),
    .A2(_2258_),
    .ZN(_2343_)
  );
  AND2_X1 _7636_ (
    .A1(divisor[22]),
    .A2(remainder[6]),
    .ZN(_2344_)
  );
  AND2_X1 _7637_ (
    .A1(divisor[23]),
    .A2(remainder[5]),
    .ZN(_2345_)
  );
  AND2_X1 _7638_ (
    .A1(divisor[24]),
    .A2(remainder[5]),
    .ZN(_2346_)
  );
  AND2_X1 _7639_ (
    .A1(_2255_),
    .A2(_2345_),
    .ZN(_2347_)
  );
  XOR2_X1 _7640_ (
    .A(_2255_),
    .B(_2345_),
    .Z(_2348_)
  );
  AND2_X1 _7641_ (
    .A1(_2344_),
    .A2(_2348_),
    .ZN(_2349_)
  );
  XOR2_X1 _7642_ (
    .A(_2344_),
    .B(_2348_),
    .Z(_2350_)
  );
  AND2_X1 _7643_ (
    .A1(_2343_),
    .A2(_2350_),
    .ZN(_2351_)
  );
  XOR2_X1 _7644_ (
    .A(_2343_),
    .B(_2350_),
    .Z(_2352_)
  );
  AND2_X1 _7645_ (
    .A1(remainder[32]),
    .A2(divisor[21]),
    .ZN(_2353_)
  );
  AND2_X1 _7646_ (
    .A1(remainder[32]),
    .A2(divisor[20]),
    .ZN(_2354_)
  );
  AND2_X1 _7647_ (
    .A1(divisor[21]),
    .A2(_2354_),
    .ZN(_2355_)
  );
  AND2_X1 _7648_ (
    .A1(_2263_),
    .A2(_2354_),
    .ZN(_2356_)
  );
  XOR2_X1 _7649_ (
    .A(_2263_),
    .B(_2354_),
    .Z(_2357_)
  );
  AND2_X1 _7650_ (
    .A1(_1337_),
    .A2(_2357_),
    .ZN(_2358_)
  );
  XOR2_X1 _7651_ (
    .A(_1337_),
    .B(_2357_),
    .Z(_2359_)
  );
  AND2_X1 _7652_ (
    .A1(_2352_),
    .A2(_2359_),
    .ZN(_2360_)
  );
  XOR2_X1 _7653_ (
    .A(_2352_),
    .B(_2359_),
    .Z(_2361_)
  );
  AND2_X1 _7654_ (
    .A1(_2342_),
    .A2(_2361_),
    .ZN(_2362_)
  );
  XOR2_X1 _7655_ (
    .A(_2342_),
    .B(_2361_),
    .Z(_2363_)
  );
  AND2_X1 _7656_ (
    .A1(_2270_),
    .A2(_2363_),
    .ZN(_2364_)
  );
  XOR2_X1 _7657_ (
    .A(_2270_),
    .B(_2363_),
    .Z(_2365_)
  );
  AND2_X1 _7658_ (
    .A1(divisor[28]),
    .A2(remainder[0]),
    .ZN(_2366_)
  );
  AND2_X1 _7659_ (
    .A1(remainder[32]),
    .A2(divisor[28]),
    .ZN(_2367_)
  );
  AND2_X1 _7660_ (
    .A1(_0541_),
    .A2(_2366_),
    .ZN(_2368_)
  );
  OR2_X1 _7661_ (
    .A1(_0542_),
    .A2(_2368_),
    .ZN(_2369_)
  );
  XOR2_X1 _7662_ (
    .A(_0541_),
    .B(_2366_),
    .Z(_2370_)
  );
  AND2_X1 _7663_ (
    .A1(_2365_),
    .A2(_2370_),
    .ZN(_2371_)
  );
  XOR2_X1 _7664_ (
    .A(_2365_),
    .B(_2370_),
    .Z(_2372_)
  );
  AND2_X1 _7665_ (
    .A1(_2330_),
    .A2(_2372_),
    .ZN(_2373_)
  );
  XOR2_X1 _7666_ (
    .A(_2330_),
    .B(_2372_),
    .Z(_2374_)
  );
  OR2_X1 _7667_ (
    .A1(_2235_),
    .A2(_2237_),
    .ZN(_2375_)
  );
  OR2_X1 _7668_ (
    .A1(_2231_),
    .A2(_2233_),
    .ZN(_2376_)
  );
  OR2_X1 _7669_ (
    .A1(_2227_),
    .A2(_2229_),
    .ZN(_2377_)
  );
  OR2_X1 _7670_ (
    .A1(_2260_),
    .A2(_2268_),
    .ZN(_2378_)
  );
  OR2_X1 _7671_ (
    .A1(_2264_),
    .A2(_2266_),
    .ZN(_2379_)
  );
  AND2_X1 _7672_ (
    .A1(_2111_),
    .A2(_2379_),
    .ZN(_2380_)
  );
  XOR2_X1 _7673_ (
    .A(_2111_),
    .B(_2379_),
    .Z(_2381_)
  );
  AND2_X1 _7674_ (
    .A1(_2225_),
    .A2(_2381_),
    .ZN(_2382_)
  );
  XOR2_X1 _7675_ (
    .A(_2225_),
    .B(_2381_),
    .Z(_2383_)
  );
  AND2_X1 _7676_ (
    .A1(_2378_),
    .A2(_2383_),
    .ZN(_2384_)
  );
  XOR2_X1 _7677_ (
    .A(_2378_),
    .B(_2383_),
    .Z(_2385_)
  );
  AND2_X1 _7678_ (
    .A1(_2377_),
    .A2(_2385_),
    .ZN(_2386_)
  );
  XOR2_X1 _7679_ (
    .A(_2377_),
    .B(_2385_),
    .Z(_2387_)
  );
  AND2_X1 _7680_ (
    .A1(_2376_),
    .A2(_2387_),
    .ZN(_2388_)
  );
  XOR2_X1 _7681_ (
    .A(_2376_),
    .B(_2387_),
    .Z(_2389_)
  );
  AND2_X1 _7682_ (
    .A1(_2025_),
    .A2(_2389_),
    .ZN(_2390_)
  );
  XOR2_X1 _7683_ (
    .A(_2025_),
    .B(_2389_),
    .Z(_2391_)
  );
  AND2_X1 _7684_ (
    .A1(_2272_),
    .A2(_2391_),
    .ZN(_2392_)
  );
  XOR2_X1 _7685_ (
    .A(_2272_),
    .B(_2391_),
    .Z(_2393_)
  );
  AND2_X1 _7686_ (
    .A1(_2375_),
    .A2(_2393_),
    .ZN(_2394_)
  );
  XOR2_X1 _7687_ (
    .A(_2375_),
    .B(_2393_),
    .Z(_2395_)
  );
  AND2_X1 _7688_ (
    .A1(_2374_),
    .A2(_2395_),
    .ZN(_2396_)
  );
  XOR2_X1 _7689_ (
    .A(_2374_),
    .B(_2395_),
    .Z(_2397_)
  );
  AND2_X1 _7690_ (
    .A1(_2329_),
    .A2(_2397_),
    .ZN(_2398_)
  );
  XOR2_X1 _7691_ (
    .A(_2329_),
    .B(_2397_),
    .Z(_2399_)
  );
  AND2_X1 _7692_ (
    .A1(_2170_),
    .A2(_2285_),
    .ZN(_2400_)
  );
  INV_X1 _7693_ (
    .A(_2400_),
    .ZN(_2401_)
  );
  OR2_X1 _7694_ (
    .A1(_2239_),
    .A2(_2241_),
    .ZN(_2402_)
  );
  AND2_X1 _7695_ (
    .A1(_2287_),
    .A2(_2402_),
    .ZN(_2403_)
  );
  XOR2_X1 _7696_ (
    .A(_2288_),
    .B(_2402_),
    .Z(_2404_)
  );
  OR2_X1 _7697_ (
    .A1(_2400_),
    .A2(_2404_),
    .ZN(_2405_)
  );
  INV_X1 _7698_ (
    .A(_2405_),
    .ZN(_2406_)
  );
  XOR2_X1 _7699_ (
    .A(_2400_),
    .B(_2404_),
    .Z(_2407_)
  );
  AND2_X1 _7700_ (
    .A1(_2399_),
    .A2(_2407_),
    .ZN(_2408_)
  );
  XOR2_X1 _7701_ (
    .A(_2399_),
    .B(_2407_),
    .Z(_2409_)
  );
  AND2_X1 _7702_ (
    .A1(_2326_),
    .A2(_2409_),
    .ZN(_2410_)
  );
  XOR2_X1 _7703_ (
    .A(_2326_),
    .B(_2409_),
    .Z(_2411_)
  );
  AND2_X1 _7704_ (
    .A1(_2325_),
    .A2(_2411_),
    .ZN(_2412_)
  );
  XOR2_X1 _7705_ (
    .A(_2325_),
    .B(_2411_),
    .Z(_2413_)
  );
  AND2_X1 _7706_ (
    .A1(_2324_),
    .A2(_2413_),
    .ZN(_2414_)
  );
  XOR2_X1 _7707_ (
    .A(_2324_),
    .B(_2413_),
    .Z(_2415_)
  );
  AND2_X1 _7708_ (
    .A1(_2299_),
    .A2(_2415_),
    .ZN(_2416_)
  );
  XOR2_X1 _7709_ (
    .A(_2299_),
    .B(_2415_),
    .Z(_2417_)
  );
  INV_X1 _7710_ (
    .A(_2417_),
    .ZN(_2418_)
  );
  OR2_X1 _7711_ (
    .A1(_2301_),
    .A2(_2307_),
    .ZN(_2419_)
  );
  AND2_X1 _7712_ (
    .A1(_2417_),
    .A2(_2419_),
    .ZN(_2420_)
  );
  XOR2_X1 _7713_ (
    .A(_2417_),
    .B(_2419_),
    .Z(_2421_)
  );
  XOR2_X1 _7714_ (
    .A(_2418_),
    .B(_2419_),
    .Z(_2422_)
  );
  AND2_X1 _7715_ (
    .A1(remainder[61]),
    .A2(_2421_),
    .ZN(_2423_)
  );
  OR2_X1 _7716_ (
    .A1(_2969_),
    .A2(_2422_),
    .ZN(_2424_)
  );
  XOR2_X1 _7717_ (
    .A(remainder[61]),
    .B(_2421_),
    .Z(_2425_)
  );
  INV_X1 _7718_ (
    .A(_2425_),
    .ZN(_2426_)
  );
  AND2_X1 _7719_ (
    .A1(_2212_),
    .A2(_2310_),
    .ZN(_2427_)
  );
  OR2_X1 _7720_ (
    .A1(_2213_),
    .A2(_2311_),
    .ZN(_2428_)
  );
  AND2_X1 _7721_ (
    .A1(_2312_),
    .A2(_2428_),
    .ZN(_2429_)
  );
  OR2_X1 _7722_ (
    .A1(_2313_),
    .A2(_2427_),
    .ZN(_2430_)
  );
  AND2_X1 _7723_ (
    .A1(_2425_),
    .A2(_2429_),
    .ZN(_2431_)
  );
  OR2_X1 _7724_ (
    .A1(_2426_),
    .A2(_2430_),
    .ZN(_2432_)
  );
  XOR2_X1 _7725_ (
    .A(_2425_),
    .B(_2429_),
    .Z(_2433_)
  );
  AND2_X1 _7726_ (
    .A1(_4613_),
    .A2(_2433_),
    .ZN(_2434_)
  );
  AND2_X1 _7727_ (
    .A1(remainder[53]),
    .A2(_4610_),
    .ZN(_2435_)
  );
  OR2_X1 _7728_ (
    .A1(_4392_),
    .A2(_4539_),
    .ZN(_2436_)
  );
  OR2_X1 _7729_ (
    .A1(remainder[52]),
    .A2(_4393_),
    .ZN(_2437_)
  );
  AND2_X1 _7730_ (
    .A1(_3678_),
    .A2(_2436_),
    .ZN(_2438_)
  );
  AND2_X1 _7731_ (
    .A1(_2437_),
    .A2(_2438_),
    .ZN(_2439_)
  );
  OR2_X1 _7732_ (
    .A1(_2434_),
    .A2(_2439_),
    .ZN(_2440_)
  );
  OR2_X1 _7733_ (
    .A1(_2435_),
    .A2(_2440_),
    .ZN(_2441_)
  );
  AND2_X1 _7734_ (
    .A1(_3911_),
    .A2(_2441_),
    .ZN(_0074_)
  );
  AND2_X1 _7735_ (
    .A1(_2424_),
    .A2(_2432_),
    .ZN(_2442_)
  );
  OR2_X1 _7736_ (
    .A1(_2423_),
    .A2(_2431_),
    .ZN(_2443_)
  );
  OR2_X1 _7737_ (
    .A1(_2416_),
    .A2(_2420_),
    .ZN(_2444_)
  );
  INV_X1 _7738_ (
    .A(_2444_),
    .ZN(_2445_)
  );
  OR2_X1 _7739_ (
    .A1(_2410_),
    .A2(_2412_),
    .ZN(_2446_)
  );
  OR2_X1 _7740_ (
    .A1(_2403_),
    .A2(_2406_),
    .ZN(_2447_)
  );
  OR2_X1 _7741_ (
    .A1(_2398_),
    .A2(_2408_),
    .ZN(_2448_)
  );
  OR2_X1 _7742_ (
    .A1(_2373_),
    .A2(_2396_),
    .ZN(_2449_)
  );
  OR2_X1 _7743_ (
    .A1(_2341_),
    .A2(_2362_),
    .ZN(_2450_)
  );
  OR2_X1 _7744_ (
    .A1(_2335_),
    .A2(_2337_),
    .ZN(_2451_)
  );
  AND2_X1 _7745_ (
    .A1(divisor[25]),
    .A2(remainder[4]),
    .ZN(_2452_)
  );
  AND2_X1 _7746_ (
    .A1(divisor[26]),
    .A2(remainder[3]),
    .ZN(_2453_)
  );
  AND2_X1 _7747_ (
    .A1(divisor[27]),
    .A2(remainder[3]),
    .ZN(_2454_)
  );
  AND2_X1 _7748_ (
    .A1(_2334_),
    .A2(_2453_),
    .ZN(_2455_)
  );
  XOR2_X1 _7749_ (
    .A(_2334_),
    .B(_2453_),
    .Z(_2456_)
  );
  AND2_X1 _7750_ (
    .A1(_2452_),
    .A2(_2456_),
    .ZN(_2457_)
  );
  XOR2_X1 _7751_ (
    .A(_2452_),
    .B(_2456_),
    .Z(_2458_)
  );
  AND2_X1 _7752_ (
    .A1(_2451_),
    .A2(_2458_),
    .ZN(_2459_)
  );
  XOR2_X1 _7753_ (
    .A(_2451_),
    .B(_2458_),
    .Z(_2460_)
  );
  AND2_X1 _7754_ (
    .A1(_2339_),
    .A2(_2460_),
    .ZN(_2461_)
  );
  XOR2_X1 _7755_ (
    .A(_2339_),
    .B(_2460_),
    .Z(_2462_)
  );
  OR2_X1 _7756_ (
    .A1(_2347_),
    .A2(_2349_),
    .ZN(_2463_)
  );
  AND2_X1 _7757_ (
    .A1(divisor[22]),
    .A2(remainder[7]),
    .ZN(_2464_)
  );
  AND2_X1 _7758_ (
    .A1(divisor[23]),
    .A2(remainder[6]),
    .ZN(_2465_)
  );
  AND2_X1 _7759_ (
    .A1(divisor[24]),
    .A2(remainder[6]),
    .ZN(_2466_)
  );
  AND2_X1 _7760_ (
    .A1(_2346_),
    .A2(_2465_),
    .ZN(_2467_)
  );
  XOR2_X1 _7761_ (
    .A(_2346_),
    .B(_2465_),
    .Z(_2468_)
  );
  AND2_X1 _7762_ (
    .A1(_2464_),
    .A2(_2468_),
    .ZN(_2469_)
  );
  XOR2_X1 _7763_ (
    .A(_2464_),
    .B(_2468_),
    .Z(_2470_)
  );
  AND2_X1 _7764_ (
    .A1(_2463_),
    .A2(_2470_),
    .ZN(_2471_)
  );
  XOR2_X1 _7765_ (
    .A(_2463_),
    .B(_2470_),
    .Z(_2472_)
  );
  MUX2_X1 _7766_ (
    .A(_2354_),
    .B(_3373_),
    .S(_2353_),
    .Z(_2473_)
  );
  AND2_X1 _7767_ (
    .A1(divisor[19]),
    .A2(_2473_),
    .ZN(_2474_)
  );
  MUX2_X1 _7768_ (
    .A(_1337_),
    .B(_3362_),
    .S(_2473_),
    .Z(_2475_)
  );
  INV_X1 _7769_ (
    .A(_2475_),
    .ZN(_2476_)
  );
  AND2_X1 _7770_ (
    .A1(_2472_),
    .A2(_2475_),
    .ZN(_2477_)
  );
  XOR2_X1 _7771_ (
    .A(_2472_),
    .B(_2475_),
    .Z(_2478_)
  );
  AND2_X1 _7772_ (
    .A1(_2462_),
    .A2(_2478_),
    .ZN(_2479_)
  );
  XOR2_X1 _7773_ (
    .A(_2462_),
    .B(_2478_),
    .Z(_2480_)
  );
  AND2_X1 _7774_ (
    .A1(_2450_),
    .A2(_2480_),
    .ZN(_2481_)
  );
  XOR2_X1 _7775_ (
    .A(_2450_),
    .B(_2480_),
    .Z(_2482_)
  );
  AND2_X1 _7776_ (
    .A1(divisor[29]),
    .A2(remainder[0]),
    .ZN(_2483_)
  );
  AND2_X1 _7777_ (
    .A1(divisor[28]),
    .A2(remainder[1]),
    .ZN(_2484_)
  );
  AND2_X1 _7778_ (
    .A1(divisor[29]),
    .A2(remainder[1]),
    .ZN(_2485_)
  );
  AND2_X1 _7779_ (
    .A1(_2366_),
    .A2(_2485_),
    .ZN(_2486_)
  );
  XOR2_X1 _7780_ (
    .A(_2483_),
    .B(_2484_),
    .Z(_2487_)
  );
  INV_X1 _7781_ (
    .A(_2487_),
    .ZN(_2488_)
  );
  XOR2_X1 _7782_ (
    .A(_2369_),
    .B(_2488_),
    .Z(_2489_)
  );
  AND2_X1 _7783_ (
    .A1(_2482_),
    .A2(_2489_),
    .ZN(_2490_)
  );
  XOR2_X1 _7784_ (
    .A(_2482_),
    .B(_2489_),
    .Z(_2491_)
  );
  AND2_X1 _7785_ (
    .A1(_2371_),
    .A2(_2491_),
    .ZN(_2492_)
  );
  XOR2_X1 _7786_ (
    .A(_2371_),
    .B(_2491_),
    .Z(_2493_)
  );
  OR2_X1 _7787_ (
    .A1(_2388_),
    .A2(_2390_),
    .ZN(_2494_)
  );
  OR2_X1 _7788_ (
    .A1(_2384_),
    .A2(_2386_),
    .ZN(_2495_)
  );
  OR2_X1 _7789_ (
    .A1(_2380_),
    .A2(_2382_),
    .ZN(_2496_)
  );
  OR2_X1 _7790_ (
    .A1(_2351_),
    .A2(_2360_),
    .ZN(_2497_)
  );
  OR2_X1 _7791_ (
    .A1(_2356_),
    .A2(_2358_),
    .ZN(_2498_)
  );
  AND2_X1 _7792_ (
    .A1(_2111_),
    .A2(_2498_),
    .ZN(_2499_)
  );
  XOR2_X1 _7793_ (
    .A(_2111_),
    .B(_2498_),
    .Z(_2500_)
  );
  AND2_X1 _7794_ (
    .A1(_2225_),
    .A2(_2500_),
    .ZN(_2501_)
  );
  XOR2_X1 _7795_ (
    .A(_2225_),
    .B(_2500_),
    .Z(_2502_)
  );
  AND2_X1 _7796_ (
    .A1(_2497_),
    .A2(_2502_),
    .ZN(_2503_)
  );
  XOR2_X1 _7797_ (
    .A(_2497_),
    .B(_2502_),
    .Z(_2504_)
  );
  AND2_X1 _7798_ (
    .A1(_2496_),
    .A2(_2504_),
    .ZN(_2505_)
  );
  XOR2_X1 _7799_ (
    .A(_2496_),
    .B(_2504_),
    .Z(_2506_)
  );
  AND2_X1 _7800_ (
    .A1(_2495_),
    .A2(_2506_),
    .ZN(_2507_)
  );
  XOR2_X1 _7801_ (
    .A(_2495_),
    .B(_2506_),
    .Z(_2508_)
  );
  AND2_X1 _7802_ (
    .A1(_2025_),
    .A2(_2508_),
    .ZN(_2509_)
  );
  XOR2_X1 _7803_ (
    .A(_2025_),
    .B(_2508_),
    .Z(_2510_)
  );
  AND2_X1 _7804_ (
    .A1(_2364_),
    .A2(_2510_),
    .ZN(_2511_)
  );
  XOR2_X1 _7805_ (
    .A(_2364_),
    .B(_2510_),
    .Z(_2512_)
  );
  AND2_X1 _7806_ (
    .A1(_2494_),
    .A2(_2512_),
    .ZN(_2513_)
  );
  XOR2_X1 _7807_ (
    .A(_2494_),
    .B(_2512_),
    .Z(_2514_)
  );
  AND2_X1 _7808_ (
    .A1(_2493_),
    .A2(_2514_),
    .ZN(_2515_)
  );
  XOR2_X1 _7809_ (
    .A(_2493_),
    .B(_2514_),
    .Z(_2516_)
  );
  AND2_X1 _7810_ (
    .A1(_2449_),
    .A2(_2516_),
    .ZN(_2517_)
  );
  XOR2_X1 _7811_ (
    .A(_2449_),
    .B(_2516_),
    .Z(_2518_)
  );
  OR2_X1 _7812_ (
    .A1(_2392_),
    .A2(_2394_),
    .ZN(_2519_)
  );
  AND2_X1 _7813_ (
    .A1(_2287_),
    .A2(_2519_),
    .ZN(_2520_)
  );
  XOR2_X1 _7814_ (
    .A(_2288_),
    .B(_2519_),
    .Z(_2521_)
  );
  OR2_X1 _7815_ (
    .A1(_2400_),
    .A2(_2521_),
    .ZN(_2522_)
  );
  INV_X1 _7816_ (
    .A(_2522_),
    .ZN(_2523_)
  );
  XOR2_X1 _7817_ (
    .A(_2400_),
    .B(_2521_),
    .Z(_2524_)
  );
  AND2_X1 _7818_ (
    .A1(_2518_),
    .A2(_2524_),
    .ZN(_2525_)
  );
  XOR2_X1 _7819_ (
    .A(_2518_),
    .B(_2524_),
    .Z(_2526_)
  );
  AND2_X1 _7820_ (
    .A1(_2448_),
    .A2(_2526_),
    .ZN(_2527_)
  );
  XOR2_X1 _7821_ (
    .A(_2448_),
    .B(_2526_),
    .Z(_2528_)
  );
  AND2_X1 _7822_ (
    .A1(_2447_),
    .A2(_2528_),
    .ZN(_2529_)
  );
  XOR2_X1 _7823_ (
    .A(_2447_),
    .B(_2528_),
    .Z(_2530_)
  );
  AND2_X1 _7824_ (
    .A1(_2446_),
    .A2(_2530_),
    .ZN(_2531_)
  );
  XOR2_X1 _7825_ (
    .A(_2446_),
    .B(_2530_),
    .Z(_2532_)
  );
  AND2_X1 _7826_ (
    .A1(_2414_),
    .A2(_2532_),
    .ZN(_2533_)
  );
  OR2_X1 _7827_ (
    .A1(_2414_),
    .A2(_2532_),
    .ZN(_2534_)
  );
  XOR2_X1 _7828_ (
    .A(_2414_),
    .B(_2532_),
    .Z(_2535_)
  );
  XOR2_X1 _7829_ (
    .A(_2445_),
    .B(_2535_),
    .Z(_2536_)
  );
  XOR2_X1 _7830_ (
    .A(_2444_),
    .B(_2535_),
    .Z(_2537_)
  );
  AND2_X1 _7831_ (
    .A1(remainder[62]),
    .A2(_2537_),
    .ZN(_2538_)
  );
  INV_X1 _7832_ (
    .A(_2538_),
    .ZN(_2539_)
  );
  AND2_X1 _7833_ (
    .A1(_2958_),
    .A2(_2536_),
    .ZN(_2540_)
  );
  INV_X1 _7834_ (
    .A(_2540_),
    .ZN(_2541_)
  );
  OR2_X1 _7835_ (
    .A1(_2538_),
    .A2(_2540_),
    .ZN(_2542_)
  );
  XOR2_X1 _7836_ (
    .A(_2443_),
    .B(_2542_),
    .Z(_2543_)
  );
  INV_X1 _7837_ (
    .A(_2543_),
    .ZN(_2544_)
  );
  AND2_X1 _7838_ (
    .A1(_4613_),
    .A2(_2544_),
    .ZN(_2545_)
  );
  AND2_X1 _7839_ (
    .A1(remainder[54]),
    .A2(_4610_),
    .ZN(_2546_)
  );
  OR2_X1 _7840_ (
    .A1(_4392_),
    .A2(_4545_),
    .ZN(_2547_)
  );
  OR2_X1 _7841_ (
    .A1(remainder[53]),
    .A2(_4393_),
    .ZN(_2548_)
  );
  AND2_X1 _7842_ (
    .A1(_3678_),
    .A2(_2547_),
    .ZN(_2549_)
  );
  AND2_X1 _7843_ (
    .A1(_2548_),
    .A2(_2549_),
    .ZN(_2550_)
  );
  OR2_X1 _7844_ (
    .A1(_2545_),
    .A2(_2550_),
    .ZN(_2551_)
  );
  OR2_X1 _7845_ (
    .A1(_2546_),
    .A2(_2551_),
    .ZN(_2552_)
  );
  AND2_X1 _7846_ (
    .A1(_3911_),
    .A2(_2552_),
    .ZN(_0075_)
  );
  OR2_X1 _7847_ (
    .A1(_2527_),
    .A2(_2529_),
    .ZN(_2553_)
  );
  OR2_X1 _7848_ (
    .A1(_2520_),
    .A2(_2523_),
    .ZN(_2554_)
  );
  OR2_X1 _7849_ (
    .A1(_2517_),
    .A2(_2525_),
    .ZN(_2555_)
  );
  OR2_X1 _7850_ (
    .A1(_2492_),
    .A2(_2515_),
    .ZN(_2556_)
  );
  AND2_X1 _7851_ (
    .A1(_2368_),
    .A2(_2488_),
    .ZN(_2557_)
  );
  OR2_X1 _7852_ (
    .A1(_2490_),
    .A2(_2557_),
    .ZN(_2558_)
  );
  OR2_X1 _7853_ (
    .A1(_2461_),
    .A2(_2479_),
    .ZN(_2559_)
  );
  OR2_X1 _7854_ (
    .A1(_2455_),
    .A2(_2457_),
    .ZN(_2560_)
  );
  AND2_X1 _7855_ (
    .A1(divisor[25]),
    .A2(remainder[5]),
    .ZN(_2561_)
  );
  AND2_X1 _7856_ (
    .A1(divisor[26]),
    .A2(remainder[4]),
    .ZN(_2562_)
  );
  AND2_X1 _7857_ (
    .A1(divisor[27]),
    .A2(remainder[4]),
    .ZN(_2563_)
  );
  AND2_X1 _7858_ (
    .A1(_2454_),
    .A2(_2562_),
    .ZN(_2564_)
  );
  XOR2_X1 _7859_ (
    .A(_2454_),
    .B(_2562_),
    .Z(_2565_)
  );
  AND2_X1 _7860_ (
    .A1(_2561_),
    .A2(_2565_),
    .ZN(_2566_)
  );
  XOR2_X1 _7861_ (
    .A(_2561_),
    .B(_2565_),
    .Z(_2567_)
  );
  AND2_X1 _7862_ (
    .A1(_2486_),
    .A2(_2567_),
    .ZN(_2568_)
  );
  XOR2_X1 _7863_ (
    .A(_2486_),
    .B(_2567_),
    .Z(_2569_)
  );
  AND2_X1 _7864_ (
    .A1(_2560_),
    .A2(_2569_),
    .ZN(_2570_)
  );
  XOR2_X1 _7865_ (
    .A(_2560_),
    .B(_2569_),
    .Z(_2571_)
  );
  AND2_X1 _7866_ (
    .A1(_2459_),
    .A2(_2571_),
    .ZN(_2572_)
  );
  XOR2_X1 _7867_ (
    .A(_2459_),
    .B(_2571_),
    .Z(_2573_)
  );
  OR2_X1 _7868_ (
    .A1(_2467_),
    .A2(_2469_),
    .ZN(_2574_)
  );
  AND2_X1 _7869_ (
    .A1(remainder[32]),
    .A2(divisor[22]),
    .ZN(_2575_)
  );
  INV_X1 _7870_ (
    .A(_2575_),
    .ZN(_2576_)
  );
  AND2_X1 _7871_ (
    .A1(divisor[23]),
    .A2(remainder[7]),
    .ZN(_2577_)
  );
  AND2_X1 _7872_ (
    .A1(divisor[24]),
    .A2(remainder[7]),
    .ZN(_2578_)
  );
  AND2_X1 _7873_ (
    .A1(_2465_),
    .A2(_2578_),
    .ZN(_2579_)
  );
  XOR2_X1 _7874_ (
    .A(_2466_),
    .B(_2577_),
    .Z(_2580_)
  );
  AND2_X1 _7875_ (
    .A1(_2575_),
    .A2(_2580_),
    .ZN(_2581_)
  );
  XOR2_X1 _7876_ (
    .A(_2575_),
    .B(_2580_),
    .Z(_2582_)
  );
  AND2_X1 _7877_ (
    .A1(_2574_),
    .A2(_2582_),
    .ZN(_2583_)
  );
  XOR2_X1 _7878_ (
    .A(_2574_),
    .B(_2582_),
    .Z(_2584_)
  );
  AND2_X1 _7879_ (
    .A1(_2475_),
    .A2(_2584_),
    .ZN(_2585_)
  );
  XOR2_X1 _7880_ (
    .A(_2475_),
    .B(_2584_),
    .Z(_2586_)
  );
  AND2_X1 _7881_ (
    .A1(_2573_),
    .A2(_2586_),
    .ZN(_2587_)
  );
  XOR2_X1 _7882_ (
    .A(_2573_),
    .B(_2586_),
    .Z(_2588_)
  );
  AND2_X1 _7883_ (
    .A1(_2559_),
    .A2(_2588_),
    .ZN(_2589_)
  );
  XOR2_X1 _7884_ (
    .A(_2559_),
    .B(_2588_),
    .Z(_2590_)
  );
  AND2_X1 _7885_ (
    .A1(divisor[28]),
    .A2(remainder[2]),
    .ZN(_2591_)
  );
  AND2_X1 _7886_ (
    .A1(divisor[30]),
    .A2(remainder[0]),
    .ZN(_2592_)
  );
  AND2_X1 _7887_ (
    .A1(divisor[30]),
    .A2(remainder[1]),
    .ZN(_2593_)
  );
  AND2_X1 _7888_ (
    .A1(_2483_),
    .A2(_2593_),
    .ZN(_2594_)
  );
  XOR2_X1 _7889_ (
    .A(_2485_),
    .B(_2592_),
    .Z(_2595_)
  );
  AND2_X1 _7890_ (
    .A1(_2591_),
    .A2(_2595_),
    .ZN(_2596_)
  );
  XOR2_X1 _7891_ (
    .A(_2591_),
    .B(_2595_),
    .Z(_2597_)
  );
  INV_X1 _7892_ (
    .A(_2597_),
    .ZN(_2598_)
  );
  AND2_X1 _7893_ (
    .A1(_0541_),
    .A2(_2488_),
    .ZN(_2599_)
  );
  XOR2_X1 _7894_ (
    .A(_2597_),
    .B(_2599_),
    .Z(_2600_)
  );
  AND2_X1 _7895_ (
    .A1(_2590_),
    .A2(_2600_),
    .ZN(_2601_)
  );
  XOR2_X1 _7896_ (
    .A(_2590_),
    .B(_2600_),
    .Z(_2602_)
  );
  AND2_X1 _7897_ (
    .A1(_2558_),
    .A2(_2602_),
    .ZN(_2603_)
  );
  XOR2_X1 _7898_ (
    .A(_2558_),
    .B(_2602_),
    .Z(_2604_)
  );
  OR2_X1 _7899_ (
    .A1(_2507_),
    .A2(_2509_),
    .ZN(_2605_)
  );
  OR2_X1 _7900_ (
    .A1(_2503_),
    .A2(_2505_),
    .ZN(_2606_)
  );
  OR2_X1 _7901_ (
    .A1(_2499_),
    .A2(_2501_),
    .ZN(_2607_)
  );
  OR2_X1 _7902_ (
    .A1(_2471_),
    .A2(_2477_),
    .ZN(_2608_)
  );
  OR2_X1 _7903_ (
    .A1(_2355_),
    .A2(_2474_),
    .ZN(_2609_)
  );
  AND2_X1 _7904_ (
    .A1(_2111_),
    .A2(_2609_),
    .ZN(_2610_)
  );
  XOR2_X1 _7905_ (
    .A(_2111_),
    .B(_2609_),
    .Z(_2611_)
  );
  AND2_X1 _7906_ (
    .A1(_2225_),
    .A2(_2611_),
    .ZN(_2612_)
  );
  XOR2_X1 _7907_ (
    .A(_2225_),
    .B(_2611_),
    .Z(_2613_)
  );
  INV_X1 _7908_ (
    .A(_2613_),
    .ZN(_2614_)
  );
  AND2_X1 _7909_ (
    .A1(_2608_),
    .A2(_2613_),
    .ZN(_2615_)
  );
  XOR2_X1 _7910_ (
    .A(_2608_),
    .B(_2613_),
    .Z(_2616_)
  );
  AND2_X1 _7911_ (
    .A1(_2607_),
    .A2(_2616_),
    .ZN(_2617_)
  );
  XOR2_X1 _7912_ (
    .A(_2607_),
    .B(_2616_),
    .Z(_2618_)
  );
  AND2_X1 _7913_ (
    .A1(_2606_),
    .A2(_2618_),
    .ZN(_2619_)
  );
  XOR2_X1 _7914_ (
    .A(_2606_),
    .B(_2618_),
    .Z(_2620_)
  );
  AND2_X1 _7915_ (
    .A1(_2025_),
    .A2(_2620_),
    .ZN(_2621_)
  );
  XOR2_X1 _7916_ (
    .A(_2025_),
    .B(_2620_),
    .Z(_2622_)
  );
  AND2_X1 _7917_ (
    .A1(_2481_),
    .A2(_2622_),
    .ZN(_2623_)
  );
  XOR2_X1 _7918_ (
    .A(_2481_),
    .B(_2622_),
    .Z(_2624_)
  );
  AND2_X1 _7919_ (
    .A1(_2605_),
    .A2(_2624_),
    .ZN(_2625_)
  );
  XOR2_X1 _7920_ (
    .A(_2605_),
    .B(_2624_),
    .Z(_2626_)
  );
  AND2_X1 _7921_ (
    .A1(_2604_),
    .A2(_2626_),
    .ZN(_2627_)
  );
  XOR2_X1 _7922_ (
    .A(_2604_),
    .B(_2626_),
    .Z(_2628_)
  );
  AND2_X1 _7923_ (
    .A1(_2556_),
    .A2(_2628_),
    .ZN(_2629_)
  );
  XOR2_X1 _7924_ (
    .A(_2556_),
    .B(_2628_),
    .Z(_2630_)
  );
  OR2_X1 _7925_ (
    .A1(_2511_),
    .A2(_2513_),
    .ZN(_2631_)
  );
  AND2_X1 _7926_ (
    .A1(_2287_),
    .A2(_2631_),
    .ZN(_2632_)
  );
  XOR2_X1 _7927_ (
    .A(_2288_),
    .B(_2631_),
    .Z(_2633_)
  );
  OR2_X1 _7928_ (
    .A1(_2400_),
    .A2(_2633_),
    .ZN(_2634_)
  );
  INV_X1 _7929_ (
    .A(_2634_),
    .ZN(_2635_)
  );
  XOR2_X1 _7930_ (
    .A(_2400_),
    .B(_2633_),
    .Z(_2636_)
  );
  AND2_X1 _7931_ (
    .A1(_2630_),
    .A2(_2636_),
    .ZN(_2637_)
  );
  XOR2_X1 _7932_ (
    .A(_2630_),
    .B(_2636_),
    .Z(_2638_)
  );
  AND2_X1 _7933_ (
    .A1(_2555_),
    .A2(_2638_),
    .ZN(_2639_)
  );
  XOR2_X1 _7934_ (
    .A(_2555_),
    .B(_2638_),
    .Z(_2640_)
  );
  AND2_X1 _7935_ (
    .A1(_2554_),
    .A2(_2640_),
    .ZN(_2641_)
  );
  XOR2_X1 _7936_ (
    .A(_2554_),
    .B(_2640_),
    .Z(_2642_)
  );
  AND2_X1 _7937_ (
    .A1(_2553_),
    .A2(_2642_),
    .ZN(_2643_)
  );
  XOR2_X1 _7938_ (
    .A(_2553_),
    .B(_2642_),
    .Z(_2644_)
  );
  AND2_X1 _7939_ (
    .A1(_2531_),
    .A2(_2644_),
    .ZN(_2645_)
  );
  XOR2_X1 _7940_ (
    .A(_2531_),
    .B(_2644_),
    .Z(_2646_)
  );
  AND2_X1 _7941_ (
    .A1(_2420_),
    .A2(_2535_),
    .ZN(_2647_)
  );
  AND2_X1 _7942_ (
    .A1(_2416_),
    .A2(_2534_),
    .ZN(_2648_)
  );
  OR2_X1 _7943_ (
    .A1(_2533_),
    .A2(_2648_),
    .ZN(_2649_)
  );
  OR2_X1 _7944_ (
    .A1(_2647_),
    .A2(_2649_),
    .ZN(_2650_)
  );
  AND2_X1 _7945_ (
    .A1(_2646_),
    .A2(_2650_),
    .ZN(_2651_)
  );
  XOR2_X1 _7946_ (
    .A(_2646_),
    .B(_2650_),
    .Z(_2652_)
  );
  AND2_X1 _7947_ (
    .A1(remainder[63]),
    .A2(_2652_),
    .ZN(_2653_)
  );
  INV_X1 _7948_ (
    .A(_2653_),
    .ZN(_2654_)
  );
  XOR2_X1 _7949_ (
    .A(remainder[63]),
    .B(_2652_),
    .Z(_2655_)
  );
  INV_X1 _7950_ (
    .A(_2655_),
    .ZN(_2656_)
  );
  AND2_X1 _7951_ (
    .A1(_2442_),
    .A2(_2539_),
    .ZN(_2657_)
  );
  OR2_X1 _7952_ (
    .A1(_2443_),
    .A2(_2538_),
    .ZN(_2658_)
  );
  AND2_X1 _7953_ (
    .A1(_2541_),
    .A2(_2658_),
    .ZN(_2659_)
  );
  OR2_X1 _7954_ (
    .A1(_2540_),
    .A2(_2657_),
    .ZN(_2660_)
  );
  AND2_X1 _7955_ (
    .A1(_2655_),
    .A2(_2659_),
    .ZN(_2661_)
  );
  OR2_X1 _7956_ (
    .A1(_2656_),
    .A2(_2660_),
    .ZN(_2662_)
  );
  OR2_X1 _7957_ (
    .A1(_2655_),
    .A2(_2659_),
    .ZN(_2663_)
  );
  AND2_X1 _7958_ (
    .A1(_4613_),
    .A2(_2663_),
    .ZN(_2664_)
  );
  AND2_X1 _7959_ (
    .A1(_2662_),
    .A2(_2664_),
    .ZN(_2665_)
  );
  AND2_X1 _7960_ (
    .A1(remainder[55]),
    .A2(_4610_),
    .ZN(_2666_)
  );
  OR2_X1 _7961_ (
    .A1(remainder[54]),
    .A2(_4393_),
    .ZN(_2667_)
  );
  OR2_X1 _7962_ (
    .A1(_4392_),
    .A2(_4550_),
    .ZN(_2668_)
  );
  AND2_X1 _7963_ (
    .A1(_3678_),
    .A2(_2668_),
    .ZN(_2669_)
  );
  AND2_X1 _7964_ (
    .A1(_2667_),
    .A2(_2669_),
    .ZN(_2670_)
  );
  OR2_X1 _7965_ (
    .A1(_2665_),
    .A2(_2670_),
    .ZN(_2671_)
  );
  OR2_X1 _7966_ (
    .A1(_2666_),
    .A2(_2671_),
    .ZN(_2672_)
  );
  AND2_X1 _7967_ (
    .A1(_3911_),
    .A2(_2672_),
    .ZN(_0076_)
  );
  AND2_X1 _7968_ (
    .A1(_2654_),
    .A2(_2662_),
    .ZN(_2673_)
  );
  OR2_X1 _7969_ (
    .A1(_2653_),
    .A2(_2661_),
    .ZN(_2674_)
  );
  OR2_X1 _7970_ (
    .A1(_2645_),
    .A2(_2651_),
    .ZN(_2675_)
  );
  OR2_X1 _7971_ (
    .A1(_2639_),
    .A2(_2641_),
    .ZN(_2676_)
  );
  OR2_X1 _7972_ (
    .A1(_2632_),
    .A2(_2635_),
    .ZN(_2677_)
  );
  OR2_X1 _7973_ (
    .A1(_2629_),
    .A2(_2637_),
    .ZN(_2678_)
  );
  OR2_X1 _7974_ (
    .A1(_2603_),
    .A2(_2627_),
    .ZN(_2679_)
  );
  AND2_X1 _7975_ (
    .A1(_0541_),
    .A2(_2598_),
    .ZN(_2680_)
  );
  AND2_X1 _7976_ (
    .A1(_2487_),
    .A2(_2680_),
    .ZN(_2681_)
  );
  OR2_X1 _7977_ (
    .A1(_2601_),
    .A2(_2681_),
    .ZN(_2682_)
  );
  OR2_X1 _7978_ (
    .A1(_2572_),
    .A2(_2587_),
    .ZN(_2683_)
  );
  OR2_X1 _7979_ (
    .A1(_2568_),
    .A2(_2570_),
    .ZN(_2684_)
  );
  OR2_X1 _7980_ (
    .A1(_2564_),
    .A2(_2566_),
    .ZN(_2685_)
  );
  OR2_X1 _7981_ (
    .A1(_2594_),
    .A2(_2596_),
    .ZN(_2686_)
  );
  AND2_X1 _7982_ (
    .A1(divisor[25]),
    .A2(remainder[6]),
    .ZN(_2687_)
  );
  AND2_X1 _7983_ (
    .A1(divisor[26]),
    .A2(remainder[5]),
    .ZN(_2688_)
  );
  AND2_X1 _7984_ (
    .A1(divisor[27]),
    .A2(remainder[5]),
    .ZN(_2689_)
  );
  AND2_X1 _7985_ (
    .A1(_2563_),
    .A2(_2688_),
    .ZN(_2690_)
  );
  XOR2_X1 _7986_ (
    .A(_2563_),
    .B(_2688_),
    .Z(_2691_)
  );
  AND2_X1 _7987_ (
    .A1(_2687_),
    .A2(_2691_),
    .ZN(_2692_)
  );
  XOR2_X1 _7988_ (
    .A(_2687_),
    .B(_2691_),
    .Z(_2693_)
  );
  AND2_X1 _7989_ (
    .A1(_2686_),
    .A2(_2693_),
    .ZN(_2694_)
  );
  XOR2_X1 _7990_ (
    .A(_2686_),
    .B(_2693_),
    .Z(_2695_)
  );
  AND2_X1 _7991_ (
    .A1(_2685_),
    .A2(_2695_),
    .ZN(_2696_)
  );
  XOR2_X1 _7992_ (
    .A(_2685_),
    .B(_2695_),
    .Z(_2697_)
  );
  AND2_X1 _7993_ (
    .A1(_2684_),
    .A2(_2697_),
    .ZN(_2698_)
  );
  XOR2_X1 _7994_ (
    .A(_2684_),
    .B(_2697_),
    .Z(_2699_)
  );
  OR2_X1 _7995_ (
    .A1(_2579_),
    .A2(_2581_),
    .ZN(_2700_)
  );
  AND2_X1 _7996_ (
    .A1(remainder[32]),
    .A2(divisor[24]),
    .ZN(_2701_)
  );
  AND2_X1 _7997_ (
    .A1(remainder[32]),
    .A2(divisor[23]),
    .ZN(_2702_)
  );
  AND2_X1 _7998_ (
    .A1(_2578_),
    .A2(_2702_),
    .ZN(_2703_)
  );
  XOR2_X1 _7999_ (
    .A(_2578_),
    .B(_2702_),
    .Z(_2704_)
  );
  AND2_X1 _8000_ (
    .A1(_2575_),
    .A2(_2704_),
    .ZN(_2705_)
  );
  XOR2_X1 _8001_ (
    .A(_2575_),
    .B(_2704_),
    .Z(_2706_)
  );
  AND2_X1 _8002_ (
    .A1(_2700_),
    .A2(_2706_),
    .ZN(_2707_)
  );
  XOR2_X1 _8003_ (
    .A(_2700_),
    .B(_2706_),
    .Z(_2708_)
  );
  AND2_X1 _8004_ (
    .A1(_2475_),
    .A2(_2708_),
    .ZN(_2709_)
  );
  XOR2_X1 _8005_ (
    .A(_2475_),
    .B(_2708_),
    .Z(_2710_)
  );
  AND2_X1 _8006_ (
    .A1(_2699_),
    .A2(_2710_),
    .ZN(_2711_)
  );
  XOR2_X1 _8007_ (
    .A(_2699_),
    .B(_2710_),
    .Z(_2712_)
  );
  AND2_X1 _8008_ (
    .A1(_2683_),
    .A2(_2712_),
    .ZN(_2713_)
  );
  XOR2_X1 _8009_ (
    .A(_2683_),
    .B(_2712_),
    .Z(_2714_)
  );
  AND2_X1 _8010_ (
    .A1(divisor[31]),
    .A2(remainder[0]),
    .ZN(_2715_)
  );
  AND2_X1 _8011_ (
    .A1(divisor[28]),
    .A2(remainder[3]),
    .ZN(_2716_)
  );
  AND2_X1 _8012_ (
    .A1(divisor[29]),
    .A2(remainder[2]),
    .ZN(_2717_)
  );
  AND2_X1 _8013_ (
    .A1(divisor[30]),
    .A2(remainder[2]),
    .ZN(_2718_)
  );
  AND2_X1 _8014_ (
    .A1(_2485_),
    .A2(_2718_),
    .ZN(_2719_)
  );
  XOR2_X1 _8015_ (
    .A(_2593_),
    .B(_2717_),
    .Z(_2720_)
  );
  AND2_X1 _8016_ (
    .A1(_2716_),
    .A2(_2720_),
    .ZN(_2721_)
  );
  XOR2_X1 _8017_ (
    .A(_2716_),
    .B(_2720_),
    .Z(_2722_)
  );
  AND2_X1 _8018_ (
    .A1(_2715_),
    .A2(_2722_),
    .ZN(_2723_)
  );
  XOR2_X1 _8019_ (
    .A(_2715_),
    .B(_2722_),
    .Z(_2724_)
  );
  INV_X1 _8020_ (
    .A(_2724_),
    .ZN(_2725_)
  );
  XOR2_X1 _8021_ (
    .A(_2680_),
    .B(_2724_),
    .Z(_2726_)
  );
  AND2_X1 _8022_ (
    .A1(_2714_),
    .A2(_2726_),
    .ZN(_2727_)
  );
  XOR2_X1 _8023_ (
    .A(_2714_),
    .B(_2726_),
    .Z(_2728_)
  );
  AND2_X1 _8024_ (
    .A1(_2682_),
    .A2(_2728_),
    .ZN(_2729_)
  );
  XOR2_X1 _8025_ (
    .A(_2682_),
    .B(_2728_),
    .Z(_2730_)
  );
  OR2_X1 _8026_ (
    .A1(_2619_),
    .A2(_2621_),
    .ZN(_2731_)
  );
  OR2_X1 _8027_ (
    .A1(_2615_),
    .A2(_2617_),
    .ZN(_2732_)
  );
  OR2_X1 _8028_ (
    .A1(_2610_),
    .A2(_2612_),
    .ZN(_2733_)
  );
  OR2_X1 _8029_ (
    .A1(_2583_),
    .A2(_2585_),
    .ZN(_2734_)
  );
  AND2_X1 _8030_ (
    .A1(_2613_),
    .A2(_2734_),
    .ZN(_2735_)
  );
  XOR2_X1 _8031_ (
    .A(_2613_),
    .B(_2734_),
    .Z(_2736_)
  );
  AND2_X1 _8032_ (
    .A1(_2733_),
    .A2(_2736_),
    .ZN(_2737_)
  );
  XOR2_X1 _8033_ (
    .A(_2733_),
    .B(_2736_),
    .Z(_2738_)
  );
  AND2_X1 _8034_ (
    .A1(_2732_),
    .A2(_2738_),
    .ZN(_2739_)
  );
  XOR2_X1 _8035_ (
    .A(_2732_),
    .B(_2738_),
    .Z(_2740_)
  );
  AND2_X1 _8036_ (
    .A1(_2025_),
    .A2(_2740_),
    .ZN(_2741_)
  );
  XOR2_X1 _8037_ (
    .A(_2025_),
    .B(_2740_),
    .Z(_2742_)
  );
  AND2_X1 _8038_ (
    .A1(_2589_),
    .A2(_2742_),
    .ZN(_2743_)
  );
  XOR2_X1 _8039_ (
    .A(_2589_),
    .B(_2742_),
    .Z(_2744_)
  );
  AND2_X1 _8040_ (
    .A1(_2731_),
    .A2(_2744_),
    .ZN(_2745_)
  );
  XOR2_X1 _8041_ (
    .A(_2731_),
    .B(_2744_),
    .Z(_2746_)
  );
  AND2_X1 _8042_ (
    .A1(_2730_),
    .A2(_2746_),
    .ZN(_2747_)
  );
  XOR2_X1 _8043_ (
    .A(_2730_),
    .B(_2746_),
    .Z(_2748_)
  );
  AND2_X1 _8044_ (
    .A1(_2679_),
    .A2(_2748_),
    .ZN(_2749_)
  );
  XOR2_X1 _8045_ (
    .A(_2679_),
    .B(_2748_),
    .Z(_2750_)
  );
  OR2_X1 _8046_ (
    .A1(_2623_),
    .A2(_2625_),
    .ZN(_2751_)
  );
  AND2_X1 _8047_ (
    .A1(_2287_),
    .A2(_2751_),
    .ZN(_2752_)
  );
  XOR2_X1 _8048_ (
    .A(_2288_),
    .B(_2751_),
    .Z(_2753_)
  );
  OR2_X1 _8049_ (
    .A1(_2400_),
    .A2(_2753_),
    .ZN(_2754_)
  );
  INV_X1 _8050_ (
    .A(_2754_),
    .ZN(_2755_)
  );
  XOR2_X1 _8051_ (
    .A(_2400_),
    .B(_2753_),
    .Z(_2756_)
  );
  AND2_X1 _8052_ (
    .A1(_2750_),
    .A2(_2756_),
    .ZN(_2757_)
  );
  XOR2_X1 _8053_ (
    .A(_2750_),
    .B(_2756_),
    .Z(_2758_)
  );
  AND2_X1 _8054_ (
    .A1(_2678_),
    .A2(_2758_),
    .ZN(_2759_)
  );
  XOR2_X1 _8055_ (
    .A(_2678_),
    .B(_2758_),
    .Z(_2760_)
  );
  AND2_X1 _8056_ (
    .A1(_2677_),
    .A2(_2760_),
    .ZN(_2761_)
  );
  XOR2_X1 _8057_ (
    .A(_2677_),
    .B(_2760_),
    .Z(_2762_)
  );
  AND2_X1 _8058_ (
    .A1(_2676_),
    .A2(_2762_),
    .ZN(_2763_)
  );
  XOR2_X1 _8059_ (
    .A(_2676_),
    .B(_2762_),
    .Z(_2764_)
  );
  AND2_X1 _8060_ (
    .A1(_2643_),
    .A2(_2764_),
    .ZN(_2765_)
  );
  OR2_X1 _8061_ (
    .A1(_2643_),
    .A2(_2764_),
    .ZN(_2766_)
  );
  XOR2_X1 _8062_ (
    .A(_2643_),
    .B(_2764_),
    .Z(_2767_)
  );
  XOR2_X1 _8063_ (
    .A(_2675_),
    .B(_2767_),
    .Z(_2768_)
  );
  AND2_X1 _8064_ (
    .A1(remainder[64]),
    .A2(_2768_),
    .ZN(_2769_)
  );
  INV_X1 _8065_ (
    .A(_2769_),
    .ZN(_2770_)
  );
  XOR2_X1 _8066_ (
    .A(remainder[64]),
    .B(_2768_),
    .Z(_2771_)
  );
  INV_X1 _8067_ (
    .A(_2771_),
    .ZN(_2772_)
  );
  AND2_X1 _8068_ (
    .A1(_2674_),
    .A2(_2771_),
    .ZN(_2773_)
  );
  OR2_X1 _8069_ (
    .A1(_2673_),
    .A2(_2772_),
    .ZN(_2774_)
  );
  OR2_X1 _8070_ (
    .A1(_2674_),
    .A2(_2771_),
    .ZN(_2775_)
  );
  AND2_X1 _8071_ (
    .A1(_4613_),
    .A2(_2775_),
    .ZN(_2776_)
  );
  AND2_X1 _8072_ (
    .A1(_2774_),
    .A2(_2776_),
    .ZN(_2777_)
  );
  AND2_X1 _8073_ (
    .A1(remainder[56]),
    .A2(_4610_),
    .ZN(_2778_)
  );
  MUX2_X1 _8074_ (
    .A(remainder[55]),
    .B(_4556_),
    .S(_4393_),
    .Z(_2779_)
  );
  AND2_X1 _8075_ (
    .A1(_3678_),
    .A2(_2779_),
    .ZN(_2780_)
  );
  OR2_X1 _8076_ (
    .A1(_2778_),
    .A2(_2780_),
    .ZN(_2781_)
  );
  OR2_X1 _8077_ (
    .A1(_2777_),
    .A2(_2781_),
    .ZN(_2782_)
  );
  AND2_X1 _8078_ (
    .A1(_3911_),
    .A2(_2782_),
    .ZN(_0077_)
  );
  AND2_X1 _8079_ (
    .A1(_2770_),
    .A2(_2774_),
    .ZN(_2783_)
  );
  OR2_X1 _8080_ (
    .A1(_2769_),
    .A2(_2773_),
    .ZN(_2784_)
  );
  OR2_X1 _8081_ (
    .A1(_2759_),
    .A2(_2761_),
    .ZN(_2785_)
  );
  OR2_X1 _8082_ (
    .A1(_2752_),
    .A2(_2755_),
    .ZN(_2786_)
  );
  OR2_X1 _8083_ (
    .A1(_2749_),
    .A2(_2757_),
    .ZN(_2787_)
  );
  OR2_X1 _8084_ (
    .A1(_2729_),
    .A2(_2747_),
    .ZN(_2788_)
  );
  AND2_X1 _8085_ (
    .A1(_0541_),
    .A2(_2725_),
    .ZN(_2789_)
  );
  AND2_X1 _8086_ (
    .A1(_2597_),
    .A2(_2789_),
    .ZN(_2790_)
  );
  OR2_X1 _8087_ (
    .A1(_2727_),
    .A2(_2790_),
    .ZN(_2791_)
  );
  OR2_X1 _8088_ (
    .A1(_2698_),
    .A2(_2711_),
    .ZN(_2792_)
  );
  OR2_X1 _8089_ (
    .A1(_2694_),
    .A2(_2696_),
    .ZN(_2793_)
  );
  OR2_X1 _8090_ (
    .A1(_2690_),
    .A2(_2692_),
    .ZN(_2794_)
  );
  OR2_X1 _8091_ (
    .A1(_2719_),
    .A2(_2721_),
    .ZN(_2795_)
  );
  AND2_X1 _8092_ (
    .A1(divisor[25]),
    .A2(remainder[7]),
    .ZN(_2796_)
  );
  AND2_X1 _8093_ (
    .A1(divisor[26]),
    .A2(remainder[6]),
    .ZN(_2797_)
  );
  AND2_X1 _8094_ (
    .A1(divisor[27]),
    .A2(remainder[6]),
    .ZN(_2798_)
  );
  AND2_X1 _8095_ (
    .A1(_2689_),
    .A2(_2797_),
    .ZN(_2799_)
  );
  XOR2_X1 _8096_ (
    .A(_2689_),
    .B(_2797_),
    .Z(_2800_)
  );
  AND2_X1 _8097_ (
    .A1(_2796_),
    .A2(_2800_),
    .ZN(_2801_)
  );
  XOR2_X1 _8098_ (
    .A(_2796_),
    .B(_2800_),
    .Z(_2802_)
  );
  AND2_X1 _8099_ (
    .A1(_2795_),
    .A2(_2802_),
    .ZN(_2803_)
  );
  XOR2_X1 _8100_ (
    .A(_2795_),
    .B(_2802_),
    .Z(_2804_)
  );
  AND2_X1 _8101_ (
    .A1(_2794_),
    .A2(_2804_),
    .ZN(_2805_)
  );
  XOR2_X1 _8102_ (
    .A(_2794_),
    .B(_2804_),
    .Z(_2806_)
  );
  AND2_X1 _8103_ (
    .A1(_2793_),
    .A2(_2806_),
    .ZN(_2807_)
  );
  XOR2_X1 _8104_ (
    .A(_2793_),
    .B(_2806_),
    .Z(_2808_)
  );
  OR2_X1 _8105_ (
    .A1(_2703_),
    .A2(_2705_),
    .ZN(_2809_)
  );
  INV_X1 _8106_ (
    .A(_2809_),
    .ZN(_2810_)
  );
  OR2_X1 _8107_ (
    .A1(_2701_),
    .A2(_2702_),
    .ZN(_2811_)
  );
  MUX2_X1 _8108_ (
    .A(_2702_),
    .B(_3384_),
    .S(_2701_),
    .Z(_2812_)
  );
  MUX2_X1 _8109_ (
    .A(_2576_),
    .B(divisor[22]),
    .S(_2812_),
    .Z(_2813_)
  );
  OR2_X1 _8110_ (
    .A1(_2810_),
    .A2(_2813_),
    .ZN(_2814_)
  );
  INV_X1 _8111_ (
    .A(_2814_),
    .ZN(_2815_)
  );
  XOR2_X1 _8112_ (
    .A(_2809_),
    .B(_2813_),
    .Z(_2816_)
  );
  OR2_X1 _8113_ (
    .A1(_2476_),
    .A2(_2816_),
    .ZN(_2817_)
  );
  XOR2_X1 _8114_ (
    .A(_2476_),
    .B(_2816_),
    .Z(_2818_)
  );
  AND2_X1 _8115_ (
    .A1(_2808_),
    .A2(_2818_),
    .ZN(_2819_)
  );
  XOR2_X1 _8116_ (
    .A(_2808_),
    .B(_2818_),
    .Z(_2820_)
  );
  AND2_X1 _8117_ (
    .A1(_2792_),
    .A2(_2820_),
    .ZN(_2821_)
  );
  XOR2_X1 _8118_ (
    .A(_2792_),
    .B(_2820_),
    .Z(_2822_)
  );
  AND2_X1 _8119_ (
    .A1(divisor[32]),
    .A2(remainder[0]),
    .ZN(_2823_)
  );
  INV_X1 _8120_ (
    .A(_2823_),
    .ZN(_2824_)
  );
  AND2_X1 _8121_ (
    .A1(divisor[31]),
    .A2(remainder[1]),
    .ZN(_2825_)
  );
  AND2_X1 _8122_ (
    .A1(divisor[32]),
    .A2(remainder[1]),
    .ZN(_2826_)
  );
  AND2_X1 _8123_ (
    .A1(_2715_),
    .A2(_2826_),
    .ZN(_2827_)
  );
  XOR2_X1 _8124_ (
    .A(_2823_),
    .B(_2825_),
    .Z(_2828_)
  );
  AND2_X1 _8125_ (
    .A1(divisor[28]),
    .A2(remainder[4]),
    .ZN(_2829_)
  );
  AND2_X1 _8126_ (
    .A1(divisor[29]),
    .A2(remainder[3]),
    .ZN(_2830_)
  );
  AND2_X1 _8127_ (
    .A1(divisor[30]),
    .A2(remainder[3]),
    .ZN(_2831_)
  );
  AND2_X1 _8128_ (
    .A1(_2718_),
    .A2(_2830_),
    .ZN(_2832_)
  );
  XOR2_X1 _8129_ (
    .A(_2718_),
    .B(_2830_),
    .Z(_2833_)
  );
  AND2_X1 _8130_ (
    .A1(_2829_),
    .A2(_2833_),
    .ZN(_2834_)
  );
  XOR2_X1 _8131_ (
    .A(_2829_),
    .B(_2833_),
    .Z(_2835_)
  );
  AND2_X1 _8132_ (
    .A1(_2828_),
    .A2(_2835_),
    .ZN(_2836_)
  );
  XOR2_X1 _8133_ (
    .A(_2828_),
    .B(_2835_),
    .Z(_2837_)
  );
  AND2_X1 _8134_ (
    .A1(_2723_),
    .A2(_2837_),
    .ZN(_2838_)
  );
  XOR2_X1 _8135_ (
    .A(_2723_),
    .B(_2837_),
    .Z(_2839_)
  );
  INV_X1 _8136_ (
    .A(_2839_),
    .ZN(_2840_)
  );
  XOR2_X1 _8137_ (
    .A(_2789_),
    .B(_2839_),
    .Z(_2841_)
  );
  AND2_X1 _8138_ (
    .A1(_2822_),
    .A2(_2841_),
    .ZN(_2842_)
  );
  XOR2_X1 _8139_ (
    .A(_2822_),
    .B(_2841_),
    .Z(_2843_)
  );
  AND2_X1 _8140_ (
    .A1(_2791_),
    .A2(_2843_),
    .ZN(_2844_)
  );
  XOR2_X1 _8141_ (
    .A(_2791_),
    .B(_2843_),
    .Z(_2845_)
  );
  OR2_X1 _8142_ (
    .A1(_2739_),
    .A2(_2741_),
    .ZN(_2846_)
  );
  OR2_X1 _8143_ (
    .A1(_2735_),
    .A2(_2737_),
    .ZN(_2847_)
  );
  OR2_X1 _8144_ (
    .A1(_2707_),
    .A2(_2709_),
    .ZN(_2848_)
  );
  AND2_X1 _8145_ (
    .A1(_2613_),
    .A2(_2848_),
    .ZN(_2849_)
  );
  XOR2_X1 _8146_ (
    .A(_2613_),
    .B(_2848_),
    .Z(_2850_)
  );
  AND2_X1 _8147_ (
    .A1(_2733_),
    .A2(_2850_),
    .ZN(_2851_)
  );
  XOR2_X1 _8148_ (
    .A(_2733_),
    .B(_2850_),
    .Z(_2852_)
  );
  AND2_X1 _8149_ (
    .A1(_2847_),
    .A2(_2852_),
    .ZN(_2853_)
  );
  XOR2_X1 _8150_ (
    .A(_2847_),
    .B(_2852_),
    .Z(_2854_)
  );
  AND2_X1 _8151_ (
    .A1(_2025_),
    .A2(_2854_),
    .ZN(_2855_)
  );
  XOR2_X1 _8152_ (
    .A(_2025_),
    .B(_2854_),
    .Z(_2856_)
  );
  AND2_X1 _8153_ (
    .A1(_2713_),
    .A2(_2856_),
    .ZN(_2857_)
  );
  XOR2_X1 _8154_ (
    .A(_2713_),
    .B(_2856_),
    .Z(_2858_)
  );
  AND2_X1 _8155_ (
    .A1(_2846_),
    .A2(_2858_),
    .ZN(_2859_)
  );
  XOR2_X1 _8156_ (
    .A(_2846_),
    .B(_2858_),
    .Z(_2860_)
  );
  AND2_X1 _8157_ (
    .A1(_2845_),
    .A2(_2860_),
    .ZN(_2861_)
  );
  XOR2_X1 _8158_ (
    .A(_2845_),
    .B(_2860_),
    .Z(_2862_)
  );
  AND2_X1 _8159_ (
    .A1(_2788_),
    .A2(_2862_),
    .ZN(_2863_)
  );
  XOR2_X1 _8160_ (
    .A(_2788_),
    .B(_2862_),
    .Z(_2864_)
  );
  OR2_X1 _8161_ (
    .A1(_2743_),
    .A2(_2745_),
    .ZN(_2865_)
  );
  AND2_X1 _8162_ (
    .A1(_2287_),
    .A2(_2865_),
    .ZN(_2866_)
  );
  XOR2_X1 _8163_ (
    .A(_2288_),
    .B(_2865_),
    .Z(_2867_)
  );
  OR2_X1 _8164_ (
    .A1(_2400_),
    .A2(_2867_),
    .ZN(_2868_)
  );
  INV_X1 _8165_ (
    .A(_2868_),
    .ZN(_2869_)
  );
  XOR2_X1 _8166_ (
    .A(_2400_),
    .B(_2867_),
    .Z(_2870_)
  );
  AND2_X1 _8167_ (
    .A1(_2864_),
    .A2(_2870_),
    .ZN(_2871_)
  );
  XOR2_X1 _8168_ (
    .A(_2864_),
    .B(_2870_),
    .Z(_2872_)
  );
  AND2_X1 _8169_ (
    .A1(_2787_),
    .A2(_2872_),
    .ZN(_2873_)
  );
  XOR2_X1 _8170_ (
    .A(_2787_),
    .B(_2872_),
    .Z(_2874_)
  );
  AND2_X1 _8171_ (
    .A1(_2786_),
    .A2(_2874_),
    .ZN(_2875_)
  );
  XOR2_X1 _8172_ (
    .A(_2786_),
    .B(_2874_),
    .Z(_2876_)
  );
  AND2_X1 _8173_ (
    .A1(_2785_),
    .A2(_2876_),
    .ZN(_2877_)
  );
  XOR2_X1 _8174_ (
    .A(_2785_),
    .B(_2876_),
    .Z(_2878_)
  );
  AND2_X1 _8175_ (
    .A1(_2763_),
    .A2(_2878_),
    .ZN(_2879_)
  );
  XOR2_X1 _8176_ (
    .A(_2763_),
    .B(_2878_),
    .Z(_2880_)
  );
  OR2_X1 _8177_ (
    .A1(_2645_),
    .A2(_2765_),
    .ZN(_2881_)
  );
  AND2_X1 _8178_ (
    .A1(_2766_),
    .A2(_2881_),
    .ZN(_2882_)
  );
  AND2_X1 _8179_ (
    .A1(_2651_),
    .A2(_2767_),
    .ZN(_2883_)
  );
  OR2_X1 _8180_ (
    .A1(_2882_),
    .A2(_2883_),
    .ZN(_2884_)
  );
  AND2_X1 _8181_ (
    .A1(_2880_),
    .A2(_2884_),
    .ZN(_2885_)
  );
  XOR2_X1 _8182_ (
    .A(_2880_),
    .B(_2884_),
    .Z(_2886_)
  );
  AND2_X1 _8183_ (
    .A1(remainder[65]),
    .A2(_2886_),
    .ZN(_2887_)
  );
  XOR2_X1 _8184_ (
    .A(remainder[65]),
    .B(_2886_),
    .Z(_2888_)
  );
  INV_X1 _8185_ (
    .A(_2888_),
    .ZN(_2889_)
  );
  AND2_X1 _8186_ (
    .A1(_2784_),
    .A2(_2888_),
    .ZN(_2890_)
  );
  OR2_X1 _8187_ (
    .A1(_2783_),
    .A2(_2889_),
    .ZN(_2891_)
  );
  OR2_X1 _8188_ (
    .A1(_2784_),
    .A2(_2888_),
    .ZN(_2892_)
  );
  AND2_X1 _8189_ (
    .A1(_4613_),
    .A2(_2892_),
    .ZN(_2893_)
  );
  AND2_X1 _8190_ (
    .A1(_2891_),
    .A2(_2893_),
    .ZN(_2894_)
  );
  AND2_X1 _8191_ (
    .A1(remainder[57]),
    .A2(_4610_),
    .ZN(_2895_)
  );
  OR2_X1 _8192_ (
    .A1(remainder[56]),
    .A2(_4393_),
    .ZN(_2896_)
  );
  OR2_X1 _8193_ (
    .A1(_4392_),
    .A2(_4561_),
    .ZN(_2897_)
  );
  AND2_X1 _8194_ (
    .A1(_3678_),
    .A2(_2897_),
    .ZN(_2898_)
  );
  AND2_X1 _8195_ (
    .A1(_2896_),
    .A2(_2898_),
    .ZN(_2899_)
  );
  OR2_X1 _8196_ (
    .A1(_2895_),
    .A2(_2899_),
    .ZN(_2900_)
  );
  OR2_X1 _8197_ (
    .A1(_2894_),
    .A2(_2900_),
    .ZN(_2901_)
  );
  AND2_X1 _8198_ (
    .A1(_3911_),
    .A2(_2901_),
    .ZN(_0078_)
  );
  OR2_X1 _8199_ (
    .A1(_2887_),
    .A2(_2890_),
    .ZN(_2902_)
  );
  OR2_X1 _8200_ (
    .A1(_2879_),
    .A2(_2885_),
    .ZN(_2903_)
  );
  OR2_X1 _8201_ (
    .A1(_2873_),
    .A2(_2875_),
    .ZN(_2904_)
  );
  OR2_X1 _8202_ (
    .A1(_2866_),
    .A2(_2869_),
    .ZN(_2905_)
  );
  OR2_X1 _8203_ (
    .A1(_2863_),
    .A2(_2871_),
    .ZN(_2906_)
  );
  OR2_X1 _8204_ (
    .A1(_2844_),
    .A2(_2861_),
    .ZN(_2907_)
  );
  AND2_X1 _8205_ (
    .A1(_0541_),
    .A2(_2840_),
    .ZN(_2908_)
  );
  AND2_X1 _8206_ (
    .A1(_2724_),
    .A2(_2908_),
    .ZN(_2909_)
  );
  OR2_X1 _8207_ (
    .A1(_2842_),
    .A2(_2909_),
    .ZN(_2910_)
  );
  OR2_X1 _8208_ (
    .A1(_2807_),
    .A2(_2819_),
    .ZN(_2911_)
  );
  OR2_X1 _8209_ (
    .A1(_2803_),
    .A2(_2805_),
    .ZN(_2912_)
  );
  OR2_X1 _8210_ (
    .A1(_2799_),
    .A2(_2801_),
    .ZN(_2913_)
  );
  OR2_X1 _8211_ (
    .A1(_2832_),
    .A2(_2834_),
    .ZN(_2914_)
  );
  AND2_X1 _8212_ (
    .A1(remainder[32]),
    .A2(divisor[25]),
    .ZN(_2915_)
  );
  AND2_X1 _8213_ (
    .A1(divisor[26]),
    .A2(remainder[7]),
    .ZN(_2916_)
  );
  AND2_X1 _8214_ (
    .A1(divisor[27]),
    .A2(remainder[7]),
    .ZN(_2917_)
  );
  AND2_X1 _8215_ (
    .A1(_2797_),
    .A2(_2917_),
    .ZN(_2918_)
  );
  XOR2_X1 _8216_ (
    .A(_2798_),
    .B(_2916_),
    .Z(_2919_)
  );
  AND2_X1 _8217_ (
    .A1(_2915_),
    .A2(_2919_),
    .ZN(_2920_)
  );
  XOR2_X1 _8218_ (
    .A(_2915_),
    .B(_2919_),
    .Z(_2921_)
  );
  AND2_X1 _8219_ (
    .A1(_2914_),
    .A2(_2921_),
    .ZN(_2922_)
  );
  XOR2_X1 _8220_ (
    .A(_2914_),
    .B(_2921_),
    .Z(_2923_)
  );
  AND2_X1 _8221_ (
    .A1(_2913_),
    .A2(_2923_),
    .ZN(_2924_)
  );
  XOR2_X1 _8222_ (
    .A(_2913_),
    .B(_2923_),
    .Z(_2925_)
  );
  AND2_X1 _8223_ (
    .A1(_2912_),
    .A2(_2925_),
    .ZN(_2926_)
  );
  XOR2_X1 _8224_ (
    .A(_2912_),
    .B(_2925_),
    .Z(_2927_)
  );
  OR2_X1 _8225_ (
    .A1(_2575_),
    .A2(_2811_),
    .ZN(_2928_)
  );
  AND2_X1 _8226_ (
    .A1(_2814_),
    .A2(_2928_),
    .ZN(_2929_)
  );
  AND2_X1 _8227_ (
    .A1(_2475_),
    .A2(_2929_),
    .ZN(_2930_)
  );
  XOR2_X1 _8228_ (
    .A(_2475_),
    .B(_2929_),
    .Z(_2931_)
  );
  INV_X1 _8229_ (
    .A(_2931_),
    .ZN(_2932_)
  );
  AND2_X1 _8230_ (
    .A1(_2927_),
    .A2(_2931_),
    .ZN(_2933_)
  );
  XOR2_X1 _8231_ (
    .A(_2927_),
    .B(_2931_),
    .Z(_2934_)
  );
  AND2_X1 _8232_ (
    .A1(_2838_),
    .A2(_2934_),
    .ZN(_2935_)
  );
  XOR2_X1 _8233_ (
    .A(_2838_),
    .B(_2934_),
    .Z(_2937_)
  );
  AND2_X1 _8234_ (
    .A1(_2911_),
    .A2(_2937_),
    .ZN(_2938_)
  );
  XOR2_X1 _8235_ (
    .A(_2911_),
    .B(_2937_),
    .Z(_2939_)
  );
  AND2_X1 _8236_ (
    .A1(divisor[31]),
    .A2(remainder[2]),
    .ZN(_2940_)
  );
  AND2_X1 _8237_ (
    .A1(remainder[1]),
    .A2(_2823_),
    .ZN(_2941_)
  );
  MUX2_X1 _8238_ (
    .A(_2826_),
    .B(_3449_),
    .S(_2823_),
    .Z(_2942_)
  );
  MUX2_X1 _8239_ (
    .A(_2824_),
    .B(remainder[0]),
    .S(_2826_),
    .Z(_2943_)
  );
  AND2_X1 _8240_ (
    .A1(_2940_),
    .A2(_2942_),
    .ZN(_2944_)
  );
  XOR2_X1 _8241_ (
    .A(_2940_),
    .B(_2942_),
    .Z(_2945_)
  );
  AND2_X1 _8242_ (
    .A1(_2827_),
    .A2(_2945_),
    .ZN(_2946_)
  );
  XOR2_X1 _8243_ (
    .A(_2827_),
    .B(_2945_),
    .Z(_2948_)
  );
  AND2_X1 _8244_ (
    .A1(divisor[28]),
    .A2(remainder[5]),
    .ZN(_2949_)
  );
  AND2_X1 _8245_ (
    .A1(divisor[29]),
    .A2(remainder[4]),
    .ZN(_2950_)
  );
  AND2_X1 _8246_ (
    .A1(divisor[30]),
    .A2(remainder[4]),
    .ZN(_2951_)
  );
  AND2_X1 _8247_ (
    .A1(_2831_),
    .A2(_2950_),
    .ZN(_2952_)
  );
  XOR2_X1 _8248_ (
    .A(_2831_),
    .B(_2950_),
    .Z(_2953_)
  );
  AND2_X1 _8249_ (
    .A1(_2949_),
    .A2(_2953_),
    .ZN(_2954_)
  );
  XOR2_X1 _8250_ (
    .A(_2949_),
    .B(_2953_),
    .Z(_2955_)
  );
  AND2_X1 _8251_ (
    .A1(_2948_),
    .A2(_2955_),
    .ZN(_2956_)
  );
  XOR2_X1 _8252_ (
    .A(_2948_),
    .B(_2955_),
    .Z(_2957_)
  );
  AND2_X1 _8253_ (
    .A1(_2836_),
    .A2(_2957_),
    .ZN(_2959_)
  );
  XOR2_X1 _8254_ (
    .A(_2836_),
    .B(_2957_),
    .Z(_2960_)
  );
  INV_X1 _8255_ (
    .A(_2960_),
    .ZN(_2961_)
  );
  XOR2_X1 _8256_ (
    .A(_2908_),
    .B(_2960_),
    .Z(_2962_)
  );
  AND2_X1 _8257_ (
    .A1(_2939_),
    .A2(_2962_),
    .ZN(_2963_)
  );
  XOR2_X1 _8258_ (
    .A(_2939_),
    .B(_2962_),
    .Z(_2964_)
  );
  AND2_X1 _8259_ (
    .A1(_2910_),
    .A2(_2964_),
    .ZN(_2965_)
  );
  XOR2_X1 _8260_ (
    .A(_2910_),
    .B(_2964_),
    .Z(_2966_)
  );
  OR2_X1 _8261_ (
    .A1(_2853_),
    .A2(_2855_),
    .ZN(_2967_)
  );
  OR2_X1 _8262_ (
    .A1(_2849_),
    .A2(_2851_),
    .ZN(_2968_)
  );
  AND2_X1 _8263_ (
    .A1(_2814_),
    .A2(_2817_),
    .ZN(_2970_)
  );
  OR2_X1 _8264_ (
    .A1(_2614_),
    .A2(_2970_),
    .ZN(_2971_)
  );
  XOR2_X1 _8265_ (
    .A(_2614_),
    .B(_2970_),
    .Z(_2972_)
  );
  AND2_X1 _8266_ (
    .A1(_2733_),
    .A2(_2972_),
    .ZN(_2973_)
  );
  INV_X1 _8267_ (
    .A(_2973_),
    .ZN(_2974_)
  );
  XOR2_X1 _8268_ (
    .A(_2733_),
    .B(_2972_),
    .Z(_2975_)
  );
  AND2_X1 _8269_ (
    .A1(_2968_),
    .A2(_2975_),
    .ZN(_2976_)
  );
  XOR2_X1 _8270_ (
    .A(_2968_),
    .B(_2975_),
    .Z(_2977_)
  );
  AND2_X1 _8271_ (
    .A1(_2025_),
    .A2(_2977_),
    .ZN(_2978_)
  );
  XOR2_X1 _8272_ (
    .A(_2025_),
    .B(_2977_),
    .Z(_2979_)
  );
  AND2_X1 _8273_ (
    .A1(_2821_),
    .A2(_2979_),
    .ZN(_2981_)
  );
  XOR2_X1 _8274_ (
    .A(_2821_),
    .B(_2979_),
    .Z(_2982_)
  );
  AND2_X1 _8275_ (
    .A1(_2967_),
    .A2(_2982_),
    .ZN(_2983_)
  );
  XOR2_X1 _8276_ (
    .A(_2967_),
    .B(_2982_),
    .Z(_2984_)
  );
  AND2_X1 _8277_ (
    .A1(_2966_),
    .A2(_2984_),
    .ZN(_2985_)
  );
  XOR2_X1 _8278_ (
    .A(_2966_),
    .B(_2984_),
    .Z(_2986_)
  );
  AND2_X1 _8279_ (
    .A1(_2907_),
    .A2(_2986_),
    .ZN(_2987_)
  );
  XOR2_X1 _8280_ (
    .A(_2907_),
    .B(_2986_),
    .Z(_2988_)
  );
  OR2_X1 _8281_ (
    .A1(_2857_),
    .A2(_2859_),
    .ZN(_2989_)
  );
  AND2_X1 _8282_ (
    .A1(_2287_),
    .A2(_2989_),
    .ZN(_2990_)
  );
  XOR2_X1 _8283_ (
    .A(_2288_),
    .B(_2989_),
    .Z(_2992_)
  );
  OR2_X1 _8284_ (
    .A1(_2400_),
    .A2(_2992_),
    .ZN(_2993_)
  );
  INV_X1 _8285_ (
    .A(_2993_),
    .ZN(_2994_)
  );
  XOR2_X1 _8286_ (
    .A(_2400_),
    .B(_2992_),
    .Z(_2995_)
  );
  AND2_X1 _8287_ (
    .A1(_2988_),
    .A2(_2995_),
    .ZN(_2996_)
  );
  XOR2_X1 _8288_ (
    .A(_2988_),
    .B(_2995_),
    .Z(_2997_)
  );
  AND2_X1 _8289_ (
    .A1(_2906_),
    .A2(_2997_),
    .ZN(_2998_)
  );
  XOR2_X1 _8290_ (
    .A(_2906_),
    .B(_2997_),
    .Z(_2999_)
  );
  AND2_X1 _8291_ (
    .A1(_2905_),
    .A2(_2999_),
    .ZN(_3000_)
  );
  XOR2_X1 _8292_ (
    .A(_2905_),
    .B(_2999_),
    .Z(_3001_)
  );
  AND2_X1 _8293_ (
    .A1(_2904_),
    .A2(_3001_),
    .ZN(_3003_)
  );
  XOR2_X1 _8294_ (
    .A(_2904_),
    .B(_3001_),
    .Z(_3004_)
  );
  AND2_X1 _8295_ (
    .A1(_2877_),
    .A2(_3004_),
    .ZN(_3005_)
  );
  XOR2_X1 _8296_ (
    .A(_2877_),
    .B(_3004_),
    .Z(_3006_)
  );
  AND2_X1 _8297_ (
    .A1(_2903_),
    .A2(_3006_),
    .ZN(_3007_)
  );
  XOR2_X1 _8298_ (
    .A(_2903_),
    .B(_3006_),
    .Z(_3008_)
  );
  AND2_X1 _8299_ (
    .A1(remainder[65]),
    .A2(_3008_),
    .ZN(_3009_)
  );
  XOR2_X1 _8300_ (
    .A(remainder[65]),
    .B(_3008_),
    .Z(_3010_)
  );
  INV_X1 _8301_ (
    .A(_3010_),
    .ZN(_3011_)
  );
  XOR2_X1 _8302_ (
    .A(_2902_),
    .B(_3010_),
    .Z(_3012_)
  );
  AND2_X1 _8303_ (
    .A1(_4613_),
    .A2(_3012_),
    .ZN(_3014_)
  );
  AND2_X1 _8304_ (
    .A1(remainder[58]),
    .A2(_4610_),
    .ZN(_3015_)
  );
  MUX2_X1 _8305_ (
    .A(remainder[57]),
    .B(_4567_),
    .S(_4393_),
    .Z(_3016_)
  );
  AND2_X1 _8306_ (
    .A1(_3678_),
    .A2(_3016_),
    .ZN(_3017_)
  );
  OR2_X1 _8307_ (
    .A1(_3015_),
    .A2(_3017_),
    .ZN(_3018_)
  );
  OR2_X1 _8308_ (
    .A1(_3014_),
    .A2(_3018_),
    .ZN(_3019_)
  );
  AND2_X1 _8309_ (
    .A1(_3911_),
    .A2(_3019_),
    .ZN(_0079_)
  );
  AND2_X1 _8310_ (
    .A1(_2890_),
    .A2(_3010_),
    .ZN(_3020_)
  );
  OR2_X1 _8311_ (
    .A1(_2891_),
    .A2(_3011_),
    .ZN(_3021_)
  );
  OR2_X1 _8312_ (
    .A1(_2887_),
    .A2(_3009_),
    .ZN(_3022_)
  );
  OR2_X1 _8313_ (
    .A1(_3020_),
    .A2(_3022_),
    .ZN(_3024_)
  );
  INV_X1 _8314_ (
    .A(_3024_),
    .ZN(_3025_)
  );
  OR2_X1 _8315_ (
    .A1(_2998_),
    .A2(_3000_),
    .ZN(_3026_)
  );
  OR2_X1 _8316_ (
    .A1(_2990_),
    .A2(_2994_),
    .ZN(_3027_)
  );
  OR2_X1 _8317_ (
    .A1(_2987_),
    .A2(_2996_),
    .ZN(_3028_)
  );
  OR2_X1 _8318_ (
    .A1(_2965_),
    .A2(_2985_),
    .ZN(_3029_)
  );
  AND2_X1 _8319_ (
    .A1(_0541_),
    .A2(_2839_),
    .ZN(_3030_)
  );
  AND2_X1 _8320_ (
    .A1(_2961_),
    .A2(_3030_),
    .ZN(_3031_)
  );
  OR2_X1 _8321_ (
    .A1(_2963_),
    .A2(_3031_),
    .ZN(_3032_)
  );
  AND2_X1 _8322_ (
    .A1(_0541_),
    .A2(_2960_),
    .ZN(_3033_)
  );
  OR2_X1 _8323_ (
    .A1(_0542_),
    .A2(_2824_),
    .ZN(_3035_)
  );
  XOR2_X1 _8324_ (
    .A(_0541_),
    .B(_2823_),
    .Z(_3036_)
  );
  OR2_X1 _8325_ (
    .A1(_2946_),
    .A2(_2956_),
    .ZN(_3037_)
  );
  OR2_X1 _8326_ (
    .A1(_2941_),
    .A2(_2944_),
    .ZN(_3038_)
  );
  AND2_X1 _8327_ (
    .A1(divisor[31]),
    .A2(remainder[3]),
    .ZN(_3039_)
  );
  AND2_X1 _8328_ (
    .A1(divisor[32]),
    .A2(remainder[2]),
    .ZN(_3040_)
  );
  INV_X1 _8329_ (
    .A(_3040_),
    .ZN(_3041_)
  );
  AND2_X1 _8330_ (
    .A1(remainder[1]),
    .A2(_3040_),
    .ZN(_3042_)
  );
  MUX2_X1 _8331_ (
    .A(_3040_),
    .B(_3460_),
    .S(_2826_),
    .Z(_3043_)
  );
  AND2_X1 _8332_ (
    .A1(_3039_),
    .A2(_3043_),
    .ZN(_3044_)
  );
  XOR2_X1 _8333_ (
    .A(_3039_),
    .B(_3043_),
    .Z(_3046_)
  );
  AND2_X1 _8334_ (
    .A1(_3038_),
    .A2(_3046_),
    .ZN(_3047_)
  );
  XOR2_X1 _8335_ (
    .A(_3038_),
    .B(_3046_),
    .Z(_3048_)
  );
  AND2_X1 _8336_ (
    .A1(divisor[28]),
    .A2(remainder[6]),
    .ZN(_3049_)
  );
  AND2_X1 _8337_ (
    .A1(divisor[29]),
    .A2(remainder[5]),
    .ZN(_3050_)
  );
  AND2_X1 _8338_ (
    .A1(divisor[30]),
    .A2(remainder[5]),
    .ZN(_3051_)
  );
  AND2_X1 _8339_ (
    .A1(_2951_),
    .A2(_3050_),
    .ZN(_3052_)
  );
  XOR2_X1 _8340_ (
    .A(_2951_),
    .B(_3050_),
    .Z(_3053_)
  );
  AND2_X1 _8341_ (
    .A1(_3049_),
    .A2(_3053_),
    .ZN(_3054_)
  );
  XOR2_X1 _8342_ (
    .A(_3049_),
    .B(_3053_),
    .Z(_3055_)
  );
  AND2_X1 _8343_ (
    .A1(_3048_),
    .A2(_3055_),
    .ZN(_3057_)
  );
  XOR2_X1 _8344_ (
    .A(_3048_),
    .B(_3055_),
    .Z(_3058_)
  );
  AND2_X1 _8345_ (
    .A1(_3037_),
    .A2(_3058_),
    .ZN(_3059_)
  );
  XOR2_X1 _8346_ (
    .A(_3037_),
    .B(_3058_),
    .Z(_3060_)
  );
  AND2_X1 _8347_ (
    .A1(_3036_),
    .A2(_3060_),
    .ZN(_3061_)
  );
  XOR2_X1 _8348_ (
    .A(_3036_),
    .B(_3060_),
    .Z(_3062_)
  );
  AND2_X1 _8349_ (
    .A1(_3033_),
    .A2(_3062_),
    .ZN(_3063_)
  );
  XOR2_X1 _8350_ (
    .A(_3033_),
    .B(_3062_),
    .Z(_3064_)
  );
  OR2_X1 _8351_ (
    .A1(_2926_),
    .A2(_2933_),
    .ZN(_3065_)
  );
  OR2_X1 _8352_ (
    .A1(_2922_),
    .A2(_2924_),
    .ZN(_3066_)
  );
  OR2_X1 _8353_ (
    .A1(_2918_),
    .A2(_2920_),
    .ZN(_3068_)
  );
  OR2_X1 _8354_ (
    .A1(_2952_),
    .A2(_2954_),
    .ZN(_3069_)
  );
  AND2_X1 _8355_ (
    .A1(remainder[32]),
    .A2(divisor[27]),
    .ZN(_3070_)
  );
  AND2_X1 _8356_ (
    .A1(remainder[32]),
    .A2(divisor[26]),
    .ZN(_3071_)
  );
  AND2_X1 _8357_ (
    .A1(divisor[27]),
    .A2(_3071_),
    .ZN(_3072_)
  );
  AND2_X1 _8358_ (
    .A1(_2917_),
    .A2(_3071_),
    .ZN(_3073_)
  );
  XOR2_X1 _8359_ (
    .A(_2917_),
    .B(_3071_),
    .Z(_3074_)
  );
  AND2_X1 _8360_ (
    .A1(_2915_),
    .A2(_3074_),
    .ZN(_3075_)
  );
  XOR2_X1 _8361_ (
    .A(_2915_),
    .B(_3074_),
    .Z(_3076_)
  );
  AND2_X1 _8362_ (
    .A1(_3069_),
    .A2(_3076_),
    .ZN(_3077_)
  );
  XOR2_X1 _8363_ (
    .A(_3069_),
    .B(_3076_),
    .Z(_3079_)
  );
  AND2_X1 _8364_ (
    .A1(_3068_),
    .A2(_3079_),
    .ZN(_3080_)
  );
  XOR2_X1 _8365_ (
    .A(_3068_),
    .B(_3079_),
    .Z(_3081_)
  );
  AND2_X1 _8366_ (
    .A1(_3066_),
    .A2(_3081_),
    .ZN(_3082_)
  );
  XOR2_X1 _8367_ (
    .A(_3066_),
    .B(_3081_),
    .Z(_3083_)
  );
  AND2_X1 _8368_ (
    .A1(_2931_),
    .A2(_3083_),
    .ZN(_3084_)
  );
  XOR2_X1 _8369_ (
    .A(_2931_),
    .B(_3083_),
    .Z(_3085_)
  );
  AND2_X1 _8370_ (
    .A1(_2959_),
    .A2(_3085_),
    .ZN(_3086_)
  );
  XOR2_X1 _8371_ (
    .A(_2959_),
    .B(_3085_),
    .Z(_3087_)
  );
  AND2_X1 _8372_ (
    .A1(_3065_),
    .A2(_3087_),
    .ZN(_3088_)
  );
  XOR2_X1 _8373_ (
    .A(_3065_),
    .B(_3087_),
    .Z(_3090_)
  );
  AND2_X1 _8374_ (
    .A1(_3064_),
    .A2(_3090_),
    .ZN(_3091_)
  );
  XOR2_X1 _8375_ (
    .A(_3064_),
    .B(_3090_),
    .Z(_3092_)
  );
  AND2_X1 _8376_ (
    .A1(_3032_),
    .A2(_3092_),
    .ZN(_3093_)
  );
  XOR2_X1 _8377_ (
    .A(_3032_),
    .B(_3092_),
    .Z(_3094_)
  );
  OR2_X1 _8378_ (
    .A1(_2976_),
    .A2(_2978_),
    .ZN(_3095_)
  );
  OR2_X1 _8379_ (
    .A1(_2935_),
    .A2(_2938_),
    .ZN(_3096_)
  );
  AND2_X1 _8380_ (
    .A1(_2971_),
    .A2(_2974_),
    .ZN(_3097_)
  );
  INV_X1 _8381_ (
    .A(_3097_),
    .ZN(_3098_)
  );
  OR2_X1 _8382_ (
    .A1(_2815_),
    .A2(_2930_),
    .ZN(_3099_)
  );
  OR2_X1 _8383_ (
    .A1(_2613_),
    .A2(_3099_),
    .ZN(_3101_)
  );
  XOR2_X1 _8384_ (
    .A(_2613_),
    .B(_3099_),
    .Z(_3102_)
  );
  XOR2_X1 _8385_ (
    .A(_2733_),
    .B(_3102_),
    .Z(_3103_)
  );
  AND2_X1 _8386_ (
    .A1(_3098_),
    .A2(_3103_),
    .ZN(_3104_)
  );
  INV_X1 _8387_ (
    .A(_3104_),
    .ZN(_3105_)
  );
  XOR2_X1 _8388_ (
    .A(_3098_),
    .B(_3103_),
    .Z(_3106_)
  );
  AND2_X1 _8389_ (
    .A1(_2025_),
    .A2(_3106_),
    .ZN(_3107_)
  );
  XOR2_X1 _8390_ (
    .A(_2025_),
    .B(_3106_),
    .Z(_3108_)
  );
  AND2_X1 _8391_ (
    .A1(_3096_),
    .A2(_3108_),
    .ZN(_3109_)
  );
  XOR2_X1 _8392_ (
    .A(_3096_),
    .B(_3108_),
    .Z(_3110_)
  );
  AND2_X1 _8393_ (
    .A1(_3095_),
    .A2(_3110_),
    .ZN(_3112_)
  );
  XOR2_X1 _8394_ (
    .A(_3095_),
    .B(_3110_),
    .Z(_3113_)
  );
  AND2_X1 _8395_ (
    .A1(_3094_),
    .A2(_3113_),
    .ZN(_3114_)
  );
  XOR2_X1 _8396_ (
    .A(_3094_),
    .B(_3113_),
    .Z(_3115_)
  );
  AND2_X1 _8397_ (
    .A1(_3029_),
    .A2(_3115_),
    .ZN(_3116_)
  );
  XOR2_X1 _8398_ (
    .A(_3029_),
    .B(_3115_),
    .Z(_3117_)
  );
  OR2_X1 _8399_ (
    .A1(_2981_),
    .A2(_2983_),
    .ZN(_3118_)
  );
  AND2_X1 _8400_ (
    .A1(_2287_),
    .A2(_3118_),
    .ZN(_3119_)
  );
  XOR2_X1 _8401_ (
    .A(_2288_),
    .B(_3118_),
    .Z(_3120_)
  );
  OR2_X1 _8402_ (
    .A1(_2400_),
    .A2(_3120_),
    .ZN(_3121_)
  );
  INV_X1 _8403_ (
    .A(_3121_),
    .ZN(_3123_)
  );
  XOR2_X1 _8404_ (
    .A(_2400_),
    .B(_3120_),
    .Z(_3124_)
  );
  AND2_X1 _8405_ (
    .A1(_3117_),
    .A2(_3124_),
    .ZN(_3125_)
  );
  XOR2_X1 _8406_ (
    .A(_3117_),
    .B(_3124_),
    .Z(_3126_)
  );
  AND2_X1 _8407_ (
    .A1(_3028_),
    .A2(_3126_),
    .ZN(_3127_)
  );
  XOR2_X1 _8408_ (
    .A(_3028_),
    .B(_3126_),
    .Z(_3128_)
  );
  AND2_X1 _8409_ (
    .A1(_3027_),
    .A2(_3128_),
    .ZN(_3129_)
  );
  XOR2_X1 _8410_ (
    .A(_3027_),
    .B(_3128_),
    .Z(_3130_)
  );
  AND2_X1 _8411_ (
    .A1(_3026_),
    .A2(_3130_),
    .ZN(_3131_)
  );
  XOR2_X1 _8412_ (
    .A(_3026_),
    .B(_3130_),
    .Z(_3132_)
  );
  AND2_X1 _8413_ (
    .A1(_3003_),
    .A2(_3132_),
    .ZN(_3134_)
  );
  XOR2_X1 _8414_ (
    .A(_3003_),
    .B(_3132_),
    .Z(_3135_)
  );
  OR2_X1 _8415_ (
    .A1(_3005_),
    .A2(_3007_),
    .ZN(_3136_)
  );
  AND2_X1 _8416_ (
    .A1(_3135_),
    .A2(_3136_),
    .ZN(_3137_)
  );
  XOR2_X1 _8417_ (
    .A(_3135_),
    .B(_3136_),
    .Z(_3138_)
  );
  AND2_X1 _8418_ (
    .A1(remainder[65]),
    .A2(_3138_),
    .ZN(_3139_)
  );
  INV_X1 _8419_ (
    .A(_3139_),
    .ZN(_3140_)
  );
  XOR2_X1 _8420_ (
    .A(remainder[65]),
    .B(_3138_),
    .Z(_3141_)
  );
  INV_X1 _8421_ (
    .A(_3141_),
    .ZN(_3142_)
  );
  OR2_X1 _8422_ (
    .A1(_3025_),
    .A2(_3142_),
    .ZN(_3143_)
  );
  INV_X1 _8423_ (
    .A(_3143_),
    .ZN(_3145_)
  );
  OR2_X1 _8424_ (
    .A1(_3024_),
    .A2(_3141_),
    .ZN(_3146_)
  );
  AND2_X1 _8425_ (
    .A1(_4613_),
    .A2(_3146_),
    .ZN(_3147_)
  );
  AND2_X1 _8426_ (
    .A1(_3143_),
    .A2(_3147_),
    .ZN(_3148_)
  );
  AND2_X1 _8427_ (
    .A1(remainder[59]),
    .A2(_4610_),
    .ZN(_3149_)
  );
  OR2_X1 _8428_ (
    .A1(remainder[58]),
    .A2(_4393_),
    .ZN(_3150_)
  );
  OR2_X1 _8429_ (
    .A1(_4392_),
    .A2(_4572_),
    .ZN(_3151_)
  );
  AND2_X1 _8430_ (
    .A1(_3678_),
    .A2(_3151_),
    .ZN(_3152_)
  );
  AND2_X1 _8431_ (
    .A1(_3150_),
    .A2(_3152_),
    .ZN(_3153_)
  );
  OR2_X1 _8432_ (
    .A1(_3149_),
    .A2(_3153_),
    .ZN(_3154_)
  );
  OR2_X1 _8433_ (
    .A1(_3148_),
    .A2(_3154_),
    .ZN(_3156_)
  );
  AND2_X1 _8434_ (
    .A1(_3911_),
    .A2(_3156_),
    .ZN(_0080_)
  );
  AND2_X1 _8435_ (
    .A1(_3140_),
    .A2(_3143_),
    .ZN(_3157_)
  );
  OR2_X1 _8436_ (
    .A1(_3139_),
    .A2(_3145_),
    .ZN(_3158_)
  );
  OR2_X1 _8437_ (
    .A1(_3134_),
    .A2(_3137_),
    .ZN(_3159_)
  );
  OR2_X1 _8438_ (
    .A1(_3127_),
    .A2(_3129_),
    .ZN(_3160_)
  );
  OR2_X1 _8439_ (
    .A1(_3119_),
    .A2(_3123_),
    .ZN(_3161_)
  );
  OR2_X1 _8440_ (
    .A1(_3116_),
    .A2(_3125_),
    .ZN(_3162_)
  );
  OR2_X1 _8441_ (
    .A1(_3093_),
    .A2(_3114_),
    .ZN(_3163_)
  );
  OR2_X1 _8442_ (
    .A1(_3063_),
    .A2(_3091_),
    .ZN(_3164_)
  );
  AND2_X1 _8443_ (
    .A1(_0541_),
    .A2(_2941_),
    .ZN(_3166_)
  );
  AND2_X1 _8444_ (
    .A1(_0541_),
    .A2(_2942_),
    .ZN(_3167_)
  );
  AND2_X1 _8445_ (
    .A1(_0542_),
    .A2(_2943_),
    .ZN(_3168_)
  );
  XOR2_X1 _8446_ (
    .A(_0541_),
    .B(_2942_),
    .Z(_3169_)
  );
  MUX2_X1 _8447_ (
    .A(_3449_),
    .B(_3169_),
    .S(_3035_),
    .Z(_3170_)
  );
  OR2_X1 _8448_ (
    .A1(_3047_),
    .A2(_3057_),
    .ZN(_3171_)
  );
  OR2_X1 _8449_ (
    .A1(_3042_),
    .A2(_3044_),
    .ZN(_3172_)
  );
  AND2_X1 _8450_ (
    .A1(divisor[31]),
    .A2(remainder[4]),
    .ZN(_3173_)
  );
  AND2_X1 _8451_ (
    .A1(divisor[32]),
    .A2(remainder[3]),
    .ZN(_3174_)
  );
  AND2_X1 _8452_ (
    .A1(remainder[3]),
    .A2(_3040_),
    .ZN(_3175_)
  );
  MUX2_X1 _8453_ (
    .A(_3040_),
    .B(_3460_),
    .S(_3174_),
    .Z(_3177_)
  );
  AND2_X1 _8454_ (
    .A1(_3173_),
    .A2(_3177_),
    .ZN(_3178_)
  );
  XOR2_X1 _8455_ (
    .A(_3173_),
    .B(_3177_),
    .Z(_3179_)
  );
  AND2_X1 _8456_ (
    .A1(_3172_),
    .A2(_3179_),
    .ZN(_3180_)
  );
  XOR2_X1 _8457_ (
    .A(_3172_),
    .B(_3179_),
    .Z(_3181_)
  );
  AND2_X1 _8458_ (
    .A1(divisor[28]),
    .A2(remainder[7]),
    .ZN(_3182_)
  );
  AND2_X1 _8459_ (
    .A1(divisor[29]),
    .A2(remainder[6]),
    .ZN(_3183_)
  );
  AND2_X1 _8460_ (
    .A1(divisor[30]),
    .A2(remainder[6]),
    .ZN(_3184_)
  );
  AND2_X1 _8461_ (
    .A1(_3051_),
    .A2(_3183_),
    .ZN(_3185_)
  );
  XOR2_X1 _8462_ (
    .A(_3051_),
    .B(_3183_),
    .Z(_3186_)
  );
  AND2_X1 _8463_ (
    .A1(_3182_),
    .A2(_3186_),
    .ZN(_3188_)
  );
  XOR2_X1 _8464_ (
    .A(_3182_),
    .B(_3186_),
    .Z(_3189_)
  );
  AND2_X1 _8465_ (
    .A1(_3181_),
    .A2(_3189_),
    .ZN(_3190_)
  );
  XOR2_X1 _8466_ (
    .A(_3181_),
    .B(_3189_),
    .Z(_3191_)
  );
  AND2_X1 _8467_ (
    .A1(_3171_),
    .A2(_3191_),
    .ZN(_3192_)
  );
  XOR2_X1 _8468_ (
    .A(_3171_),
    .B(_3191_),
    .Z(_3193_)
  );
  AND2_X1 _8469_ (
    .A1(_3170_),
    .A2(_3193_),
    .ZN(_3194_)
  );
  XOR2_X1 _8470_ (
    .A(_3170_),
    .B(_3193_),
    .Z(_3195_)
  );
  AND2_X1 _8471_ (
    .A1(_3061_),
    .A2(_3195_),
    .ZN(_3196_)
  );
  XOR2_X1 _8472_ (
    .A(_3061_),
    .B(_3195_),
    .Z(_3197_)
  );
  OR2_X1 _8473_ (
    .A1(_3082_),
    .A2(_3084_),
    .ZN(_3199_)
  );
  OR2_X1 _8474_ (
    .A1(_3077_),
    .A2(_3080_),
    .ZN(_3200_)
  );
  OR2_X1 _8475_ (
    .A1(_3073_),
    .A2(_3075_),
    .ZN(_3201_)
  );
  OR2_X1 _8476_ (
    .A1(_3052_),
    .A2(_3054_),
    .ZN(_3202_)
  );
  MUX2_X1 _8477_ (
    .A(_3071_),
    .B(_3405_),
    .S(_3070_),
    .Z(_3203_)
  );
  AND2_X1 _8478_ (
    .A1(divisor[25]),
    .A2(_3203_),
    .ZN(_3204_)
  );
  MUX2_X1 _8479_ (
    .A(_2915_),
    .B(_3394_),
    .S(_3203_),
    .Z(_3205_)
  );
  AND2_X1 _8480_ (
    .A1(_3202_),
    .A2(_3205_),
    .ZN(_3206_)
  );
  XOR2_X1 _8481_ (
    .A(_3202_),
    .B(_3205_),
    .Z(_3207_)
  );
  AND2_X1 _8482_ (
    .A1(_3201_),
    .A2(_3207_),
    .ZN(_3208_)
  );
  XOR2_X1 _8483_ (
    .A(_3201_),
    .B(_3207_),
    .Z(_3210_)
  );
  AND2_X1 _8484_ (
    .A1(_3200_),
    .A2(_3210_),
    .ZN(_3211_)
  );
  XOR2_X1 _8485_ (
    .A(_3200_),
    .B(_3210_),
    .Z(_3212_)
  );
  AND2_X1 _8486_ (
    .A1(_2931_),
    .A2(_3212_),
    .ZN(_3213_)
  );
  XOR2_X1 _8487_ (
    .A(_2931_),
    .B(_3212_),
    .Z(_3214_)
  );
  AND2_X1 _8488_ (
    .A1(_3059_),
    .A2(_3214_),
    .ZN(_3215_)
  );
  XOR2_X1 _8489_ (
    .A(_3059_),
    .B(_3214_),
    .Z(_3216_)
  );
  AND2_X1 _8490_ (
    .A1(_3199_),
    .A2(_3216_),
    .ZN(_3217_)
  );
  XOR2_X1 _8491_ (
    .A(_3199_),
    .B(_3216_),
    .Z(_3218_)
  );
  AND2_X1 _8492_ (
    .A1(_3197_),
    .A2(_3218_),
    .ZN(_3219_)
  );
  XOR2_X1 _8493_ (
    .A(_3197_),
    .B(_3218_),
    .Z(_3221_)
  );
  AND2_X1 _8494_ (
    .A1(_3164_),
    .A2(_3221_),
    .ZN(_3222_)
  );
  XOR2_X1 _8495_ (
    .A(_3164_),
    .B(_3221_),
    .Z(_3223_)
  );
  OR2_X1 _8496_ (
    .A1(_3104_),
    .A2(_3107_),
    .ZN(_3224_)
  );
  OR2_X1 _8497_ (
    .A1(_3086_),
    .A2(_3088_),
    .ZN(_3225_)
  );
  OR2_X1 _8498_ (
    .A1(_2733_),
    .A2(_3101_),
    .ZN(_3226_)
  );
  AND2_X1 _8499_ (
    .A1(_3105_),
    .A2(_3226_),
    .ZN(_3227_)
  );
  AND2_X1 _8500_ (
    .A1(_2025_),
    .A2(_3227_),
    .ZN(_3228_)
  );
  XOR2_X1 _8501_ (
    .A(_2025_),
    .B(_3227_),
    .Z(_3229_)
  );
  AND2_X1 _8502_ (
    .A1(_3225_),
    .A2(_3229_),
    .ZN(_3230_)
  );
  XOR2_X1 _8503_ (
    .A(_3225_),
    .B(_3229_),
    .Z(_3232_)
  );
  AND2_X1 _8504_ (
    .A1(_3224_),
    .A2(_3232_),
    .ZN(_3233_)
  );
  XOR2_X1 _8505_ (
    .A(_3224_),
    .B(_3232_),
    .Z(_3234_)
  );
  AND2_X1 _8506_ (
    .A1(_3223_),
    .A2(_3234_),
    .ZN(_3235_)
  );
  XOR2_X1 _8507_ (
    .A(_3223_),
    .B(_3234_),
    .Z(_3236_)
  );
  AND2_X1 _8508_ (
    .A1(_3163_),
    .A2(_3236_),
    .ZN(_3237_)
  );
  XOR2_X1 _8509_ (
    .A(_3163_),
    .B(_3236_),
    .Z(_3238_)
  );
  OR2_X1 _8510_ (
    .A1(_3109_),
    .A2(_3112_),
    .ZN(_3239_)
  );
  AND2_X1 _8511_ (
    .A1(_2287_),
    .A2(_3239_),
    .ZN(_3240_)
  );
  XOR2_X1 _8512_ (
    .A(_2287_),
    .B(_3239_),
    .Z(_3241_)
  );
  AND2_X1 _8513_ (
    .A1(_2401_),
    .A2(_3241_),
    .ZN(_3243_)
  );
  XOR2_X1 _8514_ (
    .A(_2401_),
    .B(_3241_),
    .Z(_3244_)
  );
  AND2_X1 _8515_ (
    .A1(_3238_),
    .A2(_3244_),
    .ZN(_3245_)
  );
  XOR2_X1 _8516_ (
    .A(_3238_),
    .B(_3244_),
    .Z(_3246_)
  );
  AND2_X1 _8517_ (
    .A1(_3162_),
    .A2(_3246_),
    .ZN(_3247_)
  );
  XOR2_X1 _8518_ (
    .A(_3162_),
    .B(_3246_),
    .Z(_3248_)
  );
  AND2_X1 _8519_ (
    .A1(_3161_),
    .A2(_3248_),
    .ZN(_3249_)
  );
  XOR2_X1 _8520_ (
    .A(_3161_),
    .B(_3248_),
    .Z(_3250_)
  );
  AND2_X1 _8521_ (
    .A1(_3160_),
    .A2(_3250_),
    .ZN(_3251_)
  );
  XOR2_X1 _8522_ (
    .A(_3160_),
    .B(_3250_),
    .Z(_3252_)
  );
  AND2_X1 _8523_ (
    .A1(_3131_),
    .A2(_3252_),
    .ZN(_3254_)
  );
  XOR2_X1 _8524_ (
    .A(_3131_),
    .B(_3252_),
    .Z(_3255_)
  );
  AND2_X1 _8525_ (
    .A1(_3159_),
    .A2(_3255_),
    .ZN(_3256_)
  );
  XOR2_X1 _8526_ (
    .A(_3159_),
    .B(_3255_),
    .Z(_3257_)
  );
  AND2_X1 _8527_ (
    .A1(remainder[65]),
    .A2(_3257_),
    .ZN(_3258_)
  );
  XOR2_X1 _8528_ (
    .A(remainder[65]),
    .B(_3257_),
    .Z(_3259_)
  );
  XOR2_X1 _8529_ (
    .A(_2936_),
    .B(_3257_),
    .Z(_3260_)
  );
  OR2_X1 _8530_ (
    .A1(_3158_),
    .A2(_3259_),
    .ZN(_3261_)
  );
  OR2_X1 _8531_ (
    .A1(_3157_),
    .A2(_3260_),
    .ZN(_3262_)
  );
  AND2_X1 _8532_ (
    .A1(_4613_),
    .A2(_3262_),
    .ZN(_3263_)
  );
  AND2_X1 _8533_ (
    .A1(_3261_),
    .A2(_3263_),
    .ZN(_3265_)
  );
  AND2_X1 _8534_ (
    .A1(remainder[60]),
    .A2(_4610_),
    .ZN(_3266_)
  );
  MUX2_X1 _8535_ (
    .A(remainder[59]),
    .B(_4578_),
    .S(_4393_),
    .Z(_3267_)
  );
  AND2_X1 _8536_ (
    .A1(_3678_),
    .A2(_3267_),
    .ZN(_3268_)
  );
  OR2_X1 _8537_ (
    .A1(_3266_),
    .A2(_3268_),
    .ZN(_3269_)
  );
  OR2_X1 _8538_ (
    .A1(_3265_),
    .A2(_3269_),
    .ZN(_3270_)
  );
  AND2_X1 _8539_ (
    .A1(_3911_),
    .A2(_3270_),
    .ZN(_0081_)
  );
  AND2_X1 _8540_ (
    .A1(_3020_),
    .A2(_3141_),
    .ZN(_3271_)
  );
  OR2_X1 _8541_ (
    .A1(_3021_),
    .A2(_3142_),
    .ZN(_3272_)
  );
  AND2_X1 _8542_ (
    .A1(_3259_),
    .A2(_3271_),
    .ZN(_3273_)
  );
  OR2_X1 _8543_ (
    .A1(_3260_),
    .A2(_3272_),
    .ZN(_3275_)
  );
  OR2_X1 _8544_ (
    .A1(_3022_),
    .A2(_3139_),
    .ZN(_3276_)
  );
  OR2_X1 _8545_ (
    .A1(_3258_),
    .A2(_3276_),
    .ZN(_3277_)
  );
  INV_X1 _8546_ (
    .A(_3277_),
    .ZN(_3278_)
  );
  AND2_X1 _8547_ (
    .A1(_3275_),
    .A2(_3278_),
    .ZN(_3279_)
  );
  OR2_X1 _8548_ (
    .A1(_3273_),
    .A2(_3277_),
    .ZN(_3280_)
  );
  OR2_X1 _8549_ (
    .A1(_3247_),
    .A2(_3249_),
    .ZN(_3281_)
  );
  OR2_X1 _8550_ (
    .A1(_3240_),
    .A2(_3243_),
    .ZN(_3282_)
  );
  OR2_X1 _8551_ (
    .A1(_3237_),
    .A2(_3245_),
    .ZN(_3283_)
  );
  OR2_X1 _8552_ (
    .A1(_3222_),
    .A2(_3235_),
    .ZN(_3284_)
  );
  OR2_X1 _8553_ (
    .A1(_3196_),
    .A2(_3219_),
    .ZN(_3286_)
  );
  OR2_X1 _8554_ (
    .A1(_3166_),
    .A2(_3194_),
    .ZN(_3287_)
  );
  OR2_X1 _8555_ (
    .A1(_3180_),
    .A2(_3190_),
    .ZN(_3288_)
  );
  OR2_X1 _8556_ (
    .A1(_3175_),
    .A2(_3178_),
    .ZN(_3289_)
  );
  AND2_X1 _8557_ (
    .A1(divisor[31]),
    .A2(remainder[5]),
    .ZN(_3290_)
  );
  AND2_X1 _8558_ (
    .A1(divisor[32]),
    .A2(remainder[4]),
    .ZN(_3291_)
  );
  AND2_X1 _8559_ (
    .A1(remainder[4]),
    .A2(_3174_),
    .ZN(_3292_)
  );
  MUX2_X1 _8560_ (
    .A(_3291_),
    .B(_3471_),
    .S(_3174_),
    .Z(_3293_)
  );
  AND2_X1 _8561_ (
    .A1(_3290_),
    .A2(_3293_),
    .ZN(_3294_)
  );
  XOR2_X1 _8562_ (
    .A(_3290_),
    .B(_3293_),
    .Z(_3295_)
  );
  AND2_X1 _8563_ (
    .A1(_3289_),
    .A2(_3295_),
    .ZN(_3297_)
  );
  XOR2_X1 _8564_ (
    .A(_3289_),
    .B(_3295_),
    .Z(_3298_)
  );
  AND2_X1 _8565_ (
    .A1(divisor[29]),
    .A2(remainder[7]),
    .ZN(_3299_)
  );
  AND2_X1 _8566_ (
    .A1(divisor[30]),
    .A2(remainder[7]),
    .ZN(_3300_)
  );
  AND2_X1 _8567_ (
    .A1(_3183_),
    .A2(_3300_),
    .ZN(_3301_)
  );
  XOR2_X1 _8568_ (
    .A(_3184_),
    .B(_3299_),
    .Z(_3302_)
  );
  AND2_X1 _8569_ (
    .A1(_2367_),
    .A2(_3302_),
    .ZN(_3303_)
  );
  XOR2_X1 _8570_ (
    .A(_2367_),
    .B(_3302_),
    .Z(_3304_)
  );
  AND2_X1 _8571_ (
    .A1(_3298_),
    .A2(_3304_),
    .ZN(_3305_)
  );
  XOR2_X1 _8572_ (
    .A(_3298_),
    .B(_3304_),
    .Z(_3306_)
  );
  AND2_X1 _8573_ (
    .A1(_3288_),
    .A2(_3306_),
    .ZN(_3308_)
  );
  XOR2_X1 _8574_ (
    .A(_3288_),
    .B(_3306_),
    .Z(_3309_)
  );
  AND2_X1 _8575_ (
    .A1(_2941_),
    .A2(_3040_),
    .ZN(_3310_)
  );
  AND2_X1 _8576_ (
    .A1(_2942_),
    .A2(_3040_),
    .ZN(_3311_)
  );
  XOR2_X1 _8577_ (
    .A(_2942_),
    .B(_3041_),
    .Z(_3312_)
  );
  INV_X1 _8578_ (
    .A(_3312_),
    .ZN(_3313_)
  );
  MUX2_X1 _8579_ (
    .A(_3313_),
    .B(_3041_),
    .S(_2941_),
    .Z(_3314_)
  );
  INV_X1 _8580_ (
    .A(_3314_),
    .ZN(_3315_)
  );
  AND2_X1 _8581_ (
    .A1(_0541_),
    .A2(_2943_),
    .ZN(_3316_)
  );
  XOR2_X1 _8582_ (
    .A(_3314_),
    .B(_3316_),
    .Z(_3317_)
  );
  AND2_X1 _8583_ (
    .A1(_3309_),
    .A2(_3317_),
    .ZN(_3319_)
  );
  XOR2_X1 _8584_ (
    .A(_3309_),
    .B(_3317_),
    .Z(_3320_)
  );
  AND2_X1 _8585_ (
    .A1(_3287_),
    .A2(_3320_),
    .ZN(_3321_)
  );
  XOR2_X1 _8586_ (
    .A(_3287_),
    .B(_3320_),
    .Z(_3322_)
  );
  OR2_X1 _8587_ (
    .A1(_3211_),
    .A2(_3213_),
    .ZN(_3323_)
  );
  OR2_X1 _8588_ (
    .A1(_3206_),
    .A2(_3208_),
    .ZN(_3324_)
  );
  OR2_X1 _8589_ (
    .A1(_3072_),
    .A2(_3204_),
    .ZN(_3325_)
  );
  OR2_X1 _8590_ (
    .A1(_3185_),
    .A2(_3188_),
    .ZN(_3326_)
  );
  AND2_X1 _8591_ (
    .A1(_3205_),
    .A2(_3326_),
    .ZN(_3327_)
  );
  XOR2_X1 _8592_ (
    .A(_3205_),
    .B(_3326_),
    .Z(_3328_)
  );
  AND2_X1 _8593_ (
    .A1(_3325_),
    .A2(_3328_),
    .ZN(_3330_)
  );
  XOR2_X1 _8594_ (
    .A(_3325_),
    .B(_3328_),
    .Z(_3331_)
  );
  AND2_X1 _8595_ (
    .A1(_3324_),
    .A2(_3331_),
    .ZN(_3332_)
  );
  XOR2_X1 _8596_ (
    .A(_3324_),
    .B(_3331_),
    .Z(_3333_)
  );
  AND2_X1 _8597_ (
    .A1(_2931_),
    .A2(_3333_),
    .ZN(_3334_)
  );
  XOR2_X1 _8598_ (
    .A(_2931_),
    .B(_3333_),
    .Z(_3335_)
  );
  AND2_X1 _8599_ (
    .A1(_3192_),
    .A2(_3335_),
    .ZN(_3336_)
  );
  XOR2_X1 _8600_ (
    .A(_3192_),
    .B(_3335_),
    .Z(_3337_)
  );
  AND2_X1 _8601_ (
    .A1(_3323_),
    .A2(_3337_),
    .ZN(_3338_)
  );
  XOR2_X1 _8602_ (
    .A(_3323_),
    .B(_3337_),
    .Z(_3339_)
  );
  AND2_X1 _8603_ (
    .A1(_3322_),
    .A2(_3339_),
    .ZN(_3341_)
  );
  XOR2_X1 _8604_ (
    .A(_3322_),
    .B(_3339_),
    .Z(_3342_)
  );
  AND2_X1 _8605_ (
    .A1(_3286_),
    .A2(_3342_),
    .ZN(_3343_)
  );
  XOR2_X1 _8606_ (
    .A(_3286_),
    .B(_3342_),
    .Z(_3344_)
  );
  OR2_X1 _8607_ (
    .A1(_3104_),
    .A2(_3228_),
    .ZN(_3345_)
  );
  OR2_X1 _8608_ (
    .A1(_3215_),
    .A2(_3217_),
    .ZN(_3346_)
  );
  AND2_X1 _8609_ (
    .A1(_3229_),
    .A2(_3346_),
    .ZN(_3347_)
  );
  XOR2_X1 _8610_ (
    .A(_3229_),
    .B(_3346_),
    .Z(_3348_)
  );
  AND2_X1 _8611_ (
    .A1(_3345_),
    .A2(_3348_),
    .ZN(_3349_)
  );
  XOR2_X1 _8612_ (
    .A(_3345_),
    .B(_3348_),
    .Z(_3350_)
  );
  AND2_X1 _8613_ (
    .A1(_3344_),
    .A2(_3350_),
    .ZN(_3352_)
  );
  XOR2_X1 _8614_ (
    .A(_3344_),
    .B(_3350_),
    .Z(_3353_)
  );
  AND2_X1 _8615_ (
    .A1(_3284_),
    .A2(_3353_),
    .ZN(_3354_)
  );
  XOR2_X1 _8616_ (
    .A(_3284_),
    .B(_3353_),
    .Z(_3355_)
  );
  OR2_X1 _8617_ (
    .A1(_3230_),
    .A2(_3233_),
    .ZN(_3356_)
  );
  AND2_X1 _8618_ (
    .A1(_2287_),
    .A2(_3356_),
    .ZN(_3357_)
  );
  XOR2_X1 _8619_ (
    .A(_2287_),
    .B(_3356_),
    .Z(_3358_)
  );
  AND2_X1 _8620_ (
    .A1(_2401_),
    .A2(_3358_),
    .ZN(_3359_)
  );
  XOR2_X1 _8621_ (
    .A(_2401_),
    .B(_3358_),
    .Z(_3360_)
  );
  AND2_X1 _8622_ (
    .A1(_3355_),
    .A2(_3360_),
    .ZN(_3361_)
  );
  XOR2_X1 _8623_ (
    .A(_3355_),
    .B(_3360_),
    .Z(_3363_)
  );
  AND2_X1 _8624_ (
    .A1(_3283_),
    .A2(_3363_),
    .ZN(_3364_)
  );
  XOR2_X1 _8625_ (
    .A(_3283_),
    .B(_3363_),
    .Z(_3365_)
  );
  AND2_X1 _8626_ (
    .A1(_3282_),
    .A2(_3365_),
    .ZN(_3366_)
  );
  XOR2_X1 _8627_ (
    .A(_3282_),
    .B(_3365_),
    .Z(_3367_)
  );
  AND2_X1 _8628_ (
    .A1(_3281_),
    .A2(_3367_),
    .ZN(_3368_)
  );
  XOR2_X1 _8629_ (
    .A(_3281_),
    .B(_3367_),
    .Z(_3369_)
  );
  AND2_X1 _8630_ (
    .A1(_3251_),
    .A2(_3369_),
    .ZN(_3370_)
  );
  XOR2_X1 _8631_ (
    .A(_3251_),
    .B(_3369_),
    .Z(_3371_)
  );
  OR2_X1 _8632_ (
    .A1(_3254_),
    .A2(_3256_),
    .ZN(_3372_)
  );
  AND2_X1 _8633_ (
    .A1(_3371_),
    .A2(_3372_),
    .ZN(_3374_)
  );
  XOR2_X1 _8634_ (
    .A(_3371_),
    .B(_3372_),
    .Z(_3375_)
  );
  AND2_X1 _8635_ (
    .A1(remainder[65]),
    .A2(_3375_),
    .ZN(_3376_)
  );
  INV_X1 _8636_ (
    .A(_3376_),
    .ZN(_3377_)
  );
  XOR2_X1 _8637_ (
    .A(remainder[65]),
    .B(_3375_),
    .Z(_3378_)
  );
  INV_X1 _8638_ (
    .A(_3378_),
    .ZN(_3379_)
  );
  AND2_X1 _8639_ (
    .A1(_3280_),
    .A2(_3378_),
    .ZN(_3380_)
  );
  OR2_X1 _8640_ (
    .A1(_3279_),
    .A2(_3379_),
    .ZN(_3381_)
  );
  XOR2_X1 _8641_ (
    .A(_3280_),
    .B(_3378_),
    .Z(_3382_)
  );
  AND2_X1 _8642_ (
    .A1(_4613_),
    .A2(_3382_),
    .ZN(_3383_)
  );
  AND2_X1 _8643_ (
    .A1(remainder[61]),
    .A2(_4610_),
    .ZN(_3385_)
  );
  OR2_X1 _8644_ (
    .A1(remainder[60]),
    .A2(_4393_),
    .ZN(_3386_)
  );
  OR2_X1 _8645_ (
    .A1(_4392_),
    .A2(_4583_),
    .ZN(_3387_)
  );
  AND2_X1 _8646_ (
    .A1(_3678_),
    .A2(_3387_),
    .ZN(_3388_)
  );
  AND2_X1 _8647_ (
    .A1(_3386_),
    .A2(_3388_),
    .ZN(_3389_)
  );
  OR2_X1 _8648_ (
    .A1(_3385_),
    .A2(_3389_),
    .ZN(_3390_)
  );
  OR2_X1 _8649_ (
    .A1(_3383_),
    .A2(_3390_),
    .ZN(_3391_)
  );
  AND2_X1 _8650_ (
    .A1(_3911_),
    .A2(_3391_),
    .ZN(_0082_)
  );
  OR2_X1 _8651_ (
    .A1(_3376_),
    .A2(_3380_),
    .ZN(_3392_)
  );
  OR2_X1 _8652_ (
    .A1(_3370_),
    .A2(_3374_),
    .ZN(_3393_)
  );
  OR2_X1 _8653_ (
    .A1(_3364_),
    .A2(_3366_),
    .ZN(_3395_)
  );
  OR2_X1 _8654_ (
    .A1(_3357_),
    .A2(_3359_),
    .ZN(_3396_)
  );
  OR2_X1 _8655_ (
    .A1(_3354_),
    .A2(_3361_),
    .ZN(_3397_)
  );
  OR2_X1 _8656_ (
    .A1(_3343_),
    .A2(_3352_),
    .ZN(_3398_)
  );
  OR2_X1 _8657_ (
    .A1(_3321_),
    .A2(_3341_),
    .ZN(_3399_)
  );
  AND2_X1 _8658_ (
    .A1(_3167_),
    .A2(_3315_),
    .ZN(_3400_)
  );
  OR2_X1 _8659_ (
    .A1(_3319_),
    .A2(_3400_),
    .ZN(_3401_)
  );
  AND2_X1 _8660_ (
    .A1(_0541_),
    .A2(_3314_),
    .ZN(_3402_)
  );
  OR2_X1 _8661_ (
    .A1(_2941_),
    .A2(_3311_),
    .ZN(_3403_)
  );
  AND2_X1 _8662_ (
    .A1(_3043_),
    .A2(_3174_),
    .ZN(_3404_)
  );
  XOR2_X1 _8663_ (
    .A(_3043_),
    .B(_3174_),
    .Z(_3406_)
  );
  AND2_X1 _8664_ (
    .A1(_3403_),
    .A2(_3406_),
    .ZN(_3407_)
  );
  XOR2_X1 _8665_ (
    .A(_3403_),
    .B(_3406_),
    .Z(_3408_)
  );
  AND2_X1 _8666_ (
    .A1(_3036_),
    .A2(_3408_),
    .ZN(_3409_)
  );
  XOR2_X1 _8667_ (
    .A(_3036_),
    .B(_3408_),
    .Z(_3410_)
  );
  AND2_X1 _8668_ (
    .A1(_3402_),
    .A2(_3410_),
    .ZN(_3411_)
  );
  XOR2_X1 _8669_ (
    .A(_3402_),
    .B(_3410_),
    .Z(_3412_)
  );
  OR2_X1 _8670_ (
    .A1(_3297_),
    .A2(_3305_),
    .ZN(_3413_)
  );
  OR2_X1 _8671_ (
    .A1(_3292_),
    .A2(_3294_),
    .ZN(_3414_)
  );
  AND2_X1 _8672_ (
    .A1(divisor[31]),
    .A2(remainder[6]),
    .ZN(_3415_)
  );
  AND2_X1 _8673_ (
    .A1(divisor[32]),
    .A2(remainder[5]),
    .ZN(_3417_)
  );
  AND2_X1 _8674_ (
    .A1(remainder[5]),
    .A2(_3291_),
    .ZN(_3418_)
  );
  MUX2_X1 _8675_ (
    .A(_3291_),
    .B(_3471_),
    .S(_3417_),
    .Z(_3419_)
  );
  AND2_X1 _8676_ (
    .A1(_3415_),
    .A2(_3419_),
    .ZN(_3420_)
  );
  XOR2_X1 _8677_ (
    .A(_3415_),
    .B(_3419_),
    .Z(_3421_)
  );
  AND2_X1 _8678_ (
    .A1(_3414_),
    .A2(_3421_),
    .ZN(_3422_)
  );
  XOR2_X1 _8679_ (
    .A(_3414_),
    .B(_3421_),
    .Z(_3423_)
  );
  AND2_X1 _8680_ (
    .A1(remainder[32]),
    .A2(divisor[30]),
    .ZN(_3424_)
  );
  AND2_X1 _8681_ (
    .A1(remainder[32]),
    .A2(divisor[29]),
    .ZN(_3425_)
  );
  AND2_X1 _8682_ (
    .A1(divisor[30]),
    .A2(_3425_),
    .ZN(_3426_)
  );
  AND2_X1 _8683_ (
    .A1(_3300_),
    .A2(_3425_),
    .ZN(_3428_)
  );
  XOR2_X1 _8684_ (
    .A(_3300_),
    .B(_3425_),
    .Z(_3429_)
  );
  AND2_X1 _8685_ (
    .A1(_2367_),
    .A2(_3429_),
    .ZN(_3430_)
  );
  XOR2_X1 _8686_ (
    .A(_2367_),
    .B(_3429_),
    .Z(_3431_)
  );
  AND2_X1 _8687_ (
    .A1(_3423_),
    .A2(_3431_),
    .ZN(_3432_)
  );
  XOR2_X1 _8688_ (
    .A(_3423_),
    .B(_3431_),
    .Z(_3433_)
  );
  AND2_X1 _8689_ (
    .A1(_3310_),
    .A2(_3433_),
    .ZN(_3434_)
  );
  XOR2_X1 _8690_ (
    .A(_3310_),
    .B(_3433_),
    .Z(_3435_)
  );
  AND2_X1 _8691_ (
    .A1(_3413_),
    .A2(_3435_),
    .ZN(_3436_)
  );
  XOR2_X1 _8692_ (
    .A(_3413_),
    .B(_3435_),
    .Z(_3437_)
  );
  AND2_X1 _8693_ (
    .A1(_3412_),
    .A2(_3437_),
    .ZN(_3439_)
  );
  XOR2_X1 _8694_ (
    .A(_3412_),
    .B(_3437_),
    .Z(_3440_)
  );
  AND2_X1 _8695_ (
    .A1(_3401_),
    .A2(_3440_),
    .ZN(_3441_)
  );
  XOR2_X1 _8696_ (
    .A(_3401_),
    .B(_3440_),
    .Z(_3442_)
  );
  OR2_X1 _8697_ (
    .A1(_3332_),
    .A2(_3334_),
    .ZN(_3443_)
  );
  OR2_X1 _8698_ (
    .A1(_3327_),
    .A2(_3330_),
    .ZN(_3444_)
  );
  OR2_X1 _8699_ (
    .A1(_3301_),
    .A2(_3303_),
    .ZN(_3445_)
  );
  AND2_X1 _8700_ (
    .A1(_3205_),
    .A2(_3445_),
    .ZN(_3446_)
  );
  XOR2_X1 _8701_ (
    .A(_3205_),
    .B(_3445_),
    .Z(_3447_)
  );
  AND2_X1 _8702_ (
    .A1(_3325_),
    .A2(_3447_),
    .ZN(_3448_)
  );
  XOR2_X1 _8703_ (
    .A(_3325_),
    .B(_3447_),
    .Z(_3450_)
  );
  AND2_X1 _8704_ (
    .A1(_3444_),
    .A2(_3450_),
    .ZN(_3451_)
  );
  XOR2_X1 _8705_ (
    .A(_3444_),
    .B(_3450_),
    .Z(_3452_)
  );
  AND2_X1 _8706_ (
    .A1(_2931_),
    .A2(_3452_),
    .ZN(_3453_)
  );
  XOR2_X1 _8707_ (
    .A(_2931_),
    .B(_3452_),
    .Z(_3454_)
  );
  AND2_X1 _8708_ (
    .A1(_3308_),
    .A2(_3454_),
    .ZN(_3455_)
  );
  XOR2_X1 _8709_ (
    .A(_3308_),
    .B(_3454_),
    .Z(_3456_)
  );
  AND2_X1 _8710_ (
    .A1(_3443_),
    .A2(_3456_),
    .ZN(_3457_)
  );
  XOR2_X1 _8711_ (
    .A(_3443_),
    .B(_3456_),
    .Z(_3458_)
  );
  AND2_X1 _8712_ (
    .A1(_3442_),
    .A2(_3458_),
    .ZN(_3459_)
  );
  XOR2_X1 _8713_ (
    .A(_3442_),
    .B(_3458_),
    .Z(_3461_)
  );
  AND2_X1 _8714_ (
    .A1(_3399_),
    .A2(_3461_),
    .ZN(_3462_)
  );
  XOR2_X1 _8715_ (
    .A(_3399_),
    .B(_3461_),
    .Z(_3463_)
  );
  OR2_X1 _8716_ (
    .A1(_3336_),
    .A2(_3338_),
    .ZN(_3464_)
  );
  AND2_X1 _8717_ (
    .A1(_3229_),
    .A2(_3464_),
    .ZN(_3465_)
  );
  XOR2_X1 _8718_ (
    .A(_3229_),
    .B(_3464_),
    .Z(_3466_)
  );
  AND2_X1 _8719_ (
    .A1(_3345_),
    .A2(_3466_),
    .ZN(_3467_)
  );
  XOR2_X1 _8720_ (
    .A(_3345_),
    .B(_3466_),
    .Z(_3468_)
  );
  AND2_X1 _8721_ (
    .A1(_3463_),
    .A2(_3468_),
    .ZN(_3469_)
  );
  XOR2_X1 _8722_ (
    .A(_3463_),
    .B(_3468_),
    .Z(_3470_)
  );
  AND2_X1 _8723_ (
    .A1(_3398_),
    .A2(_3470_),
    .ZN(_3472_)
  );
  XOR2_X1 _8724_ (
    .A(_3398_),
    .B(_3470_),
    .Z(_3473_)
  );
  OR2_X1 _8725_ (
    .A1(_3347_),
    .A2(_3349_),
    .ZN(_3474_)
  );
  AND2_X1 _8726_ (
    .A1(_2287_),
    .A2(_3474_),
    .ZN(_3475_)
  );
  XOR2_X1 _8727_ (
    .A(_2287_),
    .B(_3474_),
    .Z(_3476_)
  );
  AND2_X1 _8728_ (
    .A1(_2401_),
    .A2(_3476_),
    .ZN(_3477_)
  );
  XOR2_X1 _8729_ (
    .A(_2401_),
    .B(_3476_),
    .Z(_3478_)
  );
  AND2_X1 _8730_ (
    .A1(_3473_),
    .A2(_3478_),
    .ZN(_3479_)
  );
  XOR2_X1 _8731_ (
    .A(_3473_),
    .B(_3478_),
    .Z(_3480_)
  );
  AND2_X1 _8732_ (
    .A1(_3397_),
    .A2(_3480_),
    .ZN(_3481_)
  );
  XOR2_X1 _8733_ (
    .A(_3397_),
    .B(_3480_),
    .Z(_3483_)
  );
  AND2_X1 _8734_ (
    .A1(_3396_),
    .A2(_3483_),
    .ZN(_3484_)
  );
  XOR2_X1 _8735_ (
    .A(_3396_),
    .B(_3483_),
    .Z(_3485_)
  );
  AND2_X1 _8736_ (
    .A1(_3395_),
    .A2(_3485_),
    .ZN(_3486_)
  );
  XOR2_X1 _8737_ (
    .A(_3395_),
    .B(_3485_),
    .Z(_3487_)
  );
  AND2_X1 _8738_ (
    .A1(_3368_),
    .A2(_3487_),
    .ZN(_3488_)
  );
  XOR2_X1 _8739_ (
    .A(_3368_),
    .B(_3487_),
    .Z(_3489_)
  );
  INV_X1 _8740_ (
    .A(_3489_),
    .ZN(_3490_)
  );
  AND2_X1 _8741_ (
    .A1(_3393_),
    .A2(_3489_),
    .ZN(_3491_)
  );
  XOR2_X1 _8742_ (
    .A(_3393_),
    .B(_3490_),
    .Z(_3492_)
  );
  XOR2_X1 _8743_ (
    .A(_3393_),
    .B(_3489_),
    .Z(_3494_)
  );
  AND2_X1 _8744_ (
    .A1(remainder[65]),
    .A2(_3494_),
    .ZN(_3495_)
  );
  OR2_X1 _8745_ (
    .A1(_2936_),
    .A2(_3492_),
    .ZN(_3496_)
  );
  XOR2_X1 _8746_ (
    .A(_2936_),
    .B(_3492_),
    .Z(_3497_)
  );
  XOR2_X1 _8747_ (
    .A(remainder[65]),
    .B(_3492_),
    .Z(_3498_)
  );
  AND2_X1 _8748_ (
    .A1(_3392_),
    .A2(_3497_),
    .ZN(_3499_)
  );
  INV_X1 _8749_ (
    .A(_3499_),
    .ZN(_3500_)
  );
  OR2_X1 _8750_ (
    .A1(_3392_),
    .A2(_3497_),
    .ZN(_3501_)
  );
  AND2_X1 _8751_ (
    .A1(_4613_),
    .A2(_3501_),
    .ZN(_3502_)
  );
  AND2_X1 _8752_ (
    .A1(_3500_),
    .A2(_3502_),
    .ZN(_3503_)
  );
  AND2_X1 _8753_ (
    .A1(remainder[62]),
    .A2(_4610_),
    .ZN(_3505_)
  );
  OR2_X1 _8754_ (
    .A1(remainder[61]),
    .A2(_4393_),
    .ZN(_3506_)
  );
  OR2_X1 _8755_ (
    .A1(_4392_),
    .A2(_4589_),
    .ZN(_3507_)
  );
  AND2_X1 _8756_ (
    .A1(_3678_),
    .A2(_3507_),
    .ZN(_3508_)
  );
  AND2_X1 _8757_ (
    .A1(_3506_),
    .A2(_3508_),
    .ZN(_3509_)
  );
  OR2_X1 _8758_ (
    .A1(_3505_),
    .A2(_3509_),
    .ZN(_3510_)
  );
  OR2_X1 _8759_ (
    .A1(_3503_),
    .A2(_3510_),
    .ZN(_3511_)
  );
  AND2_X1 _8760_ (
    .A1(_3911_),
    .A2(_3511_),
    .ZN(_0083_)
  );
  AND2_X1 _8761_ (
    .A1(_3380_),
    .A2(_3497_),
    .ZN(_3512_)
  );
  OR2_X1 _8762_ (
    .A1(_3381_),
    .A2(_3498_),
    .ZN(_3513_)
  );
  AND2_X1 _8763_ (
    .A1(_3377_),
    .A2(_3496_),
    .ZN(_3515_)
  );
  OR2_X1 _8764_ (
    .A1(_3376_),
    .A2(_3495_),
    .ZN(_3516_)
  );
  AND2_X1 _8765_ (
    .A1(_3513_),
    .A2(_3515_),
    .ZN(_3517_)
  );
  OR2_X1 _8766_ (
    .A1(_3512_),
    .A2(_3516_),
    .ZN(_3518_)
  );
  OR2_X1 _8767_ (
    .A1(_3481_),
    .A2(_3484_),
    .ZN(_3519_)
  );
  OR2_X1 _8768_ (
    .A1(_3475_),
    .A2(_3477_),
    .ZN(_3520_)
  );
  OR2_X1 _8769_ (
    .A1(_3472_),
    .A2(_3479_),
    .ZN(_3521_)
  );
  OR2_X1 _8770_ (
    .A1(_3462_),
    .A2(_3469_),
    .ZN(_3522_)
  );
  OR2_X1 _8771_ (
    .A1(_3441_),
    .A2(_3459_),
    .ZN(_3523_)
  );
  OR2_X1 _8772_ (
    .A1(_3411_),
    .A2(_3439_),
    .ZN(_3524_)
  );
  OR2_X1 _8773_ (
    .A1(_3042_),
    .A2(_3404_),
    .ZN(_3526_)
  );
  AND2_X1 _8774_ (
    .A1(_3177_),
    .A2(_3291_),
    .ZN(_3527_)
  );
  XOR2_X1 _8775_ (
    .A(_3177_),
    .B(_3291_),
    .Z(_3528_)
  );
  AND2_X1 _8776_ (
    .A1(_3526_),
    .A2(_3528_),
    .ZN(_3529_)
  );
  XOR2_X1 _8777_ (
    .A(_3526_),
    .B(_3528_),
    .Z(_3530_)
  );
  AND2_X1 _8778_ (
    .A1(_3170_),
    .A2(_3530_),
    .ZN(_3531_)
  );
  XOR2_X1 _8779_ (
    .A(_3170_),
    .B(_3530_),
    .Z(_3532_)
  );
  AND2_X1 _8780_ (
    .A1(_3409_),
    .A2(_3532_),
    .ZN(_3533_)
  );
  XOR2_X1 _8781_ (
    .A(_3409_),
    .B(_3532_),
    .Z(_3534_)
  );
  OR2_X1 _8782_ (
    .A1(_3422_),
    .A2(_3432_),
    .ZN(_3535_)
  );
  OR2_X1 _8783_ (
    .A1(_3418_),
    .A2(_3420_),
    .ZN(_3537_)
  );
  AND2_X1 _8784_ (
    .A1(divisor[31]),
    .A2(remainder[7]),
    .ZN(_3538_)
  );
  AND2_X1 _8785_ (
    .A1(divisor[32]),
    .A2(remainder[6]),
    .ZN(_3539_)
  );
  AND2_X1 _8786_ (
    .A1(remainder[5]),
    .A2(_3539_),
    .ZN(_3540_)
  );
  MUX2_X1 _8787_ (
    .A(_3539_),
    .B(_3482_),
    .S(_3417_),
    .Z(_3541_)
  );
  AND2_X1 _8788_ (
    .A1(_3538_),
    .A2(_3541_),
    .ZN(_3542_)
  );
  XOR2_X1 _8789_ (
    .A(_3538_),
    .B(_3541_),
    .Z(_3543_)
  );
  AND2_X1 _8790_ (
    .A1(_3537_),
    .A2(_3543_),
    .ZN(_3544_)
  );
  XOR2_X1 _8791_ (
    .A(_3537_),
    .B(_3543_),
    .Z(_3545_)
  );
  MUX2_X1 _8792_ (
    .A(_3425_),
    .B(_3427_),
    .S(_3424_),
    .Z(_3546_)
  );
  AND2_X1 _8793_ (
    .A1(divisor[28]),
    .A2(_3546_),
    .ZN(_3548_)
  );
  MUX2_X1 _8794_ (
    .A(_2367_),
    .B(_3416_),
    .S(_3546_),
    .Z(_3549_)
  );
  AND2_X1 _8795_ (
    .A1(_3545_),
    .A2(_3549_),
    .ZN(_3550_)
  );
  XOR2_X1 _8796_ (
    .A(_3545_),
    .B(_3549_),
    .Z(_3551_)
  );
  AND2_X1 _8797_ (
    .A1(_3407_),
    .A2(_3551_),
    .ZN(_3552_)
  );
  XOR2_X1 _8798_ (
    .A(_3407_),
    .B(_3551_),
    .Z(_3553_)
  );
  AND2_X1 _8799_ (
    .A1(_3535_),
    .A2(_3553_),
    .ZN(_3554_)
  );
  XOR2_X1 _8800_ (
    .A(_3535_),
    .B(_3553_),
    .Z(_3555_)
  );
  AND2_X1 _8801_ (
    .A1(_3534_),
    .A2(_3555_),
    .ZN(_3556_)
  );
  XOR2_X1 _8802_ (
    .A(_3534_),
    .B(_3555_),
    .Z(_3557_)
  );
  AND2_X1 _8803_ (
    .A1(_3524_),
    .A2(_3557_),
    .ZN(_3559_)
  );
  XOR2_X1 _8804_ (
    .A(_3524_),
    .B(_3557_),
    .Z(_3560_)
  );
  OR2_X1 _8805_ (
    .A1(_3451_),
    .A2(_3453_),
    .ZN(_3561_)
  );
  OR2_X1 _8806_ (
    .A1(_3434_),
    .A2(_3436_),
    .ZN(_3562_)
  );
  OR2_X1 _8807_ (
    .A1(_3446_),
    .A2(_3448_),
    .ZN(_3563_)
  );
  OR2_X1 _8808_ (
    .A1(_3428_),
    .A2(_3430_),
    .ZN(_3564_)
  );
  AND2_X1 _8809_ (
    .A1(_3205_),
    .A2(_3564_),
    .ZN(_3565_)
  );
  XOR2_X1 _8810_ (
    .A(_3205_),
    .B(_3564_),
    .Z(_3566_)
  );
  AND2_X1 _8811_ (
    .A1(_3325_),
    .A2(_3566_),
    .ZN(_3567_)
  );
  XOR2_X1 _8812_ (
    .A(_3325_),
    .B(_3566_),
    .Z(_3568_)
  );
  AND2_X1 _8813_ (
    .A1(_3563_),
    .A2(_3568_),
    .ZN(_3570_)
  );
  XOR2_X1 _8814_ (
    .A(_3563_),
    .B(_3568_),
    .Z(_3571_)
  );
  AND2_X1 _8815_ (
    .A1(_2931_),
    .A2(_3571_),
    .ZN(_3572_)
  );
  XOR2_X1 _8816_ (
    .A(_2931_),
    .B(_3571_),
    .Z(_3573_)
  );
  AND2_X1 _8817_ (
    .A1(_3562_),
    .A2(_3573_),
    .ZN(_3574_)
  );
  XOR2_X1 _8818_ (
    .A(_3562_),
    .B(_3573_),
    .Z(_3575_)
  );
  AND2_X1 _8819_ (
    .A1(_3561_),
    .A2(_3575_),
    .ZN(_3576_)
  );
  XOR2_X1 _8820_ (
    .A(_3561_),
    .B(_3575_),
    .Z(_3577_)
  );
  AND2_X1 _8821_ (
    .A1(_3560_),
    .A2(_3577_),
    .ZN(_3578_)
  );
  XOR2_X1 _8822_ (
    .A(_3560_),
    .B(_3577_),
    .Z(_3579_)
  );
  AND2_X1 _8823_ (
    .A1(_3523_),
    .A2(_3579_),
    .ZN(_3581_)
  );
  XOR2_X1 _8824_ (
    .A(_3523_),
    .B(_3579_),
    .Z(_3582_)
  );
  OR2_X1 _8825_ (
    .A1(_3455_),
    .A2(_3457_),
    .ZN(_3583_)
  );
  AND2_X1 _8826_ (
    .A1(_3229_),
    .A2(_3583_),
    .ZN(_3584_)
  );
  XOR2_X1 _8827_ (
    .A(_3229_),
    .B(_3583_),
    .Z(_3585_)
  );
  AND2_X1 _8828_ (
    .A1(_3345_),
    .A2(_3585_),
    .ZN(_3586_)
  );
  XOR2_X1 _8829_ (
    .A(_3345_),
    .B(_3585_),
    .Z(_3587_)
  );
  AND2_X1 _8830_ (
    .A1(_3582_),
    .A2(_3587_),
    .ZN(_3588_)
  );
  XOR2_X1 _8831_ (
    .A(_3582_),
    .B(_3587_),
    .Z(_3589_)
  );
  AND2_X1 _8832_ (
    .A1(_3522_),
    .A2(_3589_),
    .ZN(_3590_)
  );
  XOR2_X1 _8833_ (
    .A(_3522_),
    .B(_3589_),
    .Z(_3592_)
  );
  OR2_X1 _8834_ (
    .A1(_3465_),
    .A2(_3467_),
    .ZN(_3593_)
  );
  AND2_X1 _8835_ (
    .A1(_2287_),
    .A2(_3593_),
    .ZN(_3594_)
  );
  XOR2_X1 _8836_ (
    .A(_2288_),
    .B(_3593_),
    .Z(_3595_)
  );
  OR2_X1 _8837_ (
    .A1(_2400_),
    .A2(_3595_),
    .ZN(_3596_)
  );
  INV_X1 _8838_ (
    .A(_3596_),
    .ZN(_3597_)
  );
  XOR2_X1 _8839_ (
    .A(_2400_),
    .B(_3595_),
    .Z(_3598_)
  );
  AND2_X1 _8840_ (
    .A1(_3592_),
    .A2(_3598_),
    .ZN(_3599_)
  );
  XOR2_X1 _8841_ (
    .A(_3592_),
    .B(_3598_),
    .Z(_3600_)
  );
  AND2_X1 _8842_ (
    .A1(_3521_),
    .A2(_3600_),
    .ZN(_3601_)
  );
  XOR2_X1 _8843_ (
    .A(_3521_),
    .B(_3600_),
    .Z(_3603_)
  );
  AND2_X1 _8844_ (
    .A1(_3520_),
    .A2(_3603_),
    .ZN(_3604_)
  );
  XOR2_X1 _8845_ (
    .A(_3520_),
    .B(_3603_),
    .Z(_3605_)
  );
  AND2_X1 _8846_ (
    .A1(_3519_),
    .A2(_3605_),
    .ZN(_3606_)
  );
  XOR2_X1 _8847_ (
    .A(_3519_),
    .B(_3605_),
    .Z(_3607_)
  );
  AND2_X1 _8848_ (
    .A1(_3486_),
    .A2(_3607_),
    .ZN(_3608_)
  );
  XOR2_X1 _8849_ (
    .A(_3486_),
    .B(_3607_),
    .Z(_3609_)
  );
  OR2_X1 _8850_ (
    .A1(_3488_),
    .A2(_3491_),
    .ZN(_3610_)
  );
  AND2_X1 _8851_ (
    .A1(_3609_),
    .A2(_3610_),
    .ZN(_3611_)
  );
  XOR2_X1 _8852_ (
    .A(_3609_),
    .B(_3610_),
    .Z(_3612_)
  );
  AND2_X1 _8853_ (
    .A1(remainder[65]),
    .A2(_3612_),
    .ZN(_3614_)
  );
  INV_X1 _8854_ (
    .A(_3614_),
    .ZN(_3615_)
  );
  XOR2_X1 _8855_ (
    .A(remainder[65]),
    .B(_3612_),
    .Z(_3616_)
  );
  XOR2_X1 _8856_ (
    .A(_2936_),
    .B(_3612_),
    .Z(_3617_)
  );
  AND2_X1 _8857_ (
    .A1(_3518_),
    .A2(_3616_),
    .ZN(_3618_)
  );
  OR2_X1 _8858_ (
    .A1(_3517_),
    .A2(_3617_),
    .ZN(_3619_)
  );
  OR2_X1 _8859_ (
    .A1(_3518_),
    .A2(_3616_),
    .ZN(_3620_)
  );
  AND2_X1 _8860_ (
    .A1(_4613_),
    .A2(_3620_),
    .ZN(_3621_)
  );
  AND2_X1 _8861_ (
    .A1(_3619_),
    .A2(_3621_),
    .ZN(_3622_)
  );
  AND2_X1 _8862_ (
    .A1(remainder[63]),
    .A2(_4610_),
    .ZN(_3623_)
  );
  OR2_X1 _8863_ (
    .A1(remainder[62]),
    .A2(_4393_),
    .ZN(_3625_)
  );
  OR2_X1 _8864_ (
    .A1(_4392_),
    .A2(_4594_),
    .ZN(_3626_)
  );
  AND2_X1 _8865_ (
    .A1(_3678_),
    .A2(_3626_),
    .ZN(_3627_)
  );
  AND2_X1 _8866_ (
    .A1(_3625_),
    .A2(_3627_),
    .ZN(_3628_)
  );
  OR2_X1 _8867_ (
    .A1(_3623_),
    .A2(_3628_),
    .ZN(_3629_)
  );
  OR2_X1 _8868_ (
    .A1(_3622_),
    .A2(_3629_),
    .ZN(_3630_)
  );
  AND2_X1 _8869_ (
    .A1(_3911_),
    .A2(_3630_),
    .ZN(_0084_)
  );
  AND2_X1 _8870_ (
    .A1(_3615_),
    .A2(_3619_),
    .ZN(_3631_)
  );
  OR2_X1 _8871_ (
    .A1(_3614_),
    .A2(_3618_),
    .ZN(_3632_)
  );
  OR2_X1 _8872_ (
    .A1(_3608_),
    .A2(_3611_),
    .ZN(_3633_)
  );
  OR2_X1 _8873_ (
    .A1(_3601_),
    .A2(_3604_),
    .ZN(_3635_)
  );
  OR2_X1 _8874_ (
    .A1(_3594_),
    .A2(_3597_),
    .ZN(_3636_)
  );
  OR2_X1 _8875_ (
    .A1(_3590_),
    .A2(_3599_),
    .ZN(_3637_)
  );
  OR2_X1 _8876_ (
    .A1(_3581_),
    .A2(_3588_),
    .ZN(_3638_)
  );
  OR2_X1 _8877_ (
    .A1(_3559_),
    .A2(_3578_),
    .ZN(_3639_)
  );
  OR2_X1 _8878_ (
    .A1(_3533_),
    .A2(_3556_),
    .ZN(_3640_)
  );
  OR2_X1 _8879_ (
    .A1(_3166_),
    .A2(_3531_),
    .ZN(_3641_)
  );
  AND2_X1 _8880_ (
    .A1(_3167_),
    .A2(_3314_),
    .ZN(_3642_)
  );
  MUX2_X1 _8881_ (
    .A(_3168_),
    .B(_3169_),
    .S(_3041_),
    .Z(_3643_)
  );
  OR2_X1 _8882_ (
    .A1(_3642_),
    .A2(_3643_),
    .ZN(_3644_)
  );
  OR2_X1 _8883_ (
    .A1(_3175_),
    .A2(_3527_),
    .ZN(_3646_)
  );
  AND2_X1 _8884_ (
    .A1(_3293_),
    .A2(_3417_),
    .ZN(_3647_)
  );
  XOR2_X1 _8885_ (
    .A(_3293_),
    .B(_3417_),
    .Z(_3648_)
  );
  AND2_X1 _8886_ (
    .A1(_2941_),
    .A2(_3648_),
    .ZN(_3649_)
  );
  XOR2_X1 _8887_ (
    .A(_2941_),
    .B(_3648_),
    .Z(_3650_)
  );
  AND2_X1 _8888_ (
    .A1(_3646_),
    .A2(_3650_),
    .ZN(_3651_)
  );
  XOR2_X1 _8889_ (
    .A(_3646_),
    .B(_3650_),
    .Z(_3652_)
  );
  AND2_X1 _8890_ (
    .A1(_3644_),
    .A2(_3652_),
    .ZN(_3653_)
  );
  XOR2_X1 _8891_ (
    .A(_3644_),
    .B(_3652_),
    .Z(_3654_)
  );
  AND2_X1 _8892_ (
    .A1(_3641_),
    .A2(_3654_),
    .ZN(_3655_)
  );
  XOR2_X1 _8893_ (
    .A(_3641_),
    .B(_3654_),
    .Z(_3657_)
  );
  OR2_X1 _8894_ (
    .A1(_3544_),
    .A2(_3550_),
    .ZN(_3658_)
  );
  OR2_X1 _8895_ (
    .A1(_3540_),
    .A2(_3542_),
    .ZN(_3659_)
  );
  AND2_X1 _8896_ (
    .A1(remainder[32]),
    .A2(divisor[31]),
    .ZN(_3660_)
  );
  AND2_X1 _8897_ (
    .A1(divisor[32]),
    .A2(remainder[7]),
    .ZN(_3661_)
  );
  AND2_X1 _8898_ (
    .A1(remainder[7]),
    .A2(_3539_),
    .ZN(_3662_)
  );
  MUX2_X1 _8899_ (
    .A(_3539_),
    .B(_3482_),
    .S(_3661_),
    .Z(_3663_)
  );
  AND2_X1 _8900_ (
    .A1(_3660_),
    .A2(_3663_),
    .ZN(_3664_)
  );
  XOR2_X1 _8901_ (
    .A(_3660_),
    .B(_3663_),
    .Z(_3665_)
  );
  AND2_X1 _8902_ (
    .A1(_3659_),
    .A2(_3665_),
    .ZN(_3666_)
  );
  XOR2_X1 _8903_ (
    .A(_3659_),
    .B(_3665_),
    .Z(_3668_)
  );
  AND2_X1 _8904_ (
    .A1(_3549_),
    .A2(_3668_),
    .ZN(_3669_)
  );
  XOR2_X1 _8905_ (
    .A(_3549_),
    .B(_3668_),
    .Z(_3670_)
  );
  AND2_X1 _8906_ (
    .A1(_3529_),
    .A2(_3670_),
    .ZN(_3671_)
  );
  XOR2_X1 _8907_ (
    .A(_3529_),
    .B(_3670_),
    .Z(_3672_)
  );
  AND2_X1 _8908_ (
    .A1(_3658_),
    .A2(_3672_),
    .ZN(_3673_)
  );
  XOR2_X1 _8909_ (
    .A(_3658_),
    .B(_3672_),
    .Z(_3674_)
  );
  AND2_X1 _8910_ (
    .A1(_3657_),
    .A2(_3674_),
    .ZN(_3675_)
  );
  XOR2_X1 _8911_ (
    .A(_3657_),
    .B(_3674_),
    .Z(_3676_)
  );
  AND2_X1 _8912_ (
    .A1(_3640_),
    .A2(_3676_),
    .ZN(_3677_)
  );
  XOR2_X1 _8913_ (
    .A(_3640_),
    .B(_3676_),
    .Z(_3679_)
  );
  OR2_X1 _8914_ (
    .A1(_3570_),
    .A2(_3572_),
    .ZN(_3680_)
  );
  OR2_X1 _8915_ (
    .A1(_3552_),
    .A2(_3554_),
    .ZN(_3681_)
  );
  OR2_X1 _8916_ (
    .A1(_3565_),
    .A2(_3567_),
    .ZN(_3682_)
  );
  INV_X1 _8917_ (
    .A(_3682_),
    .ZN(_3683_)
  );
  OR2_X1 _8918_ (
    .A1(_3426_),
    .A2(_3548_),
    .ZN(_3684_)
  );
  INV_X1 _8919_ (
    .A(_3684_),
    .ZN(_3685_)
  );
  OR2_X1 _8920_ (
    .A1(_3205_),
    .A2(_3684_),
    .ZN(_3686_)
  );
  XOR2_X1 _8921_ (
    .A(_3205_),
    .B(_3685_),
    .Z(_3687_)
  );
  XOR2_X1 _8922_ (
    .A(_3325_),
    .B(_3687_),
    .Z(_3688_)
  );
  OR2_X1 _8923_ (
    .A1(_3683_),
    .A2(_3688_),
    .ZN(_3690_)
  );
  XOR2_X1 _8924_ (
    .A(_3682_),
    .B(_3688_),
    .Z(_3691_)
  );
  OR2_X1 _8925_ (
    .A1(_2932_),
    .A2(_3691_),
    .ZN(_3692_)
  );
  XOR2_X1 _8926_ (
    .A(_2932_),
    .B(_3691_),
    .Z(_3693_)
  );
  AND2_X1 _8927_ (
    .A1(_3681_),
    .A2(_3693_),
    .ZN(_3694_)
  );
  XOR2_X1 _8928_ (
    .A(_3681_),
    .B(_3693_),
    .Z(_3695_)
  );
  AND2_X1 _8929_ (
    .A1(_3680_),
    .A2(_3695_),
    .ZN(_3696_)
  );
  XOR2_X1 _8930_ (
    .A(_3680_),
    .B(_3695_),
    .Z(_3697_)
  );
  AND2_X1 _8931_ (
    .A1(_3679_),
    .A2(_3697_),
    .ZN(_3698_)
  );
  XOR2_X1 _8932_ (
    .A(_3679_),
    .B(_3697_),
    .Z(_3699_)
  );
  AND2_X1 _8933_ (
    .A1(_3639_),
    .A2(_3699_),
    .ZN(_3701_)
  );
  XOR2_X1 _8934_ (
    .A(_3639_),
    .B(_3699_),
    .Z(_3702_)
  );
  OR2_X1 _8935_ (
    .A1(_3574_),
    .A2(_3576_),
    .ZN(_3703_)
  );
  AND2_X1 _8936_ (
    .A1(_3229_),
    .A2(_3703_),
    .ZN(_3704_)
  );
  XOR2_X1 _8937_ (
    .A(_3229_),
    .B(_3703_),
    .Z(_3705_)
  );
  AND2_X1 _8938_ (
    .A1(_3345_),
    .A2(_3705_),
    .ZN(_3706_)
  );
  XOR2_X1 _8939_ (
    .A(_3345_),
    .B(_3705_),
    .Z(_3707_)
  );
  AND2_X1 _8940_ (
    .A1(_3702_),
    .A2(_3707_),
    .ZN(_3708_)
  );
  XOR2_X1 _8941_ (
    .A(_3702_),
    .B(_3707_),
    .Z(_3709_)
  );
  AND2_X1 _8942_ (
    .A1(_3638_),
    .A2(_3709_),
    .ZN(_3710_)
  );
  XOR2_X1 _8943_ (
    .A(_3638_),
    .B(_3709_),
    .Z(_3712_)
  );
  OR2_X1 _8944_ (
    .A1(_3584_),
    .A2(_3586_),
    .ZN(_3713_)
  );
  AND2_X1 _8945_ (
    .A1(_2287_),
    .A2(_3713_),
    .ZN(_3714_)
  );
  INV_X1 _8946_ (
    .A(_3714_),
    .ZN(_3715_)
  );
  XOR2_X1 _8947_ (
    .A(_2288_),
    .B(_3713_),
    .Z(_3716_)
  );
  OR2_X1 _8948_ (
    .A1(_2400_),
    .A2(_3716_),
    .ZN(_3717_)
  );
  XOR2_X1 _8949_ (
    .A(_2400_),
    .B(_3716_),
    .Z(_3718_)
  );
  AND2_X1 _8950_ (
    .A1(_3712_),
    .A2(_3718_),
    .ZN(_3719_)
  );
  XOR2_X1 _8951_ (
    .A(_3712_),
    .B(_3718_),
    .Z(_3720_)
  );
  AND2_X1 _8952_ (
    .A1(_3637_),
    .A2(_3720_),
    .ZN(_3721_)
  );
  XOR2_X1 _8953_ (
    .A(_3637_),
    .B(_3720_),
    .Z(_3723_)
  );
  AND2_X1 _8954_ (
    .A1(_3636_),
    .A2(_3723_),
    .ZN(_3724_)
  );
  XOR2_X1 _8955_ (
    .A(_3636_),
    .B(_3723_),
    .Z(_3725_)
  );
  AND2_X1 _8956_ (
    .A1(_3635_),
    .A2(_3725_),
    .ZN(_3726_)
  );
  XOR2_X1 _8957_ (
    .A(_3635_),
    .B(_3725_),
    .Z(_3727_)
  );
  AND2_X1 _8958_ (
    .A1(_3606_),
    .A2(_3727_),
    .ZN(_3728_)
  );
  XOR2_X1 _8959_ (
    .A(_3606_),
    .B(_3727_),
    .Z(_3729_)
  );
  AND2_X1 _8960_ (
    .A1(_3633_),
    .A2(_3729_),
    .ZN(_3730_)
  );
  XOR2_X1 _8961_ (
    .A(_3633_),
    .B(_3729_),
    .Z(_3731_)
  );
  AND2_X1 _8962_ (
    .A1(remainder[65]),
    .A2(_3731_),
    .ZN(_3732_)
  );
  XOR2_X1 _8963_ (
    .A(remainder[65]),
    .B(_3731_),
    .Z(_3734_)
  );
  XOR2_X1 _8964_ (
    .A(_2936_),
    .B(_3731_),
    .Z(_3735_)
  );
  OR2_X1 _8965_ (
    .A1(_3632_),
    .A2(_3734_),
    .ZN(_3736_)
  );
  OR2_X1 _8966_ (
    .A1(_3631_),
    .A2(_3735_),
    .ZN(_3737_)
  );
  AND2_X1 _8967_ (
    .A1(_4613_),
    .A2(_3737_),
    .ZN(_3738_)
  );
  AND2_X1 _8968_ (
    .A1(_3736_),
    .A2(_3738_),
    .ZN(_3739_)
  );
  AND2_X1 _8969_ (
    .A1(remainder[64]),
    .A2(_4610_),
    .ZN(_3740_)
  );
  OR2_X1 _8970_ (
    .A1(_4392_),
    .A2(_4600_),
    .ZN(_3741_)
  );
  OR2_X1 _8971_ (
    .A1(remainder[63]),
    .A2(_4393_),
    .ZN(_3742_)
  );
  AND2_X1 _8972_ (
    .A1(_3678_),
    .A2(_3741_),
    .ZN(_3743_)
  );
  AND2_X1 _8973_ (
    .A1(_3742_),
    .A2(_3743_),
    .ZN(_3745_)
  );
  OR2_X1 _8974_ (
    .A1(_3740_),
    .A2(_3745_),
    .ZN(_3746_)
  );
  OR2_X1 _8975_ (
    .A1(_3739_),
    .A2(_3746_),
    .ZN(_3747_)
  );
  AND2_X1 _8976_ (
    .A1(_3911_),
    .A2(_3747_),
    .ZN(_0085_)
  );
  AND2_X1 _8977_ (
    .A1(_3512_),
    .A2(_3616_),
    .ZN(_3748_)
  );
  AND2_X1 _8978_ (
    .A1(_3734_),
    .A2(_3748_),
    .ZN(_3749_)
  );
  OR2_X1 _8979_ (
    .A1(_3516_),
    .A2(_3614_),
    .ZN(_3750_)
  );
  OR2_X1 _8980_ (
    .A1(_3732_),
    .A2(_3750_),
    .ZN(_3751_)
  );
  OR2_X1 _8981_ (
    .A1(_3749_),
    .A2(_3751_),
    .ZN(_3752_)
  );
  OR2_X1 _8982_ (
    .A1(_3728_),
    .A2(_3730_),
    .ZN(_3753_)
  );
  OR2_X1 _8983_ (
    .A1(_3721_),
    .A2(_3724_),
    .ZN(_3755_)
  );
  AND2_X1 _8984_ (
    .A1(_3715_),
    .A2(_3717_),
    .ZN(_3756_)
  );
  OR2_X1 _8985_ (
    .A1(_3710_),
    .A2(_3719_),
    .ZN(_3757_)
  );
  OR2_X1 _8986_ (
    .A1(_3677_),
    .A2(_3698_),
    .ZN(_3758_)
  );
  OR2_X1 _8987_ (
    .A1(_3655_),
    .A2(_3675_),
    .ZN(_3759_)
  );
  AND2_X1 _8988_ (
    .A1(_3690_),
    .A2(_3692_),
    .ZN(_3760_)
  );
  XOR2_X1 _8989_ (
    .A(_3759_),
    .B(_3760_),
    .Z(_3761_)
  );
  OR2_X1 _8990_ (
    .A1(_3400_),
    .A2(_3653_),
    .ZN(_3762_)
  );
  OR2_X1 _8991_ (
    .A1(_3666_),
    .A2(_3669_),
    .ZN(_3763_)
  );
  OR2_X1 _8992_ (
    .A1(_3325_),
    .A2(_3686_),
    .ZN(_3764_)
  );
  AND2_X1 _8993_ (
    .A1(_3690_),
    .A2(_3764_),
    .ZN(_3766_)
  );
  XOR2_X1 _8994_ (
    .A(_2931_),
    .B(_3763_),
    .Z(_3767_)
  );
  XOR2_X1 _8995_ (
    .A(_3762_),
    .B(_3767_),
    .Z(_3768_)
  );
  XOR2_X1 _8996_ (
    .A(_3766_),
    .B(_3768_),
    .Z(_3769_)
  );
  OR2_X1 _8997_ (
    .A1(_3671_),
    .A2(_3673_),
    .ZN(_3770_)
  );
  OR2_X1 _8998_ (
    .A1(_0542_),
    .A2(_3312_),
    .ZN(_3771_)
  );
  OR2_X1 _8999_ (
    .A1(_3292_),
    .A2(_3647_),
    .ZN(_3772_)
  );
  XOR2_X1 _9000_ (
    .A(_3771_),
    .B(_3772_),
    .Z(_3773_)
  );
  OR2_X1 _9001_ (
    .A1(_3649_),
    .A2(_3651_),
    .ZN(_3774_)
  );
  XOR2_X1 _9002_ (
    .A(_3773_),
    .B(_3774_),
    .Z(_3775_)
  );
  XOR2_X1 _9003_ (
    .A(_3419_),
    .B(_3539_),
    .Z(_3777_)
  );
  XOR2_X1 _9004_ (
    .A(_3406_),
    .B(_3777_),
    .Z(_3778_)
  );
  XOR2_X1 _9005_ (
    .A(_3036_),
    .B(_3403_),
    .Z(_3779_)
  );
  XOR2_X1 _9006_ (
    .A(_3778_),
    .B(_3779_),
    .Z(_3780_)
  );
  OR2_X1 _9007_ (
    .A1(_3662_),
    .A2(_3664_),
    .ZN(_3781_)
  );
  XOR2_X1 _9008_ (
    .A(remainder[32]),
    .B(remainder[7]),
    .Z(_3782_)
  );
  AND2_X1 _9009_ (
    .A1(divisor[32]),
    .A2(_3782_),
    .ZN(_3783_)
  );
  XOR2_X1 _9010_ (
    .A(_3781_),
    .B(_3783_),
    .Z(_3784_)
  );
  XOR2_X1 _9011_ (
    .A(_3549_),
    .B(_3660_),
    .Z(_3785_)
  );
  XOR2_X1 _9012_ (
    .A(_3784_),
    .B(_3785_),
    .Z(_3786_)
  );
  XOR2_X1 _9013_ (
    .A(_3780_),
    .B(_3786_),
    .Z(_3788_)
  );
  XOR2_X1 _9014_ (
    .A(_3775_),
    .B(_3788_),
    .Z(_3789_)
  );
  XOR2_X1 _9015_ (
    .A(_3770_),
    .B(_3789_),
    .Z(_3790_)
  );
  XOR2_X1 _9016_ (
    .A(_3769_),
    .B(_3790_),
    .Z(_3791_)
  );
  XOR2_X1 _9017_ (
    .A(_3761_),
    .B(_3791_),
    .Z(_3792_)
  );
  XOR2_X1 _9018_ (
    .A(_3758_),
    .B(_3792_),
    .Z(_3793_)
  );
  OR2_X1 _9019_ (
    .A1(_3694_),
    .A2(_3696_),
    .ZN(_3794_)
  );
  XOR2_X1 _9020_ (
    .A(_3229_),
    .B(_3794_),
    .Z(_3795_)
  );
  XOR2_X1 _9021_ (
    .A(_3345_),
    .B(_3795_),
    .Z(_3796_)
  );
  XOR2_X1 _9022_ (
    .A(_3793_),
    .B(_3796_),
    .Z(_3797_)
  );
  MUX2_X1 _9023_ (
    .A(_0512_),
    .B(_2286_),
    .S(_2170_),
    .Z(_3799_)
  );
  XOR2_X1 _9024_ (
    .A(_3797_),
    .B(_3799_),
    .Z(_3800_)
  );
  OR2_X1 _9025_ (
    .A1(_3701_),
    .A2(_3708_),
    .ZN(_3801_)
  );
  OR2_X1 _9026_ (
    .A1(_3704_),
    .A2(_3706_),
    .ZN(_3802_)
  );
  XOR2_X1 _9027_ (
    .A(_3801_),
    .B(_3802_),
    .Z(_3803_)
  );
  XOR2_X1 _9028_ (
    .A(_3800_),
    .B(_3803_),
    .Z(_3804_)
  );
  XOR2_X1 _9029_ (
    .A(_3757_),
    .B(_3804_),
    .Z(_3805_)
  );
  XOR2_X1 _9030_ (
    .A(_3756_),
    .B(_3805_),
    .Z(_3806_)
  );
  XOR2_X1 _9031_ (
    .A(_3755_),
    .B(_3806_),
    .Z(_3807_)
  );
  XOR2_X1 _9032_ (
    .A(remainder[65]),
    .B(_3726_),
    .Z(_3808_)
  );
  XOR2_X1 _9033_ (
    .A(_3807_),
    .B(_3808_),
    .Z(_3810_)
  );
  XOR2_X1 _9034_ (
    .A(_3753_),
    .B(_3810_),
    .Z(_3811_)
  );
  XOR2_X1 _9035_ (
    .A(_3752_),
    .B(_3811_),
    .Z(_3812_)
  );
  OR2_X1 _9036_ (
    .A1(_3829_),
    .A2(_3812_),
    .ZN(_3813_)
  );
  AND2_X1 _9037_ (
    .A1(_3829_),
    .A2(_4609_),
    .ZN(_3814_)
  );
  AND2_X1 _9038_ (
    .A1(_3689_),
    .A2(_3911_),
    .ZN(_3815_)
  );
  AND2_X1 _9039_ (
    .A1(remainder[65]),
    .A2(_4608_),
    .ZN(_3816_)
  );
  OR2_X1 _9040_ (
    .A1(_3819_),
    .A2(_3816_),
    .ZN(_3817_)
  );
  AND2_X1 _9041_ (
    .A1(_3815_),
    .A2(_3817_),
    .ZN(_3818_)
  );
  AND2_X1 _9042_ (
    .A1(_3813_),
    .A2(_3818_),
    .ZN(_0086_)
  );
  AND2_X1 _9043_ (
    .A1(remainder[8]),
    .A2(_3819_),
    .ZN(_3820_)
  );
  MUX2_X1 _9044_ (
    .A(remainder[0]),
    .B(remainder[33]),
    .S(resHi),
    .Z(io_resp_bits_data[0])
  );
  AND2_X1 _9045_ (
    .A1(_3814_),
    .A2(io_resp_bits_data[0]),
    .ZN(_3821_)
  );
  OR2_X1 _9046_ (
    .A1(_3820_),
    .A2(_3821_),
    .ZN(_3822_)
  );
  MUX2_X1 _9047_ (
    .A(_4393_),
    .B(_3822_),
    .S(_3689_),
    .Z(_3823_)
  );
  AND2_X1 _9048_ (
    .A1(_3911_),
    .A2(_3823_),
    .ZN(_3824_)
  );
  AND2_X1 _9049_ (
    .A1(io_req_bits_in1[0]),
    .A2(_3902_),
    .ZN(_3825_)
  );
  AND2_X1 _9050_ (
    .A1(_3911_),
    .A2(_4610_),
    .ZN(_3826_)
  );
  AND2_X1 _9051_ (
    .A1(remainder[0]),
    .A2(_3826_),
    .ZN(_3827_)
  );
  OR2_X1 _9052_ (
    .A1(_3825_),
    .A2(_3827_),
    .ZN(_3828_)
  );
  OR2_X1 _9053_ (
    .A1(_3824_),
    .A2(_3828_),
    .ZN(_0087_)
  );
  AND2_X1 _9054_ (
    .A1(remainder[1]),
    .A2(_3826_),
    .ZN(_3830_)
  );
  MUX2_X1 _9055_ (
    .A(remainder[1]),
    .B(remainder[34]),
    .S(resHi),
    .Z(io_resp_bits_data[1])
  );
  OR2_X1 _9056_ (
    .A1(io_resp_bits_data[0]),
    .A2(io_resp_bits_data[1]),
    .ZN(_3831_)
  );
  XOR2_X1 _9057_ (
    .A(io_resp_bits_data[0]),
    .B(io_resp_bits_data[1]),
    .Z(_3832_)
  );
  AND2_X1 _9058_ (
    .A1(_3814_),
    .A2(_3832_),
    .ZN(_3833_)
  );
  AND2_X1 _9059_ (
    .A1(remainder[9]),
    .A2(_3819_),
    .ZN(_3834_)
  );
  OR2_X1 _9060_ (
    .A1(_3833_),
    .A2(_3834_),
    .ZN(_3835_)
  );
  MUX2_X1 _9061_ (
    .A(remainder[0]),
    .B(_3835_),
    .S(_3689_),
    .Z(_3836_)
  );
  MUX2_X1 _9062_ (
    .A(io_req_bits_in1[1]),
    .B(_3836_),
    .S(_3911_),
    .Z(_3837_)
  );
  OR2_X1 _9063_ (
    .A1(_3830_),
    .A2(_3837_),
    .ZN(_0088_)
  );
  AND2_X1 _9064_ (
    .A1(remainder[2]),
    .A2(_3826_),
    .ZN(_3839_)
  );
  AND2_X1 _9065_ (
    .A1(remainder[10]),
    .A2(_3819_),
    .ZN(_3840_)
  );
  OR2_X1 _9066_ (
    .A1(_3678_),
    .A2(_3840_),
    .ZN(_3841_)
  );
  MUX2_X1 _9067_ (
    .A(remainder[2]),
    .B(remainder[35]),
    .S(resHi),
    .Z(io_resp_bits_data[2])
  );
  OR2_X1 _9068_ (
    .A1(_3831_),
    .A2(io_resp_bits_data[2]),
    .ZN(_3842_)
  );
  XOR2_X1 _9069_ (
    .A(_3831_),
    .B(io_resp_bits_data[2]),
    .Z(_3843_)
  );
  AND2_X1 _9070_ (
    .A1(_3814_),
    .A2(_3843_),
    .ZN(_3844_)
  );
  OR2_X1 _9071_ (
    .A1(_3841_),
    .A2(_3844_),
    .ZN(_3845_)
  );
  OR2_X1 _9072_ (
    .A1(remainder[1]),
    .A2(_3689_),
    .ZN(_3846_)
  );
  AND2_X1 _9073_ (
    .A1(_3845_),
    .A2(_3846_),
    .ZN(_3848_)
  );
  MUX2_X1 _9074_ (
    .A(io_req_bits_in1[2]),
    .B(_3848_),
    .S(_3911_),
    .Z(_3849_)
  );
  OR2_X1 _9075_ (
    .A1(_3839_),
    .A2(_3849_),
    .ZN(_0089_)
  );
  AND2_X1 _9076_ (
    .A1(remainder[3]),
    .A2(_3826_),
    .ZN(_3850_)
  );
  AND2_X1 _9077_ (
    .A1(remainder[11]),
    .A2(_3819_),
    .ZN(_3851_)
  );
  OR2_X1 _9078_ (
    .A1(_3678_),
    .A2(_3851_),
    .ZN(_3852_)
  );
  MUX2_X1 _9079_ (
    .A(remainder[3]),
    .B(remainder[36]),
    .S(resHi),
    .Z(io_resp_bits_data[3])
  );
  OR2_X1 _9080_ (
    .A1(_3842_),
    .A2(io_resp_bits_data[3]),
    .ZN(_3853_)
  );
  XOR2_X1 _9081_ (
    .A(_3842_),
    .B(io_resp_bits_data[3]),
    .Z(_3854_)
  );
  AND2_X1 _9082_ (
    .A1(_3814_),
    .A2(_3854_),
    .ZN(_3855_)
  );
  OR2_X1 _9083_ (
    .A1(_3852_),
    .A2(_3855_),
    .ZN(_3857_)
  );
  OR2_X1 _9084_ (
    .A1(remainder[2]),
    .A2(_3689_),
    .ZN(_3858_)
  );
  AND2_X1 _9085_ (
    .A1(_3857_),
    .A2(_3858_),
    .ZN(_3859_)
  );
  MUX2_X1 _9086_ (
    .A(io_req_bits_in1[3]),
    .B(_3859_),
    .S(_3911_),
    .Z(_3860_)
  );
  OR2_X1 _9087_ (
    .A1(_3850_),
    .A2(_3860_),
    .ZN(_0090_)
  );
  AND2_X1 _9088_ (
    .A1(remainder[4]),
    .A2(_3826_),
    .ZN(_3861_)
  );
  AND2_X1 _9089_ (
    .A1(remainder[12]),
    .A2(_3819_),
    .ZN(_3862_)
  );
  OR2_X1 _9090_ (
    .A1(_3678_),
    .A2(_3862_),
    .ZN(_3863_)
  );
  MUX2_X1 _9091_ (
    .A(remainder[4]),
    .B(remainder[37]),
    .S(resHi),
    .Z(io_resp_bits_data[4])
  );
  OR2_X1 _9092_ (
    .A1(_3853_),
    .A2(io_resp_bits_data[4]),
    .ZN(_3864_)
  );
  XOR2_X1 _9093_ (
    .A(_3853_),
    .B(io_resp_bits_data[4]),
    .Z(_3866_)
  );
  AND2_X1 _9094_ (
    .A1(_3814_),
    .A2(_3866_),
    .ZN(_3867_)
  );
  OR2_X1 _9095_ (
    .A1(_3863_),
    .A2(_3867_),
    .ZN(_3868_)
  );
  OR2_X1 _9096_ (
    .A1(remainder[3]),
    .A2(_3689_),
    .ZN(_3869_)
  );
  AND2_X1 _9097_ (
    .A1(_3868_),
    .A2(_3869_),
    .ZN(_3870_)
  );
  MUX2_X1 _9098_ (
    .A(io_req_bits_in1[4]),
    .B(_3870_),
    .S(_3911_),
    .Z(_3871_)
  );
  OR2_X1 _9099_ (
    .A1(_3861_),
    .A2(_3871_),
    .ZN(_0091_)
  );
  AND2_X1 _9100_ (
    .A1(remainder[5]),
    .A2(_3826_),
    .ZN(_3872_)
  );
  OR2_X1 _9101_ (
    .A1(remainder[4]),
    .A2(_3689_),
    .ZN(_3873_)
  );
  AND2_X1 _9102_ (
    .A1(remainder[13]),
    .A2(_3819_),
    .ZN(_3874_)
  );
  OR2_X1 _9103_ (
    .A1(_3678_),
    .A2(_3874_),
    .ZN(_3876_)
  );
  MUX2_X1 _9104_ (
    .A(remainder[5]),
    .B(remainder[38]),
    .S(resHi),
    .Z(io_resp_bits_data[5])
  );
  OR2_X1 _9105_ (
    .A1(_3864_),
    .A2(io_resp_bits_data[5]),
    .ZN(_3877_)
  );
  XOR2_X1 _9106_ (
    .A(_3864_),
    .B(io_resp_bits_data[5]),
    .Z(_3878_)
  );
  AND2_X1 _9107_ (
    .A1(_3814_),
    .A2(_3878_),
    .ZN(_3879_)
  );
  OR2_X1 _9108_ (
    .A1(_3876_),
    .A2(_3879_),
    .ZN(_3880_)
  );
  AND2_X1 _9109_ (
    .A1(_3873_),
    .A2(_3880_),
    .ZN(_3881_)
  );
  MUX2_X1 _9110_ (
    .A(io_req_bits_in1[5]),
    .B(_3881_),
    .S(_3911_),
    .Z(_3882_)
  );
  OR2_X1 _9111_ (
    .A1(_3872_),
    .A2(_3882_),
    .ZN(_0092_)
  );
  AND2_X1 _9112_ (
    .A1(remainder[6]),
    .A2(_3826_),
    .ZN(_3883_)
  );
  AND2_X1 _9113_ (
    .A1(remainder[14]),
    .A2(_3819_),
    .ZN(_3885_)
  );
  OR2_X1 _9114_ (
    .A1(_3678_),
    .A2(_3885_),
    .ZN(_3886_)
  );
  MUX2_X1 _9115_ (
    .A(remainder[6]),
    .B(remainder[39]),
    .S(resHi),
    .Z(io_resp_bits_data[6])
  );
  OR2_X1 _9116_ (
    .A1(_3877_),
    .A2(io_resp_bits_data[6]),
    .ZN(_3887_)
  );
  XOR2_X1 _9117_ (
    .A(_3877_),
    .B(io_resp_bits_data[6]),
    .Z(_3888_)
  );
  AND2_X1 _9118_ (
    .A1(_3814_),
    .A2(_3888_),
    .ZN(_3889_)
  );
  OR2_X1 _9119_ (
    .A1(_3886_),
    .A2(_3889_),
    .ZN(_3890_)
  );
  OR2_X1 _9120_ (
    .A1(remainder[5]),
    .A2(_3689_),
    .ZN(_3891_)
  );
  AND2_X1 _9121_ (
    .A1(_3890_),
    .A2(_3891_),
    .ZN(_3892_)
  );
  MUX2_X1 _9122_ (
    .A(io_req_bits_in1[6]),
    .B(_3892_),
    .S(_3911_),
    .Z(_3893_)
  );
  OR2_X1 _9123_ (
    .A1(_3883_),
    .A2(_3893_),
    .ZN(_0093_)
  );
  AND2_X1 _9124_ (
    .A1(remainder[15]),
    .A2(_3819_),
    .ZN(_3894_)
  );
  OR2_X1 _9125_ (
    .A1(_3678_),
    .A2(_3894_),
    .ZN(_3895_)
  );
  MUX2_X1 _9126_ (
    .A(remainder[7]),
    .B(remainder[40]),
    .S(resHi),
    .Z(io_resp_bits_data[7])
  );
  OR2_X1 _9127_ (
    .A1(_3887_),
    .A2(io_resp_bits_data[7]),
    .ZN(_3896_)
  );
  XOR2_X1 _9128_ (
    .A(_3887_),
    .B(io_resp_bits_data[7]),
    .Z(_3897_)
  );
  AND2_X1 _9129_ (
    .A1(_3814_),
    .A2(_3897_),
    .ZN(_3898_)
  );
  OR2_X1 _9130_ (
    .A1(_3895_),
    .A2(_3898_),
    .ZN(_3899_)
  );
  OR2_X1 _9131_ (
    .A1(remainder[6]),
    .A2(_3689_),
    .ZN(_3900_)
  );
  AND2_X1 _9132_ (
    .A1(_3911_),
    .A2(_3900_),
    .ZN(_3901_)
  );
  AND2_X1 _9133_ (
    .A1(_3899_),
    .A2(_3901_),
    .ZN(_3903_)
  );
  AND2_X1 _9134_ (
    .A1(remainder[7]),
    .A2(_3826_),
    .ZN(_3904_)
  );
  AND2_X1 _9135_ (
    .A1(io_req_bits_in1[7]),
    .A2(_3902_),
    .ZN(_3905_)
  );
  OR2_X1 _9136_ (
    .A1(_3904_),
    .A2(_3905_),
    .ZN(_3906_)
  );
  OR2_X1 _9137_ (
    .A1(_3903_),
    .A2(_3906_),
    .ZN(_0094_)
  );
  AND2_X1 _9138_ (
    .A1(remainder[16]),
    .A2(_3819_),
    .ZN(_3907_)
  );
  OR2_X1 _9139_ (
    .A1(_3678_),
    .A2(_3907_),
    .ZN(_3908_)
  );
  MUX2_X1 _9140_ (
    .A(remainder[8]),
    .B(remainder[41]),
    .S(resHi),
    .Z(io_resp_bits_data[8])
  );
  OR2_X1 _9141_ (
    .A1(_3896_),
    .A2(io_resp_bits_data[8]),
    .ZN(_3909_)
  );
  XOR2_X1 _9142_ (
    .A(_3896_),
    .B(io_resp_bits_data[8]),
    .Z(_3910_)
  );
  AND2_X1 _9143_ (
    .A1(_3814_),
    .A2(_3910_),
    .ZN(_3912_)
  );
  OR2_X1 _9144_ (
    .A1(_3908_),
    .A2(_3912_),
    .ZN(_3913_)
  );
  OR2_X1 _9145_ (
    .A1(remainder[7]),
    .A2(_3689_),
    .ZN(_3914_)
  );
  AND2_X1 _9146_ (
    .A1(_3911_),
    .A2(_3914_),
    .ZN(_3915_)
  );
  AND2_X1 _9147_ (
    .A1(_3913_),
    .A2(_3915_),
    .ZN(_3916_)
  );
  AND2_X1 _9148_ (
    .A1(remainder[8]),
    .A2(_3826_),
    .ZN(_3917_)
  );
  AND2_X1 _9149_ (
    .A1(io_req_bits_in1[8]),
    .A2(_3902_),
    .ZN(_3918_)
  );
  OR2_X1 _9150_ (
    .A1(_3917_),
    .A2(_3918_),
    .ZN(_3919_)
  );
  OR2_X1 _9151_ (
    .A1(_3916_),
    .A2(_3919_),
    .ZN(_0095_)
  );
  AND2_X1 _9152_ (
    .A1(remainder[17]),
    .A2(_3819_),
    .ZN(_3920_)
  );
  OR2_X1 _9153_ (
    .A1(_3678_),
    .A2(_3920_),
    .ZN(_3922_)
  );
  MUX2_X1 _9154_ (
    .A(remainder[9]),
    .B(remainder[42]),
    .S(resHi),
    .Z(io_resp_bits_data[9])
  );
  OR2_X1 _9155_ (
    .A1(_3909_),
    .A2(io_resp_bits_data[9]),
    .ZN(_3923_)
  );
  XOR2_X1 _9156_ (
    .A(_3909_),
    .B(io_resp_bits_data[9]),
    .Z(_3924_)
  );
  AND2_X1 _9157_ (
    .A1(_3814_),
    .A2(_3924_),
    .ZN(_3925_)
  );
  OR2_X1 _9158_ (
    .A1(_3922_),
    .A2(_3925_),
    .ZN(_3926_)
  );
  OR2_X1 _9159_ (
    .A1(remainder[8]),
    .A2(_3689_),
    .ZN(_3927_)
  );
  AND2_X1 _9160_ (
    .A1(_3911_),
    .A2(_3927_),
    .ZN(_3928_)
  );
  AND2_X1 _9161_ (
    .A1(_3926_),
    .A2(_3928_),
    .ZN(_3929_)
  );
  AND2_X1 _9162_ (
    .A1(remainder[9]),
    .A2(_3826_),
    .ZN(_3930_)
  );
  AND2_X1 _9163_ (
    .A1(io_req_bits_in1[9]),
    .A2(_3902_),
    .ZN(_3932_)
  );
  OR2_X1 _9164_ (
    .A1(_3930_),
    .A2(_3932_),
    .ZN(_3933_)
  );
  OR2_X1 _9165_ (
    .A1(_3929_),
    .A2(_3933_),
    .ZN(_0096_)
  );
  AND2_X1 _9166_ (
    .A1(remainder[18]),
    .A2(_3819_),
    .ZN(_3934_)
  );
  OR2_X1 _9167_ (
    .A1(_3678_),
    .A2(_3934_),
    .ZN(_3935_)
  );
  MUX2_X1 _9168_ (
    .A(remainder[10]),
    .B(remainder[43]),
    .S(resHi),
    .Z(io_resp_bits_data[10])
  );
  OR2_X1 _9169_ (
    .A1(_3923_),
    .A2(io_resp_bits_data[10]),
    .ZN(_3936_)
  );
  XOR2_X1 _9170_ (
    .A(_3923_),
    .B(io_resp_bits_data[10]),
    .Z(_3937_)
  );
  AND2_X1 _9171_ (
    .A1(_3814_),
    .A2(_3937_),
    .ZN(_3938_)
  );
  OR2_X1 _9172_ (
    .A1(_3935_),
    .A2(_3938_),
    .ZN(_3939_)
  );
  OR2_X1 _9173_ (
    .A1(remainder[9]),
    .A2(_3689_),
    .ZN(_3941_)
  );
  AND2_X1 _9174_ (
    .A1(_3911_),
    .A2(_3941_),
    .ZN(_3942_)
  );
  AND2_X1 _9175_ (
    .A1(_3939_),
    .A2(_3942_),
    .ZN(_3943_)
  );
  AND2_X1 _9176_ (
    .A1(remainder[10]),
    .A2(_3826_),
    .ZN(_3944_)
  );
  AND2_X1 _9177_ (
    .A1(io_req_bits_in1[10]),
    .A2(_3902_),
    .ZN(_3945_)
  );
  OR2_X1 _9178_ (
    .A1(_3944_),
    .A2(_3945_),
    .ZN(_3946_)
  );
  OR2_X1 _9179_ (
    .A1(_3943_),
    .A2(_3946_),
    .ZN(_0097_)
  );
  AND2_X1 _9180_ (
    .A1(remainder[19]),
    .A2(_3819_),
    .ZN(_3947_)
  );
  OR2_X1 _9181_ (
    .A1(_3678_),
    .A2(_3947_),
    .ZN(_3948_)
  );
  MUX2_X1 _9182_ (
    .A(remainder[11]),
    .B(remainder[44]),
    .S(resHi),
    .Z(io_resp_bits_data[11])
  );
  OR2_X1 _9183_ (
    .A1(_3936_),
    .A2(io_resp_bits_data[11]),
    .ZN(_3950_)
  );
  XOR2_X1 _9184_ (
    .A(_3936_),
    .B(io_resp_bits_data[11]),
    .Z(_3951_)
  );
  AND2_X1 _9185_ (
    .A1(_3814_),
    .A2(_3951_),
    .ZN(_3952_)
  );
  OR2_X1 _9186_ (
    .A1(_3948_),
    .A2(_3952_),
    .ZN(_3953_)
  );
  OR2_X1 _9187_ (
    .A1(remainder[10]),
    .A2(_3689_),
    .ZN(_3954_)
  );
  AND2_X1 _9188_ (
    .A1(_3911_),
    .A2(_3954_),
    .ZN(_3955_)
  );
  AND2_X1 _9189_ (
    .A1(_3953_),
    .A2(_3955_),
    .ZN(_3956_)
  );
  AND2_X1 _9190_ (
    .A1(remainder[11]),
    .A2(_3826_),
    .ZN(_3957_)
  );
  AND2_X1 _9191_ (
    .A1(io_req_bits_in1[11]),
    .A2(_3902_),
    .ZN(_3958_)
  );
  OR2_X1 _9192_ (
    .A1(_3957_),
    .A2(_3958_),
    .ZN(_3959_)
  );
  OR2_X1 _9193_ (
    .A1(_3956_),
    .A2(_3959_),
    .ZN(_0098_)
  );
  AND2_X1 _9194_ (
    .A1(remainder[20]),
    .A2(_3819_),
    .ZN(_3961_)
  );
  OR2_X1 _9195_ (
    .A1(_3678_),
    .A2(_3961_),
    .ZN(_3962_)
  );
  MUX2_X1 _9196_ (
    .A(remainder[12]),
    .B(remainder[45]),
    .S(resHi),
    .Z(io_resp_bits_data[12])
  );
  OR2_X1 _9197_ (
    .A1(_3950_),
    .A2(io_resp_bits_data[12]),
    .ZN(_3963_)
  );
  XOR2_X1 _9198_ (
    .A(_3950_),
    .B(io_resp_bits_data[12]),
    .Z(_3964_)
  );
  AND2_X1 _9199_ (
    .A1(_3814_),
    .A2(_3964_),
    .ZN(_3965_)
  );
  OR2_X1 _9200_ (
    .A1(_3962_),
    .A2(_3965_),
    .ZN(_3966_)
  );
  OR2_X1 _9201_ (
    .A1(remainder[11]),
    .A2(_3689_),
    .ZN(_3967_)
  );
  AND2_X1 _9202_ (
    .A1(_3911_),
    .A2(_3967_),
    .ZN(_3968_)
  );
  AND2_X1 _9203_ (
    .A1(_3966_),
    .A2(_3968_),
    .ZN(_3970_)
  );
  AND2_X1 _9204_ (
    .A1(remainder[12]),
    .A2(_3826_),
    .ZN(_3971_)
  );
  AND2_X1 _9205_ (
    .A1(io_req_bits_in1[12]),
    .A2(_3902_),
    .ZN(_3972_)
  );
  OR2_X1 _9206_ (
    .A1(_3971_),
    .A2(_3972_),
    .ZN(_3973_)
  );
  OR2_X1 _9207_ (
    .A1(_3970_),
    .A2(_3973_),
    .ZN(_0099_)
  );
  AND2_X1 _9208_ (
    .A1(remainder[21]),
    .A2(_3819_),
    .ZN(_3974_)
  );
  OR2_X1 _9209_ (
    .A1(_3678_),
    .A2(_3974_),
    .ZN(_3975_)
  );
  MUX2_X1 _9210_ (
    .A(remainder[13]),
    .B(remainder[46]),
    .S(resHi),
    .Z(io_resp_bits_data[13])
  );
  OR2_X1 _9211_ (
    .A1(_3963_),
    .A2(io_resp_bits_data[13]),
    .ZN(_3976_)
  );
  XOR2_X1 _9212_ (
    .A(_3963_),
    .B(io_resp_bits_data[13]),
    .Z(_3977_)
  );
  AND2_X1 _9213_ (
    .A1(_3814_),
    .A2(_3977_),
    .ZN(_3979_)
  );
  OR2_X1 _9214_ (
    .A1(_3975_),
    .A2(_3979_),
    .ZN(_3980_)
  );
  OR2_X1 _9215_ (
    .A1(remainder[12]),
    .A2(_3689_),
    .ZN(_3981_)
  );
  AND2_X1 _9216_ (
    .A1(_3911_),
    .A2(_3981_),
    .ZN(_3982_)
  );
  AND2_X1 _9217_ (
    .A1(_3980_),
    .A2(_3982_),
    .ZN(_3983_)
  );
  AND2_X1 _9218_ (
    .A1(remainder[13]),
    .A2(_3826_),
    .ZN(_3984_)
  );
  AND2_X1 _9219_ (
    .A1(io_req_bits_in1[13]),
    .A2(_3902_),
    .ZN(_3985_)
  );
  OR2_X1 _9220_ (
    .A1(_3984_),
    .A2(_3985_),
    .ZN(_3986_)
  );
  OR2_X1 _9221_ (
    .A1(_3983_),
    .A2(_3986_),
    .ZN(_0100_)
  );
  AND2_X1 _9222_ (
    .A1(remainder[22]),
    .A2(_3819_),
    .ZN(_3987_)
  );
  OR2_X1 _9223_ (
    .A1(_3678_),
    .A2(_3987_),
    .ZN(_3989_)
  );
  MUX2_X1 _9224_ (
    .A(remainder[14]),
    .B(remainder[47]),
    .S(resHi),
    .Z(io_resp_bits_data[14])
  );
  OR2_X1 _9225_ (
    .A1(_3976_),
    .A2(io_resp_bits_data[14]),
    .ZN(_3990_)
  );
  XOR2_X1 _9226_ (
    .A(_3976_),
    .B(io_resp_bits_data[14]),
    .Z(_3991_)
  );
  AND2_X1 _9227_ (
    .A1(_3814_),
    .A2(_3991_),
    .ZN(_3992_)
  );
  OR2_X1 _9228_ (
    .A1(_3989_),
    .A2(_3992_),
    .ZN(_3993_)
  );
  OR2_X1 _9229_ (
    .A1(remainder[13]),
    .A2(_3689_),
    .ZN(_3994_)
  );
  AND2_X1 _9230_ (
    .A1(_3911_),
    .A2(_3994_),
    .ZN(_3995_)
  );
  AND2_X1 _9231_ (
    .A1(_3993_),
    .A2(_3995_),
    .ZN(_3996_)
  );
  AND2_X1 _9232_ (
    .A1(remainder[14]),
    .A2(_3826_),
    .ZN(_3997_)
  );
  AND2_X1 _9233_ (
    .A1(io_req_bits_in1[14]),
    .A2(_3902_),
    .ZN(_3998_)
  );
  OR2_X1 _9234_ (
    .A1(_3997_),
    .A2(_3998_),
    .ZN(_3999_)
  );
  OR2_X1 _9235_ (
    .A1(_3996_),
    .A2(_3999_),
    .ZN(_0101_)
  );
  AND2_X1 _9236_ (
    .A1(remainder[23]),
    .A2(_3819_),
    .ZN(_4000_)
  );
  OR2_X1 _9237_ (
    .A1(_3678_),
    .A2(_4000_),
    .ZN(_4001_)
  );
  MUX2_X1 _9238_ (
    .A(remainder[15]),
    .B(remainder[48]),
    .S(resHi),
    .Z(io_resp_bits_data[15])
  );
  OR2_X1 _9239_ (
    .A1(_3990_),
    .A2(io_resp_bits_data[15]),
    .ZN(_4002_)
  );
  XOR2_X1 _9240_ (
    .A(_3990_),
    .B(io_resp_bits_data[15]),
    .Z(_4003_)
  );
  AND2_X1 _9241_ (
    .A1(_3814_),
    .A2(_4003_),
    .ZN(_4004_)
  );
  OR2_X1 _9242_ (
    .A1(_4001_),
    .A2(_4004_),
    .ZN(_4005_)
  );
  OR2_X1 _9243_ (
    .A1(remainder[14]),
    .A2(_3689_),
    .ZN(_4007_)
  );
  AND2_X1 _9244_ (
    .A1(_3911_),
    .A2(_4007_),
    .ZN(_4008_)
  );
  AND2_X1 _9245_ (
    .A1(_4005_),
    .A2(_4008_),
    .ZN(_4009_)
  );
  AND2_X1 _9246_ (
    .A1(remainder[15]),
    .A2(_3826_),
    .ZN(_4010_)
  );
  AND2_X1 _9247_ (
    .A1(io_req_bits_in1[15]),
    .A2(_3902_),
    .ZN(_4011_)
  );
  OR2_X1 _9248_ (
    .A1(_4010_),
    .A2(_4011_),
    .ZN(_4012_)
  );
  OR2_X1 _9249_ (
    .A1(_4009_),
    .A2(_4012_),
    .ZN(_0102_)
  );
  AND2_X1 _9250_ (
    .A1(remainder[24]),
    .A2(_3819_),
    .ZN(_4013_)
  );
  OR2_X1 _9251_ (
    .A1(_3678_),
    .A2(_4013_),
    .ZN(_4014_)
  );
  MUX2_X1 _9252_ (
    .A(remainder[16]),
    .B(remainder[49]),
    .S(resHi),
    .Z(io_resp_bits_data[16])
  );
  OR2_X1 _9253_ (
    .A1(_4002_),
    .A2(io_resp_bits_data[16]),
    .ZN(_4016_)
  );
  XOR2_X1 _9254_ (
    .A(_4002_),
    .B(io_resp_bits_data[16]),
    .Z(_4017_)
  );
  AND2_X1 _9255_ (
    .A1(_3814_),
    .A2(_4017_),
    .ZN(_4018_)
  );
  OR2_X1 _9256_ (
    .A1(_4014_),
    .A2(_4018_),
    .ZN(_4019_)
  );
  OR2_X1 _9257_ (
    .A1(remainder[15]),
    .A2(_3689_),
    .ZN(_4020_)
  );
  AND2_X1 _9258_ (
    .A1(_3911_),
    .A2(_4020_),
    .ZN(_4021_)
  );
  AND2_X1 _9259_ (
    .A1(_4019_),
    .A2(_4021_),
    .ZN(_4022_)
  );
  AND2_X1 _9260_ (
    .A1(remainder[16]),
    .A2(_3826_),
    .ZN(_4023_)
  );
  AND2_X1 _9261_ (
    .A1(io_req_bits_in1[16]),
    .A2(_3902_),
    .ZN(_4024_)
  );
  OR2_X1 _9262_ (
    .A1(_4023_),
    .A2(_4024_),
    .ZN(_4025_)
  );
  OR2_X1 _9263_ (
    .A1(_4022_),
    .A2(_4025_),
    .ZN(_0103_)
  );
  AND2_X1 _9264_ (
    .A1(remainder[25]),
    .A2(_3819_),
    .ZN(_4027_)
  );
  OR2_X1 _9265_ (
    .A1(_3678_),
    .A2(_4027_),
    .ZN(_4028_)
  );
  MUX2_X1 _9266_ (
    .A(remainder[17]),
    .B(remainder[50]),
    .S(resHi),
    .Z(io_resp_bits_data[17])
  );
  OR2_X1 _9267_ (
    .A1(_4016_),
    .A2(io_resp_bits_data[17]),
    .ZN(_4029_)
  );
  XOR2_X1 _9268_ (
    .A(_4016_),
    .B(io_resp_bits_data[17]),
    .Z(_4030_)
  );
  AND2_X1 _9269_ (
    .A1(_3814_),
    .A2(_4030_),
    .ZN(_4031_)
  );
  OR2_X1 _9270_ (
    .A1(_4028_),
    .A2(_4031_),
    .ZN(_4032_)
  );
  OR2_X1 _9271_ (
    .A1(remainder[16]),
    .A2(_3689_),
    .ZN(_4033_)
  );
  AND2_X1 _9272_ (
    .A1(_3911_),
    .A2(_4033_),
    .ZN(_4034_)
  );
  AND2_X1 _9273_ (
    .A1(_4032_),
    .A2(_4034_),
    .ZN(_4036_)
  );
  AND2_X1 _9274_ (
    .A1(remainder[17]),
    .A2(_3826_),
    .ZN(_4037_)
  );
  AND2_X1 _9275_ (
    .A1(io_req_bits_in1[17]),
    .A2(_3902_),
    .ZN(_4038_)
  );
  OR2_X1 _9276_ (
    .A1(_4037_),
    .A2(_4038_),
    .ZN(_4039_)
  );
  OR2_X1 _9277_ (
    .A1(_4036_),
    .A2(_4039_),
    .ZN(_0104_)
  );
  AND2_X1 _9278_ (
    .A1(remainder[26]),
    .A2(_3819_),
    .ZN(_4040_)
  );
  OR2_X1 _9279_ (
    .A1(_3678_),
    .A2(_4040_),
    .ZN(_4041_)
  );
  MUX2_X1 _9280_ (
    .A(remainder[18]),
    .B(remainder[51]),
    .S(resHi),
    .Z(io_resp_bits_data[18])
  );
  OR2_X1 _9281_ (
    .A1(_4029_),
    .A2(io_resp_bits_data[18]),
    .ZN(_4042_)
  );
  XOR2_X1 _9282_ (
    .A(_4029_),
    .B(io_resp_bits_data[18]),
    .Z(_4043_)
  );
  AND2_X1 _9283_ (
    .A1(_3814_),
    .A2(_4043_),
    .ZN(_4045_)
  );
  OR2_X1 _9284_ (
    .A1(_4041_),
    .A2(_4045_),
    .ZN(_4046_)
  );
  OR2_X1 _9285_ (
    .A1(remainder[17]),
    .A2(_3689_),
    .ZN(_4047_)
  );
  AND2_X1 _9286_ (
    .A1(_3911_),
    .A2(_4047_),
    .ZN(_4048_)
  );
  AND2_X1 _9287_ (
    .A1(_4046_),
    .A2(_4048_),
    .ZN(_4049_)
  );
  AND2_X1 _9288_ (
    .A1(remainder[18]),
    .A2(_3826_),
    .ZN(_4050_)
  );
  AND2_X1 _9289_ (
    .A1(io_req_bits_in1[18]),
    .A2(_3902_),
    .ZN(_4051_)
  );
  OR2_X1 _9290_ (
    .A1(_4050_),
    .A2(_4051_),
    .ZN(_4052_)
  );
  OR2_X1 _9291_ (
    .A1(_4049_),
    .A2(_4052_),
    .ZN(_0105_)
  );
  AND2_X1 _9292_ (
    .A1(remainder[27]),
    .A2(_3819_),
    .ZN(_4053_)
  );
  OR2_X1 _9293_ (
    .A1(_3678_),
    .A2(_4053_),
    .ZN(_4055_)
  );
  MUX2_X1 _9294_ (
    .A(remainder[19]),
    .B(remainder[52]),
    .S(resHi),
    .Z(io_resp_bits_data[19])
  );
  OR2_X1 _9295_ (
    .A1(_4042_),
    .A2(io_resp_bits_data[19]),
    .ZN(_4056_)
  );
  XOR2_X1 _9296_ (
    .A(_4042_),
    .B(io_resp_bits_data[19]),
    .Z(_4057_)
  );
  AND2_X1 _9297_ (
    .A1(_3814_),
    .A2(_4057_),
    .ZN(_4058_)
  );
  OR2_X1 _9298_ (
    .A1(_4055_),
    .A2(_4058_),
    .ZN(_4059_)
  );
  OR2_X1 _9299_ (
    .A1(remainder[18]),
    .A2(_3689_),
    .ZN(_4060_)
  );
  AND2_X1 _9300_ (
    .A1(_3911_),
    .A2(_4060_),
    .ZN(_4061_)
  );
  AND2_X1 _9301_ (
    .A1(_4059_),
    .A2(_4061_),
    .ZN(_4062_)
  );
  AND2_X1 _9302_ (
    .A1(remainder[19]),
    .A2(_3826_),
    .ZN(_4063_)
  );
  AND2_X1 _9303_ (
    .A1(io_req_bits_in1[19]),
    .A2(_3902_),
    .ZN(_4065_)
  );
  OR2_X1 _9304_ (
    .A1(_4063_),
    .A2(_4065_),
    .ZN(_4066_)
  );
  OR2_X1 _9305_ (
    .A1(_4062_),
    .A2(_4066_),
    .ZN(_0106_)
  );
  AND2_X1 _9306_ (
    .A1(remainder[28]),
    .A2(_3819_),
    .ZN(_4067_)
  );
  OR2_X1 _9307_ (
    .A1(_3678_),
    .A2(_4067_),
    .ZN(_4068_)
  );
  MUX2_X1 _9308_ (
    .A(remainder[20]),
    .B(remainder[53]),
    .S(resHi),
    .Z(io_resp_bits_data[20])
  );
  OR2_X1 _9309_ (
    .A1(_4056_),
    .A2(io_resp_bits_data[20]),
    .ZN(_4069_)
  );
  XOR2_X1 _9310_ (
    .A(_4056_),
    .B(io_resp_bits_data[20]),
    .Z(_4070_)
  );
  AND2_X1 _9311_ (
    .A1(_3814_),
    .A2(_4070_),
    .ZN(_4071_)
  );
  OR2_X1 _9312_ (
    .A1(_4068_),
    .A2(_4071_),
    .ZN(_4072_)
  );
  OR2_X1 _9313_ (
    .A1(remainder[19]),
    .A2(_3689_),
    .ZN(_4074_)
  );
  AND2_X1 _9314_ (
    .A1(_3911_),
    .A2(_4074_),
    .ZN(_4075_)
  );
  AND2_X1 _9315_ (
    .A1(_4072_),
    .A2(_4075_),
    .ZN(_4076_)
  );
  AND2_X1 _9316_ (
    .A1(remainder[20]),
    .A2(_3826_),
    .ZN(_4077_)
  );
  AND2_X1 _9317_ (
    .A1(io_req_bits_in1[20]),
    .A2(_3902_),
    .ZN(_4078_)
  );
  OR2_X1 _9318_ (
    .A1(_4077_),
    .A2(_4078_),
    .ZN(_4079_)
  );
  OR2_X1 _9319_ (
    .A1(_4076_),
    .A2(_4079_),
    .ZN(_0107_)
  );
  AND2_X1 _9320_ (
    .A1(remainder[29]),
    .A2(_3819_),
    .ZN(_4080_)
  );
  OR2_X1 _9321_ (
    .A1(_3678_),
    .A2(_4080_),
    .ZN(_4081_)
  );
  MUX2_X1 _9322_ (
    .A(remainder[21]),
    .B(remainder[54]),
    .S(resHi),
    .Z(io_resp_bits_data[21])
  );
  OR2_X1 _9323_ (
    .A1(_4069_),
    .A2(io_resp_bits_data[21]),
    .ZN(_4082_)
  );
  XOR2_X1 _9324_ (
    .A(_4069_),
    .B(io_resp_bits_data[21]),
    .Z(_4083_)
  );
  AND2_X1 _9325_ (
    .A1(_3814_),
    .A2(_4083_),
    .ZN(_4084_)
  );
  OR2_X1 _9326_ (
    .A1(_4081_),
    .A2(_4084_),
    .ZN(_4085_)
  );
  OR2_X1 _9327_ (
    .A1(remainder[20]),
    .A2(_3689_),
    .ZN(_4086_)
  );
  AND2_X1 _9328_ (
    .A1(_3911_),
    .A2(_4086_),
    .ZN(_4087_)
  );
  AND2_X1 _9329_ (
    .A1(_4085_),
    .A2(_4087_),
    .ZN(_4088_)
  );
  AND2_X1 _9330_ (
    .A1(remainder[21]),
    .A2(_3826_),
    .ZN(_4089_)
  );
  AND2_X1 _9331_ (
    .A1(io_req_bits_in1[21]),
    .A2(_3902_),
    .ZN(_4090_)
  );
  OR2_X1 _9332_ (
    .A1(_4089_),
    .A2(_4090_),
    .ZN(_4091_)
  );
  OR2_X1 _9333_ (
    .A1(_4088_),
    .A2(_4091_),
    .ZN(_0108_)
  );
  AND2_X1 _9334_ (
    .A1(remainder[30]),
    .A2(_3819_),
    .ZN(_4093_)
  );
  OR2_X1 _9335_ (
    .A1(_3678_),
    .A2(_4093_),
    .ZN(_4094_)
  );
  MUX2_X1 _9336_ (
    .A(remainder[22]),
    .B(remainder[55]),
    .S(resHi),
    .Z(io_resp_bits_data[22])
  );
  OR2_X1 _9337_ (
    .A1(_4082_),
    .A2(io_resp_bits_data[22]),
    .ZN(_4095_)
  );
  INV_X1 _9338_ (
    .A(_4095_),
    .ZN(_4096_)
  );
  XOR2_X1 _9339_ (
    .A(_4082_),
    .B(io_resp_bits_data[22]),
    .Z(_4097_)
  );
  AND2_X1 _9340_ (
    .A1(_3814_),
    .A2(_4097_),
    .ZN(_4098_)
  );
  OR2_X1 _9341_ (
    .A1(_4094_),
    .A2(_4098_),
    .ZN(_4099_)
  );
  OR2_X1 _9342_ (
    .A1(remainder[21]),
    .A2(_3689_),
    .ZN(_4100_)
  );
  AND2_X1 _9343_ (
    .A1(_3911_),
    .A2(_4100_),
    .ZN(_4102_)
  );
  AND2_X1 _9344_ (
    .A1(_4099_),
    .A2(_4102_),
    .ZN(_4103_)
  );
  AND2_X1 _9345_ (
    .A1(remainder[22]),
    .A2(_3826_),
    .ZN(_4104_)
  );
  AND2_X1 _9346_ (
    .A1(io_req_bits_in1[22]),
    .A2(_3902_),
    .ZN(_4105_)
  );
  OR2_X1 _9347_ (
    .A1(_4104_),
    .A2(_4105_),
    .ZN(_4106_)
  );
  OR2_X1 _9348_ (
    .A1(_4103_),
    .A2(_4106_),
    .ZN(_0109_)
  );
  AND2_X1 _9349_ (
    .A1(remainder[31]),
    .A2(_3819_),
    .ZN(_4107_)
  );
  OR2_X1 _9350_ (
    .A1(_3678_),
    .A2(_4107_),
    .ZN(_4108_)
  );
  MUX2_X1 _9351_ (
    .A(remainder[23]),
    .B(remainder[56]),
    .S(resHi),
    .Z(io_resp_bits_data[23])
  );
  INV_X1 _9352_ (
    .A(io_resp_bits_data[23]),
    .ZN(_4109_)
  );
  AND2_X1 _9353_ (
    .A1(_4096_),
    .A2(_4109_),
    .ZN(_4111_)
  );
  INV_X1 _9354_ (
    .A(_4111_),
    .ZN(_4112_)
  );
  XOR2_X1 _9355_ (
    .A(_4095_),
    .B(io_resp_bits_data[23]),
    .Z(_4113_)
  );
  AND2_X1 _9356_ (
    .A1(_3814_),
    .A2(_4113_),
    .ZN(_4114_)
  );
  OR2_X1 _9357_ (
    .A1(_4108_),
    .A2(_4114_),
    .ZN(_4115_)
  );
  OR2_X1 _9358_ (
    .A1(remainder[22]),
    .A2(_3689_),
    .ZN(_4116_)
  );
  AND2_X1 _9359_ (
    .A1(_3911_),
    .A2(_4116_),
    .ZN(_4117_)
  );
  AND2_X1 _9360_ (
    .A1(_4115_),
    .A2(_4117_),
    .ZN(_4118_)
  );
  AND2_X1 _9361_ (
    .A1(remainder[23]),
    .A2(_3826_),
    .ZN(_4119_)
  );
  AND2_X1 _9362_ (
    .A1(io_req_bits_in1[23]),
    .A2(_3902_),
    .ZN(_4120_)
  );
  OR2_X1 _9363_ (
    .A1(_4119_),
    .A2(_4120_),
    .ZN(_4122_)
  );
  OR2_X1 _9364_ (
    .A1(_4118_),
    .A2(_4122_),
    .ZN(_0110_)
  );
  MUX2_X1 _9365_ (
    .A(_3493_),
    .B(_3013_),
    .S(resHi),
    .Z(_4123_)
  );
  INV_X1 _9366_ (
    .A(_4123_),
    .ZN(io_resp_bits_data[24])
  );
  OR2_X1 _9367_ (
    .A1(_4111_),
    .A2(_4123_),
    .ZN(_4124_)
  );
  OR2_X1 _9368_ (
    .A1(_4112_),
    .A2(io_resp_bits_data[24]),
    .ZN(_4125_)
  );
  AND2_X1 _9369_ (
    .A1(_3814_),
    .A2(_4124_),
    .ZN(_4126_)
  );
  AND2_X1 _9370_ (
    .A1(_4125_),
    .A2(_4126_),
    .ZN(_4127_)
  );
  OR2_X1 _9371_ (
    .A1(remainder[33]),
    .A2(_0186_),
    .ZN(_4128_)
  );
  AND2_X1 _9372_ (
    .A1(_3819_),
    .A2(_4128_),
    .ZN(_4129_)
  );
  AND2_X1 _9373_ (
    .A1(_0232_),
    .A2(_4129_),
    .ZN(_4131_)
  );
  OR2_X1 _9374_ (
    .A1(_3678_),
    .A2(_4131_),
    .ZN(_4132_)
  );
  OR2_X1 _9375_ (
    .A1(_4127_),
    .A2(_4132_),
    .ZN(_4133_)
  );
  OR2_X1 _9376_ (
    .A1(remainder[23]),
    .A2(_3689_),
    .ZN(_4134_)
  );
  AND2_X1 _9377_ (
    .A1(_3911_),
    .A2(_4134_),
    .ZN(_4135_)
  );
  AND2_X1 _9378_ (
    .A1(_4133_),
    .A2(_4135_),
    .ZN(_4136_)
  );
  AND2_X1 _9379_ (
    .A1(remainder[24]),
    .A2(_3826_),
    .ZN(_4137_)
  );
  AND2_X1 _9380_ (
    .A1(io_req_bits_in1[24]),
    .A2(_3902_),
    .ZN(_4138_)
  );
  OR2_X1 _9381_ (
    .A1(_4137_),
    .A2(_4138_),
    .ZN(_4139_)
  );
  OR2_X1 _9382_ (
    .A1(_4136_),
    .A2(_4139_),
    .ZN(_0111_)
  );
  MUX2_X1 _9383_ (
    .A(remainder[25]),
    .B(remainder[58]),
    .S(resHi),
    .Z(io_resp_bits_data[25])
  );
  AND2_X1 _9384_ (
    .A1(_4125_),
    .A2(io_resp_bits_data[25]),
    .ZN(_4141_)
  );
  INV_X1 _9385_ (
    .A(_4141_),
    .ZN(_4142_)
  );
  OR2_X1 _9386_ (
    .A1(_4125_),
    .A2(io_resp_bits_data[25]),
    .ZN(_4143_)
  );
  AND2_X1 _9387_ (
    .A1(_3814_),
    .A2(_4143_),
    .ZN(_4144_)
  );
  AND2_X1 _9388_ (
    .A1(_4142_),
    .A2(_4144_),
    .ZN(_4145_)
  );
  OR2_X1 _9389_ (
    .A1(_0231_),
    .A2(_0233_),
    .ZN(_4146_)
  );
  AND2_X1 _9390_ (
    .A1(_3819_),
    .A2(_4146_),
    .ZN(_4147_)
  );
  AND2_X1 _9391_ (
    .A1(_0235_),
    .A2(_4147_),
    .ZN(_4148_)
  );
  OR2_X1 _9392_ (
    .A1(_3678_),
    .A2(_4148_),
    .ZN(_4149_)
  );
  OR2_X1 _9393_ (
    .A1(_4145_),
    .A2(_4149_),
    .ZN(_4151_)
  );
  OR2_X1 _9394_ (
    .A1(remainder[24]),
    .A2(_3689_),
    .ZN(_4152_)
  );
  AND2_X1 _9395_ (
    .A1(_3911_),
    .A2(_4152_),
    .ZN(_4153_)
  );
  AND2_X1 _9396_ (
    .A1(_4151_),
    .A2(_4153_),
    .ZN(_4154_)
  );
  AND2_X1 _9397_ (
    .A1(remainder[25]),
    .A2(_3826_),
    .ZN(_4155_)
  );
  AND2_X1 _9398_ (
    .A1(io_req_bits_in1[25]),
    .A2(_3902_),
    .ZN(_4156_)
  );
  OR2_X1 _9399_ (
    .A1(_4155_),
    .A2(_4156_),
    .ZN(_4157_)
  );
  OR2_X1 _9400_ (
    .A1(_4154_),
    .A2(_4157_),
    .ZN(_0112_)
  );
  MUX2_X1 _9401_ (
    .A(remainder[26]),
    .B(remainder[59]),
    .S(resHi),
    .Z(io_resp_bits_data[26])
  );
  OR2_X1 _9402_ (
    .A1(_4143_),
    .A2(io_resp_bits_data[26]),
    .ZN(_4158_)
  );
  XOR2_X1 _9403_ (
    .A(_4143_),
    .B(io_resp_bits_data[26]),
    .Z(_4159_)
  );
  AND2_X1 _9404_ (
    .A1(_3814_),
    .A2(_4159_),
    .ZN(_4160_)
  );
  OR2_X1 _9405_ (
    .A1(_0236_),
    .A2(_0238_),
    .ZN(_4161_)
  );
  AND2_X1 _9406_ (
    .A1(_3819_),
    .A2(_4161_),
    .ZN(_4162_)
  );
  AND2_X1 _9407_ (
    .A1(_0241_),
    .A2(_4162_),
    .ZN(_4163_)
  );
  OR2_X1 _9408_ (
    .A1(_3678_),
    .A2(_4163_),
    .ZN(_4164_)
  );
  OR2_X1 _9409_ (
    .A1(_4160_),
    .A2(_4164_),
    .ZN(_4165_)
  );
  OR2_X1 _9410_ (
    .A1(remainder[25]),
    .A2(_3689_),
    .ZN(_4166_)
  );
  AND2_X1 _9411_ (
    .A1(_3911_),
    .A2(_4166_),
    .ZN(_4167_)
  );
  AND2_X1 _9412_ (
    .A1(_4165_),
    .A2(_4167_),
    .ZN(_4168_)
  );
  AND2_X1 _9413_ (
    .A1(remainder[26]),
    .A2(_3826_),
    .ZN(_4170_)
  );
  AND2_X1 _9414_ (
    .A1(io_req_bits_in1[26]),
    .A2(_3902_),
    .ZN(_4171_)
  );
  OR2_X1 _9415_ (
    .A1(_4170_),
    .A2(_4171_),
    .ZN(_4172_)
  );
  OR2_X1 _9416_ (
    .A1(_4168_),
    .A2(_4172_),
    .ZN(_0113_)
  );
  MUX2_X1 _9417_ (
    .A(remainder[27]),
    .B(remainder[60]),
    .S(resHi),
    .Z(io_resp_bits_data[27])
  );
  AND2_X1 _9418_ (
    .A1(_4158_),
    .A2(io_resp_bits_data[27]),
    .ZN(_4173_)
  );
  INV_X1 _9419_ (
    .A(_4173_),
    .ZN(_4174_)
  );
  OR2_X1 _9420_ (
    .A1(_4158_),
    .A2(io_resp_bits_data[27]),
    .ZN(_4175_)
  );
  AND2_X1 _9421_ (
    .A1(_3814_),
    .A2(_4175_),
    .ZN(_4176_)
  );
  AND2_X1 _9422_ (
    .A1(_4174_),
    .A2(_4176_),
    .ZN(_4177_)
  );
  AND2_X1 _9423_ (
    .A1(_0223_),
    .A2(_0225_),
    .ZN(_4179_)
  );
  OR2_X1 _9424_ (
    .A1(_0222_),
    .A2(_0224_),
    .ZN(_4180_)
  );
  OR2_X1 _9425_ (
    .A1(_0242_),
    .A2(_4180_),
    .ZN(_4181_)
  );
  OR2_X1 _9426_ (
    .A1(_0243_),
    .A2(_4179_),
    .ZN(_4182_)
  );
  AND2_X1 _9427_ (
    .A1(_3819_),
    .A2(_4181_),
    .ZN(_4183_)
  );
  AND2_X1 _9428_ (
    .A1(_4182_),
    .A2(_4183_),
    .ZN(_4184_)
  );
  OR2_X1 _9429_ (
    .A1(_3678_),
    .A2(_4184_),
    .ZN(_4185_)
  );
  OR2_X1 _9430_ (
    .A1(_4177_),
    .A2(_4185_),
    .ZN(_4186_)
  );
  OR2_X1 _9431_ (
    .A1(remainder[26]),
    .A2(_3689_),
    .ZN(_4187_)
  );
  AND2_X1 _9432_ (
    .A1(_3911_),
    .A2(_4187_),
    .ZN(_4188_)
  );
  AND2_X1 _9433_ (
    .A1(_4186_),
    .A2(_4188_),
    .ZN(_4190_)
  );
  AND2_X1 _9434_ (
    .A1(remainder[27]),
    .A2(_3826_),
    .ZN(_4191_)
  );
  AND2_X1 _9435_ (
    .A1(io_req_bits_in1[27]),
    .A2(_3902_),
    .ZN(_4192_)
  );
  OR2_X1 _9436_ (
    .A1(_4191_),
    .A2(_4192_),
    .ZN(_4193_)
  );
  OR2_X1 _9437_ (
    .A1(_4190_),
    .A2(_4193_),
    .ZN(_0114_)
  );
  MUX2_X1 _9438_ (
    .A(remainder[28]),
    .B(remainder[61]),
    .S(resHi),
    .Z(io_resp_bits_data[28])
  );
  AND2_X1 _9439_ (
    .A1(_4175_),
    .A2(io_resp_bits_data[28]),
    .ZN(_4194_)
  );
  INV_X1 _9440_ (
    .A(_4194_),
    .ZN(_4195_)
  );
  OR2_X1 _9441_ (
    .A1(_4175_),
    .A2(io_resp_bits_data[28]),
    .ZN(_4196_)
  );
  AND2_X1 _9442_ (
    .A1(_3814_),
    .A2(_4196_),
    .ZN(_4197_)
  );
  AND2_X1 _9443_ (
    .A1(_4195_),
    .A2(_4197_),
    .ZN(_4199_)
  );
  OR2_X1 _9444_ (
    .A1(_0218_),
    .A2(_0247_),
    .ZN(_4200_)
  );
  AND2_X1 _9445_ (
    .A1(_3819_),
    .A2(_4200_),
    .ZN(_4201_)
  );
  AND2_X1 _9446_ (
    .A1(_0249_),
    .A2(_4201_),
    .ZN(_4202_)
  );
  OR2_X1 _9447_ (
    .A1(_3678_),
    .A2(_4202_),
    .ZN(_4203_)
  );
  OR2_X1 _9448_ (
    .A1(_4199_),
    .A2(_4203_),
    .ZN(_4204_)
  );
  OR2_X1 _9449_ (
    .A1(remainder[27]),
    .A2(_3689_),
    .ZN(_4205_)
  );
  AND2_X1 _9450_ (
    .A1(_3911_),
    .A2(_4205_),
    .ZN(_4206_)
  );
  AND2_X1 _9451_ (
    .A1(_4204_),
    .A2(_4206_),
    .ZN(_4207_)
  );
  AND2_X1 _9452_ (
    .A1(remainder[28]),
    .A2(_3826_),
    .ZN(_4208_)
  );
  AND2_X1 _9453_ (
    .A1(io_req_bits_in1[28]),
    .A2(_3902_),
    .ZN(_4210_)
  );
  OR2_X1 _9454_ (
    .A1(_4208_),
    .A2(_4210_),
    .ZN(_4211_)
  );
  OR2_X1 _9455_ (
    .A1(_4207_),
    .A2(_4211_),
    .ZN(_0115_)
  );
  MUX2_X1 _9456_ (
    .A(remainder[29]),
    .B(remainder[62]),
    .S(resHi),
    .Z(io_resp_bits_data[29])
  );
  OR2_X1 _9457_ (
    .A1(_4196_),
    .A2(io_resp_bits_data[29]),
    .ZN(_4212_)
  );
  XOR2_X1 _9458_ (
    .A(_4196_),
    .B(io_resp_bits_data[29]),
    .Z(_4213_)
  );
  AND2_X1 _9459_ (
    .A1(_3814_),
    .A2(_4213_),
    .ZN(_4214_)
  );
  OR2_X1 _9460_ (
    .A1(_0213_),
    .A2(_0251_),
    .ZN(_4215_)
  );
  AND2_X1 _9461_ (
    .A1(_3819_),
    .A2(_0253_),
    .ZN(_4216_)
  );
  AND2_X1 _9462_ (
    .A1(_4215_),
    .A2(_4216_),
    .ZN(_4217_)
  );
  OR2_X1 _9463_ (
    .A1(_3678_),
    .A2(_4217_),
    .ZN(_4219_)
  );
  OR2_X1 _9464_ (
    .A1(_4214_),
    .A2(_4219_),
    .ZN(_4220_)
  );
  OR2_X1 _9465_ (
    .A1(remainder[28]),
    .A2(_3689_),
    .ZN(_4221_)
  );
  AND2_X1 _9466_ (
    .A1(_3911_),
    .A2(_4221_),
    .ZN(_4222_)
  );
  AND2_X1 _9467_ (
    .A1(_4220_),
    .A2(_4222_),
    .ZN(_4223_)
  );
  AND2_X1 _9468_ (
    .A1(remainder[29]),
    .A2(_3826_),
    .ZN(_4224_)
  );
  AND2_X1 _9469_ (
    .A1(io_req_bits_in1[29]),
    .A2(_3902_),
    .ZN(_4225_)
  );
  OR2_X1 _9470_ (
    .A1(_4224_),
    .A2(_4225_),
    .ZN(_4226_)
  );
  OR2_X1 _9471_ (
    .A1(_4223_),
    .A2(_4226_),
    .ZN(_0116_)
  );
  MUX2_X1 _9472_ (
    .A(remainder[30]),
    .B(remainder[63]),
    .S(resHi),
    .Z(io_resp_bits_data[30])
  );
  OR2_X1 _9473_ (
    .A1(_4212_),
    .A2(io_resp_bits_data[30]),
    .ZN(_4228_)
  );
  XOR2_X1 _9474_ (
    .A(_4212_),
    .B(io_resp_bits_data[30]),
    .Z(_4229_)
  );
  AND2_X1 _9475_ (
    .A1(_3814_),
    .A2(_4229_),
    .ZN(_4230_)
  );
  OR2_X1 _9476_ (
    .A1(_0255_),
    .A2(_0256_),
    .ZN(_4231_)
  );
  AND2_X1 _9477_ (
    .A1(_3819_),
    .A2(_0259_),
    .ZN(_4232_)
  );
  AND2_X1 _9478_ (
    .A1(_4231_),
    .A2(_4232_),
    .ZN(_4233_)
  );
  OR2_X1 _9479_ (
    .A1(_3678_),
    .A2(_4233_),
    .ZN(_4234_)
  );
  OR2_X1 _9480_ (
    .A1(_4230_),
    .A2(_4234_),
    .ZN(_4235_)
  );
  OR2_X1 _9481_ (
    .A1(remainder[29]),
    .A2(_3689_),
    .ZN(_4236_)
  );
  AND2_X1 _9482_ (
    .A1(_3911_),
    .A2(_4236_),
    .ZN(_4237_)
  );
  AND2_X1 _9483_ (
    .A1(_4235_),
    .A2(_4237_),
    .ZN(_4239_)
  );
  AND2_X1 _9484_ (
    .A1(remainder[30]),
    .A2(_3826_),
    .ZN(_4240_)
  );
  AND2_X1 _9485_ (
    .A1(io_req_bits_in1[30]),
    .A2(_3902_),
    .ZN(_4241_)
  );
  OR2_X1 _9486_ (
    .A1(_4240_),
    .A2(_4241_),
    .ZN(_4242_)
  );
  OR2_X1 _9487_ (
    .A1(_4239_),
    .A2(_4242_),
    .ZN(_0117_)
  );
  MUX2_X1 _9488_ (
    .A(remainder[31]),
    .B(remainder[64]),
    .S(resHi),
    .Z(io_resp_bits_data[31])
  );
  XOR2_X1 _9489_ (
    .A(_4228_),
    .B(io_resp_bits_data[31]),
    .Z(_4243_)
  );
  AND2_X1 _9490_ (
    .A1(_3814_),
    .A2(_4243_),
    .ZN(_4244_)
  );
  OR2_X1 _9491_ (
    .A1(_0261_),
    .A2(_0262_),
    .ZN(_4245_)
  );
  AND2_X1 _9492_ (
    .A1(_3819_),
    .A2(_4245_),
    .ZN(_4246_)
  );
  AND2_X1 _9493_ (
    .A1(_0265_),
    .A2(_4246_),
    .ZN(_4248_)
  );
  OR2_X1 _9494_ (
    .A1(_3678_),
    .A2(_4248_),
    .ZN(_4249_)
  );
  OR2_X1 _9495_ (
    .A1(_4244_),
    .A2(_4249_),
    .ZN(_4250_)
  );
  OR2_X1 _9496_ (
    .A1(remainder[30]),
    .A2(_3689_),
    .ZN(_4251_)
  );
  AND2_X1 _9497_ (
    .A1(_3911_),
    .A2(_4251_),
    .ZN(_4252_)
  );
  AND2_X1 _9498_ (
    .A1(_4250_),
    .A2(_4252_),
    .ZN(_4253_)
  );
  AND2_X1 _9499_ (
    .A1(remainder[31]),
    .A2(_3826_),
    .ZN(_4254_)
  );
  AND2_X1 _9500_ (
    .A1(io_req_bits_in1[31]),
    .A2(_3902_),
    .ZN(_4255_)
  );
  OR2_X1 _9501_ (
    .A1(_4254_),
    .A2(_4255_),
    .ZN(_4256_)
  );
  OR2_X1 _9502_ (
    .A1(_4253_),
    .A2(_4256_),
    .ZN(_0118_)
  );
  OR2_X1 _9503_ (
    .A1(state[2]),
    .A2(_3978_),
    .ZN(_4258_)
  );
  AND2_X1 _9504_ (
    .A1(_3253_),
    .A2(_4110_),
    .ZN(_4259_)
  );
  AND2_X1 _9505_ (
    .A1(_4258_),
    .A2(_4259_),
    .ZN(_0119_)
  );
  MUX2_X1 _9506_ (
    .A(_4401_),
    .B(isHi),
    .S(_3911_),
    .Z(_0120_)
  );
  DFF_X1 \count[0]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0014_),
    .Q(count[0]),
    .QN(_count_T_1[0])
  );
  DFF_X1 \count[1]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0015_),
    .Q(count[1]),
    .QN(_0002_)
  );
  DFF_X1 \count[2]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0016_),
    .Q(count[2]),
    .QN(_4769_)
  );
  DFF_X1 \count[3]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0017_),
    .Q(count[3]),
    .QN(_4768_)
  );
  DFF_X1 \count[4]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0018_),
    .Q(count[4]),
    .QN(_4767_)
  );
  DFF_X1 \count[5]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0019_),
    .Q(count[5]),
    .QN(_0001_)
  );
  DFF_X1 \divisor[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_0020_),
    .Q(divisor[0]),
    .QN(_4776_[0])
  );
  DFF_X1 \divisor[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_0030_),
    .Q(divisor[10]),
    .QN(_4776_[10])
  );
  DFF_X1 \divisor[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_0031_),
    .Q(divisor[11]),
    .QN(_4776_[11])
  );
  DFF_X1 \divisor[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_0032_),
    .Q(divisor[12]),
    .QN(_4776_[12])
  );
  DFF_X1 \divisor[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_0033_),
    .Q(divisor[13]),
    .QN(_4776_[13])
  );
  DFF_X1 \divisor[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_0034_),
    .Q(divisor[14]),
    .QN(_4776_[14])
  );
  DFF_X1 \divisor[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_0035_),
    .Q(divisor[15]),
    .QN(_4776_[15])
  );
  DFF_X1 \divisor[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_0036_),
    .Q(divisor[16]),
    .QN(_4776_[16])
  );
  DFF_X1 \divisor[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_0037_),
    .Q(divisor[17]),
    .QN(_4776_[17])
  );
  DFF_X1 \divisor[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_0038_),
    .Q(divisor[18]),
    .QN(_4776_[18])
  );
  DFF_X1 \divisor[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_0039_),
    .Q(divisor[19]),
    .QN(_4776_[19])
  );
  DFF_X1 \divisor[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_0021_),
    .Q(divisor[1]),
    .QN(_4776_[1])
  );
  DFF_X1 \divisor[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_0040_),
    .Q(divisor[20]),
    .QN(_4776_[20])
  );
  DFF_X1 \divisor[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_0041_),
    .Q(divisor[21]),
    .QN(_4776_[21])
  );
  DFF_X1 \divisor[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_0042_),
    .Q(divisor[22]),
    .QN(_4776_[22])
  );
  DFF_X1 \divisor[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_0043_),
    .Q(divisor[23]),
    .QN(_4776_[23])
  );
  DFF_X1 \divisor[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_0044_),
    .Q(divisor[24]),
    .QN(_4776_[24])
  );
  DFF_X1 \divisor[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_0045_),
    .Q(divisor[25]),
    .QN(_4776_[25])
  );
  DFF_X1 \divisor[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_0046_),
    .Q(divisor[26]),
    .QN(_4776_[26])
  );
  DFF_X1 \divisor[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_0047_),
    .Q(divisor[27]),
    .QN(_4776_[27])
  );
  DFF_X1 \divisor[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_0048_),
    .Q(divisor[28]),
    .QN(_4776_[28])
  );
  DFF_X1 \divisor[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_0049_),
    .Q(divisor[29]),
    .QN(_4776_[29])
  );
  DFF_X1 \divisor[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_0022_),
    .Q(divisor[2]),
    .QN(_4776_[2])
  );
  DFF_X1 \divisor[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_0050_),
    .Q(divisor[30]),
    .QN(_4776_[30])
  );
  DFF_X1 \divisor[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_0051_),
    .Q(divisor[31]),
    .QN(_4776_[31])
  );
  DFF_X1 \divisor[32]$_DFFE_PP_  (
    .CK(clock),
    .D(_0052_),
    .Q(divisor[32]),
    .QN(_4776_[32])
  );
  DFF_X1 \divisor[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_0023_),
    .Q(divisor[3]),
    .QN(_4776_[3])
  );
  DFF_X1 \divisor[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_0024_),
    .Q(divisor[4]),
    .QN(_4776_[4])
  );
  DFF_X1 \divisor[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_0025_),
    .Q(divisor[5]),
    .QN(_4776_[5])
  );
  DFF_X1 \divisor[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_0026_),
    .Q(divisor[6]),
    .QN(_4776_[6])
  );
  DFF_X1 \divisor[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_0027_),
    .Q(divisor[7]),
    .QN(_4776_[7])
  );
  DFF_X1 \divisor[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_0028_),
    .Q(divisor[8]),
    .QN(_4776_[8])
  );
  DFF_X1 \divisor[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_0029_),
    .Q(divisor[9]),
    .QN(_4776_[9])
  );
  DFF_X1 \isHi$_DFFE_PP_  (
    .CK(clock),
    .D(_0120_),
    .Q(isHi),
    .QN(_eOut_T_4)
  );
  DFF_X1 \neg_out$_DFFE_PP_  (
    .CK(clock),
    .D(_0008_),
    .Q(neg_out),
    .QN(_state_T[1])
  );
  DFF_X1 \remainder[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_0087_),
    .Q(remainder[0]),
    .QN(_4732_)
  );
  DFF_X1 \remainder[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_0097_),
    .Q(remainder[10]),
    .QN(_4722_)
  );
  DFF_X1 \remainder[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_0098_),
    .Q(remainder[11]),
    .QN(_4721_)
  );
  DFF_X1 \remainder[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_0099_),
    .Q(remainder[12]),
    .QN(_4720_)
  );
  DFF_X1 \remainder[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_0100_),
    .Q(remainder[13]),
    .QN(_4719_)
  );
  DFF_X1 \remainder[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_0101_),
    .Q(remainder[14]),
    .QN(_4718_)
  );
  DFF_X1 \remainder[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_0102_),
    .Q(remainder[15]),
    .QN(_4717_)
  );
  DFF_X1 \remainder[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_0103_),
    .Q(remainder[16]),
    .QN(_4716_)
  );
  DFF_X1 \remainder[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_0104_),
    .Q(remainder[17]),
    .QN(_4715_)
  );
  DFF_X1 \remainder[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_0105_),
    .Q(remainder[18]),
    .QN(_4714_)
  );
  DFF_X1 \remainder[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_0106_),
    .Q(remainder[19]),
    .QN(_4713_)
  );
  DFF_X1 \remainder[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_0088_),
    .Q(remainder[1]),
    .QN(_4731_)
  );
  DFF_X1 \remainder[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_0107_),
    .Q(remainder[20]),
    .QN(_4712_)
  );
  DFF_X1 \remainder[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_0108_),
    .Q(remainder[21]),
    .QN(_4711_)
  );
  DFF_X1 \remainder[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_0109_),
    .Q(remainder[22]),
    .QN(_4710_)
  );
  DFF_X1 \remainder[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_0110_),
    .Q(remainder[23]),
    .QN(_4709_)
  );
  DFF_X1 \remainder[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_0111_),
    .Q(remainder[24]),
    .QN(_4708_)
  );
  DFF_X1 \remainder[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_0112_),
    .Q(remainder[25]),
    .QN(_4707_)
  );
  DFF_X1 \remainder[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_0113_),
    .Q(remainder[26]),
    .QN(_4706_)
  );
  DFF_X1 \remainder[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_0114_),
    .Q(remainder[27]),
    .QN(_4705_)
  );
  DFF_X1 \remainder[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_0115_),
    .Q(remainder[28]),
    .QN(_4704_)
  );
  DFF_X1 \remainder[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_0116_),
    .Q(remainder[29]),
    .QN(_4703_)
  );
  DFF_X1 \remainder[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_0089_),
    .Q(remainder[2]),
    .QN(_4730_)
  );
  DFF_X1 \remainder[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_0117_),
    .Q(remainder[30]),
    .QN(_4702_)
  );
  DFF_X1 \remainder[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_0118_),
    .Q(remainder[31]),
    .QN(_4701_)
  );
  DFF_X1 \remainder[32]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0053_),
    .Q(remainder[32]),
    .QN(_4766_)
  );
  DFF_X1 \remainder[33]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0054_),
    .Q(remainder[33]),
    .QN(_4765_)
  );
  DFF_X1 \remainder[34]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0055_),
    .Q(remainder[34]),
    .QN(_4764_)
  );
  DFF_X1 \remainder[35]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0056_),
    .Q(remainder[35]),
    .QN(_4763_)
  );
  DFF_X1 \remainder[36]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0057_),
    .Q(remainder[36]),
    .QN(_4762_)
  );
  DFF_X1 \remainder[37]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0058_),
    .Q(remainder[37]),
    .QN(_4761_)
  );
  DFF_X1 \remainder[38]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0059_),
    .Q(remainder[38]),
    .QN(_4760_)
  );
  DFF_X1 \remainder[39]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0060_),
    .Q(remainder[39]),
    .QN(_4759_)
  );
  DFF_X1 \remainder[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_0090_),
    .Q(remainder[3]),
    .QN(_4729_)
  );
  DFF_X1 \remainder[40]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0061_),
    .Q(remainder[40]),
    .QN(_4758_)
  );
  DFF_X1 \remainder[41]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0062_),
    .Q(remainder[41]),
    .QN(_4757_)
  );
  DFF_X1 \remainder[42]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0063_),
    .Q(remainder[42]),
    .QN(_4756_)
  );
  DFF_X1 \remainder[43]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0064_),
    .Q(remainder[43]),
    .QN(_4755_)
  );
  DFF_X1 \remainder[44]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0065_),
    .Q(remainder[44]),
    .QN(_4754_)
  );
  DFF_X1 \remainder[45]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0066_),
    .Q(remainder[45]),
    .QN(_4753_)
  );
  DFF_X1 \remainder[46]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0067_),
    .Q(remainder[46]),
    .QN(_4752_)
  );
  DFF_X1 \remainder[47]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0068_),
    .Q(remainder[47]),
    .QN(_4751_)
  );
  DFF_X1 \remainder[48]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0069_),
    .Q(remainder[48]),
    .QN(_4750_)
  );
  DFF_X1 \remainder[49]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0070_),
    .Q(remainder[49]),
    .QN(_4749_)
  );
  DFF_X1 \remainder[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_0091_),
    .Q(remainder[4]),
    .QN(_4728_)
  );
  DFF_X1 \remainder[50]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0071_),
    .Q(remainder[50]),
    .QN(_4748_)
  );
  DFF_X1 \remainder[51]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0072_),
    .Q(remainder[51]),
    .QN(_4747_)
  );
  DFF_X1 \remainder[52]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0073_),
    .Q(remainder[52]),
    .QN(_4746_)
  );
  DFF_X1 \remainder[53]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0074_),
    .Q(remainder[53]),
    .QN(_4745_)
  );
  DFF_X1 \remainder[54]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0075_),
    .Q(remainder[54]),
    .QN(_4744_)
  );
  DFF_X1 \remainder[55]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0076_),
    .Q(remainder[55]),
    .QN(_4743_)
  );
  DFF_X1 \remainder[56]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0077_),
    .Q(remainder[56]),
    .QN(_4742_)
  );
  DFF_X1 \remainder[57]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0078_),
    .Q(remainder[57]),
    .QN(_4741_)
  );
  DFF_X1 \remainder[58]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0079_),
    .Q(remainder[58]),
    .QN(_4740_)
  );
  DFF_X1 \remainder[59]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0080_),
    .Q(remainder[59]),
    .QN(_4739_)
  );
  DFF_X1 \remainder[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_0092_),
    .Q(remainder[5]),
    .QN(_4727_)
  );
  DFF_X1 \remainder[60]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0081_),
    .Q(remainder[60]),
    .QN(_4738_)
  );
  DFF_X1 \remainder[61]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0082_),
    .Q(remainder[61]),
    .QN(_4737_)
  );
  DFF_X1 \remainder[62]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0083_),
    .Q(remainder[62]),
    .QN(_4736_)
  );
  DFF_X1 \remainder[63]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0084_),
    .Q(remainder[63]),
    .QN(_4735_)
  );
  DFF_X1 \remainder[64]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0085_),
    .Q(remainder[64]),
    .QN(_4734_)
  );
  DFF_X1 \remainder[65]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_0086_),
    .Q(remainder[65]),
    .QN(_4733_)
  );
  DFF_X1 \remainder[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_0093_),
    .Q(remainder[6]),
    .QN(_4726_)
  );
  DFF_X1 \remainder[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_0094_),
    .Q(remainder[7]),
    .QN(_4725_)
  );
  DFF_X1 \remainder[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_0095_),
    .Q(remainder[8]),
    .QN(_4724_)
  );
  DFF_X1 \remainder[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_0096_),
    .Q(remainder[9]),
    .QN(_4723_)
  );
  DFF_X1 \req_tag[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_0009_),
    .Q(req_tag[0]),
    .QN(_4774_)
  );
  DFF_X1 \req_tag[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_0010_),
    .Q(req_tag[1]),
    .QN(_4773_)
  );
  DFF_X1 \req_tag[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_0011_),
    .Q(req_tag[2]),
    .QN(_4772_)
  );
  DFF_X1 \req_tag[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_0012_),
    .Q(req_tag[3]),
    .QN(_4771_)
  );
  DFF_X1 \req_tag[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_0013_),
    .Q(req_tag[4]),
    .QN(_4770_)
  );
  DFF_X1 \resHi$_SDFF_PP0_  (
    .CK(clock),
    .D(_0005_),
    .Q(resHi),
    .QN(_4775_)
  );
  DFF_X1 \state[0]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0006_),
    .Q(state[0]),
    .QN(_0004_)
  );
  DFF_X1 \state[1]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0007_),
    .Q(state[1]),
    .QN(_0003_)
  );
  DFF_X1 \state[2]$_SDFF_PP0_  (
    .CK(clock),
    .D(_0119_),
    .Q(state[2]),
    .QN(_0000_)
  );
  assign _GEN_0[64:32] = { _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65], _GEN_0[65] };
  assign _GEN_2[64:32] = { _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65], _GEN_2[65] };
  assign _GEN_35 = { remainder[65], remainder[65], remainder[65], remainder[65], remainder[65], remainder[65], remainder[65], remainder[65], remainder[65], remainder[65:33] };
  assign _decoded_T_4[1] = io_req_bits_fn[0];
  assign _decoded_T_6 = io_req_bits_fn[1];
  assign _decoded_T_7[0] = io_req_bits_fn[2];
  assign _decoded_orMatrixOutputs_T_4[0] = io_req_bits_fn[1];
  assign _divisor_T[31:0] = io_req_bits_in2;
  assign _prod_T_2 = { remainder[32], remainder[7:0] };
  assign _remainder_T_2[23:0] = remainder[31:8];
  assign { _state_T[2], _state_T[0] } = 2'h3;
  assign accum = remainder[65:33];
  assign decoded_andMatrixInput_0_3 = io_req_bits_fn[0];
  assign decoded_andMatrixInput_0_4 = io_req_bits_fn[1];
  assign decoded_andMatrixInput_1_2 = io_req_bits_fn[2];
  assign decoded_plaInput = io_req_bits_fn[2:0];
  assign hi = io_req_bits_in1[31:16];
  assign hi_1 = io_req_bits_in2[31:16];
  assign io_resp_bits_tag = req_tag;
  assign lhs_in = io_req_bits_in1;
  assign loOut = io_resp_bits_data[15:0];
  assign mplier = remainder[31:0];
  assign mplierSign = remainder[32];
  assign mulReg = { remainder[65:33], remainder[31:0] };
  assign negated_remainder[0] = io_resp_bits_data[0];
  assign nextMplierSign = _remainder_T_2[32];
  assign nextMulReg[64:0] = { _remainder_T_2[65:33], _remainder_T_2[31:24], remainder[31:8] };
  assign nextMulReg1 = { _remainder_T_2[65:33], _remainder_T_2[31:24], remainder[31:8] };
  assign nextMulReg_hi = { nextMulReg[65], _remainder_T_2[65:33], _remainder_T_2[31:24] };
  assign result = io_resp_bits_data;
  assign rhs_sign = _divisor_T[32];
  assign unrolls_0[32:1] = remainder[31:0];
endmodule
module PlusArgTimeout(clock, reset, io_count);
  input clock;
  wire clock;
  input [31:0] io_count;
  wire [31:0] io_count;
  input reset;
  wire reset;
endmodule
module RVCExpander(io_in, io_out_bits, io_out_rd, io_out_rs1, io_out_rs2, io_rvc);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire [30:0] _GEN_0;
  wire [30:0] _GEN_1;
  wire [31:0] _io_out_T_10_bits;
  wire [4:0] _io_out_T_10_rd;
  wire [4:0] _io_out_T_10_rs1;
  wire [31:0] _io_out_T_12_bits;
  wire [4:0] _io_out_T_12_rd;
  wire [4:0] _io_out_T_12_rs1;
  wire [31:0] _io_out_T_14_bits;
  wire [4:0] _io_out_T_14_rd;
  wire [4:0] _io_out_T_14_rs1;
  wire [31:0] _io_out_T_16_bits;
  wire [4:0] _io_out_T_16_rd;
  wire [4:0] _io_out_T_16_rs1;
  wire [31:0] _io_out_T_18_bits;
  wire [4:0] _io_out_T_18_rd;
  wire [4:0] _io_out_T_18_rs1;
  wire [4:0] _io_out_T_18_rs2;
  wire [4:0] _io_out_T_2;
  wire [31:0] _io_out_T_20_bits;
  wire [4:0] _io_out_T_20_rs2;
  wire [31:0] _io_out_T_22_bits;
  wire [4:0] _io_out_T_22_rs2;
  wire [31:0] _io_out_T_24_bits;
  wire [4:0] _io_out_T_24_rs2;
  wire [31:0] _io_out_T_26_bits;
  wire [4:0] _io_out_T_26_rs2;
  wire [31:0] _io_out_T_28_bits;
  wire [4:0] _io_out_T_28_rs2;
  wire [31:0] _io_out_T_30_bits;
  wire [4:0] _io_out_T_30_rs2;
  wire [31:0] _io_out_T_32_bits;
  wire [4:0] _io_out_T_32_rs2;
  wire [31:0] _io_out_T_34_bits;
  wire [31:0] _io_out_T_36_bits;
  wire [31:0] _io_out_T_38_bits;
  wire [31:0] _io_out_T_40_bits;
  wire [31:0] _io_out_T_42_bits;
  wire [31:0] _io_out_T_44_bits;
  wire [31:0] _io_out_T_46_bits;
  wire [31:0] _io_out_T_48_bits;
  wire [31:0] _io_out_T_4_bits;
  wire [4:0] _io_out_T_4_rd;
  wire [4:0] _io_out_T_4_rs1;
  wire [31:0] _io_out_T_6_bits;
  wire [4:0] _io_out_T_6_rd;
  wire [4:0] _io_out_T_6_rs1;
  wire [31:0] _io_out_T_8_bits;
  wire [4:0] _io_out_T_8_rd;
  wire [4:0] _io_out_T_8_rs1;
  wire [26:0] _io_out_s_T_116;
  wire [26:0] _io_out_s_T_138;
  wire [6:0] _io_out_s_T_148;
  wire [7:0] _io_out_s_T_15;
  wire [11:0] _io_out_s_T_150;
  wire [9:0] _io_out_s_T_161;
  wire [20:0] _io_out_s_T_169;
  wire [4:0] _io_out_s_T_17;
  wire [27:0] _io_out_s_T_20;
  wire [2:0] _io_out_s_T_230;
  wire [25:0] _io_out_s_T_251;
  wire [30:0] _io_out_s_T_260;
  wire [31:0] _io_out_s_T_270;
  wire [24:0] _io_out_s_T_277;
  wire [30:0] _io_out_s_T_278;
  wire [30:0] _io_out_s_T_281;
  wire [31:0] _io_out_s_T_283;
  wire [6:0] _io_out_s_T_31;
  wire [4:0] _io_out_s_T_349;
  wire [12:0] _io_out_s_T_354;
  wire [26:0] _io_out_s_T_36;
  wire [25:0] _io_out_s_T_438;
  wire [28:0] _io_out_s_T_448;
  wire [27:0] _io_out_s_T_457;
  wire [27:0] _io_out_s_T_466;
  wire [8:0] _io_out_s_T_473;
  wire [28:0] _io_out_s_T_480;
  wire [7:0] _io_out_s_T_486;
  wire [27:0] _io_out_s_T_493;
  wire [27:0] _io_out_s_T_506;
  wire [26:0] _io_out_s_T_52;
  wire [4:0] _io_out_s_T_6;
  wire [29:0] _io_out_s_T_7;
  wire [26:0] _io_out_s_T_74;
  wire [27:0] _io_out_s_T_94;
  wire [24:0] _io_out_s_add_T_3;
  wire [24:0] _io_out_s_ebreak_T_1;
  wire [2:0] _io_out_s_funct_T_2;
  wire [2:0] _io_out_s_funct_T_4;
  wire [2:0] _io_out_s_funct_T_6;
  wire [24:0] _io_out_s_jalr_ebreak_T_2;
  wire [24:0] _io_out_s_jr_reserved_T_2;
  wire _io_out_s_load_opc_T_1;
  wire [14:0] _io_out_s_me_T_2;
  wire [31:0] _io_out_s_me_T_4;
  wire [24:0] _io_out_s_mv_T_2;
  input [31:0] io_in;
  wire [31:0] io_in;
  output [31:0] io_out_bits;
  wire [31:0] io_out_bits;
  output [4:0] io_out_rd;
  wire [4:0] io_out_rd;
  output [4:0] io_out_rs1;
  wire [4:0] io_out_rs1;
  output [4:0] io_out_rs2;
  wire [4:0] io_out_rs2;
  wire [31:0] io_out_s_0_bits;
  wire [31:0] io_out_s_10_bits;
  wire [31:0] io_out_s_11_bits;
  wire [4:0] io_out_s_11_rd;
  wire [4:0] io_out_s_11_rs2;
  wire [31:0] io_out_s_12_bits;
  wire [31:0] io_out_s_13_bits;
  wire [31:0] io_out_s_14_bits;
  wire [31:0] io_out_s_15_bits;
  wire [31:0] io_out_s_16_bits;
  wire [31:0] io_out_s_17_bits;
  wire [31:0] io_out_s_18_bits;
  wire [31:0] io_out_s_19_bits;
  wire [31:0] io_out_s_1_bits;
  wire [31:0] io_out_s_20_bits;
  wire [4:0] io_out_s_20_rd;
  wire [4:0] io_out_s_20_rs1;
  wire [4:0] io_out_s_20_rs2;
  wire [31:0] io_out_s_21_bits;
  wire [31:0] io_out_s_22_bits;
  wire [31:0] io_out_s_23_bits;
  wire [4:0] io_out_s_24_rs1;
  wire [4:0] io_out_s_24_rs2;
  wire [31:0] io_out_s_2_bits;
  wire [31:0] io_out_s_3_bits;
  wire [31:0] io_out_s_4_bits;
  wire [31:0] io_out_s_5_bits;
  wire [31:0] io_out_s_6_bits;
  wire [31:0] io_out_s_7_bits;
  wire [31:0] io_out_s_8_bits;
  wire [31:0] io_out_s_9_bits;
  wire [31:0] io_out_s_add_bits;
  wire [24:0] io_out_s_ebreak;
  wire [2:0] io_out_s_funct;
  wire [24:0] io_out_s_jalr;
  wire [31:0] io_out_s_jalr_add_bits;
  wire [4:0] io_out_s_jalr_add_rd;
  wire [4:0] io_out_s_jalr_add_rs1;
  wire [31:0] io_out_s_jalr_ebreak_bits;
  wire [24:0] io_out_s_jr;
  wire [31:0] io_out_s_jr_mv_bits;
  wire [4:0] io_out_s_jr_mv_rd;
  wire [4:0] io_out_s_jr_mv_rs1;
  wire [4:0] io_out_s_jr_mv_rs2;
  wire [31:0] io_out_s_jr_reserved_bits;
  wire [6:0] io_out_s_load_opc;
  wire [31:0] io_out_s_me_bits;
  wire [31:0] io_out_s_mv_bits;
  wire [6:0] io_out_s_opc;
  wire [6:0] io_out_s_opc_1;
  wire [6:0] io_out_s_opc_2;
  wire [6:0] io_out_s_opc_3;
  wire [31:0] io_out_s_res_bits;
  wire [24:0] io_out_s_reserved;
  wire [30:0] io_out_s_sub;
  output io_rvc;
  wire io_rvc;
  INV_X1 _0618_ (
    .A(io_in[12]),
    .ZN(_0601_)
  );
  INV_X1 _0619_ (
    .A(io_in[8]),
    .ZN(_0602_)
  );
  INV_X1 _0620_ (
    .A(io_in[11]),
    .ZN(_0603_)
  );
  INV_X1 _0621_ (
    .A(io_in[10]),
    .ZN(_0604_)
  );
  INV_X1 _0622_ (
    .A(io_in[0]),
    .ZN(_0605_)
  );
  INV_X1 _0623_ (
    .A(io_in[14]),
    .ZN(_0606_)
  );
  INV_X1 _0624_ (
    .A(io_in[13]),
    .ZN(_0607_)
  );
  INV_X1 _0625_ (
    .A(io_in[1]),
    .ZN(_0608_)
  );
  INV_X1 _0626_ (
    .A(io_in[15]),
    .ZN(_0609_)
  );
  AND2_X1 _0627_ (
    .A1(io_in[0]),
    .A2(io_in[1]),
    .ZN(_0610_)
  );
  INV_X1 _0628_ (
    .A(_0610_),
    .ZN(io_rvc)
  );
  OR2_X1 _0629_ (
    .A1(io_in[2]),
    .A2(io_rvc),
    .ZN(_0611_)
  );
  OR2_X1 _0630_ (
    .A1(io_in[6]),
    .A2(io_in[5]),
    .ZN(_0612_)
  );
  INV_X1 _0631_ (
    .A(_0612_),
    .ZN(_0613_)
  );
  OR2_X1 _0632_ (
    .A1(io_in[2]),
    .A2(io_in[3]),
    .ZN(_0614_)
  );
  OR2_X1 _0633_ (
    .A1(io_in[4]),
    .A2(_0614_),
    .ZN(_0615_)
  );
  INV_X1 _0634_ (
    .A(_0615_),
    .ZN(_0616_)
  );
  AND2_X1 _0635_ (
    .A1(_0613_),
    .A2(_0616_),
    .ZN(_0617_)
  );
  OR2_X1 _0636_ (
    .A1(_0612_),
    .A2(_0615_),
    .ZN(_0000_)
  );
  AND2_X1 _0637_ (
    .A1(_0601_),
    .A2(_0617_),
    .ZN(_0001_)
  );
  OR2_X1 _0638_ (
    .A1(io_in[12]),
    .A2(_0000_),
    .ZN(_0002_)
  );
  OR2_X1 _0639_ (
    .A1(io_in[11]),
    .A2(io_in[10]),
    .ZN(_0003_)
  );
  INV_X1 _0640_ (
    .A(_0003_),
    .ZN(_0004_)
  );
  OR2_X1 _0641_ (
    .A1(io_in[7]),
    .A2(io_in[9]),
    .ZN(_0005_)
  );
  INV_X1 _0642_ (
    .A(_0005_),
    .ZN(_0006_)
  );
  AND2_X1 _0643_ (
    .A1(_0004_),
    .A2(_0006_),
    .ZN(_0007_)
  );
  OR2_X1 _0644_ (
    .A1(_0003_),
    .A2(_0005_),
    .ZN(_0008_)
  );
  AND2_X1 _0645_ (
    .A1(_0602_),
    .A2(_0007_),
    .ZN(_0009_)
  );
  OR2_X1 _0646_ (
    .A1(io_in[8]),
    .A2(_0008_),
    .ZN(_0010_)
  );
  AND2_X1 _0647_ (
    .A1(_0617_),
    .A2(_0010_),
    .ZN(_0011_)
  );
  AND2_X1 _0648_ (
    .A1(_0606_),
    .A2(_0607_),
    .ZN(_0012_)
  );
  OR2_X1 _0649_ (
    .A1(io_in[14]),
    .A2(io_in[13]),
    .ZN(_0013_)
  );
  AND2_X1 _0650_ (
    .A1(_0605_),
    .A2(io_in[15]),
    .ZN(_0014_)
  );
  OR2_X1 _0651_ (
    .A1(io_in[0]),
    .A2(_0609_),
    .ZN(_0015_)
  );
  AND2_X1 _0652_ (
    .A1(io_in[1]),
    .A2(_0014_),
    .ZN(_0016_)
  );
  OR2_X1 _0653_ (
    .A1(_0608_),
    .A2(_0015_),
    .ZN(_0017_)
  );
  AND2_X1 _0654_ (
    .A1(io_in[1]),
    .A2(_0012_),
    .ZN(_0018_)
  );
  AND2_X1 _0655_ (
    .A1(_0012_),
    .A2(_0016_),
    .ZN(_0019_)
  );
  OR2_X1 _0656_ (
    .A1(_0013_),
    .A2(_0017_),
    .ZN(_0020_)
  );
  OR2_X1 _0657_ (
    .A1(_0011_),
    .A2(_0020_),
    .ZN(_0021_)
  );
  INV_X1 _0658_ (
    .A(_0021_),
    .ZN(_0022_)
  );
  OR2_X1 _0659_ (
    .A1(_0001_),
    .A2(_0021_),
    .ZN(_0023_)
  );
  OR2_X1 _0660_ (
    .A1(io_in[0]),
    .A2(io_in[15]),
    .ZN(_0024_)
  );
  INV_X1 _0661_ (
    .A(_0024_),
    .ZN(_0025_)
  );
  AND2_X1 _0662_ (
    .A1(io_in[1]),
    .A2(_0025_),
    .ZN(_0026_)
  );
  OR2_X1 _0663_ (
    .A1(_0608_),
    .A2(_0024_),
    .ZN(_0027_)
  );
  AND2_X1 _0664_ (
    .A1(io_in[14]),
    .A2(io_in[1]),
    .ZN(_0028_)
  );
  AND2_X1 _0665_ (
    .A1(_0025_),
    .A2(_0028_),
    .ZN(_0029_)
  );
  OR2_X1 _0666_ (
    .A1(_0606_),
    .A2(io_in[13]),
    .ZN(_0030_)
  );
  OR2_X1 _0667_ (
    .A1(_0027_),
    .A2(_0030_),
    .ZN(_0031_)
  );
  INV_X1 _0668_ (
    .A(_0031_),
    .ZN(_0032_)
  );
  AND2_X1 _0669_ (
    .A1(_0608_),
    .A2(_0014_),
    .ZN(_0033_)
  );
  OR2_X1 _0670_ (
    .A1(io_in[1]),
    .A2(_0015_),
    .ZN(_0034_)
  );
  OR2_X1 _0671_ (
    .A1(_0606_),
    .A2(_0034_),
    .ZN(_0035_)
  );
  AND2_X1 _0672_ (
    .A1(io_in[14]),
    .A2(io_in[13]),
    .ZN(_0036_)
  );
  OR2_X1 _0673_ (
    .A1(_0606_),
    .A2(_0607_),
    .ZN(_0037_)
  );
  OR2_X1 _0674_ (
    .A1(_0034_),
    .A2(_0037_),
    .ZN(_0038_)
  );
  AND2_X1 _0675_ (
    .A1(_0606_),
    .A2(io_in[13]),
    .ZN(_0039_)
  );
  OR2_X1 _0676_ (
    .A1(io_in[14]),
    .A2(_0607_),
    .ZN(_0040_)
  );
  AND2_X1 _0677_ (
    .A1(_0608_),
    .A2(_0039_),
    .ZN(_0041_)
  );
  OR2_X1 _0678_ (
    .A1(io_in[1]),
    .A2(_0040_),
    .ZN(_0042_)
  );
  AND2_X1 _0679_ (
    .A1(_0025_),
    .A2(_0041_),
    .ZN(_0043_)
  );
  OR2_X1 _0680_ (
    .A1(_0024_),
    .A2(_0042_),
    .ZN(_0044_)
  );
  OR2_X1 _0681_ (
    .A1(io_in[12]),
    .A2(_0010_),
    .ZN(_0045_)
  );
  INV_X1 _0682_ (
    .A(_0045_),
    .ZN(_0046_)
  );
  AND2_X1 _0683_ (
    .A1(_0613_),
    .A2(_0046_),
    .ZN(_0047_)
  );
  OR2_X1 _0684_ (
    .A1(_0043_),
    .A2(_0047_),
    .ZN(_0048_)
  );
  OR2_X1 _0685_ (
    .A1(io_in[1]),
    .A2(_0030_),
    .ZN(_0049_)
  );
  INV_X1 _0686_ (
    .A(_0049_),
    .ZN(_0050_)
  );
  OR2_X1 _0687_ (
    .A1(_0024_),
    .A2(_0049_),
    .ZN(_0051_)
  );
  AND2_X1 _0688_ (
    .A1(_0048_),
    .A2(_0051_),
    .ZN(_0052_)
  );
  OR2_X1 _0689_ (
    .A1(_0024_),
    .A2(_0037_),
    .ZN(_0053_)
  );
  OR2_X1 _0690_ (
    .A1(io_in[14]),
    .A2(_0015_),
    .ZN(_0054_)
  );
  AND2_X1 _0691_ (
    .A1(_0053_),
    .A2(_0054_),
    .ZN(_0055_)
  );
  OR2_X1 _0692_ (
    .A1(io_in[1]),
    .A2(_0055_),
    .ZN(_0056_)
  );
  INV_X1 _0693_ (
    .A(_0056_),
    .ZN(_0057_)
  );
  OR2_X1 _0694_ (
    .A1(_0052_),
    .A2(_0057_),
    .ZN(_0058_)
  );
  MUX2_X1 _0695_ (
    .A(io_in[13]),
    .B(_0058_),
    .S(_0035_),
    .Z(_0059_)
  );
  AND2_X1 _0696_ (
    .A1(_0608_),
    .A2(_0036_),
    .ZN(_0060_)
  );
  AND2_X1 _0697_ (
    .A1(io_in[0]),
    .A2(_0609_),
    .ZN(_0061_)
  );
  OR2_X1 _0698_ (
    .A1(_0605_),
    .A2(io_in[15]),
    .ZN(_0062_)
  );
  OR2_X1 _0699_ (
    .A1(_0037_),
    .A2(_0062_),
    .ZN(_0063_)
  );
  AND2_X1 _0700_ (
    .A1(_0060_),
    .A2(_0061_),
    .ZN(_0064_)
  );
  OR2_X1 _0701_ (
    .A1(io_in[1]),
    .A2(_0063_),
    .ZN(_0065_)
  );
  AND2_X1 _0702_ (
    .A1(_0050_),
    .A2(_0061_),
    .ZN(_0066_)
  );
  OR2_X1 _0703_ (
    .A1(_0049_),
    .A2(_0062_),
    .ZN(_0067_)
  );
  AND2_X1 _0704_ (
    .A1(_0065_),
    .A2(_0067_),
    .ZN(_0068_)
  );
  OR2_X1 _0705_ (
    .A1(_0064_),
    .A2(_0066_),
    .ZN(_0069_)
  );
  OR2_X1 _0706_ (
    .A1(io_in[1]),
    .A2(_0013_),
    .ZN(_0070_)
  );
  INV_X1 _0707_ (
    .A(_0070_),
    .ZN(_0071_)
  );
  AND2_X1 _0708_ (
    .A1(_0061_),
    .A2(_0071_),
    .ZN(_0072_)
  );
  OR2_X1 _0709_ (
    .A1(_0062_),
    .A2(_0070_),
    .ZN(_0073_)
  );
  OR2_X1 _0710_ (
    .A1(_0066_),
    .A2(_0072_),
    .ZN(_0074_)
  );
  AND2_X1 _0711_ (
    .A1(_0068_),
    .A2(_0073_),
    .ZN(_0075_)
  );
  AND2_X1 _0712_ (
    .A1(_0059_),
    .A2(_0075_),
    .ZN(_0076_)
  );
  AND2_X1 _0713_ (
    .A1(_0008_),
    .A2(_0064_),
    .ZN(_0077_)
  );
  AND2_X1 _0714_ (
    .A1(_0001_),
    .A2(_0064_),
    .ZN(_0078_)
  );
  AND2_X1 _0715_ (
    .A1(io_in[0]),
    .A2(_0041_),
    .ZN(_0079_)
  );
  OR2_X1 _0716_ (
    .A1(_0605_),
    .A2(_0042_),
    .ZN(_0080_)
  );
  AND2_X1 _0717_ (
    .A1(_0041_),
    .A2(_0061_),
    .ZN(_0081_)
  );
  OR2_X1 _0718_ (
    .A1(_0042_),
    .A2(_0062_),
    .ZN(_0082_)
  );
  OR2_X1 _0719_ (
    .A1(_0078_),
    .A2(_0081_),
    .ZN(_0083_)
  );
  OR2_X1 _0720_ (
    .A1(_0077_),
    .A2(_0083_),
    .ZN(_0084_)
  );
  OR2_X1 _0721_ (
    .A1(_0076_),
    .A2(_0084_),
    .ZN(_0085_)
  );
  AND2_X1 _0722_ (
    .A1(_0012_),
    .A2(_0026_),
    .ZN(_0086_)
  );
  INV_X1 _0723_ (
    .A(_0086_),
    .ZN(_0087_)
  );
  AND2_X1 _0724_ (
    .A1(io_in[0]),
    .A2(_0608_),
    .ZN(_0088_)
  );
  OR2_X1 _0725_ (
    .A1(_0605_),
    .A2(io_in[1]),
    .ZN(_0089_)
  );
  AND2_X1 _0726_ (
    .A1(io_in[15]),
    .A2(_0088_),
    .ZN(_0090_)
  );
  OR2_X1 _0727_ (
    .A1(_0609_),
    .A2(_0089_),
    .ZN(_0091_)
  );
  AND2_X1 _0728_ (
    .A1(io_in[0]),
    .A2(io_in[15]),
    .ZN(_0092_)
  );
  AND2_X1 _0729_ (
    .A1(_0050_),
    .A2(_0092_),
    .ZN(_0093_)
  );
  OR2_X1 _0730_ (
    .A1(_0037_),
    .A2(_0091_),
    .ZN(_0094_)
  );
  OR2_X1 _0731_ (
    .A1(_0606_),
    .A2(_0091_),
    .ZN(_0095_)
  );
  AND2_X1 _0732_ (
    .A1(io_in[14]),
    .A2(_0090_),
    .ZN(_0096_)
  );
  AND2_X1 _0733_ (
    .A1(_0012_),
    .A2(_0090_),
    .ZN(_0097_)
  );
  OR2_X1 _0734_ (
    .A1(_0013_),
    .A2(_0091_),
    .ZN(_0098_)
  );
  OR2_X1 _0735_ (
    .A1(_0039_),
    .A2(_0091_),
    .ZN(_0099_)
  );
  INV_X1 _0736_ (
    .A(_0099_),
    .ZN(_0100_)
  );
  OR2_X1 _0737_ (
    .A1(_0086_),
    .A2(_0097_),
    .ZN(_0101_)
  );
  AND2_X1 _0738_ (
    .A1(_0087_),
    .A2(_0095_),
    .ZN(_0102_)
  );
  OR2_X1 _0739_ (
    .A1(_0086_),
    .A2(_0100_),
    .ZN(_0103_)
  );
  INV_X1 _0740_ (
    .A(_0103_),
    .ZN(_0104_)
  );
  AND2_X1 _0741_ (
    .A1(_0085_),
    .A2(_0104_),
    .ZN(_0105_)
  );
  OR2_X1 _0742_ (
    .A1(io_in[14]),
    .A2(_0027_),
    .ZN(_0106_)
  );
  AND2_X1 _0743_ (
    .A1(_0026_),
    .A2(_0039_),
    .ZN(_0107_)
  );
  AND2_X1 _0744_ (
    .A1(_0039_),
    .A2(_0092_),
    .ZN(_0108_)
  );
  AND2_X1 _0745_ (
    .A1(_0039_),
    .A2(_0090_),
    .ZN(_0109_)
  );
  OR2_X1 _0746_ (
    .A1(_0040_),
    .A2(_0091_),
    .ZN(_0110_)
  );
  OR2_X1 _0747_ (
    .A1(_0107_),
    .A2(_0109_),
    .ZN(_0111_)
  );
  OR2_X1 _0748_ (
    .A1(_0105_),
    .A2(_0111_),
    .ZN(_0112_)
  );
  OR2_X1 _0749_ (
    .A1(_0027_),
    .A2(_0037_),
    .ZN(_0113_)
  );
  AND2_X1 _0750_ (
    .A1(_0020_),
    .A2(_0113_),
    .ZN(_0114_)
  );
  INV_X1 _0751_ (
    .A(_0114_),
    .ZN(_0115_)
  );
  AND2_X1 _0752_ (
    .A1(_0009_),
    .A2(_0032_),
    .ZN(_0116_)
  );
  MUX2_X1 _0753_ (
    .A(_0009_),
    .B(_0112_),
    .S(_0031_),
    .Z(_0117_)
  );
  OR2_X1 _0754_ (
    .A1(_0115_),
    .A2(_0117_),
    .ZN(_0118_)
  );
  AND2_X1 _0755_ (
    .A1(_0023_),
    .A2(_0118_),
    .ZN(_0119_)
  );
  AND2_X1 _0756_ (
    .A1(_0014_),
    .A2(_0039_),
    .ZN(_0120_)
  );
  AND2_X1 _0757_ (
    .A1(_0016_),
    .A2(_0039_),
    .ZN(_0121_)
  );
  OR2_X1 _0758_ (
    .A1(_0119_),
    .A2(_0121_),
    .ZN(_0122_)
  );
  OR2_X1 _0759_ (
    .A1(_0017_),
    .A2(_0030_),
    .ZN(_0123_)
  );
  AND2_X1 _0760_ (
    .A1(_0122_),
    .A2(_0123_),
    .ZN(_0124_)
  );
  AND2_X1 _0761_ (
    .A1(_0016_),
    .A2(_0036_),
    .ZN(_0125_)
  );
  OR2_X1 _0762_ (
    .A1(_0610_),
    .A2(_0125_),
    .ZN(_0126_)
  );
  OR2_X1 _0763_ (
    .A1(_0124_),
    .A2(_0126_),
    .ZN(_0127_)
  );
  AND2_X1 _0764_ (
    .A1(_0611_),
    .A2(_0127_),
    .ZN(io_out_bits[2])
  );
  AND2_X1 _0765_ (
    .A1(io_in[3]),
    .A2(_0610_),
    .ZN(_0128_)
  );
  AND2_X1 _0766_ (
    .A1(_0027_),
    .A2(_0094_),
    .ZN(_0129_)
  );
  AND2_X1 _0767_ (
    .A1(_0027_),
    .A2(_0095_),
    .ZN(_0130_)
  );
  INV_X1 _0768_ (
    .A(_0130_),
    .ZN(_0131_)
  );
  OR2_X1 _0769_ (
    .A1(_0012_),
    .A2(_0024_),
    .ZN(_0132_)
  );
  OR2_X1 _0770_ (
    .A1(io_in[1]),
    .A2(_0132_),
    .ZN(_0133_)
  );
  INV_X1 _0771_ (
    .A(_0133_),
    .ZN(_0134_)
  );
  AND2_X1 _0772_ (
    .A1(_0047_),
    .A2(_0133_),
    .ZN(_0135_)
  );
  AND2_X1 _0773_ (
    .A1(_0012_),
    .A2(_0033_),
    .ZN(_0136_)
  );
  OR2_X1 _0774_ (
    .A1(_0135_),
    .A2(_0136_),
    .ZN(_0137_)
  );
  OR2_X1 _0775_ (
    .A1(_0015_),
    .A2(_0042_),
    .ZN(_0138_)
  );
  INV_X1 _0776_ (
    .A(_0138_),
    .ZN(_0139_)
  );
  AND2_X1 _0777_ (
    .A1(_0035_),
    .A2(_0138_),
    .ZN(_0140_)
  );
  AND2_X1 _0778_ (
    .A1(_0075_),
    .A2(_0140_),
    .ZN(_0141_)
  );
  AND2_X1 _0779_ (
    .A1(_0035_),
    .A2(_0073_),
    .ZN(_0142_)
  );
  AND2_X1 _0780_ (
    .A1(_0137_),
    .A2(_0141_),
    .ZN(_0143_)
  );
  OR2_X1 _0781_ (
    .A1(_0083_),
    .A2(_0143_),
    .ZN(_0144_)
  );
  AND2_X1 _0782_ (
    .A1(_0098_),
    .A2(_0144_),
    .ZN(_0145_)
  );
  AND2_X1 _0783_ (
    .A1(io_in[11]),
    .A2(io_in[10]),
    .ZN(_0146_)
  );
  OR2_X1 _0784_ (
    .A1(_0603_),
    .A2(_0604_),
    .ZN(_0147_)
  );
  AND2_X1 _0785_ (
    .A1(_0097_),
    .A2(_0146_),
    .ZN(_0148_)
  );
  INV_X1 _0786_ (
    .A(_0148_),
    .ZN(_0149_)
  );
  AND2_X1 _0787_ (
    .A1(io_in[12]),
    .A2(_0148_),
    .ZN(_0150_)
  );
  OR2_X1 _0788_ (
    .A1(_0109_),
    .A2(_0150_),
    .ZN(_0151_)
  );
  OR2_X1 _0789_ (
    .A1(_0145_),
    .A2(_0151_),
    .ZN(_0152_)
  );
  AND2_X1 _0790_ (
    .A1(_0130_),
    .A2(_0152_),
    .ZN(_0153_)
  );
  OR2_X1 _0791_ (
    .A1(_0019_),
    .A2(_0116_),
    .ZN(_0154_)
  );
  OR2_X1 _0792_ (
    .A1(_0153_),
    .A2(_0154_),
    .ZN(_0155_)
  );
  AND2_X1 _0793_ (
    .A1(_0009_),
    .A2(_0012_),
    .ZN(_0156_)
  );
  OR2_X1 _0794_ (
    .A1(_0010_),
    .A2(_0013_),
    .ZN(_0157_)
  );
  AND2_X1 _0795_ (
    .A1(_0617_),
    .A2(_0009_),
    .ZN(_0158_)
  );
  AND2_X1 _0796_ (
    .A1(_0001_),
    .A2(_0156_),
    .ZN(_0159_)
  );
  OR2_X1 _0797_ (
    .A1(_0002_),
    .A2(_0157_),
    .ZN(_0160_)
  );
  AND2_X1 _0798_ (
    .A1(_0016_),
    .A2(_0160_),
    .ZN(_0161_)
  );
  OR2_X1 _0799_ (
    .A1(_0017_),
    .A2(_0159_),
    .ZN(_0162_)
  );
  AND2_X1 _0800_ (
    .A1(io_rvc),
    .A2(_0162_),
    .ZN(_0163_)
  );
  AND2_X1 _0801_ (
    .A1(_0155_),
    .A2(_0163_),
    .ZN(_0164_)
  );
  OR2_X1 _0802_ (
    .A1(_0128_),
    .A2(_0164_),
    .ZN(io_out_bits[3])
  );
  AND2_X1 _0803_ (
    .A1(io_in[4]),
    .A2(_0610_),
    .ZN(_0165_)
  );
  AND2_X1 _0804_ (
    .A1(io_in[1]),
    .A2(_0013_),
    .ZN(_0166_)
  );
  AND2_X1 _0805_ (
    .A1(_0014_),
    .A2(_0166_),
    .ZN(_0167_)
  );
  INV_X1 _0806_ (
    .A(_0167_),
    .ZN(_0168_)
  );
  AND2_X1 _0807_ (
    .A1(io_in[1]),
    .A2(_0108_),
    .ZN(_0169_)
  );
  AND2_X1 _0808_ (
    .A1(_0018_),
    .A2(_0092_),
    .ZN(_0170_)
  );
  OR2_X1 _0809_ (
    .A1(_0169_),
    .A2(_0170_),
    .ZN(_0171_)
  );
  AND2_X1 _0810_ (
    .A1(_0028_),
    .A2(_0092_),
    .ZN(_0172_)
  );
  AND2_X1 _0811_ (
    .A1(io_in[15]),
    .A2(_0610_),
    .ZN(_0173_)
  );
  AND2_X1 _0812_ (
    .A1(_0018_),
    .A2(_0061_),
    .ZN(_0174_)
  );
  AND2_X1 _0813_ (
    .A1(_0609_),
    .A2(_0610_),
    .ZN(_0175_)
  );
  AND2_X1 _0814_ (
    .A1(io_rvc),
    .A2(_0168_),
    .ZN(_0176_)
  );
  OR2_X1 _0815_ (
    .A1(_0610_),
    .A2(_0167_),
    .ZN(_0177_)
  );
  AND2_X1 _0816_ (
    .A1(_0030_),
    .A2(_0040_),
    .ZN(_0178_)
  );
  OR2_X1 _0817_ (
    .A1(_0034_),
    .A2(_0178_),
    .ZN(_0179_)
  );
  OR2_X1 _0818_ (
    .A1(_0033_),
    .A2(_0134_),
    .ZN(_0180_)
  );
  AND2_X1 _0819_ (
    .A1(_0133_),
    .A2(_0179_),
    .ZN(_0181_)
  );
  AND2_X1 _0820_ (
    .A1(_0038_),
    .A2(_0181_),
    .ZN(_0182_)
  );
  OR2_X1 _0821_ (
    .A1(_0091_),
    .A2(_0178_),
    .ZN(_0183_)
  );
  OR2_X1 _0822_ (
    .A1(_0012_),
    .A2(_0091_),
    .ZN(_0184_)
  );
  AND2_X1 _0823_ (
    .A1(_0013_),
    .A2(_0090_),
    .ZN(_0185_)
  );
  OR2_X1 _0824_ (
    .A1(_0081_),
    .A2(_0185_),
    .ZN(_0186_)
  );
  INV_X1 _0825_ (
    .A(_0186_),
    .ZN(_0187_)
  );
  AND2_X1 _0826_ (
    .A1(_0025_),
    .A2(_0166_),
    .ZN(_0188_)
  );
  OR2_X1 _0827_ (
    .A1(_0012_),
    .A2(_0027_),
    .ZN(_0189_)
  );
  OR2_X1 _0828_ (
    .A1(_0036_),
    .A2(_0189_),
    .ZN(_0190_)
  );
  AND2_X1 _0829_ (
    .A1(_0182_),
    .A2(_0187_),
    .ZN(_0191_)
  );
  AND2_X1 _0830_ (
    .A1(_0190_),
    .A2(_0191_),
    .ZN(_0192_)
  );
  OR2_X1 _0831_ (
    .A1(_0116_),
    .A2(_0192_),
    .ZN(_0193_)
  );
  AND2_X1 _0832_ (
    .A1(_0114_),
    .A2(_0193_),
    .ZN(_0194_)
  );
  OR2_X1 _0833_ (
    .A1(_0022_),
    .A2(_0194_),
    .ZN(_0195_)
  );
  AND2_X1 _0834_ (
    .A1(_0176_),
    .A2(_0195_),
    .ZN(_0196_)
  );
  OR2_X1 _0835_ (
    .A1(_0165_),
    .A2(_0196_),
    .ZN(io_out_bits[4])
  );
  OR2_X1 _0836_ (
    .A1(_0148_),
    .A2(_0186_),
    .ZN(_0197_)
  );
  AND2_X1 _0837_ (
    .A1(io_in[5]),
    .A2(_0610_),
    .ZN(_0198_)
  );
  OR2_X1 _0838_ (
    .A1(_0033_),
    .A2(_0198_),
    .ZN(_0199_)
  );
  OR2_X1 _0839_ (
    .A1(_0077_),
    .A2(_0199_),
    .ZN(_0200_)
  );
  OR2_X1 _0840_ (
    .A1(_0197_),
    .A2(_0200_),
    .ZN(_0201_)
  );
  OR2_X1 _0841_ (
    .A1(_0161_),
    .A2(_0201_),
    .ZN(io_out_bits[5])
  );
  AND2_X1 _0842_ (
    .A1(_0617_),
    .A2(_0019_),
    .ZN(_0202_)
  );
  AND2_X1 _0843_ (
    .A1(_0045_),
    .A2(_0202_),
    .ZN(_0203_)
  );
  AND2_X1 _0844_ (
    .A1(io_in[6]),
    .A2(_0610_),
    .ZN(_0204_)
  );
  OR2_X1 _0845_ (
    .A1(_0186_),
    .A2(_0204_),
    .ZN(_0205_)
  );
  OR2_X1 _0846_ (
    .A1(_0203_),
    .A2(_0205_),
    .ZN(io_out_bits[6])
  );
  AND2_X1 _0847_ (
    .A1(io_in[7]),
    .A2(_0610_),
    .ZN(_0206_)
  );
  AND2_X1 _0848_ (
    .A1(io_in[7]),
    .A2(_0072_),
    .ZN(_0207_)
  );
  OR2_X1 _0849_ (
    .A1(_0081_),
    .A2(_0207_),
    .ZN(_0208_)
  );
  AND2_X1 _0850_ (
    .A1(_0034_),
    .A2(_0073_),
    .ZN(_0209_)
  );
  OR2_X1 _0851_ (
    .A1(_0033_),
    .A2(_0072_),
    .ZN(_0210_)
  );
  AND2_X1 _0852_ (
    .A1(io_in[2]),
    .A2(_0209_),
    .ZN(_0211_)
  );
  OR2_X1 _0853_ (
    .A1(_0208_),
    .A2(_0211_),
    .ZN(_0212_)
  );
  AND2_X1 _0854_ (
    .A1(_0068_),
    .A2(_0098_),
    .ZN(_0213_)
  );
  OR2_X1 _0855_ (
    .A1(_0069_),
    .A2(_0097_),
    .ZN(_0214_)
  );
  MUX2_X1 _0856_ (
    .A(io_in[7]),
    .B(_0212_),
    .S(_0213_),
    .Z(_0215_)
  );
  AND2_X1 _0857_ (
    .A1(_0184_),
    .A2(_0215_),
    .ZN(_0216_)
  );
  AND2_X1 _0858_ (
    .A1(io_in[12]),
    .A2(_0096_),
    .ZN(_0217_)
  );
  OR2_X1 _0859_ (
    .A1(_0216_),
    .A2(_0217_),
    .ZN(_0218_)
  );
  AND2_X1 _0860_ (
    .A1(_0027_),
    .A2(_0218_),
    .ZN(_0219_)
  );
  AND2_X1 _0861_ (
    .A1(io_in[7]),
    .A2(_0026_),
    .ZN(_0220_)
  );
  OR2_X1 _0862_ (
    .A1(_0019_),
    .A2(_0220_),
    .ZN(_0221_)
  );
  OR2_X1 _0863_ (
    .A1(_0219_),
    .A2(_0221_),
    .ZN(_0222_)
  );
  AND2_X1 _0864_ (
    .A1(io_in[12]),
    .A2(_0011_),
    .ZN(_0223_)
  );
  AND2_X1 _0865_ (
    .A1(io_in[7]),
    .A2(_0000_),
    .ZN(_0224_)
  );
  OR2_X1 _0866_ (
    .A1(_0020_),
    .A2(_0224_),
    .ZN(_0225_)
  );
  OR2_X1 _0867_ (
    .A1(_0223_),
    .A2(_0225_),
    .ZN(_0226_)
  );
  AND2_X1 _0868_ (
    .A1(_0176_),
    .A2(_0226_),
    .ZN(_0227_)
  );
  AND2_X1 _0869_ (
    .A1(_0222_),
    .A2(_0227_),
    .ZN(_0228_)
  );
  OR2_X1 _0870_ (
    .A1(_0206_),
    .A2(_0228_),
    .ZN(io_out_bits[7])
  );
  AND2_X1 _0871_ (
    .A1(io_in[8]),
    .A2(_0610_),
    .ZN(_0229_)
  );
  AND2_X1 _0872_ (
    .A1(_0000_),
    .A2(_0019_),
    .ZN(_0230_)
  );
  AND2_X1 _0873_ (
    .A1(io_in[8]),
    .A2(_0230_),
    .ZN(_0231_)
  );
  AND2_X1 _0874_ (
    .A1(io_in[8]),
    .A2(_0026_),
    .ZN(_0232_)
  );
  AND2_X1 _0875_ (
    .A1(io_in[8]),
    .A2(_0214_),
    .ZN(_0233_)
  );
  AND2_X1 _0876_ (
    .A1(io_in[8]),
    .A2(_0072_),
    .ZN(_0234_)
  );
  AND2_X1 _0877_ (
    .A1(io_in[3]),
    .A2(_0209_),
    .ZN(_0235_)
  );
  OR2_X1 _0878_ (
    .A1(_0234_),
    .A2(_0235_),
    .ZN(_0236_)
  );
  AND2_X1 _0879_ (
    .A1(_0082_),
    .A2(_0213_),
    .ZN(_0237_)
  );
  OR2_X1 _0880_ (
    .A1(_0064_),
    .A2(_0081_),
    .ZN(_0238_)
  );
  AND2_X1 _0881_ (
    .A1(_0236_),
    .A2(_0237_),
    .ZN(_0239_)
  );
  OR2_X1 _0882_ (
    .A1(_0233_),
    .A2(_0239_),
    .ZN(_0240_)
  );
  AND2_X1 _0883_ (
    .A1(_0027_),
    .A2(_0110_),
    .ZN(_0241_)
  );
  AND2_X1 _0884_ (
    .A1(_0240_),
    .A2(_0241_),
    .ZN(_0242_)
  );
  OR2_X1 _0885_ (
    .A1(_0232_),
    .A2(_0242_),
    .ZN(_0243_)
  );
  AND2_X1 _0886_ (
    .A1(_0020_),
    .A2(_0243_),
    .ZN(_0244_)
  );
  OR2_X1 _0887_ (
    .A1(_0231_),
    .A2(_0244_),
    .ZN(_0245_)
  );
  AND2_X1 _0888_ (
    .A1(_0176_),
    .A2(_0245_),
    .ZN(_0246_)
  );
  OR2_X1 _0889_ (
    .A1(_0229_),
    .A2(_0246_),
    .ZN(io_out_bits[8])
  );
  AND2_X1 _0890_ (
    .A1(io_in[9]),
    .A2(_0026_),
    .ZN(_0247_)
  );
  AND2_X1 _0891_ (
    .A1(io_in[9]),
    .A2(_0214_),
    .ZN(_0248_)
  );
  OR2_X1 _0892_ (
    .A1(io_in[6]),
    .A2(_0039_),
    .ZN(_0249_)
  );
  MUX2_X1 _0893_ (
    .A(io_in[4]),
    .B(_0249_),
    .S(_0033_),
    .Z(_0250_)
  );
  AND2_X1 _0894_ (
    .A1(_0138_),
    .A2(_0250_),
    .ZN(_0251_)
  );
  MUX2_X1 _0895_ (
    .A(io_in[9]),
    .B(_0251_),
    .S(_0073_),
    .Z(_0252_)
  );
  AND2_X1 _0896_ (
    .A1(_0237_),
    .A2(_0252_),
    .ZN(_0253_)
  );
  OR2_X1 _0897_ (
    .A1(_0248_),
    .A2(_0253_),
    .ZN(_0254_)
  );
  AND2_X1 _0898_ (
    .A1(_0241_),
    .A2(_0254_),
    .ZN(_0255_)
  );
  OR2_X1 _0899_ (
    .A1(_0247_),
    .A2(_0255_),
    .ZN(_0256_)
  );
  AND2_X1 _0900_ (
    .A1(io_rvc),
    .A2(_0017_),
    .ZN(_0257_)
  );
  AND2_X1 _0901_ (
    .A1(_0256_),
    .A2(_0257_),
    .ZN(_0258_)
  );
  AND2_X1 _0902_ (
    .A1(io_in[15]),
    .A2(_0028_),
    .ZN(_0259_)
  );
  OR2_X1 _0903_ (
    .A1(_0610_),
    .A2(_0259_),
    .ZN(_0260_)
  );
  INV_X1 _0904_ (
    .A(_0260_),
    .ZN(_0261_)
  );
  OR2_X1 _0905_ (
    .A1(_0230_),
    .A2(_0260_),
    .ZN(_0262_)
  );
  AND2_X1 _0906_ (
    .A1(io_in[9]),
    .A2(_0262_),
    .ZN(_0263_)
  );
  OR2_X1 _0907_ (
    .A1(_0258_),
    .A2(_0263_),
    .ZN(io_out_bits[9])
  );
  AND2_X1 _0908_ (
    .A1(_0067_),
    .A2(_0209_),
    .ZN(_0264_)
  );
  OR2_X1 _0909_ (
    .A1(_0066_),
    .A2(_0210_),
    .ZN(_0265_)
  );
  AND2_X1 _0910_ (
    .A1(_0130_),
    .A2(_0264_),
    .ZN(_0266_)
  );
  AND2_X1 _0911_ (
    .A1(_0176_),
    .A2(_0266_),
    .ZN(_0267_)
  );
  OR2_X1 _0912_ (
    .A1(io_in[10]),
    .A2(_0267_),
    .ZN(_0268_)
  );
  MUX2_X1 _0913_ (
    .A(io_in[10]),
    .B(_0082_),
    .S(_0065_),
    .Z(_0269_)
  );
  AND2_X1 _0914_ (
    .A1(_0110_),
    .A2(_0269_),
    .ZN(_0270_)
  );
  AND2_X1 _0915_ (
    .A1(_0020_),
    .A2(_0270_),
    .ZN(_0271_)
  );
  AND2_X1 _0916_ (
    .A1(io_in[10]),
    .A2(_0230_),
    .ZN(_0272_)
  );
  OR2_X1 _0917_ (
    .A1(_0271_),
    .A2(_0272_),
    .ZN(_0273_)
  );
  AND2_X1 _0918_ (
    .A1(_0268_),
    .A2(_0273_),
    .ZN(io_out_bits[10])
  );
  AND2_X1 _0919_ (
    .A1(_0068_),
    .A2(_0209_),
    .ZN(_0274_)
  );
  INV_X1 _0920_ (
    .A(_0274_),
    .ZN(_0275_)
  );
  OR2_X1 _0921_ (
    .A1(_0177_),
    .A2(_0230_),
    .ZN(_0276_)
  );
  OR2_X1 _0922_ (
    .A1(_0131_),
    .A2(_0276_),
    .ZN(_0277_)
  );
  OR2_X1 _0923_ (
    .A1(_0275_),
    .A2(_0277_),
    .ZN(_0278_)
  );
  AND2_X1 _0924_ (
    .A1(io_in[11]),
    .A2(_0278_),
    .ZN(io_out_bits[11])
  );
  AND2_X1 _0925_ (
    .A1(io_in[6]),
    .A2(io_in[5]),
    .ZN(_0279_)
  );
  OR2_X1 _0926_ (
    .A1(_0147_),
    .A2(_0279_),
    .ZN(_0280_)
  );
  AND2_X1 _0927_ (
    .A1(_0097_),
    .A2(_0280_),
    .ZN(_0281_)
  );
  OR2_X1 _0928_ (
    .A1(_0043_),
    .A2(_0120_),
    .ZN(_0282_)
  );
  AND2_X1 _0929_ (
    .A1(_0094_),
    .A2(_0106_),
    .ZN(_0283_)
  );
  INV_X1 _0930_ (
    .A(_0283_),
    .ZN(_0284_)
  );
  OR2_X1 _0931_ (
    .A1(_0282_),
    .A2(_0284_),
    .ZN(_0285_)
  );
  AND2_X1 _0932_ (
    .A1(io_in[2]),
    .A2(_0077_),
    .ZN(_0286_)
  );
  OR2_X1 _0933_ (
    .A1(_0285_),
    .A2(_0286_),
    .ZN(_0287_)
  );
  AND2_X1 _0934_ (
    .A1(io_in[12]),
    .A2(_0610_),
    .ZN(_0288_)
  );
  AND2_X1 _0935_ (
    .A1(io_in[12]),
    .A2(_0079_),
    .ZN(_0289_)
  );
  OR2_X1 _0936_ (
    .A1(_0281_),
    .A2(_0289_),
    .ZN(_0290_)
  );
  OR2_X1 _0937_ (
    .A1(_0288_),
    .A2(_0290_),
    .ZN(_0291_)
  );
  OR2_X1 _0938_ (
    .A1(_0287_),
    .A2(_0291_),
    .ZN(io_out_bits[12])
  );
  AND2_X1 _0939_ (
    .A1(io_in[3]),
    .A2(_0077_),
    .ZN(_0292_)
  );
  OR2_X1 _0940_ (
    .A1(_0180_),
    .A2(_0289_),
    .ZN(_0293_)
  );
  AND2_X1 _0941_ (
    .A1(io_in[11]),
    .A2(_0604_),
    .ZN(_0294_)
  );
  AND2_X1 _0942_ (
    .A1(io_in[6]),
    .A2(io_in[11]),
    .ZN(_0295_)
  );
  OR2_X1 _0943_ (
    .A1(_0294_),
    .A2(_0295_),
    .ZN(_0296_)
  );
  AND2_X1 _0944_ (
    .A1(_0097_),
    .A2(_0296_),
    .ZN(_0297_)
  );
  OR2_X1 _0945_ (
    .A1(_0605_),
    .A2(io_in[13]),
    .ZN(_0298_)
  );
  AND2_X1 _0946_ (
    .A1(_0166_),
    .A2(_0298_),
    .ZN(_0299_)
  );
  OR2_X1 _0947_ (
    .A1(_0297_),
    .A2(_0299_),
    .ZN(_0300_)
  );
  OR2_X1 _0948_ (
    .A1(_0292_),
    .A2(_0300_),
    .ZN(_0301_)
  );
  OR2_X1 _0949_ (
    .A1(_0293_),
    .A2(_0301_),
    .ZN(io_out_bits[13])
  );
  AND2_X1 _0950_ (
    .A1(io_in[4]),
    .A2(_0077_),
    .ZN(_0302_)
  );
  AND2_X1 _0951_ (
    .A1(_0601_),
    .A2(_0612_),
    .ZN(_0303_)
  );
  OR2_X1 _0952_ (
    .A1(_0147_),
    .A2(_0303_),
    .ZN(_0304_)
  );
  AND2_X1 _0953_ (
    .A1(_0097_),
    .A2(_0304_),
    .ZN(_0305_)
  );
  AND2_X1 _0954_ (
    .A1(io_in[14]),
    .A2(_0610_),
    .ZN(_0306_)
  );
  OR2_X1 _0955_ (
    .A1(_0305_),
    .A2(_0306_),
    .ZN(_0307_)
  );
  OR2_X1 _0956_ (
    .A1(_0289_),
    .A2(_0307_),
    .ZN(_0308_)
  );
  OR2_X1 _0957_ (
    .A1(_0302_),
    .A2(_0308_),
    .ZN(io_out_bits[14])
  );
  AND2_X1 _0958_ (
    .A1(_0133_),
    .A2(_0209_),
    .ZN(_0309_)
  );
  OR2_X1 _0959_ (
    .A1(_0134_),
    .A2(_0210_),
    .ZN(_0310_)
  );
  AND2_X1 _0960_ (
    .A1(io_in[7]),
    .A2(_0310_),
    .ZN(_0311_)
  );
  OR2_X1 _0961_ (
    .A1(io_in[12]),
    .A2(_0617_),
    .ZN(_0312_)
  );
  AND2_X1 _0962_ (
    .A1(io_in[7]),
    .A2(_0019_),
    .ZN(_0313_)
  );
  AND2_X1 _0963_ (
    .A1(_0312_),
    .A2(_0313_),
    .ZN(_0314_)
  );
  OR2_X1 _0964_ (
    .A1(_0173_),
    .A2(_0314_),
    .ZN(_0315_)
  );
  OR2_X1 _0965_ (
    .A1(_0311_),
    .A2(_0315_),
    .ZN(_0316_)
  );
  AND2_X1 _0966_ (
    .A1(io_in[7]),
    .A2(_0103_),
    .ZN(_0317_)
  );
  AND2_X1 _0967_ (
    .A1(io_in[5]),
    .A2(_0077_),
    .ZN(_0318_)
  );
  OR2_X1 _0968_ (
    .A1(_0289_),
    .A2(_0318_),
    .ZN(_0319_)
  );
  OR2_X1 _0969_ (
    .A1(_0317_),
    .A2(_0319_),
    .ZN(_0320_)
  );
  OR2_X1 _0970_ (
    .A1(_0316_),
    .A2(_0320_),
    .ZN(io_out_bits[15])
  );
  AND2_X1 _0971_ (
    .A1(io_in[16]),
    .A2(_0610_),
    .ZN(_0321_)
  );
  AND2_X1 _0972_ (
    .A1(_0019_),
    .A2(_0312_),
    .ZN(_0322_)
  );
  AND2_X1 _0973_ (
    .A1(io_in[8]),
    .A2(_0322_),
    .ZN(_0323_)
  );
  OR2_X1 _0974_ (
    .A1(_0321_),
    .A2(_0323_),
    .ZN(_0324_)
  );
  OR2_X1 _0975_ (
    .A1(io_in[6]),
    .A2(_0007_),
    .ZN(_0325_)
  );
  AND2_X1 _0976_ (
    .A1(_0010_),
    .A2(_0064_),
    .ZN(_0326_)
  );
  AND2_X1 _0977_ (
    .A1(_0325_),
    .A2(_0326_),
    .ZN(_0327_)
  );
  AND2_X1 _0978_ (
    .A1(io_in[8]),
    .A2(_0097_),
    .ZN(_0328_)
  );
  OR2_X1 _0979_ (
    .A1(io_in[8]),
    .A2(_0309_),
    .ZN(_0329_)
  );
  MUX2_X1 _0980_ (
    .A(io_in[12]),
    .B(_0329_),
    .S(_0082_),
    .Z(_0330_)
  );
  AND2_X1 _0981_ (
    .A1(_0213_),
    .A2(_0330_),
    .ZN(_0331_)
  );
  OR2_X1 _0982_ (
    .A1(_0328_),
    .A2(_0331_),
    .ZN(_0332_)
  );
  OR2_X1 _0983_ (
    .A1(_0327_),
    .A2(_0332_),
    .ZN(_0333_)
  );
  OR2_X1 _0984_ (
    .A1(io_in[8]),
    .A2(_0102_),
    .ZN(_0334_)
  );
  OR2_X1 _0985_ (
    .A1(io_in[12]),
    .A2(_0110_),
    .ZN(_0335_)
  );
  AND2_X1 _0986_ (
    .A1(io_rvc),
    .A2(_0020_),
    .ZN(_0336_)
  );
  AND2_X1 _0987_ (
    .A1(_0335_),
    .A2(_0336_),
    .ZN(_0337_)
  );
  AND2_X1 _0988_ (
    .A1(_0334_),
    .A2(_0337_),
    .ZN(_0338_)
  );
  AND2_X1 _0989_ (
    .A1(_0333_),
    .A2(_0338_),
    .ZN(_0339_)
  );
  OR2_X1 _0990_ (
    .A1(_0324_),
    .A2(_0339_),
    .ZN(io_out_bits[16])
  );
  OR2_X1 _0991_ (
    .A1(_0310_),
    .A2(_0322_),
    .ZN(_0340_)
  );
  AND2_X1 _0992_ (
    .A1(io_in[9]),
    .A2(_0340_),
    .ZN(_0341_)
  );
  AND2_X1 _0993_ (
    .A1(io_in[17]),
    .A2(_0610_),
    .ZN(_0342_)
  );
  OR2_X1 _0994_ (
    .A1(_0341_),
    .A2(_0342_),
    .ZN(_0343_)
  );
  AND2_X1 _0995_ (
    .A1(io_in[9]),
    .A2(_0103_),
    .ZN(_0344_)
  );
  AND2_X1 _0996_ (
    .A1(io_in[12]),
    .A2(_0064_),
    .ZN(_0345_)
  );
  OR2_X1 _0997_ (
    .A1(io_in[12]),
    .A2(_0007_),
    .ZN(_0346_)
  );
  AND2_X1 _0998_ (
    .A1(_0064_),
    .A2(_0346_),
    .ZN(_0347_)
  );
  AND2_X1 _0999_ (
    .A1(io_in[12]),
    .A2(_0077_),
    .ZN(_0348_)
  );
  OR2_X1 _1000_ (
    .A1(_0289_),
    .A2(_0348_),
    .ZN(_0349_)
  );
  OR2_X1 _1001_ (
    .A1(_0344_),
    .A2(_0349_),
    .ZN(_0350_)
  );
  OR2_X1 _1002_ (
    .A1(_0343_),
    .A2(_0350_),
    .ZN(io_out_bits[17])
  );
  AND2_X1 _1003_ (
    .A1(io_in[10]),
    .A2(_0086_),
    .ZN(_0351_)
  );
  OR2_X1 _1004_ (
    .A1(_0171_),
    .A2(_0175_),
    .ZN(_0352_)
  );
  AND2_X1 _1005_ (
    .A1(io_in[18]),
    .A2(_0352_),
    .ZN(_0353_)
  );
  OR2_X1 _1006_ (
    .A1(_0351_),
    .A2(_0353_),
    .ZN(_0354_)
  );
  AND2_X1 _1007_ (
    .A1(io_in[10]),
    .A2(_0322_),
    .ZN(_0355_)
  );
  OR2_X1 _1008_ (
    .A1(_0100_),
    .A2(_0355_),
    .ZN(_0356_)
  );
  AND2_X1 _1009_ (
    .A1(io_in[10]),
    .A2(_0072_),
    .ZN(_0357_)
  );
  AND2_X1 _1010_ (
    .A1(io_in[18]),
    .A2(_0172_),
    .ZN(_0358_)
  );
  OR2_X1 _1011_ (
    .A1(_0357_),
    .A2(_0358_),
    .ZN(_0359_)
  );
  OR2_X1 _1012_ (
    .A1(_0293_),
    .A2(_0359_),
    .ZN(_0360_)
  );
  OR2_X1 _1013_ (
    .A1(_0348_),
    .A2(_0360_),
    .ZN(_0361_)
  );
  OR2_X1 _1014_ (
    .A1(_0356_),
    .A2(_0361_),
    .ZN(_0362_)
  );
  OR2_X1 _1015_ (
    .A1(_0354_),
    .A2(_0362_),
    .ZN(io_out_bits[18])
  );
  AND2_X1 _1016_ (
    .A1(io_in[11]),
    .A2(_0072_),
    .ZN(_0363_)
  );
  AND2_X1 _1017_ (
    .A1(io_in[19]),
    .A2(_0172_),
    .ZN(_0364_)
  );
  OR2_X1 _1018_ (
    .A1(_0363_),
    .A2(_0364_),
    .ZN(_0365_)
  );
  AND2_X1 _1019_ (
    .A1(io_in[11]),
    .A2(_0086_),
    .ZN(_0366_)
  );
  AND2_X1 _1020_ (
    .A1(io_in[19]),
    .A2(_0352_),
    .ZN(_0367_)
  );
  OR2_X1 _1021_ (
    .A1(_0366_),
    .A2(_0367_),
    .ZN(_0368_)
  );
  AND2_X1 _1022_ (
    .A1(io_in[11]),
    .A2(_0322_),
    .ZN(_0369_)
  );
  OR2_X1 _1023_ (
    .A1(_0349_),
    .A2(_0369_),
    .ZN(_0370_)
  );
  OR2_X1 _1024_ (
    .A1(_0368_),
    .A2(_0370_),
    .ZN(_0371_)
  );
  OR2_X1 _1025_ (
    .A1(_0365_),
    .A2(_0371_),
    .ZN(io_out_bits[19])
  );
  OR2_X1 _1026_ (
    .A1(_0101_),
    .A2(_0167_),
    .ZN(_0372_)
  );
  OR2_X1 _1027_ (
    .A1(_0265_),
    .A2(_0372_),
    .ZN(_0373_)
  );
  AND2_X1 _1028_ (
    .A1(io_in[2]),
    .A2(_0373_),
    .ZN(_0374_)
  );
  AND2_X1 _1029_ (
    .A1(io_in[12]),
    .A2(_0158_),
    .ZN(_0375_)
  );
  OR2_X1 _1030_ (
    .A1(io_in[2]),
    .A2(_0375_),
    .ZN(_0376_)
  );
  AND2_X1 _1031_ (
    .A1(_0019_),
    .A2(_0376_),
    .ZN(_0377_)
  );
  AND2_X1 _1032_ (
    .A1(io_in[20]),
    .A2(_0610_),
    .ZN(_0378_)
  );
  OR2_X1 _1033_ (
    .A1(_0349_),
    .A2(_0378_),
    .ZN(_0379_)
  );
  OR2_X1 _1034_ (
    .A1(_0377_),
    .A2(_0379_),
    .ZN(_0380_)
  );
  OR2_X1 _1035_ (
    .A1(_0374_),
    .A2(_0380_),
    .ZN(io_out_bits[20])
  );
  OR2_X1 _1036_ (
    .A1(_0081_),
    .A2(_0265_),
    .ZN(_0381_)
  );
  AND2_X1 _1037_ (
    .A1(_0606_),
    .A2(_0090_),
    .ZN(_0382_)
  );
  OR2_X1 _1038_ (
    .A1(_0016_),
    .A2(_0086_),
    .ZN(_0383_)
  );
  OR2_X1 _1039_ (
    .A1(_0382_),
    .A2(_0383_),
    .ZN(_0384_)
  );
  OR2_X1 _1040_ (
    .A1(_0381_),
    .A2(_0384_),
    .ZN(_0385_)
  );
  AND2_X1 _1041_ (
    .A1(io_in[3]),
    .A2(_0385_),
    .ZN(_0386_)
  );
  AND2_X1 _1042_ (
    .A1(io_in[21]),
    .A2(_0610_),
    .ZN(_0387_)
  );
  OR2_X1 _1043_ (
    .A1(_0348_),
    .A2(_0387_),
    .ZN(_0388_)
  );
  OR2_X1 _1044_ (
    .A1(_0386_),
    .A2(_0388_),
    .ZN(io_out_bits[21])
  );
  AND2_X1 _1045_ (
    .A1(_0013_),
    .A2(_0175_),
    .ZN(_0389_)
  );
  OR2_X1 _1046_ (
    .A1(_0173_),
    .A2(_0389_),
    .ZN(_0390_)
  );
  INV_X1 _1047_ (
    .A(_0390_),
    .ZN(_0391_)
  );
  AND2_X1 _1048_ (
    .A1(io_in[22]),
    .A2(_0610_),
    .ZN(_0392_)
  );
  AND2_X1 _1049_ (
    .A1(_0605_),
    .A2(io_in[1]),
    .ZN(_0393_)
  );
  OR2_X1 _1050_ (
    .A1(_0016_),
    .A2(_0029_),
    .ZN(_0394_)
  );
  AND2_X1 _1051_ (
    .A1(io_in[4]),
    .A2(_0394_),
    .ZN(_0395_)
  );
  AND2_X1 _1052_ (
    .A1(io_in[4]),
    .A2(_0086_),
    .ZN(_0396_)
  );
  AND2_X1 _1053_ (
    .A1(io_in[6]),
    .A2(_0044_),
    .ZN(_0397_)
  );
  MUX2_X1 _1054_ (
    .A(_0397_),
    .B(io_in[4]),
    .S(_0381_),
    .Z(_0398_)
  );
  AND2_X1 _1055_ (
    .A1(_0065_),
    .A2(_0398_),
    .ZN(_0399_)
  );
  OR2_X1 _1056_ (
    .A1(_0348_),
    .A2(_0382_),
    .ZN(_0400_)
  );
  OR2_X1 _1057_ (
    .A1(_0399_),
    .A2(_0400_),
    .ZN(_0401_)
  );
  OR2_X1 _1058_ (
    .A1(_0086_),
    .A2(_0090_),
    .ZN(_0402_)
  );
  INV_X1 _1059_ (
    .A(_0402_),
    .ZN(_0403_)
  );
  AND2_X1 _1060_ (
    .A1(io_in[4]),
    .A2(_0102_),
    .ZN(_0404_)
  );
  OR2_X1 _1061_ (
    .A1(_0403_),
    .A2(_0404_),
    .ZN(_0405_)
  );
  AND2_X1 _1062_ (
    .A1(_0401_),
    .A2(_0405_),
    .ZN(_0406_)
  );
  OR2_X1 _1063_ (
    .A1(_0396_),
    .A2(_0406_),
    .ZN(_0407_)
  );
  AND2_X1 _1064_ (
    .A1(_0017_),
    .A2(_0189_),
    .ZN(_0408_)
  );
  AND2_X1 _1065_ (
    .A1(_0407_),
    .A2(_0408_),
    .ZN(_0409_)
  );
  OR2_X1 _1066_ (
    .A1(_0395_),
    .A2(_0409_),
    .ZN(_0410_)
  );
  MUX2_X1 _1067_ (
    .A(io_in[22]),
    .B(_0410_),
    .S(io_rvc),
    .Z(io_out_bits[22])
  );
  AND2_X1 _1068_ (
    .A1(io_rvc),
    .A2(_0095_),
    .ZN(_0411_)
  );
  AND2_X1 _1069_ (
    .A1(_0065_),
    .A2(_0133_),
    .ZN(_0412_)
  );
  AND2_X1 _1070_ (
    .A1(io_in[5]),
    .A2(_0412_),
    .ZN(_0413_)
  );
  OR2_X1 _1071_ (
    .A1(_0098_),
    .A2(_0146_),
    .ZN(_0414_)
  );
  OR2_X1 _1072_ (
    .A1(io_in[10]),
    .A2(_0033_),
    .ZN(_0415_)
  );
  AND2_X1 _1073_ (
    .A1(_0180_),
    .A2(_0415_),
    .ZN(_0416_)
  );
  OR2_X1 _1074_ (
    .A1(_0097_),
    .A2(_0348_),
    .ZN(_0417_)
  );
  OR2_X1 _1075_ (
    .A1(_0416_),
    .A2(_0417_),
    .ZN(_0418_)
  );
  AND2_X1 _1076_ (
    .A1(_0414_),
    .A2(_0418_),
    .ZN(_0419_)
  );
  OR2_X1 _1077_ (
    .A1(_0413_),
    .A2(_0419_),
    .ZN(_0420_)
  );
  AND2_X1 _1078_ (
    .A1(_0411_),
    .A2(_0420_),
    .ZN(_0421_)
  );
  AND2_X1 _1079_ (
    .A1(io_in[23]),
    .A2(_0610_),
    .ZN(_0422_)
  );
  OR2_X1 _1080_ (
    .A1(_0421_),
    .A2(_0422_),
    .ZN(io_out_bits[23])
  );
  AND2_X1 _1081_ (
    .A1(io_in[24]),
    .A2(_0610_),
    .ZN(_0423_)
  );
  AND2_X1 _1082_ (
    .A1(io_in[11]),
    .A2(_0274_),
    .ZN(_0424_)
  );
  OR2_X1 _1083_ (
    .A1(_0348_),
    .A2(_0424_),
    .ZN(_0425_)
  );
  AND2_X1 _1084_ (
    .A1(_0098_),
    .A2(_0425_),
    .ZN(_0426_)
  );
  OR2_X1 _1085_ (
    .A1(_0075_),
    .A2(_0077_),
    .ZN(_0427_)
  );
  INV_X1 _1086_ (
    .A(_0427_),
    .ZN(_0428_)
  );
  OR2_X1 _1087_ (
    .A1(_0097_),
    .A2(_0428_),
    .ZN(_0429_)
  );
  AND2_X1 _1088_ (
    .A1(io_in[6]),
    .A2(_0429_),
    .ZN(_0430_)
  );
  OR2_X1 _1089_ (
    .A1(_0426_),
    .A2(_0430_),
    .ZN(_0431_)
  );
  AND2_X1 _1090_ (
    .A1(_0017_),
    .A2(_0130_),
    .ZN(_0432_)
  );
  AND2_X1 _1091_ (
    .A1(_0149_),
    .A2(_0432_),
    .ZN(_0433_)
  );
  AND2_X1 _1092_ (
    .A1(_0431_),
    .A2(_0433_),
    .ZN(_0434_)
  );
  AND2_X1 _1093_ (
    .A1(io_in[6]),
    .A2(_0393_),
    .ZN(_0435_)
  );
  OR2_X1 _1094_ (
    .A1(_0434_),
    .A2(_0435_),
    .ZN(_0436_)
  );
  OR2_X1 _1095_ (
    .A1(_0423_),
    .A2(_0435_),
    .ZN(io_out_rs2[4])
  );
  MUX2_X1 _1096_ (
    .A(io_in[24]),
    .B(_0436_),
    .S(io_rvc),
    .Z(io_out_bits[24])
  );
  AND2_X1 _1097_ (
    .A1(io_in[25]),
    .A2(_0610_),
    .ZN(_0437_)
  );
  MUX2_X1 _1098_ (
    .A(_0146_),
    .B(_0238_),
    .S(_0098_),
    .Z(_0438_)
  );
  INV_X1 _1099_ (
    .A(_0438_),
    .ZN(_0439_)
  );
  AND2_X1 _1100_ (
    .A1(io_in[12]),
    .A2(_0439_),
    .ZN(_0440_)
  );
  OR2_X1 _1101_ (
    .A1(_0348_),
    .A2(_0440_),
    .ZN(_0441_)
  );
  AND2_X1 _1102_ (
    .A1(_0184_),
    .A2(_0441_),
    .ZN(_0442_)
  );
  OR2_X1 _1103_ (
    .A1(_0081_),
    .A2(_0347_),
    .ZN(_0443_)
  );
  OR2_X1 _1104_ (
    .A1(_0185_),
    .A2(_0443_),
    .ZN(_0444_)
  );
  AND2_X1 _1105_ (
    .A1(io_in[2]),
    .A2(_0444_),
    .ZN(_0445_)
  );
  OR2_X1 _1106_ (
    .A1(_0442_),
    .A2(_0445_),
    .ZN(_0446_)
  );
  AND2_X1 _1107_ (
    .A1(_0336_),
    .A2(_0446_),
    .ZN(_0447_)
  );
  OR2_X1 _1108_ (
    .A1(_0437_),
    .A2(_0447_),
    .ZN(io_out_bits[25])
  );
  AND2_X1 _1109_ (
    .A1(io_in[26]),
    .A2(_0610_),
    .ZN(_0448_)
  );
  AND2_X1 _1110_ (
    .A1(io_in[2]),
    .A2(_0188_),
    .ZN(_0449_)
  );
  AND2_X1 _1111_ (
    .A1(_0133_),
    .A2(_0264_),
    .ZN(_0450_)
  );
  AND2_X1 _1112_ (
    .A1(io_in[7]),
    .A2(_0450_),
    .ZN(_0451_)
  );
  AND2_X1 _1113_ (
    .A1(io_in[12]),
    .A2(_0072_),
    .ZN(_0452_)
  );
  AND2_X1 _1114_ (
    .A1(io_in[12]),
    .A2(_0074_),
    .ZN(_0453_)
  );
  OR2_X1 _1115_ (
    .A1(_0451_),
    .A2(_0453_),
    .ZN(_0454_)
  );
  AND2_X1 _1116_ (
    .A1(_0065_),
    .A2(_0454_),
    .ZN(_0455_)
  );
  OR2_X1 _1117_ (
    .A1(_0064_),
    .A2(_0180_),
    .ZN(_0456_)
  );
  AND2_X1 _1118_ (
    .A1(io_in[5]),
    .A2(_0456_),
    .ZN(_0457_)
  );
  MUX2_X1 _1119_ (
    .A(_0457_),
    .B(io_in[12]),
    .S(_0077_),
    .Z(_0458_)
  );
  OR2_X1 _1120_ (
    .A1(_0455_),
    .A2(_0458_),
    .ZN(_0459_)
  );
  AND2_X1 _1121_ (
    .A1(_0099_),
    .A2(_0459_),
    .ZN(_0460_)
  );
  AND2_X1 _1122_ (
    .A1(io_in[5]),
    .A2(_0096_),
    .ZN(_0461_)
  );
  AND2_X1 _1123_ (
    .A1(io_in[12]),
    .A2(_0294_),
    .ZN(_0462_)
  );
  AND2_X1 _1124_ (
    .A1(_0097_),
    .A2(_0462_),
    .ZN(_0463_)
  );
  OR2_X1 _1125_ (
    .A1(_0461_),
    .A2(_0463_),
    .ZN(_0464_)
  );
  OR2_X1 _1126_ (
    .A1(_0460_),
    .A2(_0464_),
    .ZN(_0465_)
  );
  AND2_X1 _1127_ (
    .A1(_0027_),
    .A2(_0465_),
    .ZN(_0466_)
  );
  OR2_X1 _1128_ (
    .A1(_0449_),
    .A2(_0466_),
    .ZN(_0467_)
  );
  AND2_X1 _1129_ (
    .A1(_0336_),
    .A2(_0467_),
    .ZN(_0468_)
  );
  OR2_X1 _1130_ (
    .A1(_0448_),
    .A2(_0468_),
    .ZN(io_out_bits[26])
  );
  AND2_X1 _1131_ (
    .A1(io_in[27]),
    .A2(_0610_),
    .ZN(_0469_)
  );
  AND2_X1 _1132_ (
    .A1(io_in[3]),
    .A2(_0188_),
    .ZN(_0470_)
  );
  OR2_X1 _1133_ (
    .A1(io_in[3]),
    .A2(_0008_),
    .ZN(_0471_)
  );
  AND2_X1 _1134_ (
    .A1(_0347_),
    .A2(_0471_),
    .ZN(_0472_)
  );
  AND2_X1 _1135_ (
    .A1(io_in[6]),
    .A2(_0139_),
    .ZN(_0473_)
  );
  MUX2_X1 _1136_ (
    .A(io_in[6]),
    .B(io_in[8]),
    .S(_0044_),
    .Z(_0474_)
  );
  AND2_X1 _1137_ (
    .A1(_0056_),
    .A2(_0474_),
    .ZN(_0475_)
  );
  AND2_X1 _1138_ (
    .A1(_0051_),
    .A2(_0475_),
    .ZN(_0476_)
  );
  OR2_X1 _1139_ (
    .A1(_0473_),
    .A2(_0476_),
    .ZN(_0477_)
  );
  AND2_X1 _1140_ (
    .A1(_0142_),
    .A2(_0477_),
    .ZN(_0478_)
  );
  OR2_X1 _1141_ (
    .A1(_0081_),
    .A2(_0452_),
    .ZN(_0479_)
  );
  OR2_X1 _1142_ (
    .A1(_0478_),
    .A2(_0479_),
    .ZN(_0480_)
  );
  OR2_X1 _1143_ (
    .A1(io_in[6]),
    .A2(_0082_),
    .ZN(_0481_)
  );
  AND2_X1 _1144_ (
    .A1(_0480_),
    .A2(_0481_),
    .ZN(_0482_)
  );
  MUX2_X1 _1145_ (
    .A(io_in[12]),
    .B(_0482_),
    .S(_0067_),
    .Z(_0483_)
  );
  AND2_X1 _1146_ (
    .A1(_0065_),
    .A2(_0483_),
    .ZN(_0484_)
  );
  OR2_X1 _1147_ (
    .A1(_0472_),
    .A2(_0484_),
    .ZN(_0485_)
  );
  MUX2_X1 _1148_ (
    .A(_0013_),
    .B(_0485_),
    .S(_0091_),
    .Z(_0486_)
  );
  OR2_X1 _1149_ (
    .A1(_0463_),
    .A2(_0486_),
    .ZN(_0487_)
  );
  OR2_X1 _1150_ (
    .A1(io_in[6]),
    .A2(_0184_),
    .ZN(_0488_)
  );
  AND2_X1 _1151_ (
    .A1(_0027_),
    .A2(_0488_),
    .ZN(_0489_)
  );
  AND2_X1 _1152_ (
    .A1(_0487_),
    .A2(_0489_),
    .ZN(_0490_)
  );
  OR2_X1 _1153_ (
    .A1(_0470_),
    .A2(_0490_),
    .ZN(_0491_)
  );
  AND2_X1 _1154_ (
    .A1(_0336_),
    .A2(_0491_),
    .ZN(_0492_)
  );
  OR2_X1 _1155_ (
    .A1(_0469_),
    .A2(_0492_),
    .ZN(io_out_bits[27])
  );
  AND2_X1 _1156_ (
    .A1(io_in[28]),
    .A2(_0610_),
    .ZN(_0493_)
  );
  AND2_X1 _1157_ (
    .A1(io_in[4]),
    .A2(_0107_),
    .ZN(_0494_)
  );
  AND2_X1 _1158_ (
    .A1(io_in[9]),
    .A2(_0450_),
    .ZN(_0495_)
  );
  OR2_X1 _1159_ (
    .A1(_0453_),
    .A2(_0495_),
    .ZN(_0496_)
  );
  AND2_X1 _1160_ (
    .A1(_0065_),
    .A2(_0496_),
    .ZN(_0497_)
  );
  OR2_X1 _1161_ (
    .A1(io_in[4]),
    .A2(_0008_),
    .ZN(_0498_)
  );
  AND2_X1 _1162_ (
    .A1(_0347_),
    .A2(_0498_),
    .ZN(_0499_)
  );
  OR2_X1 _1163_ (
    .A1(_0497_),
    .A2(_0499_),
    .ZN(_0500_)
  );
  AND2_X1 _1164_ (
    .A1(_0099_),
    .A2(_0500_),
    .ZN(_0501_)
  );
  OR2_X1 _1165_ (
    .A1(_0217_),
    .A2(_0463_),
    .ZN(_0502_)
  );
  OR2_X1 _1166_ (
    .A1(_0501_),
    .A2(_0502_),
    .ZN(_0503_)
  );
  AND2_X1 _1167_ (
    .A1(_0106_),
    .A2(_0503_),
    .ZN(_0504_)
  );
  OR2_X1 _1168_ (
    .A1(_0494_),
    .A2(_0504_),
    .ZN(_0505_)
  );
  AND2_X1 _1169_ (
    .A1(_0031_),
    .A2(_0261_),
    .ZN(_0506_)
  );
  AND2_X1 _1170_ (
    .A1(_0114_),
    .A2(_0506_),
    .ZN(_0507_)
  );
  AND2_X1 _1171_ (
    .A1(_0505_),
    .A2(_0507_),
    .ZN(_0508_)
  );
  OR2_X1 _1172_ (
    .A1(_0493_),
    .A2(_0508_),
    .ZN(io_out_bits[28])
  );
  AND2_X1 _1173_ (
    .A1(io_in[29]),
    .A2(_0610_),
    .ZN(_0509_)
  );
  AND2_X1 _1174_ (
    .A1(io_in[10]),
    .A2(_0450_),
    .ZN(_0510_)
  );
  OR2_X1 _1175_ (
    .A1(_0345_),
    .A2(_0453_),
    .ZN(_0511_)
  );
  OR2_X1 _1176_ (
    .A1(_0463_),
    .A2(_0511_),
    .ZN(_0512_)
  );
  OR2_X1 _1177_ (
    .A1(_0510_),
    .A2(_0512_),
    .ZN(_0513_)
  );
  OR2_X1 _1178_ (
    .A1(_0099_),
    .A2(_0463_),
    .ZN(_0514_)
  );
  OR2_X1 _1179_ (
    .A1(io_in[12]),
    .A2(_0065_),
    .ZN(_0515_)
  );
  AND2_X1 _1180_ (
    .A1(_0514_),
    .A2(_0515_),
    .ZN(_0516_)
  );
  AND2_X1 _1181_ (
    .A1(_0513_),
    .A2(_0516_),
    .ZN(_0517_)
  );
  OR2_X1 _1182_ (
    .A1(_0217_),
    .A2(_0517_),
    .ZN(_0518_)
  );
  AND2_X1 _1183_ (
    .A1(_0608_),
    .A2(_0518_),
    .ZN(_0519_)
  );
  OR2_X1 _1184_ (
    .A1(_0509_),
    .A2(_0519_),
    .ZN(io_out_bits[29])
  );
  AND2_X1 _1185_ (
    .A1(io_in[30]),
    .A2(_0610_),
    .ZN(_0520_)
  );
  OR2_X1 _1186_ (
    .A1(_0217_),
    .A2(_0520_),
    .ZN(_0521_)
  );
  AND2_X1 _1187_ (
    .A1(io_in[11]),
    .A2(_0612_),
    .ZN(_0522_)
  );
  INV_X1 _1188_ (
    .A(_0522_),
    .ZN(_0523_)
  );
  AND2_X1 _1189_ (
    .A1(io_in[10]),
    .A2(_0523_),
    .ZN(_0524_)
  );
  AND2_X1 _1190_ (
    .A1(_0097_),
    .A2(_0524_),
    .ZN(_0525_)
  );
  AND2_X1 _1191_ (
    .A1(io_in[8]),
    .A2(_0079_),
    .ZN(_0526_)
  );
  OR2_X1 _1192_ (
    .A1(_0525_),
    .A2(_0526_),
    .ZN(_0527_)
  );
  OR2_X1 _1193_ (
    .A1(_0521_),
    .A2(_0527_),
    .ZN(_0528_)
  );
  OR2_X1 _1194_ (
    .A1(_0512_),
    .A2(_0528_),
    .ZN(io_out_bits[30])
  );
  AND2_X1 _1195_ (
    .A1(io_in[31]),
    .A2(_0610_),
    .ZN(_0529_)
  );
  OR2_X1 _1196_ (
    .A1(_0289_),
    .A2(_0529_),
    .ZN(_0530_)
  );
  OR2_X1 _1197_ (
    .A1(_0502_),
    .A2(_0530_),
    .ZN(_0531_)
  );
  OR2_X1 _1198_ (
    .A1(_0511_),
    .A2(_0531_),
    .ZN(io_out_bits[31])
  );
  OR2_X1 _1199_ (
    .A1(io_in[7]),
    .A2(_0176_),
    .ZN(_0532_)
  );
  AND2_X1 _1200_ (
    .A1(io_in[7]),
    .A2(_0093_),
    .ZN(_0533_)
  );
  AND2_X1 _1201_ (
    .A1(io_in[2]),
    .A2(_0073_),
    .ZN(_0534_)
  );
  OR2_X1 _1202_ (
    .A1(_0208_),
    .A2(_0534_),
    .ZN(_0535_)
  );
  MUX2_X1 _1203_ (
    .A(io_in[7]),
    .B(_0535_),
    .S(_0213_),
    .Z(_0536_)
  );
  AND2_X1 _1204_ (
    .A1(_0183_),
    .A2(_0536_),
    .ZN(_0537_)
  );
  OR2_X1 _1205_ (
    .A1(_0533_),
    .A2(_0537_),
    .ZN(_0538_)
  );
  AND2_X1 _1206_ (
    .A1(_0129_),
    .A2(_0538_),
    .ZN(_0539_)
  );
  OR2_X1 _1207_ (
    .A1(_0220_),
    .A2(_0539_),
    .ZN(_0540_)
  );
  AND2_X1 _1208_ (
    .A1(_0020_),
    .A2(_0540_),
    .ZN(_0541_)
  );
  OR2_X1 _1209_ (
    .A1(_0202_),
    .A2(_0313_),
    .ZN(_0542_)
  );
  AND2_X1 _1210_ (
    .A1(_0002_),
    .A2(_0542_),
    .ZN(_0543_)
  );
  OR2_X1 _1211_ (
    .A1(_0177_),
    .A2(_0543_),
    .ZN(_0544_)
  );
  OR2_X1 _1212_ (
    .A1(_0541_),
    .A2(_0544_),
    .ZN(_0545_)
  );
  AND2_X1 _1213_ (
    .A1(_0532_),
    .A2(_0545_),
    .ZN(io_out_rd[0])
  );
  AND2_X1 _1214_ (
    .A1(io_in[8]),
    .A2(_0276_),
    .ZN(_0546_)
  );
  AND2_X1 _1215_ (
    .A1(io_in[8]),
    .A2(_0093_),
    .ZN(_0547_)
  );
  MUX2_X1 _1216_ (
    .A(io_in[8]),
    .B(io_in[3]),
    .S(_0073_),
    .Z(_0548_)
  );
  AND2_X1 _1217_ (
    .A1(_0237_),
    .A2(_0548_),
    .ZN(_0549_)
  );
  OR2_X1 _1218_ (
    .A1(_0233_),
    .A2(_0549_),
    .ZN(_0550_)
  );
  AND2_X1 _1219_ (
    .A1(_0183_),
    .A2(_0550_),
    .ZN(_0551_)
  );
  OR2_X1 _1220_ (
    .A1(_0547_),
    .A2(_0551_),
    .ZN(_0552_)
  );
  AND2_X1 _1221_ (
    .A1(_0129_),
    .A2(_0552_),
    .ZN(_0553_)
  );
  OR2_X1 _1222_ (
    .A1(_0232_),
    .A2(_0553_),
    .ZN(_0554_)
  );
  AND2_X1 _1223_ (
    .A1(_0257_),
    .A2(_0554_),
    .ZN(_0555_)
  );
  OR2_X1 _1224_ (
    .A1(_0546_),
    .A2(_0555_),
    .ZN(io_out_rd[1])
  );
  AND2_X1 _1225_ (
    .A1(io_in[9]),
    .A2(_0276_),
    .ZN(_0556_)
  );
  AND2_X1 _1226_ (
    .A1(io_in[9]),
    .A2(_0093_),
    .ZN(_0557_)
  );
  MUX2_X1 _1227_ (
    .A(io_in[9]),
    .B(io_in[4]),
    .S(_0073_),
    .Z(_0558_)
  );
  AND2_X1 _1228_ (
    .A1(_0237_),
    .A2(_0558_),
    .ZN(_0559_)
  );
  OR2_X1 _1229_ (
    .A1(_0248_),
    .A2(_0559_),
    .ZN(_0560_)
  );
  AND2_X1 _1230_ (
    .A1(_0183_),
    .A2(_0560_),
    .ZN(_0561_)
  );
  OR2_X1 _1231_ (
    .A1(_0557_),
    .A2(_0561_),
    .ZN(_0562_)
  );
  AND2_X1 _1232_ (
    .A1(_0129_),
    .A2(_0562_),
    .ZN(_0563_)
  );
  OR2_X1 _1233_ (
    .A1(_0247_),
    .A2(_0563_),
    .ZN(_0564_)
  );
  AND2_X1 _1234_ (
    .A1(_0257_),
    .A2(_0564_),
    .ZN(_0565_)
  );
  OR2_X1 _1235_ (
    .A1(_0556_),
    .A2(_0565_),
    .ZN(io_out_rd[2])
  );
  AND2_X1 _1236_ (
    .A1(_0080_),
    .A2(_0094_),
    .ZN(_0566_)
  );
  AND2_X1 _1237_ (
    .A1(_0020_),
    .A2(_0566_),
    .ZN(_0567_)
  );
  OR2_X1 _1238_ (
    .A1(_0272_),
    .A2(_0567_),
    .ZN(_0568_)
  );
  OR2_X1 _1239_ (
    .A1(_0026_),
    .A2(_0072_),
    .ZN(_0569_)
  );
  AND2_X1 _1240_ (
    .A1(_0027_),
    .A2(_0075_),
    .ZN(_0570_)
  );
  OR2_X1 _1241_ (
    .A1(_0069_),
    .A2(_0569_),
    .ZN(_0571_)
  );
  AND2_X1 _1242_ (
    .A1(_0176_),
    .A2(_0570_),
    .ZN(_0572_)
  );
  OR2_X1 _1243_ (
    .A1(io_in[10]),
    .A2(_0572_),
    .ZN(_0573_)
  );
  AND2_X1 _1244_ (
    .A1(_0568_),
    .A2(_0573_),
    .ZN(io_out_rd[3])
  );
  OR2_X1 _1245_ (
    .A1(_0276_),
    .A2(_0571_),
    .ZN(_0574_)
  );
  AND2_X1 _1246_ (
    .A1(io_in[11]),
    .A2(_0574_),
    .ZN(io_out_rd[4])
  );
  OR2_X1 _1247_ (
    .A1(_0064_),
    .A2(_0402_),
    .ZN(_0575_)
  );
  OR2_X1 _1248_ (
    .A1(_0238_),
    .A2(_0402_),
    .ZN(_0576_)
  );
  AND2_X1 _1249_ (
    .A1(io_in[7]),
    .A2(_0576_),
    .ZN(_0577_)
  );
  OR2_X1 _1250_ (
    .A1(_0316_),
    .A2(_0577_),
    .ZN(io_out_rs1[0])
  );
  MUX2_X1 _1251_ (
    .A(io_in[8]),
    .B(_0329_),
    .S(_0082_),
    .Z(_0578_)
  );
  AND2_X1 _1252_ (
    .A1(io_in[8]),
    .A2(_0575_),
    .ZN(_0579_)
  );
  AND2_X1 _1253_ (
    .A1(_0068_),
    .A2(_0403_),
    .ZN(_0580_)
  );
  OR2_X1 _1254_ (
    .A1(_0579_),
    .A2(_0580_),
    .ZN(_0581_)
  );
  AND2_X1 _1255_ (
    .A1(_0578_),
    .A2(_0581_),
    .ZN(_0582_)
  );
  AND2_X1 _1256_ (
    .A1(_0336_),
    .A2(_0582_),
    .ZN(_0583_)
  );
  OR2_X1 _1257_ (
    .A1(_0324_),
    .A2(_0583_),
    .ZN(io_out_rs1[1])
  );
  AND2_X1 _1258_ (
    .A1(io_in[9]),
    .A2(_0576_),
    .ZN(_0584_)
  );
  OR2_X1 _1259_ (
    .A1(_0343_),
    .A2(_0584_),
    .ZN(io_out_rs1[2])
  );
  AND2_X1 _1260_ (
    .A1(io_in[10]),
    .A2(_0238_),
    .ZN(_0585_)
  );
  OR2_X1 _1261_ (
    .A1(_0109_),
    .A2(_0180_),
    .ZN(_0586_)
  );
  OR2_X1 _1262_ (
    .A1(_0359_),
    .A2(_0586_),
    .ZN(_0587_)
  );
  OR2_X1 _1263_ (
    .A1(_0585_),
    .A2(_0587_),
    .ZN(_0588_)
  );
  OR2_X1 _1264_ (
    .A1(_0356_),
    .A2(_0588_),
    .ZN(_0589_)
  );
  OR2_X1 _1265_ (
    .A1(_0354_),
    .A2(_0589_),
    .ZN(io_out_rs1[3])
  );
  OR2_X1 _1266_ (
    .A1(_0365_),
    .A2(_0368_),
    .ZN(_0590_)
  );
  AND2_X1 _1267_ (
    .A1(io_in[11]),
    .A2(_0238_),
    .ZN(_0591_)
  );
  OR2_X1 _1268_ (
    .A1(_0369_),
    .A2(_0591_),
    .ZN(_0592_)
  );
  OR2_X1 _1269_ (
    .A1(_0590_),
    .A2(_0592_),
    .ZN(io_out_rs1[4])
  );
  AND2_X1 _1270_ (
    .A1(io_in[2]),
    .A2(_0411_),
    .ZN(_0593_)
  );
  OR2_X1 _1271_ (
    .A1(_0378_),
    .A2(_0593_),
    .ZN(io_out_rs2[0])
  );
  AND2_X1 _1272_ (
    .A1(io_in[3]),
    .A2(_0411_),
    .ZN(_0594_)
  );
  OR2_X1 _1273_ (
    .A1(_0387_),
    .A2(_0594_),
    .ZN(io_out_rs2[1])
  );
  OR2_X1 _1274_ (
    .A1(io_in[22]),
    .A2(_0391_),
    .ZN(_0595_)
  );
  OR2_X1 _1275_ (
    .A1(_0096_),
    .A2(_0174_),
    .ZN(_0596_)
  );
  INV_X1 _1276_ (
    .A(_0596_),
    .ZN(_0597_)
  );
  AND2_X1 _1277_ (
    .A1(io_in[4]),
    .A2(_0597_),
    .ZN(_0598_)
  );
  AND2_X1 _1278_ (
    .A1(_0595_),
    .A2(_0598_),
    .ZN(_0599_)
  );
  OR2_X1 _1279_ (
    .A1(_0392_),
    .A2(_0599_),
    .ZN(io_out_rs2[2])
  );
  MUX2_X1 _1280_ (
    .A(_0095_),
    .B(io_in[5]),
    .S(_0393_),
    .Z(_0600_)
  );
  MUX2_X1 _1281_ (
    .A(io_in[23]),
    .B(_0600_),
    .S(io_rvc),
    .Z(io_out_rs2[3])
  );
  assign _GEN_0 = { 5'h00, io_in[12], io_in[6:2], 2'h1, io_in[9:7], 5'h15, io_in[9:7], 7'h13 };
  assign { _GEN_1[30:15], _GEN_1[11:0] } = { 8'h01, io_in[4:2], 2'h1, io_in[9:7], 2'h1, io_in[9:7], 3'h3, io_in[12], 3'h3 };
  assign { _io_out_T_10_bits[31:30], _io_out_T_10_bits[25], _io_out_T_10_bits[19], _io_out_T_10_bits[14:13], _io_out_T_10_bits[6], _io_out_T_10_bits[1:0] } = { 2'h0, io_in[12], 2'h0, _io_out_T_10_bits[18], 3'h3 };
  assign _io_out_T_10_rd = { 2'h1, io_in[4:2] };
  assign _io_out_T_10_rs1 = { 1'h0, _io_out_T_10_bits[18:15] };
  assign { _io_out_T_12_bits[31:30], _io_out_T_12_bits[25], _io_out_T_12_bits[19], _io_out_T_12_bits[14:13], _io_out_T_12_bits[6], _io_out_T_12_bits[1:0] } = { 2'h0, io_in[12], 2'h0, _io_out_T_12_bits[18], 3'h3 };
  assign _io_out_T_12_rd = { 2'h1, io_in[4:2] };
  assign _io_out_T_12_rs1 = { 1'h0, _io_out_T_12_bits[18:15] };
  assign { _io_out_T_14_bits[31:30], _io_out_T_14_bits[25], _io_out_T_14_bits[19], _io_out_T_14_bits[14:13], _io_out_T_14_bits[6], _io_out_T_14_bits[1:0] } = { 2'h0, io_in[12], 2'h0, _io_out_T_14_bits[18], 3'h3 };
  assign _io_out_T_14_rd = { 2'h1, io_in[4:2] };
  assign _io_out_T_14_rs1 = { 1'h0, _io_out_T_14_bits[18:15] };
  assign { _io_out_T_16_bits[31:30], _io_out_T_16_bits[25], _io_out_T_16_bits[19], _io_out_T_16_bits[14:13], _io_out_T_16_bits[6], _io_out_T_16_bits[1:0] } = { 2'h0, io_in[12], 2'h0, _io_out_T_16_bits[18], 3'h3 };
  assign _io_out_T_16_rd = { 2'h1, io_in[4:2] };
  assign _io_out_T_16_rs1 = { 1'h0, _io_out_T_16_bits[18:15] };
  assign { _io_out_T_18_bits[30], _io_out_T_18_bits[25], _io_out_T_18_bits[14], _io_out_T_18_bits[6], _io_out_T_18_bits[1:0] } = { _io_out_T_18_bits[31], io_in[12], 4'h3 };
  assign _io_out_T_18_rd[4] = _io_out_T_18_bits[19];
  assign _io_out_T_18_rs1 = _io_out_T_18_bits[19:15];
  assign _io_out_T_18_rs2 = { 2'h1, io_in[4:2] };
  assign _io_out_T_2 = { io_in[1:0], io_in[15:13] };
  assign _io_out_T_20_bits[1:0] = 2'h3;
  assign _io_out_T_20_rs2 = { 2'h1, io_in[4:2] };
  assign _io_out_T_22_bits[1:0] = 2'h3;
  assign _io_out_T_22_rs2 = { 2'h1, io_in[4:2] };
  assign _io_out_T_24_bits[1:0] = 2'h3;
  assign _io_out_T_24_rs2 = { 2'h1, io_in[4:2] };
  assign _io_out_T_26_bits[1:0] = 2'h3;
  assign _io_out_T_26_rs2 = { 2'h1, io_in[4:2] };
  assign _io_out_T_28_bits[1:0] = 2'h3;
  assign _io_out_T_28_rs2 = { 2'h1, io_in[4:2] };
  assign _io_out_T_30_bits[1:0] = 2'h3;
  assign _io_out_T_30_rs2[4] = 1'h0;
  assign _io_out_T_32_bits[1:0] = 2'h3;
  assign _io_out_T_32_rs2[4] = 1'h0;
  assign _io_out_T_34_bits[1:0] = 2'h3;
  assign _io_out_T_36_bits[1:0] = 2'h3;
  assign _io_out_T_38_bits[1:0] = 2'h3;
  assign _io_out_T_40_bits[1:0] = 2'h3;
  assign _io_out_T_42_bits[1:0] = 2'h3;
  assign _io_out_T_44_bits[1:0] = 2'h3;
  assign _io_out_T_46_bits[1:0] = 2'h3;
  assign _io_out_T_48_bits[1:0] = 2'h3;
  assign { _io_out_T_4_bits[31:30], _io_out_T_4_bits[25:24], _io_out_T_4_bits[21:19], _io_out_T_4_bits[14:5], _io_out_T_4_bits[1:0] } = { 2'h0, io_in[12:11], 4'h0, _io_out_T_4_bits[18], _io_out_T_4_bits[18], 2'h1, io_in[4:2], 4'h3 };
  assign _io_out_T_4_rd = { 2'h1, io_in[4:2] };
  assign _io_out_T_4_rs1 = { 1'h0, _io_out_T_4_bits[18:15] };
  assign { _io_out_T_6_bits[31:30], _io_out_T_6_bits[25:24], _io_out_T_6_bits[21:19], _io_out_T_6_bits[14:13], _io_out_T_6_bits[11:5], _io_out_T_6_bits[1:0] } = { 2'h0, io_in[12:11], 4'h0, _io_out_T_6_bits[18], 2'h1, io_in[4:2], 4'h3 };
  assign _io_out_T_6_rd = { 2'h1, io_in[4:2] };
  assign _io_out_T_6_rs1 = { 1'h0, _io_out_T_6_bits[18:15] };
  assign { _io_out_T_8_bits[31:30], _io_out_T_8_bits[25:24], _io_out_T_8_bits[21:19], _io_out_T_8_bits[14:13], _io_out_T_8_bits[11:5], _io_out_T_8_bits[1:0] } = { 2'h0, io_in[12:11], 4'h0, _io_out_T_8_bits[18], 2'h1, io_in[4:2], 4'h3 };
  assign _io_out_T_8_rd = { 2'h1, io_in[4:2] };
  assign _io_out_T_8_rs1 = { 1'h0, _io_out_T_8_bits[18:15] };
  assign _io_out_s_T_116 = { io_in[5], io_in[12], 2'h1, io_in[4:2], 2'h1, io_in[9:7], 3'h2, io_in[11:10], io_in[6], 9'h023 };
  assign _io_out_s_T_138 = { io_in[5], io_in[12], 2'h1, io_in[4:2], 2'h1, io_in[9:7], 3'h2, io_in[11:10], io_in[6], 9'h027 };
  assign _io_out_s_T_148 = { io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12] };
  assign _io_out_s_T_15 = { io_in[6:5], io_in[12:10], 3'h0 };
  assign _io_out_s_T_150 = { io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[6:2] };
  assign _io_out_s_T_161 = { io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12] };
  assign _io_out_s_T_169 = { io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[8], io_in[10:9], io_in[6], io_in[7], io_in[2], io_in[11], io_in[5:3], 1'h0 };
  assign _io_out_s_T_17 = { 2'h1, io_in[9:7] };
  assign _io_out_s_T_20 = { io_in[6:5], io_in[12:10], 5'h01, io_in[9:7], 5'h0d, io_in[4:2], 7'h07 };
  assign _io_out_s_T_230 = { io_in[12], io_in[12], io_in[12] };
  assign _io_out_s_T_251 = { io_in[12], io_in[6:2], 2'h1, io_in[9:7], 5'h15, io_in[9:7], 7'h13 };
  assign _io_out_s_T_260 = { 5'h10, io_in[12], io_in[6:2], 2'h1, io_in[9:7], 5'h15, io_in[9:7], 7'h13 };
  assign _io_out_s_T_270 = { io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[6:2], 2'h1, io_in[9:7], 5'h1d, io_in[9:7], 7'h13 };
  assign _io_out_s_T_277 = { 2'h1, io_in[4:2], 2'h1, io_in[9:7], _GEN_1[14:12], 2'h1, io_in[9:7], 3'h3, io_in[12], 3'h3 };
  assign _io_out_s_T_278[29:0] = { 7'h01, io_in[4:2], 2'h1, io_in[9:7], _GEN_1[14:12], 2'h1, io_in[9:7], 3'h3, io_in[12], 3'h3 };
  assign _io_out_s_T_281[29:0] = { 4'h0, io_in[12], io_in[6:2], 2'h1, io_in[9:7], 5'h15, io_in[9:7], 7'h13 };
  assign { _io_out_s_T_283[29:14], _io_out_s_T_283[12:0] } = { _io_out_s_T_283[31], _io_out_s_T_283[31], _io_out_s_T_283[31], _io_out_s_T_283[31], io_in[12], io_in[6:2], 2'h1, io_in[9:7], 4'hd, io_in[9:7], 7'h13 };
  assign _io_out_s_T_31 = { io_in[5], io_in[12:10], io_in[6], 2'h0 };
  assign _io_out_s_T_349 = { io_in[12], io_in[12], io_in[12], io_in[12], io_in[12] };
  assign _io_out_s_T_354 = { io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[6:5], io_in[2], io_in[11:10], io_in[4:3], 1'h0 };
  assign _io_out_s_T_36 = { io_in[5], io_in[12:10], io_in[6], 4'h1, io_in[9:7], 5'h09, io_in[4:2], 7'h03 };
  assign _io_out_s_T_438 = { io_in[12], io_in[6:2], io_in[11:7], 3'h1, io_in[11:7], 7'h13 };
  assign _io_out_s_T_448 = { io_in[4:2], io_in[12], io_in[6:5], 11'h013, io_in[11:7], 7'h07 };
  assign { _io_out_s_T_457[27:5], _io_out_s_T_457[3:0] } = { io_in[3:2], io_in[12], io_in[6:4], 10'h012, io_in[11:7], 2'h0, _io_out_s_T_457[4], _io_out_s_T_457[4], 2'h3 };
  assign _io_out_s_T_466 = { io_in[3:2], io_in[12], io_in[6:4], 10'h012, io_in[11:7], 7'h07 };
  assign _io_out_s_T_473 = { io_in[9:7], io_in[12:10], 3'h0 };
  assign _io_out_s_T_480 = { io_in[9:7], io_in[12], io_in[6:2], 8'h13, io_in[11:10], 10'h027 };
  assign _io_out_s_T_486 = { io_in[8:7], io_in[12:9], 2'h0 };
  assign _io_out_s_T_493 = { io_in[8:7], io_in[12], io_in[6:2], 8'h12, io_in[11:9], 9'h023 };
  assign _io_out_s_T_506 = { io_in[8:7], io_in[12], io_in[6:2], 8'h12, io_in[11:9], 9'h027 };
  assign _io_out_s_T_52 = { io_in[5], io_in[12:10], io_in[6], 4'h1, io_in[9:7], 5'h09, io_in[4:2], 7'h07 };
  assign _io_out_s_T_6 = { 2'h1, io_in[4:2] };
  assign { _io_out_s_T_7[29:4], _io_out_s_T_7[2:0] } = { io_in[10:7], io_in[12:11], io_in[5], io_in[6], 12'h041, io_in[4:2], 3'h1, _io_out_s_T_7[3], 2'h3 };
  assign _io_out_s_T_74 = { io_in[5], io_in[12], 2'h1, io_in[4:2], 2'h1, io_in[9:7], 3'h2, io_in[11:10], io_in[6], 9'h03f };
  assign _io_out_s_T_94 = { io_in[6:5], io_in[12], 2'h1, io_in[4:2], 2'h1, io_in[9:7], 3'h3, io_in[11:10], 10'h027 };
  assign _io_out_s_add_T_3 = { io_in[6:2], io_in[11:7], 3'h0, io_in[11:7], 7'h33 };
  assign _io_out_s_ebreak_T_1 = { io_in[6:2], io_in[11:7], 15'h0073 };
  assign _io_out_s_funct_T_2 = { io_in[12], io_in[6:5] };
  assign _io_out_s_funct_T_4[1:0] = 2'h0;
  assign _io_out_s_funct_T_6[0] = 1'h0;
  assign { _io_out_s_jalr_ebreak_T_2[24:21], _io_out_s_jalr_ebreak_T_2[19:8], _io_out_s_jalr_ebreak_T_2[6:0] } = { io_in[6:3], io_in[11:7], 9'h003, _io_out_s_T_457[4], 1'h0, _io_out_s_jalr_ebreak_T_2[7], 2'h3 };
  assign _io_out_s_jr_reserved_T_2 = { io_in[6:2], io_in[11:7], 8'h00, _io_out_s_jalr_ebreak_T_2[7], _io_out_s_jalr_ebreak_T_2[7], _io_out_s_T_457[4], _io_out_s_T_457[4], 3'h7 };
  assign _io_out_s_load_opc_T_1 = _io_out_s_jalr_ebreak_T_2[7];
  assign _io_out_s_me_T_2 = { io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12] };
  assign _io_out_s_me_T_4 = { io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[6:2], 12'h000 };
  assign _io_out_s_mv_T_2 = { io_in[6:2], 8'h00, io_in[11:7], 7'h33 };
  assign io_out_bits[1:0] = 2'h3;
  assign io_out_s_0_bits = { 2'h0, io_in[10:7], io_in[12:11], io_in[5], io_in[6], 12'h041, io_in[4:2], 3'h1, _io_out_s_T_7[3], _io_out_s_T_7[3], 2'h3 };
  assign io_out_s_10_bits = { io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[6:2], 8'h00, io_in[11:7], 7'h13 };
  assign { io_out_s_11_bits[31:29], io_out_s_11_bits[22:20], io_out_s_11_bits[11:6], io_out_s_11_bits[4], io_out_s_11_bits[1:0] } = { io_in[12], io_in[12], io_in[12], io_out_s_11_bits[23], io_out_s_11_bits[23], io_out_s_11_bits[23], io_in[11:7], 4'h7 };
  assign io_out_s_11_rd = io_in[11:7];
  assign io_out_s_11_rs2 = { 2'h1, io_in[4:2] };
  assign { io_out_s_12_bits[29:26], io_out_s_12_bits[22:15], io_out_s_12_bits[11:6], io_out_s_12_bits[4], io_out_s_12_bits[2:0] } = { io_out_s_12_bits[31], io_out_s_12_bits[31], io_out_s_12_bits[31], io_out_s_12_bits[31], io_in[4:2], 2'h1, io_in[9:7], 2'h1, io_in[9:7], 5'h0b };
  assign io_out_s_13_bits = { io_in[12], io_in[8], io_in[10:9], io_in[6], io_in[7], io_in[2], io_in[11], io_in[5:3], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], 12'h06f };
  assign io_out_s_14_bits = { io_in[12], io_in[12], io_in[12], io_in[12], io_in[6:5], io_in[2], 7'h01, io_in[9:7], 3'h0, io_in[11:10], io_in[4:3], io_in[12], 7'h63 };
  assign io_out_s_15_bits = { io_in[12], io_in[12], io_in[12], io_in[12], io_in[6:5], io_in[2], 7'h01, io_in[9:7], 3'h1, io_in[11:10], io_in[4:3], io_in[12], 7'h63 };
  assign io_out_s_16_bits = { 6'h00, io_in[12], io_in[6:2], io_in[11:7], 3'h1, io_in[11:7], 7'h13 };
  assign io_out_s_17_bits = { 3'h0, io_in[4:2], io_in[12], io_in[6:5], 11'h013, io_in[11:7], 7'h07 };
  assign io_out_s_18_bits = { 4'h0, io_in[3:2], io_in[12], io_in[6:4], 10'h012, io_in[11:7], 2'h0, _io_out_s_T_457[4], _io_out_s_T_457[4], _io_out_s_T_457[4], 2'h3 };
  assign io_out_s_19_bits = { 4'h0, io_in[3:2], io_in[12], io_in[6:4], 10'h012, io_in[11:7], 7'h07 };
  assign io_out_s_1_bits = { 4'h0, io_in[6:5], io_in[12:10], 5'h01, io_in[9:7], 5'h0d, io_in[4:2], 7'h07 };
  assign { io_out_s_20_bits[31:21], io_out_s_20_bits[14:12], io_out_s_20_bits[1:0] } = { 7'h00, io_in[6:3], 5'h03 };
  assign io_out_s_20_rd[4:1] = io_out_s_20_bits[11:8];
  assign io_out_s_20_rs1 = io_out_s_20_bits[19:15];
  assign io_out_s_20_rs2 = io_in[6:2];
  assign io_out_s_21_bits = { 3'h0, io_in[9:7], io_in[12], io_in[6:2], 8'h13, io_in[11:10], 10'h027 };
  assign io_out_s_22_bits = { 4'h0, io_in[8:7], io_in[12], io_in[6:2], 8'h12, io_in[11:9], 9'h023 };
  assign io_out_s_23_bits = { 4'h0, io_in[8:7], io_in[12], io_in[6:2], 8'h12, io_in[11:9], 9'h027 };
  assign io_out_s_24_rs1 = io_in[19:15];
  assign io_out_s_24_rs2 = io_in[24:20];
  assign io_out_s_2_bits = { 5'h00, io_in[5], io_in[12:10], io_in[6], 4'h1, io_in[9:7], 5'h09, io_in[4:2], 7'h03 };
  assign io_out_s_3_bits = { 5'h00, io_in[5], io_in[12:10], io_in[6], 4'h1, io_in[9:7], 5'h09, io_in[4:2], 7'h07 };
  assign io_out_s_4_bits = { 5'h00, io_in[5], io_in[12], 2'h1, io_in[4:2], 2'h1, io_in[9:7], 3'h2, io_in[11:10], io_in[6], 9'h03f };
  assign io_out_s_5_bits = { 4'h0, io_in[6:5], io_in[12], 2'h1, io_in[4:2], 2'h1, io_in[9:7], 3'h3, io_in[11:10], 10'h027 };
  assign io_out_s_6_bits = { 5'h00, io_in[5], io_in[12], 2'h1, io_in[4:2], 2'h1, io_in[9:7], 3'h2, io_in[11:10], io_in[6], 9'h023 };
  assign io_out_s_7_bits = { 5'h00, io_in[5], io_in[12], 2'h1, io_in[4:2], 2'h1, io_in[9:7], 3'h2, io_in[11:10], io_in[6], 9'h027 };
  assign io_out_s_8_bits = { io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[6:2], io_in[11:7], 3'h0, io_in[11:7], 7'h13 };
  assign io_out_s_9_bits = { io_in[12], io_in[8], io_in[10:9], io_in[6], io_in[7], io_in[2], io_in[11], io_in[5:3], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], 12'h0ef };
  assign io_out_s_add_bits = { 7'h00, io_in[6:2], io_in[11:7], 3'h0, io_in[11:7], 7'h33 };
  assign io_out_s_ebreak = { io_in[6:3], 1'h1, io_in[11:7], 15'h0073 };
  assign io_out_s_funct = _GEN_1[14:12];
  assign io_out_s_jalr = { io_in[6:2], io_in[11:7], 15'h00e7 };
  assign { io_out_s_jalr_add_bits[31:21], io_out_s_jalr_add_bits[19:8], io_out_s_jalr_add_bits[5:3], io_out_s_jalr_add_bits[1:0] } = { 7'h00, io_in[6:3], io_in[11:7], 3'h0, io_out_s_20_bits[11:8], 1'h1, io_out_s_20_bits[4], 3'h3 };
  assign io_out_s_jalr_add_rd[4:1] = io_out_s_20_bits[11:8];
  assign io_out_s_jalr_add_rs1 = io_in[11:7];
  assign io_out_s_jalr_ebreak_bits = { 7'h00, io_in[6:3], _io_out_s_jalr_ebreak_T_2[20], io_in[11:7], 7'h00, _io_out_s_jalr_ebreak_T_2[7], 2'h3, _io_out_s_T_457[4], 1'h0, _io_out_s_jalr_ebreak_T_2[7], 2'h3 };
  assign io_out_s_jr = { io_in[6:2], io_in[11:7], 15'h0067 };
  assign { io_out_s_jr_mv_bits[31:20], io_out_s_jr_mv_bits[14:8], io_out_s_jr_mv_bits[6], io_out_s_jr_mv_bits[4], io_out_s_jr_mv_bits[2:0] } = { 7'h00, io_in[6:2], 3'h0, io_out_s_20_bits[11:8], io_out_s_jalr_add_bits[2], io_out_s_20_bits[4], io_out_s_jalr_add_bits[6], 2'h3 };
  assign io_out_s_jr_mv_rd = { io_out_s_20_bits[11:8], io_out_s_jr_mv_bits[7] };
  assign io_out_s_jr_mv_rs1 = io_out_s_jr_mv_bits[19:15];
  assign io_out_s_jr_mv_rs2 = io_in[6:2];
  assign io_out_s_jr_reserved_bits = { 7'h00, io_in[6:2], io_in[11:7], 8'h00, _io_out_s_jalr_ebreak_T_2[7], _io_out_s_jalr_ebreak_T_2[7], _io_out_s_T_457[4], _io_out_s_T_457[4], 3'h7 };
  assign io_out_s_load_opc = { 2'h0, _io_out_s_T_457[4], _io_out_s_T_457[4], _io_out_s_T_457[4], 2'h3 };
  assign io_out_s_me_bits = { io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[12], io_in[6:2], io_in[11:7], 3'h3, io_out_s_11_bits[3], 3'h7 };
  assign io_out_s_mv_bits = { 7'h00, io_in[6:2], 8'h00, io_in[11:7], 7'h33 };
  assign io_out_s_opc = { 3'h1, _io_out_s_T_7[3], _io_out_s_T_7[3], 2'h3 };
  assign io_out_s_opc_1 = { 3'h3, io_out_s_11_bits[3], 3'h7 };
  assign io_out_s_opc_2 = { 3'h1, io_out_s_11_bits[3], io_out_s_11_bits[3], 2'h3 };
  assign io_out_s_opc_3 = { 3'h3, io_in[12], 3'h3 };
  assign io_out_s_res_bits = { io_in[12], io_in[12], io_in[12], io_in[4:3], io_in[5], io_in[2], io_in[6], 4'h0, io_in[11:7], 3'h0, io_in[11:7], 3'h1, io_out_s_11_bits[3], io_out_s_11_bits[3], 2'h3 };
  assign io_out_s_reserved = { io_in[6:2], io_in[11:7], 15'h001f };
  assign io_out_s_sub = { _io_out_s_T_278[30], 30'h00000000 };
endmodule
module Rocket(clock, reset, io_hartid, io_interrupts_debug, io_interrupts_mtip, io_interrupts_msip, io_interrupts_meip, io_imem_might_request, io_imem_req_valid, io_imem_req_bits_pc, io_imem_req_bits_speculative, io_imem_resp_ready, io_imem_resp_valid, io_imem_resp_bits_pc, io_imem_resp_bits_data, io_imem_resp_bits_xcpt_ae_inst, io_imem_resp_bits_replay, io_imem_btb_update_valid, io_imem_bht_update_valid, io_imem_flush_icache, io_dmem_req_ready
, io_dmem_req_valid, io_dmem_req_bits_addr, io_dmem_req_bits_tag, io_dmem_req_bits_cmd, io_dmem_req_bits_size, io_dmem_req_bits_signed, io_dmem_req_bits_dv, io_dmem_s1_kill, io_dmem_s1_data_data, io_dmem_s2_nack, io_dmem_resp_valid, io_dmem_resp_bits_tag, io_dmem_resp_bits_data, io_dmem_resp_bits_replay, io_dmem_resp_bits_has_data, io_dmem_resp_bits_data_word_bypass, io_dmem_replay_next, io_dmem_s2_xcpt_ma_ld, io_dmem_s2_xcpt_ma_st, io_dmem_s2_xcpt_pf_ld, io_dmem_s2_xcpt_pf_st
, io_dmem_s2_xcpt_ae_ld, io_dmem_s2_xcpt_ae_st, io_dmem_ordered, io_dmem_perf_grant, io_ptw_status_debug, io_ptw_pmp_0_cfg_l, io_ptw_pmp_0_cfg_a, io_ptw_pmp_0_cfg_x, io_ptw_pmp_0_cfg_w, io_ptw_pmp_0_cfg_r, io_ptw_pmp_0_addr, io_ptw_pmp_0_mask, io_ptw_pmp_1_cfg_l, io_ptw_pmp_1_cfg_a, io_ptw_pmp_1_cfg_x, io_ptw_pmp_1_cfg_w, io_ptw_pmp_1_cfg_r, io_ptw_pmp_1_addr, io_ptw_pmp_1_mask, io_ptw_pmp_2_cfg_l, io_ptw_pmp_2_cfg_a
, io_ptw_pmp_2_cfg_x, io_ptw_pmp_2_cfg_w, io_ptw_pmp_2_cfg_r, io_ptw_pmp_2_addr, io_ptw_pmp_2_mask, io_ptw_pmp_3_cfg_l, io_ptw_pmp_3_cfg_a, io_ptw_pmp_3_cfg_x, io_ptw_pmp_3_cfg_w, io_ptw_pmp_3_cfg_r, io_ptw_pmp_3_addr, io_ptw_pmp_3_mask, io_ptw_pmp_4_cfg_l, io_ptw_pmp_4_cfg_a, io_ptw_pmp_4_cfg_x, io_ptw_pmp_4_cfg_w, io_ptw_pmp_4_cfg_r, io_ptw_pmp_4_addr, io_ptw_pmp_4_mask, io_ptw_pmp_5_cfg_l, io_ptw_pmp_5_cfg_a
, io_ptw_pmp_5_cfg_x, io_ptw_pmp_5_cfg_w, io_ptw_pmp_5_cfg_r, io_ptw_pmp_5_addr, io_ptw_pmp_5_mask, io_ptw_pmp_6_cfg_l, io_ptw_pmp_6_cfg_a, io_ptw_pmp_6_cfg_x, io_ptw_pmp_6_cfg_w, io_ptw_pmp_6_cfg_r, io_ptw_pmp_6_addr, io_ptw_pmp_6_mask, io_ptw_pmp_7_cfg_l, io_ptw_pmp_7_cfg_a, io_ptw_pmp_7_cfg_x, io_ptw_pmp_7_cfg_w, io_ptw_pmp_7_cfg_r, io_ptw_pmp_7_addr, io_ptw_pmp_7_mask, io_ptw_customCSRs_csrs_0_value, io_rocc_cmd_valid
, io_wfi);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire [1:0] _10441_;
  wire [1:0] _10442_;
  wire PlusArgTimeout_clock;
  wire [31:0] PlusArgTimeout_io_count;
  wire PlusArgTimeout_reset;
  wire [4:0] _T_11;
  wire [2:0] _T_113;
  wire [2:0] _T_114;
  wire [2:0] _T_115;
  wire [4:0] _T_116;
  wire [4:0] _T_118;
  wire [4:0] _T_119;
  wire [4:0] _T_12;
  wire [4:0] _T_13;
  wire [31:0] _T_143;
  wire [2:0] _T_35;
  wire [2:0] _T_37;
  wire _T_40;
  wire _T_41;
  wire _T_42;
  wire [3:0] _T_74;
  wire _T_93;
  wire [1:0] _bypass_src_T;
  wire [1:0] _bypass_src_T_2;
  wire [15:0] _csr_io_inst_0_T_3;
  wire [2:0] _csr_io_rw_cmd_T;
  wire [2:0] _csr_io_rw_cmd_T_1;
  wire _ctrl_stalld_T_15;
  wire _ex_imm_b11_T_5;
  wire _ex_imm_b11_T_8;
  wire [7:0] _ex_imm_b19_12_T_4;
  wire [10:0] _ex_imm_b30_20_T_2;
  wire _ex_imm_sign_T_2;
  wire [31:0] _ex_op1_T;
  wire [31:0] _ex_op2_T;
  wire [3:0] _ex_op2_T_1;
  wire _ex_reg_valid_T;
  wire [31:0] _ex_rs_T_13;
  wire [31:0] _ex_rs_T_6;
  wire [7:0] _id_ctrl_decoder_decoded_T;
  wire [8:0] _id_ctrl_decoder_decoded_T_10;
  wire [8:0] _id_ctrl_decoder_decoded_T_100;
  wire [8:0] _id_ctrl_decoder_decoded_T_102;
  wire [9:0] _id_ctrl_decoder_decoded_T_104;
  wire [13:0] _id_ctrl_decoder_decoded_T_106;
  wire [14:0] _id_ctrl_decoder_decoded_T_108;
  wire [14:0] _id_ctrl_decoder_decoded_T_110;
  wire [13:0] _id_ctrl_decoder_decoded_T_112;
  wire [16:0] _id_ctrl_decoder_decoded_T_114;
  wire [19:0] _id_ctrl_decoder_decoded_T_116;
  wire [27:0] _id_ctrl_decoder_decoded_T_118;
  wire [5:0] _id_ctrl_decoder_decoded_T_12;
  wire [30:0] _id_ctrl_decoder_decoded_T_120;
  wire [14:0] _id_ctrl_decoder_decoded_T_122;
  wire [12:0] _id_ctrl_decoder_decoded_T_124;
  wire [27:0] _id_ctrl_decoder_decoded_T_126;
  wire [31:0] _id_ctrl_decoder_decoded_T_128;
  wire [16:0] _id_ctrl_decoder_decoded_T_130;
  wire [12:0] _id_ctrl_decoder_decoded_T_132;
  wire [15:0] _id_ctrl_decoder_decoded_T_134;
  wire [27:0] _id_ctrl_decoder_decoded_T_136;
  wire [31:0] _id_ctrl_decoder_decoded_T_138;
  wire [6:0] _id_ctrl_decoder_decoded_T_14;
  wire [12:0] _id_ctrl_decoder_decoded_T_140;
  wire [8:0] _id_ctrl_decoder_decoded_T_16;
  wire [7:0] _id_ctrl_decoder_decoded_T_18;
  wire [7:0] _id_ctrl_decoder_decoded_T_2;
  wire [8:0] _id_ctrl_decoder_decoded_T_20;
  wire [15:0] _id_ctrl_decoder_decoded_T_22;
  wire [12:0] _id_ctrl_decoder_decoded_T_24;
  wire [7:0] _id_ctrl_decoder_decoded_T_26;
  wire [8:0] _id_ctrl_decoder_decoded_T_28;
  wire [8:0] _id_ctrl_decoder_decoded_T_30;
  wire [9:0] _id_ctrl_decoder_decoded_T_32;
  wire [6:0] _id_ctrl_decoder_decoded_T_34;
  wire [27:0] _id_ctrl_decoder_decoded_T_36;
  wire [30:0] _id_ctrl_decoder_decoded_T_38;
  wire [7:0] _id_ctrl_decoder_decoded_T_4;
  wire [9:0] _id_ctrl_decoder_decoded_T_40;
  wire [14:0] _id_ctrl_decoder_decoded_T_42;
  wire [15:0] _id_ctrl_decoder_decoded_T_44;
  wire [7:0] _id_ctrl_decoder_decoded_T_46;
  wire [8:0] _id_ctrl_decoder_decoded_T_48;
  wire [8:0] _id_ctrl_decoder_decoded_T_50;
  wire [7:0] _id_ctrl_decoder_decoded_T_52;
  wire [7:0] _id_ctrl_decoder_decoded_T_54;
  wire [8:0] _id_ctrl_decoder_decoded_T_56;
  wire [11:0] _id_ctrl_decoder_decoded_T_58;
  wire [7:0] _id_ctrl_decoder_decoded_T_6;
  wire [14:0] _id_ctrl_decoder_decoded_T_60;
  wire [15:0] _id_ctrl_decoder_decoded_T_62;
  wire [7:0] _id_ctrl_decoder_decoded_T_64;
  wire [8:0] _id_ctrl_decoder_decoded_T_66;
  wire [8:0] _id_ctrl_decoder_decoded_T_68;
  wire [14:0] _id_ctrl_decoder_decoded_T_70;
  wire [8:0] _id_ctrl_decoder_decoded_T_72;
  wire [13:0] _id_ctrl_decoder_decoded_T_74;
  wire [7:0] _id_ctrl_decoder_decoded_T_76;
  wire [14:0] _id_ctrl_decoder_decoded_T_78;
  wire [7:0] _id_ctrl_decoder_decoded_T_8;
  wire [15:0] _id_ctrl_decoder_decoded_T_80;
  wire [15:0] _id_ctrl_decoder_decoded_T_82;
  wire [15:0] _id_ctrl_decoder_decoded_T_84;
  wire [14:0] _id_ctrl_decoder_decoded_T_86;
  wire [7:0] _id_ctrl_decoder_decoded_T_88;
  wire [8:0] _id_ctrl_decoder_decoded_T_90;
  wire [8:0] _id_ctrl_decoder_decoded_T_92;
  wire [8:0] _id_ctrl_decoder_decoded_T_94;
  wire [14:0] _id_ctrl_decoder_decoded_T_96;
  wire [7:0] _id_ctrl_decoder_decoded_T_98;
  wire _id_illegal_insn_T_11;
  wire _id_illegal_insn_T_15;
  wire _id_illegal_insn_T_33;
  wire [31:0] _io_fpu_time_T;
  wire [31:0] _mem_br_target_T_3;
  wire [31:0] _mem_br_target_T_5;
  wire [3:0] _mem_br_target_T_6;
  wire [31:0] _mem_br_target_T_7;
  wire [31:0] _mem_br_target_T_8;
  wire _mem_reg_load_T_1;
  wire [31:0] _mem_reg_rs2_T_3;
  wire [31:0] _mem_reg_rs2_T_6;
  wire [31:0] _mem_reg_rs2_T_7;
  wire _mem_reg_valid_T;
  wire [31:0] _mem_reg_wdata_T;
  wire [31:0] _r;
  wire _take_pc_mem_T;
  wire _wb_reg_replay_T;
  wire _wb_reg_valid_T;
  wire [31:0] alu_io_adder_out;
  wire alu_io_cmp_out;
  wire [3:0] alu_io_fn;
  wire [31:0] alu_io_in1;
  wire [31:0] alu_io_in2;
  wire [31:0] alu_io_out;
  wire blocked;
  wire [31:0] bpu_io_bp_0_address;
  wire bpu_io_bp_0_control_action;
  wire bpu_io_bp_0_control_r;
  wire [1:0] bpu_io_bp_0_control_tmatch;
  wire bpu_io_bp_0_control_w;
  wire bpu_io_bp_0_control_x;
  wire bpu_io_debug_if;
  wire bpu_io_debug_ld;
  wire bpu_io_debug_st;
  wire [31:0] bpu_io_ea;
  wire [31:0] bpu_io_pc;
  wire bpu_io_status_debug;
  wire bpu_io_xcpt_if;
  wire bpu_io_xcpt_ld;
  wire bpu_io_xcpt_st;
  input clock;
  wire clock;
  wire [31:0] coreMonitorBundle_inst;
  wire [31:0] coreMonitorBundle_pc;
  wire csr_clock;
  wire [31:0] csr_io_bp_0_address;
  wire csr_io_bp_0_control_action;
  wire csr_io_bp_0_control_r;
  wire [1:0] csr_io_bp_0_control_tmatch;
  wire csr_io_bp_0_control_w;
  wire csr_io_bp_0_control_x;
  wire [31:0] csr_io_cause;
  wire csr_io_csr_stall;
  wire [31:0] csr_io_customCSRs_0_value;
  wire csr_io_decode_0_fp_csr;
  wire csr_io_decode_0_fp_illegal;
  wire [31:0] csr_io_decode_0_inst;
  wire csr_io_decode_0_read_illegal;
  wire csr_io_decode_0_rocc_illegal;
  wire csr_io_decode_0_system_illegal;
  wire csr_io_decode_0_write_flush;
  wire csr_io_decode_0_write_illegal;
  wire csr_io_eret;
  wire [31:0] csr_io_evec;
  wire csr_io_exception;
  wire csr_io_gva;
  wire csr_io_hartid;
  wire csr_io_inhibit_cycle;
  wire [31:0] csr_io_inst_0;
  wire csr_io_interrupt;
  wire [31:0] csr_io_interrupt_cause;
  wire csr_io_interrupts_debug;
  wire csr_io_interrupts_meip;
  wire csr_io_interrupts_msip;
  wire csr_io_interrupts_mtip;
  wire [31:0] csr_io_pc;
  wire [29:0] csr_io_pmp_0_addr;
  wire [1:0] csr_io_pmp_0_cfg_a;
  wire csr_io_pmp_0_cfg_l;
  wire csr_io_pmp_0_cfg_r;
  wire csr_io_pmp_0_cfg_w;
  wire csr_io_pmp_0_cfg_x;
  wire [31:0] csr_io_pmp_0_mask;
  wire [29:0] csr_io_pmp_1_addr;
  wire [1:0] csr_io_pmp_1_cfg_a;
  wire csr_io_pmp_1_cfg_l;
  wire csr_io_pmp_1_cfg_r;
  wire csr_io_pmp_1_cfg_w;
  wire csr_io_pmp_1_cfg_x;
  wire [31:0] csr_io_pmp_1_mask;
  wire [29:0] csr_io_pmp_2_addr;
  wire [1:0] csr_io_pmp_2_cfg_a;
  wire csr_io_pmp_2_cfg_l;
  wire csr_io_pmp_2_cfg_r;
  wire csr_io_pmp_2_cfg_w;
  wire csr_io_pmp_2_cfg_x;
  wire [31:0] csr_io_pmp_2_mask;
  wire [29:0] csr_io_pmp_3_addr;
  wire [1:0] csr_io_pmp_3_cfg_a;
  wire csr_io_pmp_3_cfg_l;
  wire csr_io_pmp_3_cfg_r;
  wire csr_io_pmp_3_cfg_w;
  wire csr_io_pmp_3_cfg_x;
  wire [31:0] csr_io_pmp_3_mask;
  wire [29:0] csr_io_pmp_4_addr;
  wire [1:0] csr_io_pmp_4_cfg_a;
  wire csr_io_pmp_4_cfg_l;
  wire csr_io_pmp_4_cfg_r;
  wire csr_io_pmp_4_cfg_w;
  wire csr_io_pmp_4_cfg_x;
  wire [31:0] csr_io_pmp_4_mask;
  wire [29:0] csr_io_pmp_5_addr;
  wire [1:0] csr_io_pmp_5_cfg_a;
  wire csr_io_pmp_5_cfg_l;
  wire csr_io_pmp_5_cfg_r;
  wire csr_io_pmp_5_cfg_w;
  wire csr_io_pmp_5_cfg_x;
  wire [31:0] csr_io_pmp_5_mask;
  wire [29:0] csr_io_pmp_6_addr;
  wire [1:0] csr_io_pmp_6_cfg_a;
  wire csr_io_pmp_6_cfg_l;
  wire csr_io_pmp_6_cfg_r;
  wire csr_io_pmp_6_cfg_w;
  wire csr_io_pmp_6_cfg_x;
  wire [31:0] csr_io_pmp_6_mask;
  wire [29:0] csr_io_pmp_7_addr;
  wire [1:0] csr_io_pmp_7_cfg_a;
  wire csr_io_pmp_7_cfg_l;
  wire csr_io_pmp_7_cfg_r;
  wire csr_io_pmp_7_cfg_w;
  wire csr_io_pmp_7_cfg_x;
  wire [31:0] csr_io_pmp_7_mask;
  wire csr_io_retire;
  wire [11:0] csr_io_rw_addr;
  wire [2:0] csr_io_rw_cmd;
  wire [31:0] csr_io_rw_rdata;
  wire [31:0] csr_io_rw_wdata;
  wire csr_io_singleStep;
  wire csr_io_status_cease;
  wire csr_io_status_debug;
  wire [1:0] csr_io_status_dprv;
  wire csr_io_status_dv;
  wire [1:0] csr_io_status_fs;
  wire csr_io_status_gva;
  wire csr_io_status_hie;
  wire [31:0] csr_io_status_isa;
  wire csr_io_status_mbe;
  wire csr_io_status_mie;
  wire csr_io_status_mpie;
  wire [1:0] csr_io_status_mpp;
  wire csr_io_status_mprv;
  wire csr_io_status_mpv;
  wire csr_io_status_mxr;
  wire [1:0] csr_io_status_prv;
  wire csr_io_status_sbe;
  wire csr_io_status_sd;
  wire csr_io_status_sd_rv32;
  wire csr_io_status_sie;
  wire csr_io_status_spie;
  wire csr_io_status_spp;
  wire csr_io_status_sum;
  wire [1:0] csr_io_status_sxl;
  wire csr_io_status_tsr;
  wire csr_io_status_tvm;
  wire csr_io_status_tw;
  wire csr_io_status_ube;
  wire csr_io_status_uie;
  wire csr_io_status_upie;
  wire [1:0] csr_io_status_uxl;
  wire csr_io_status_v;
  wire [1:0] csr_io_status_vs;
  wire csr_io_status_wfi;
  wire [1:0] csr_io_status_xs;
  wire [7:0] csr_io_status_zero1;
  wire [22:0] csr_io_status_zero2;
  wire [31:0] csr_io_time;
  wire csr_io_trace_0_exception;
  wire [31:0] csr_io_trace_0_iaddr;
  wire [31:0] csr_io_trace_0_insn;
  wire csr_io_trace_0_valid;
  wire [31:0] csr_io_tval;
  wire csr_io_ungated_clock;
  wire csr_reset;
  wire div_clock;
  wire div_io_kill;
  wire div_io_kill_REG;
  wire [3:0] div_io_req_bits_fn;
  wire [31:0] div_io_req_bits_in1;
  wire [31:0] div_io_req_bits_in2;
  wire [4:0] div_io_req_bits_tag;
  wire div_io_req_ready;
  wire div_io_req_valid;
  wire [31:0] div_io_resp_bits_data;
  wire [4:0] div_io_resp_bits_tag;
  wire div_io_resp_ready;
  wire div_io_resp_valid;
  wire div_reset;
  wire [4:0] dmem_resp_waddr;
  wire [3:0] ex_ctrl_alu_fn;
  wire ex_ctrl_branch;
  wire [2:0] ex_ctrl_csr;
  wire ex_ctrl_div;
  wire ex_ctrl_fence_i;
  wire ex_ctrl_fp;
  wire ex_ctrl_jal;
  wire ex_ctrl_jalr;
  wire ex_ctrl_mem;
  wire [4:0] ex_ctrl_mem_cmd;
  wire ex_ctrl_mul;
  wire ex_ctrl_rfs1;
  wire ex_ctrl_rfs2;
  wire ex_ctrl_rocc;
  wire ex_ctrl_rxs2;
  wire [1:0] ex_ctrl_sel_alu1;
  wire [1:0] ex_ctrl_sel_alu2;
  wire [2:0] ex_ctrl_sel_imm;
  wire ex_ctrl_wfd;
  wire ex_ctrl_wxd;
  wire [5:0] ex_dcache_tag;
  wire [31:0] ex_reg_cause;
  wire ex_reg_flush_pipe;
  wire [31:0] ex_reg_inst;
  wire ex_reg_load_use;
  wire [1:0] ex_reg_mem_size;
  wire [31:0] ex_reg_pc;
  wire [31:0] ex_reg_raw_inst;
  wire ex_reg_replay;
  wire ex_reg_rs_bypass_0;
  wire ex_reg_rs_bypass_1;
  wire [1:0] ex_reg_rs_lsb_0;
  wire [1:0] ex_reg_rs_lsb_1;
  wire [29:0] ex_reg_rs_msb_0;
  wire [29:0] ex_reg_rs_msb_1;
  wire ex_reg_rvc;
  wire ex_reg_valid;
  wire ex_reg_xcpt;
  wire ex_reg_xcpt_interrupt;
  wire [31:0] ex_rs_1;
  wire [4:0] ex_waddr;
  wire ibuf_clock;
  wire [31:0] ibuf_io_imem_bits_data;
  wire [31:0] ibuf_io_imem_bits_pc;
  wire ibuf_io_imem_bits_replay;
  wire ibuf_io_imem_bits_xcpt_ae_inst;
  wire ibuf_io_imem_ready;
  wire ibuf_io_imem_valid;
  wire [31:0] ibuf_io_inst_0_bits_inst_bits;
  wire [4:0] ibuf_io_inst_0_bits_inst_rd;
  wire [4:0] ibuf_io_inst_0_bits_inst_rs1;
  wire [4:0] ibuf_io_inst_0_bits_inst_rs2;
  wire [31:0] ibuf_io_inst_0_bits_raw;
  wire ibuf_io_inst_0_bits_replay;
  wire ibuf_io_inst_0_bits_rvc;
  wire ibuf_io_inst_0_bits_xcpt0_ae_inst;
  wire ibuf_io_inst_0_bits_xcpt1_ae_inst;
  wire ibuf_io_inst_0_bits_xcpt1_gf_inst;
  wire ibuf_io_inst_0_bits_xcpt1_pf_inst;
  wire ibuf_io_inst_0_ready;
  wire ibuf_io_inst_0_valid;
  wire ibuf_io_kill;
  wire [31:0] ibuf_io_pc;
  wire ibuf_reset;
  wire id_amo_aq;
  wire id_amo_rl;
  wire id_ctrl_decoder_1;
  wire [4:0] id_ctrl_decoder_15;
  wire id_ctrl_decoder_16;
  wire id_ctrl_decoder_17;
  wire id_ctrl_decoder_19;
  wire id_ctrl_decoder_2;
  wire id_ctrl_decoder_20;
  wire id_ctrl_decoder_27;
  wire id_ctrl_decoder_8;
  wire id_ctrl_decoder_decoded_andMatrixInput_0;
  wire id_ctrl_decoder_decoded_andMatrixInput_1;
  wire id_ctrl_decoder_decoded_andMatrixInput_10;
  wire id_ctrl_decoder_decoded_andMatrixInput_10_20;
  wire id_ctrl_decoder_decoded_andMatrixInput_11;
  wire id_ctrl_decoder_decoded_andMatrixInput_11_1;
  wire id_ctrl_decoder_decoded_andMatrixInput_12;
  wire id_ctrl_decoder_decoded_andMatrixInput_12_2;
  wire id_ctrl_decoder_decoded_andMatrixInput_12_25;
  wire id_ctrl_decoder_decoded_andMatrixInput_12_33;
  wire id_ctrl_decoder_decoded_andMatrixInput_13;
  wire id_ctrl_decoder_decoded_andMatrixInput_13_1;
  wire id_ctrl_decoder_decoded_andMatrixInput_13_19;
  wire id_ctrl_decoder_decoded_andMatrixInput_14;
  wire id_ctrl_decoder_decoded_andMatrixInput_14_1;
  wire id_ctrl_decoder_decoded_andMatrixInput_15;
  wire id_ctrl_decoder_decoded_andMatrixInput_15_1;
  wire id_ctrl_decoder_decoded_andMatrixInput_15_14;
  wire id_ctrl_decoder_decoded_andMatrixInput_16;
  wire id_ctrl_decoder_decoded_andMatrixInput_17;
  wire id_ctrl_decoder_decoded_andMatrixInput_17_3;
  wire id_ctrl_decoder_decoded_andMatrixInput_17_5;
  wire id_ctrl_decoder_decoded_andMatrixInput_18;
  wire id_ctrl_decoder_decoded_andMatrixInput_19;
  wire id_ctrl_decoder_decoded_andMatrixInput_19_3;
  wire id_ctrl_decoder_decoded_andMatrixInput_2;
  wire id_ctrl_decoder_decoded_andMatrixInput_20;
  wire id_ctrl_decoder_decoded_andMatrixInput_20_6;
  wire id_ctrl_decoder_decoded_andMatrixInput_2_5;
  wire id_ctrl_decoder_decoded_andMatrixInput_3;
  wire id_ctrl_decoder_decoded_andMatrixInput_3_5;
  wire id_ctrl_decoder_decoded_andMatrixInput_4;
  wire id_ctrl_decoder_decoded_andMatrixInput_4_18;
  wire id_ctrl_decoder_decoded_andMatrixInput_4_6;
  wire id_ctrl_decoder_decoded_andMatrixInput_5;
  wire id_ctrl_decoder_decoded_andMatrixInput_5_18;
  wire id_ctrl_decoder_decoded_andMatrixInput_5_8;
  wire id_ctrl_decoder_decoded_andMatrixInput_6;
  wire id_ctrl_decoder_decoded_andMatrixInput_6_1;
  wire id_ctrl_decoder_decoded_andMatrixInput_6_12;
  wire id_ctrl_decoder_decoded_andMatrixInput_6_17;
  wire id_ctrl_decoder_decoded_andMatrixInput_7;
  wire id_ctrl_decoder_decoded_andMatrixInput_7_15;
  wire id_ctrl_decoder_decoded_andMatrixInput_7_17;
  wire id_ctrl_decoder_decoded_andMatrixInput_7_2;
  wire id_ctrl_decoder_decoded_andMatrixInput_7_24;
  wire id_ctrl_decoder_decoded_andMatrixInput_7_50;
  wire id_ctrl_decoder_decoded_andMatrixInput_7_54;
  wire id_ctrl_decoder_decoded_andMatrixInput_8_22;
  wire id_ctrl_decoder_decoded_andMatrixInput_8_8;
  wire [9:0] id_ctrl_decoder_decoded_hi_58;
  wire [6:0] id_ctrl_decoder_decoded_hi_lo_17;
  wire [7:0] id_ctrl_decoder_decoded_hi_lo_18;
  wire [6:0] id_ctrl_decoder_decoded_hi_lo_62;
  wire [31:0] id_ctrl_decoder_decoded_invInputs;
  wire [40:0] id_ctrl_decoder_decoded_invMatrixOutputs;
  wire [4:0] id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_lo;
  wire [9:0] id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi;
  wire [9:0] id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo;
  wire [7:0] id_ctrl_decoder_decoded_lo_11;
  wire [5:0] id_ctrl_decoder_decoded_lo_12;
  wire [13:0] id_ctrl_decoder_decoded_lo_18;
  wire [14:0] id_ctrl_decoder_decoded_lo_19;
  wire [7:0] id_ctrl_decoder_decoded_lo_22;
  wire [5:0] id_ctrl_decoder_decoded_lo_29;
  wire [7:0] id_ctrl_decoder_decoded_lo_31;
  wire [6:0] id_ctrl_decoder_decoded_lo_35;
  wire [6:0] id_ctrl_decoder_decoded_lo_37;
  wire [6:0] id_ctrl_decoder_decoded_lo_39;
  wire [7:0] id_ctrl_decoder_decoded_lo_40;
  wire [7:0] id_ctrl_decoder_decoded_lo_41;
  wire [6:0] id_ctrl_decoder_decoded_lo_53;
  wire [6:0] id_ctrl_decoder_decoded_lo_56;
  wire [7:0] id_ctrl_decoder_decoded_lo_57;
  wire [9:0] id_ctrl_decoder_decoded_lo_58;
  wire [13:0] id_ctrl_decoder_decoded_lo_59;
  wire [14:0] id_ctrl_decoder_decoded_lo_60;
  wire [6:0] id_ctrl_decoder_decoded_lo_61;
  wire [5:0] id_ctrl_decoder_decoded_lo_62;
  wire [13:0] id_ctrl_decoder_decoded_lo_63;
  wire [15:0] id_ctrl_decoder_decoded_lo_64;
  wire [7:0] id_ctrl_decoder_decoded_lo_65;
  wire [5:0] id_ctrl_decoder_decoded_lo_66;
  wire [7:0] id_ctrl_decoder_decoded_lo_67;
  wire [13:0] id_ctrl_decoder_decoded_lo_68;
  wire [15:0] id_ctrl_decoder_decoded_lo_69;
  wire [5:0] id_ctrl_decoder_decoded_lo_70;
  wire [6:0] id_ctrl_decoder_decoded_lo_lo_15;
  wire [6:0] id_ctrl_decoder_decoded_lo_lo_56;
  wire [6:0] id_ctrl_decoder_decoded_lo_lo_60;
  wire [7:0] id_ctrl_decoder_decoded_lo_lo_61;
  wire [6:0] id_ctrl_decoder_decoded_lo_lo_65;
  wire [7:0] id_ctrl_decoder_decoded_lo_lo_66;
  wire [40:0] id_ctrl_decoder_decoded_orMatrixOutputs;
  wire [4:0] id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_6;
  wire [19:0] id_ctrl_decoder_decoded_orMatrixOutputs_lo_17;
  wire [9:0] id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_10;
  wire [31:0] id_ctrl_decoder_decoded_plaInput;
  wire [3:0] id_fence_succ;
  wire [4:0] id_raddr1;
  wire [4:0] id_raddr2;
  wire id_reg_fence;
  wire id_reg_pause;
  wire [4:0] id_waddr;
  wire imem_might_request_reg;
  wire [31:0] inst;
  input io_dmem_ordered;
  wire io_dmem_ordered;
  input io_dmem_perf_grant;
  wire io_dmem_perf_grant;
  input io_dmem_replay_next;
  wire io_dmem_replay_next;
  output [31:0] io_dmem_req_bits_addr;
  wire [31:0] io_dmem_req_bits_addr;
  output [4:0] io_dmem_req_bits_cmd;
  wire [4:0] io_dmem_req_bits_cmd;
  output io_dmem_req_bits_dv;
  wire io_dmem_req_bits_dv;
  output io_dmem_req_bits_signed;
  wire io_dmem_req_bits_signed;
  output [1:0] io_dmem_req_bits_size;
  wire [1:0] io_dmem_req_bits_size;
  output [6:0] io_dmem_req_bits_tag;
  wire [6:0] io_dmem_req_bits_tag;
  input io_dmem_req_ready;
  wire io_dmem_req_ready;
  output io_dmem_req_valid;
  wire io_dmem_req_valid;
  input [31:0] io_dmem_resp_bits_data;
  wire [31:0] io_dmem_resp_bits_data;
  input [31:0] io_dmem_resp_bits_data_word_bypass;
  wire [31:0] io_dmem_resp_bits_data_word_bypass;
  input io_dmem_resp_bits_has_data;
  wire io_dmem_resp_bits_has_data;
  input io_dmem_resp_bits_replay;
  wire io_dmem_resp_bits_replay;
  input [6:0] io_dmem_resp_bits_tag;
  wire [6:0] io_dmem_resp_bits_tag;
  input io_dmem_resp_valid;
  wire io_dmem_resp_valid;
  output [31:0] io_dmem_s1_data_data;
  wire [31:0] io_dmem_s1_data_data;
  output io_dmem_s1_kill;
  wire io_dmem_s1_kill;
  input io_dmem_s2_nack;
  wire io_dmem_s2_nack;
  input io_dmem_s2_xcpt_ae_ld;
  wire io_dmem_s2_xcpt_ae_ld;
  input io_dmem_s2_xcpt_ae_st;
  wire io_dmem_s2_xcpt_ae_st;
  input io_dmem_s2_xcpt_ma_ld;
  wire io_dmem_s2_xcpt_ma_ld;
  input io_dmem_s2_xcpt_ma_st;
  wire io_dmem_s2_xcpt_ma_st;
  input io_dmem_s2_xcpt_pf_ld;
  wire io_dmem_s2_xcpt_pf_ld;
  input io_dmem_s2_xcpt_pf_st;
  wire io_dmem_s2_xcpt_pf_st;
  input io_hartid;
  wire io_hartid;
  output io_imem_bht_update_valid;
  wire io_imem_bht_update_valid;
  output io_imem_btb_update_valid;
  wire io_imem_btb_update_valid;
  output io_imem_flush_icache;
  wire io_imem_flush_icache;
  output io_imem_might_request;
  wire io_imem_might_request;
  output [31:0] io_imem_req_bits_pc;
  wire [31:0] io_imem_req_bits_pc;
  output io_imem_req_bits_speculative;
  wire io_imem_req_bits_speculative;
  output io_imem_req_valid;
  wire io_imem_req_valid;
  input [31:0] io_imem_resp_bits_data;
  wire [31:0] io_imem_resp_bits_data;
  input [31:0] io_imem_resp_bits_pc;
  wire [31:0] io_imem_resp_bits_pc;
  input io_imem_resp_bits_replay;
  wire io_imem_resp_bits_replay;
  input io_imem_resp_bits_xcpt_ae_inst;
  wire io_imem_resp_bits_xcpt_ae_inst;
  output io_imem_resp_ready;
  wire io_imem_resp_ready;
  input io_imem_resp_valid;
  wire io_imem_resp_valid;
  input io_interrupts_debug;
  wire io_interrupts_debug;
  input io_interrupts_meip;
  wire io_interrupts_meip;
  input io_interrupts_msip;
  wire io_interrupts_msip;
  input io_interrupts_mtip;
  wire io_interrupts_mtip;
  output [31:0] io_ptw_customCSRs_csrs_0_value;
  wire [31:0] io_ptw_customCSRs_csrs_0_value;
  output [29:0] io_ptw_pmp_0_addr;
  wire [29:0] io_ptw_pmp_0_addr;
  output [1:0] io_ptw_pmp_0_cfg_a;
  wire [1:0] io_ptw_pmp_0_cfg_a;
  output io_ptw_pmp_0_cfg_l;
  wire io_ptw_pmp_0_cfg_l;
  output io_ptw_pmp_0_cfg_r;
  wire io_ptw_pmp_0_cfg_r;
  output io_ptw_pmp_0_cfg_w;
  wire io_ptw_pmp_0_cfg_w;
  output io_ptw_pmp_0_cfg_x;
  wire io_ptw_pmp_0_cfg_x;
  output [31:0] io_ptw_pmp_0_mask;
  wire [31:0] io_ptw_pmp_0_mask;
  output [29:0] io_ptw_pmp_1_addr;
  wire [29:0] io_ptw_pmp_1_addr;
  output [1:0] io_ptw_pmp_1_cfg_a;
  wire [1:0] io_ptw_pmp_1_cfg_a;
  output io_ptw_pmp_1_cfg_l;
  wire io_ptw_pmp_1_cfg_l;
  output io_ptw_pmp_1_cfg_r;
  wire io_ptw_pmp_1_cfg_r;
  output io_ptw_pmp_1_cfg_w;
  wire io_ptw_pmp_1_cfg_w;
  output io_ptw_pmp_1_cfg_x;
  wire io_ptw_pmp_1_cfg_x;
  output [31:0] io_ptw_pmp_1_mask;
  wire [31:0] io_ptw_pmp_1_mask;
  output [29:0] io_ptw_pmp_2_addr;
  wire [29:0] io_ptw_pmp_2_addr;
  output [1:0] io_ptw_pmp_2_cfg_a;
  wire [1:0] io_ptw_pmp_2_cfg_a;
  output io_ptw_pmp_2_cfg_l;
  wire io_ptw_pmp_2_cfg_l;
  output io_ptw_pmp_2_cfg_r;
  wire io_ptw_pmp_2_cfg_r;
  output io_ptw_pmp_2_cfg_w;
  wire io_ptw_pmp_2_cfg_w;
  output io_ptw_pmp_2_cfg_x;
  wire io_ptw_pmp_2_cfg_x;
  output [31:0] io_ptw_pmp_2_mask;
  wire [31:0] io_ptw_pmp_2_mask;
  output [29:0] io_ptw_pmp_3_addr;
  wire [29:0] io_ptw_pmp_3_addr;
  output [1:0] io_ptw_pmp_3_cfg_a;
  wire [1:0] io_ptw_pmp_3_cfg_a;
  output io_ptw_pmp_3_cfg_l;
  wire io_ptw_pmp_3_cfg_l;
  output io_ptw_pmp_3_cfg_r;
  wire io_ptw_pmp_3_cfg_r;
  output io_ptw_pmp_3_cfg_w;
  wire io_ptw_pmp_3_cfg_w;
  output io_ptw_pmp_3_cfg_x;
  wire io_ptw_pmp_3_cfg_x;
  output [31:0] io_ptw_pmp_3_mask;
  wire [31:0] io_ptw_pmp_3_mask;
  output [29:0] io_ptw_pmp_4_addr;
  wire [29:0] io_ptw_pmp_4_addr;
  output [1:0] io_ptw_pmp_4_cfg_a;
  wire [1:0] io_ptw_pmp_4_cfg_a;
  output io_ptw_pmp_4_cfg_l;
  wire io_ptw_pmp_4_cfg_l;
  output io_ptw_pmp_4_cfg_r;
  wire io_ptw_pmp_4_cfg_r;
  output io_ptw_pmp_4_cfg_w;
  wire io_ptw_pmp_4_cfg_w;
  output io_ptw_pmp_4_cfg_x;
  wire io_ptw_pmp_4_cfg_x;
  output [31:0] io_ptw_pmp_4_mask;
  wire [31:0] io_ptw_pmp_4_mask;
  output [29:0] io_ptw_pmp_5_addr;
  wire [29:0] io_ptw_pmp_5_addr;
  output [1:0] io_ptw_pmp_5_cfg_a;
  wire [1:0] io_ptw_pmp_5_cfg_a;
  output io_ptw_pmp_5_cfg_l;
  wire io_ptw_pmp_5_cfg_l;
  output io_ptw_pmp_5_cfg_r;
  wire io_ptw_pmp_5_cfg_r;
  output io_ptw_pmp_5_cfg_w;
  wire io_ptw_pmp_5_cfg_w;
  output io_ptw_pmp_5_cfg_x;
  wire io_ptw_pmp_5_cfg_x;
  output [31:0] io_ptw_pmp_5_mask;
  wire [31:0] io_ptw_pmp_5_mask;
  output [29:0] io_ptw_pmp_6_addr;
  wire [29:0] io_ptw_pmp_6_addr;
  output [1:0] io_ptw_pmp_6_cfg_a;
  wire [1:0] io_ptw_pmp_6_cfg_a;
  output io_ptw_pmp_6_cfg_l;
  wire io_ptw_pmp_6_cfg_l;
  output io_ptw_pmp_6_cfg_r;
  wire io_ptw_pmp_6_cfg_r;
  output io_ptw_pmp_6_cfg_w;
  wire io_ptw_pmp_6_cfg_w;
  output io_ptw_pmp_6_cfg_x;
  wire io_ptw_pmp_6_cfg_x;
  output [31:0] io_ptw_pmp_6_mask;
  wire [31:0] io_ptw_pmp_6_mask;
  output [29:0] io_ptw_pmp_7_addr;
  wire [29:0] io_ptw_pmp_7_addr;
  output [1:0] io_ptw_pmp_7_cfg_a;
  wire [1:0] io_ptw_pmp_7_cfg_a;
  output io_ptw_pmp_7_cfg_l;
  wire io_ptw_pmp_7_cfg_l;
  output io_ptw_pmp_7_cfg_r;
  wire io_ptw_pmp_7_cfg_r;
  output io_ptw_pmp_7_cfg_w;
  wire io_ptw_pmp_7_cfg_w;
  output io_ptw_pmp_7_cfg_x;
  wire io_ptw_pmp_7_cfg_x;
  output [31:0] io_ptw_pmp_7_mask;
  wire [31:0] io_ptw_pmp_7_mask;
  output io_ptw_status_debug;
  wire io_ptw_status_debug;
  output io_rocc_cmd_valid;
  wire io_rocc_cmd_valid;
  output io_wfi;
  wire io_wfi;
  wire [31:0] ll_wdata;
  wire mem_br_taken;
  wire [31:0] mem_br_target;
  wire [5:0] mem_br_target_b10_5;
  wire [3:0] mem_br_target_b4_1;
  wire mem_br_target_hi_hi_hi;
  wire [10:0] mem_br_target_hi_hi_lo;
  wire [7:0] mem_br_target_hi_lo_hi;
  wire [7:0] mem_br_target_hi_lo_hi_1;
  wire mem_br_target_hi_lo_lo;
  wire mem_br_target_hi_lo_lo_1;
  wire mem_br_target_sign;
  wire mem_ctrl_branch;
  wire [2:0] mem_ctrl_csr;
  wire mem_ctrl_div;
  wire mem_ctrl_fence_i;
  wire mem_ctrl_fp;
  wire mem_ctrl_jal;
  wire mem_ctrl_jalr;
  wire mem_ctrl_mem;
  wire mem_ctrl_mul;
  wire mem_ctrl_rocc;
  wire mem_ctrl_wxd;
  wire [3:0] mem_ldst_cause;
  wire [31:0] mem_npc;
  wire [31:0] mem_reg_cause;
  wire mem_reg_flush_pipe;
  wire mem_reg_hls_or_dv;
  wire [31:0] mem_reg_inst;
  wire mem_reg_load;
  wire [31:0] mem_reg_pc;
  wire [31:0] mem_reg_raw_inst;
  wire mem_reg_replay;
  wire [31:0] mem_reg_rs2;
  wire mem_reg_rvc;
  wire mem_reg_slow_bypass;
  wire mem_reg_store;
  wire mem_reg_valid;
  wire [31:0] mem_reg_wdata;
  wire mem_reg_xcpt;
  wire mem_reg_xcpt_interrupt;
  wire [4:0] mem_waddr;
  wire [31:0] r;
  wire replay_wb_rocc;
  input reset;
  wire reset;
  wire [31:0] \rf[0] ;
  wire [31:0] \rf[10] ;
  wire [31:0] \rf[11] ;
  wire [31:0] \rf[12] ;
  wire [31:0] \rf[13] ;
  wire [31:0] \rf[14] ;
  wire [31:0] \rf[15] ;
  wire [31:0] \rf[16] ;
  wire [31:0] \rf[17] ;
  wire [31:0] \rf[18] ;
  wire [31:0] \rf[19] ;
  wire [31:0] \rf[1] ;
  wire [31:0] \rf[20] ;
  wire [31:0] \rf[21] ;
  wire [31:0] \rf[22] ;
  wire [31:0] \rf[23] ;
  wire [31:0] \rf[24] ;
  wire [31:0] \rf[25] ;
  wire [31:0] \rf[26] ;
  wire [31:0] \rf[27] ;
  wire [31:0] \rf[28] ;
  wire [31:0] \rf[29] ;
  wire [31:0] \rf[2] ;
  wire [31:0] \rf[30] ;
  wire [31:0] \rf[3] ;
  wire [31:0] \rf[4] ;
  wire [31:0] \rf[5] ;
  wire [31:0] \rf[6] ;
  wire [31:0] \rf[7] ;
  wire [31:0] \rf[8] ;
  wire [31:0] \rf[9] ;
  wire rf_MPORT_mask;
  wire rf_id_rs_MPORT_1_en;
  wire rf_id_rs_MPORT_en;
  wire [1:0] size;
  wire take_pc_mem_wb;
  wire tval_dmem_addr;
  wire [2:0] wb_ctrl_csr;
  wire wb_ctrl_div;
  wire wb_ctrl_fence_i;
  wire wb_ctrl_mem;
  wire wb_ctrl_rocc;
  wire wb_ctrl_wxd;
  wire [31:0] wb_reg_cause;
  wire wb_reg_flush_pipe;
  wire wb_reg_hls_or_dv;
  wire [31:0] wb_reg_inst;
  wire [31:0] wb_reg_pc;
  wire [31:0] wb_reg_raw_inst;
  wire wb_reg_replay;
  wire wb_reg_valid;
  wire [31:0] wb_reg_wdata;
  wire wb_reg_xcpt;
  wire wb_valid;
  wire [4:0] wb_waddr;
  wire wb_xcpt;
  INV_X1 _10443_ (
    .A(csr_io_interrupt),
    .ZN(_02978_)
  );
  INV_X1 _10444_ (
    .A(reset),
    .ZN(_02979_)
  );
  INV_X1 _10445_ (
    .A(ex_reg_rs_lsb_0[0]),
    .ZN(_02980_)
  );
  INV_X1 _10446_ (
    .A(mem_reg_wdata[28]),
    .ZN(_02981_)
  );
  INV_X1 _10447_ (
    .A(mem_reg_inst[7]),
    .ZN(_02982_)
  );
  INV_X1 _10448_ (
    .A(ex_reg_inst[7]),
    .ZN(_02983_)
  );
  INV_X1 _10449_ (
    .A(mem_reg_inst[8]),
    .ZN(_02984_)
  );
  INV_X1 _10450_ (
    .A(ex_reg_inst[8]),
    .ZN(_02985_)
  );
  INV_X1 _10451_ (
    .A(mem_reg_inst[9]),
    .ZN(_02986_)
  );
  INV_X1 _10452_ (
    .A(mem_reg_inst[10]),
    .ZN(_02987_)
  );
  INV_X1 _10453_ (
    .A(ex_reg_inst[10]),
    .ZN(_02988_)
  );
  INV_X1 _10454_ (
    .A(mem_reg_inst[11]),
    .ZN(_02989_)
  );
  INV_X1 _10455_ (
    .A(ex_reg_inst[11]),
    .ZN(_02990_)
  );
  INV_X1 _10456_ (
    .A(ex_reg_pc[4]),
    .ZN(_02991_)
  );
  INV_X1 _10457_ (
    .A(ex_reg_pc[10]),
    .ZN(_02992_)
  );
  INV_X1 _10458_ (
    .A(ex_reg_pc[11]),
    .ZN(_02993_)
  );
  INV_X1 _10459_ (
    .A(ex_reg_pc[12]),
    .ZN(_02994_)
  );
  INV_X1 _10460_ (
    .A(ex_reg_pc[13]),
    .ZN(_02995_)
  );
  INV_X1 _10461_ (
    .A(ex_reg_pc[14]),
    .ZN(_02996_)
  );
  INV_X1 _10462_ (
    .A(ex_reg_pc[15]),
    .ZN(_02997_)
  );
  INV_X1 _10463_ (
    .A(ex_reg_pc[16]),
    .ZN(_02998_)
  );
  INV_X1 _10464_ (
    .A(ex_reg_pc[17]),
    .ZN(_02999_)
  );
  INV_X1 _10465_ (
    .A(csr_io_decode_0_inst[12]),
    .ZN(_03000_)
  );
  INV_X1 _10466_ (
    .A(csr_io_decode_0_inst[13]),
    .ZN(_03001_)
  );
  INV_X1 _10467_ (
    .A(csr_io_decode_0_inst[14]),
    .ZN(_03002_)
  );
  INV_X1 _10468_ (
    .A(csr_io_decode_0_inst[23]),
    .ZN(_03003_)
  );
  INV_X1 _10469_ (
    .A(csr_io_decode_0_inst[25]),
    .ZN(_03004_)
  );
  INV_X1 _10470_ (
    .A(csr_io_decode_0_inst[26]),
    .ZN(_03005_)
  );
  INV_X1 _10471_ (
    .A(csr_io_decode_0_inst[27]),
    .ZN(_03006_)
  );
  INV_X1 _10472_ (
    .A(csr_io_decode_0_inst[28]),
    .ZN(_03007_)
  );
  INV_X1 _10473_ (
    .A(csr_io_decode_0_inst[29]),
    .ZN(_03008_)
  );
  INV_X1 _10474_ (
    .A(csr_io_decode_0_inst[31]),
    .ZN(_03009_)
  );
  INV_X1 _10475_ (
    .A(ex_reg_mem_size[1]),
    .ZN(_03010_)
  );
  INV_X1 _10476_ (
    .A(bpu_io_pc[3]),
    .ZN(_03011_)
  );
  INV_X1 _10477_ (
    .A(bpu_io_pc[4]),
    .ZN(_03012_)
  );
  INV_X1 _10478_ (
    .A(bpu_io_pc[5]),
    .ZN(_03013_)
  );
  INV_X1 _10479_ (
    .A(bpu_io_pc[6]),
    .ZN(_03014_)
  );
  INV_X1 _10480_ (
    .A(bpu_io_pc[7]),
    .ZN(_03015_)
  );
  INV_X1 _10481_ (
    .A(bpu_io_pc[8]),
    .ZN(_03016_)
  );
  INV_X1 _10482_ (
    .A(bpu_io_pc[9]),
    .ZN(_03017_)
  );
  INV_X1 _10483_ (
    .A(bpu_io_pc[10]),
    .ZN(_03018_)
  );
  INV_X1 _10484_ (
    .A(bpu_io_pc[11]),
    .ZN(_03019_)
  );
  INV_X1 _10485_ (
    .A(bpu_io_pc[12]),
    .ZN(_03020_)
  );
  INV_X1 _10486_ (
    .A(bpu_io_pc[13]),
    .ZN(_03021_)
  );
  INV_X1 _10487_ (
    .A(bpu_io_pc[14]),
    .ZN(_03022_)
  );
  INV_X1 _10488_ (
    .A(bpu_io_pc[17]),
    .ZN(_03023_)
  );
  INV_X1 _10489_ (
    .A(bpu_io_pc[28]),
    .ZN(_03024_)
  );
  INV_X1 _10490_ (
    .A(wb_ctrl_wxd),
    .ZN(_03025_)
  );
  INV_X1 _10491_ (
    .A(wb_reg_inst[8]),
    .ZN(_03026_)
  );
  INV_X1 _10492_ (
    .A(wb_reg_inst[9]),
    .ZN(_03027_)
  );
  INV_X1 _10493_ (
    .A(wb_reg_inst[10]),
    .ZN(_03028_)
  );
  INV_X1 _10494_ (
    .A(wb_reg_inst[11]),
    .ZN(_03029_)
  );
  INV_X1 _10495_ (
    .A(mem_ctrl_jalr),
    .ZN(_03030_)
  );
  INV_X1 _10496_ (
    .A(mem_ctrl_branch),
    .ZN(_03031_)
  );
  INV_X1 _10497_ (
    .A(ex_ctrl_mem_cmd[0]),
    .ZN(_03032_)
  );
  INV_X1 _10498_ (
    .A(ex_ctrl_sel_alu1[0]),
    .ZN(_03033_)
  );
  INV_X1 _10499_ (
    .A(ex_ctrl_rxs2),
    .ZN(_03034_)
  );
  INV_X1 _10500_ (
    .A(ex_reg_rs_lsb_1[0]),
    .ZN(_03035_)
  );
  INV_X1 _10501_ (
    .A(csr_io_decode_0_inst[6]),
    .ZN(_03036_)
  );
  INV_X1 _10502_ (
    .A(csr_io_decode_0_inst[2]),
    .ZN(_03037_)
  );
  INV_X1 _10503_ (
    .A(csr_io_decode_0_inst[5]),
    .ZN(_03038_)
  );
  INV_X1 _10504_ (
    .A(csr_io_decode_0_inst[4]),
    .ZN(_03039_)
  );
  INV_X1 _10505_ (
    .A(csr_io_decode_0_inst[3]),
    .ZN(_03040_)
  );
  INV_X1 _10506_ (
    .A(_00021_),
    .ZN(_03041_)
  );
  INV_X1 _10507_ (
    .A(_00012_),
    .ZN(_03042_)
  );
  INV_X1 _10508_ (
    .A(_00018_),
    .ZN(_03043_)
  );
  INV_X1 _10509_ (
    .A(ibuf_io_inst_0_bits_inst_rs1[0]),
    .ZN(_03044_)
  );
  INV_X1 _10510_ (
    .A(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_03045_)
  );
  INV_X1 _10511_ (
    .A(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_03046_)
  );
  INV_X1 _10512_ (
    .A(ibuf_io_inst_0_bits_inst_rs1[3]),
    .ZN(_03047_)
  );
  INV_X1 _10513_ (
    .A(ibuf_io_inst_0_bits_inst_rs2[0]),
    .ZN(_03048_)
  );
  INV_X1 _10514_ (
    .A(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_03049_)
  );
  INV_X1 _10515_ (
    .A(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03050_)
  );
  INV_X1 _10516_ (
    .A(ibuf_io_inst_0_bits_inst_rs2[3]),
    .ZN(_03051_)
  );
  INV_X1 _10517_ (
    .A(ibuf_io_inst_0_bits_inst_rd[0]),
    .ZN(_03052_)
  );
  INV_X1 _10518_ (
    .A(ibuf_io_inst_0_bits_inst_rd[1]),
    .ZN(_03053_)
  );
  INV_X1 _10519_ (
    .A(ibuf_io_inst_0_bits_inst_rd[2]),
    .ZN(_03054_)
  );
  INV_X1 _10520_ (
    .A(ibuf_io_inst_0_bits_inst_rd[3]),
    .ZN(_03055_)
  );
  INV_X1 _10521_ (
    .A(_00027_),
    .ZN(_03056_)
  );
  INV_X1 _10522_ (
    .A(_00026_),
    .ZN(_03057_)
  );
  INV_X1 _10523_ (
    .A(_10441_[0]),
    .ZN(_03058_)
  );
  INV_X1 _10524_ (
    .A(_00019_),
    .ZN(_03059_)
  );
  INV_X1 _10525_ (
    .A(ibuf_io_inst_0_bits_xcpt1_gf_inst),
    .ZN(_03060_)
  );
  INV_X1 _10526_ (
    .A(_00031_),
    .ZN(_03061_)
  );
  INV_X1 _10527_ (
    .A(_00035_),
    .ZN(_03062_)
  );
  INV_X1 _10528_ (
    .A(ibuf_io_inst_0_bits_inst_rs1[4]),
    .ZN(_03063_)
  );
  INV_X1 _10529_ (
    .A(ibuf_io_inst_0_bits_inst_rs2[4]),
    .ZN(_03064_)
  );
  INV_X1 _10530_ (
    .A(ibuf_io_inst_0_bits_rvc),
    .ZN(_03065_)
  );
  INV_X1 _10531_ (
    .A(ibuf_io_inst_0_bits_xcpt0_ae_inst),
    .ZN(_03066_)
  );
  INV_X1 _10532_ (
    .A(bpu_io_xcpt_if),
    .ZN(_03067_)
  );
  INV_X1 _10533_ (
    .A(div_io_resp_bits_tag[0]),
    .ZN(_03068_)
  );
  INV_X1 _10534_ (
    .A(io_dmem_resp_bits_tag[1]),
    .ZN(_03069_)
  );
  INV_X1 _10535_ (
    .A(div_io_resp_bits_tag[1]),
    .ZN(_03070_)
  );
  INV_X1 _10536_ (
    .A(io_dmem_resp_bits_tag[2]),
    .ZN(_03071_)
  );
  INV_X1 _10537_ (
    .A(div_io_resp_bits_tag[2]),
    .ZN(_03072_)
  );
  INV_X1 _10538_ (
    .A(io_dmem_resp_bits_tag[3]),
    .ZN(_03073_)
  );
  INV_X1 _10539_ (
    .A(div_io_resp_bits_tag[3]),
    .ZN(_03074_)
  );
  INV_X1 _10540_ (
    .A(io_dmem_resp_bits_tag[4]),
    .ZN(_03075_)
  );
  INV_X1 _10541_ (
    .A(wb_reg_xcpt),
    .ZN(_03076_)
  );
  INV_X1 _10542_ (
    .A(csr_io_status_isa[12]),
    .ZN(_03077_)
  );
  INV_X1 _10543_ (
    .A(csr_io_status_isa[0]),
    .ZN(_03078_)
  );
  INV_X1 _10544_ (
    .A(csr_io_status_isa[2]),
    .ZN(_03079_)
  );
  INV_X1 _10545_ (
    .A(io_dmem_ordered),
    .ZN(_03080_)
  );
  INV_X1 _10546_ (
    .A(io_dmem_resp_valid),
    .ZN(_03081_)
  );
  INV_X1 _10547_ (
    .A(io_dmem_resp_bits_tag[0]),
    .ZN(_03082_)
  );
  INV_X1 _10548_ (
    .A(io_dmem_perf_grant),
    .ZN(_03083_)
  );
  INV_X1 _10549_ (
    .A(div_io_req_ready),
    .ZN(_03084_)
  );
  INV_X1 _10550_ (
    .A(io_dmem_req_ready),
    .ZN(_03085_)
  );
  INV_X1 _10551_ (
    .A(io_dmem_s2_nack),
    .ZN(_03086_)
  );
  INV_X1 _10552_ (
    .A(wb_reg_replay),
    .ZN(_03087_)
  );
  INV_X1 _10553_ (
    .A(wb_reg_valid),
    .ZN(_03088_)
  );
  INV_X1 _10554_ (
    .A(io_dmem_s2_xcpt_ae_ld),
    .ZN(_03089_)
  );
  INV_X1 _10555_ (
    .A(csr_io_eret),
    .ZN(_03090_)
  );
  INV_X1 _10556_ (
    .A(_take_pc_mem_T),
    .ZN(_03091_)
  );
  INV_X1 _10557_ (
    .A(_00028_),
    .ZN(_03092_)
  );
  INV_X1 _10558_ (
    .A(div_io_resp_valid),
    .ZN(_03093_)
  );
  INV_X1 _10559_ (
    .A(mem_reg_xcpt_interrupt),
    .ZN(_03094_)
  );
  INV_X1 _10560_ (
    .A(csr_io_inhibit_cycle),
    .ZN(_03095_)
  );
  AND2_X1 _10561_ (
    .A1(io_dmem_resp_valid),
    .A2(io_dmem_resp_bits_has_data),
    .ZN(_03096_)
  );
  AND2_X1 _10562_ (
    .A1(_03082_),
    .A2(_03096_),
    .ZN(_03097_)
  );
  AND2_X1 _10563_ (
    .A1(io_dmem_resp_bits_replay),
    .A2(_03097_),
    .ZN(_03098_)
  );
  INV_X1 _10564_ (
    .A(_03098_),
    .ZN(_03099_)
  );
  MUX2_X1 _10565_ (
    .A(_03068_),
    .B(_03069_),
    .S(_03098_),
    .Z(_03100_)
  );
  MUX2_X1 _10566_ (
    .A(div_io_resp_bits_tag[0]),
    .B(io_dmem_resp_bits_tag[1]),
    .S(_03098_),
    .Z(_03101_)
  );
  MUX2_X1 _10567_ (
    .A(_03070_),
    .B(_03071_),
    .S(_03098_),
    .Z(_03102_)
  );
  MUX2_X1 _10568_ (
    .A(div_io_resp_bits_tag[1]),
    .B(io_dmem_resp_bits_tag[2]),
    .S(_03098_),
    .Z(_03103_)
  );
  OR2_X1 _10569_ (
    .A1(_03100_),
    .A2(_03103_),
    .ZN(_03104_)
  );
  MUX2_X1 _10570_ (
    .A(_03072_),
    .B(_03073_),
    .S(_03098_),
    .Z(_03105_)
  );
  MUX2_X1 _10571_ (
    .A(div_io_resp_bits_tag[2]),
    .B(io_dmem_resp_bits_tag[3]),
    .S(_03098_),
    .Z(_03106_)
  );
  OR2_X1 _10572_ (
    .A1(_03104_),
    .A2(_03106_),
    .ZN(_03107_)
  );
  MUX2_X1 _10573_ (
    .A(_03074_),
    .B(_03075_),
    .S(_03098_),
    .Z(_03108_)
  );
  MUX2_X1 _10574_ (
    .A(div_io_resp_bits_tag[3]),
    .B(io_dmem_resp_bits_tag[4]),
    .S(_03098_),
    .Z(_03109_)
  );
  MUX2_X1 _10575_ (
    .A(div_io_resp_bits_tag[4]),
    .B(io_dmem_resp_bits_tag[5]),
    .S(_03098_),
    .Z(_03110_)
  );
  INV_X1 _10576_ (
    .A(_03110_),
    .ZN(_03111_)
  );
  AND2_X1 _10577_ (
    .A1(wb_ctrl_wxd),
    .A2(wb_reg_valid),
    .ZN(_03112_)
  );
  OR2_X1 _10578_ (
    .A1(_03025_),
    .A2(_03088_),
    .ZN(_03113_)
  );
  OR2_X1 _10579_ (
    .A1(_03093_),
    .A2(_03112_),
    .ZN(_03114_)
  );
  INV_X1 _10580_ (
    .A(_03114_),
    .ZN(_03115_)
  );
  AND2_X1 _10581_ (
    .A1(_03099_),
    .A2(_03114_),
    .ZN(_03116_)
  );
  OR2_X1 _10582_ (
    .A1(_03098_),
    .A2(_03115_),
    .ZN(_03117_)
  );
  OR2_X1 _10583_ (
    .A1(_03110_),
    .A2(_03116_),
    .ZN(_03118_)
  );
  OR2_X1 _10584_ (
    .A1(_03109_),
    .A2(_03118_),
    .ZN(_03119_)
  );
  OR2_X1 _10585_ (
    .A1(_03107_),
    .A2(_03119_),
    .ZN(_03120_)
  );
  AND2_X1 _10586_ (
    .A1(_r[1]),
    .A2(_03120_),
    .ZN(_03121_)
  );
  AND2_X1 _10587_ (
    .A1(wb_reg_inst[7]),
    .A2(_03026_),
    .ZN(_03122_)
  );
  AND2_X1 _10588_ (
    .A1(_03027_),
    .A2(_03122_),
    .ZN(_03123_)
  );
  AND2_X1 _10589_ (
    .A1(_03028_),
    .A2(_03123_),
    .ZN(_03124_)
  );
  AND2_X1 _10590_ (
    .A1(wb_ctrl_mem),
    .A2(_03081_),
    .ZN(_03125_)
  );
  OR2_X1 _10591_ (
    .A1(wb_ctrl_div),
    .A2(_03125_),
    .ZN(_03126_)
  );
  AND2_X1 _10592_ (
    .A1(wb_ctrl_mem),
    .A2(wb_reg_valid),
    .ZN(_03127_)
  );
  AND2_X1 _10593_ (
    .A1(io_dmem_s2_xcpt_pf_st),
    .A2(_03127_),
    .ZN(_03128_)
  );
  AND2_X1 _10594_ (
    .A1(io_dmem_s2_xcpt_pf_ld),
    .A2(_03127_),
    .ZN(_03129_)
  );
  OR2_X1 _10595_ (
    .A1(wb_reg_xcpt),
    .A2(_03129_),
    .ZN(_03130_)
  );
  INV_X1 _10596_ (
    .A(_03130_),
    .ZN(_03131_)
  );
  OR2_X1 _10597_ (
    .A1(_03128_),
    .A2(_03130_),
    .ZN(_03132_)
  );
  AND2_X1 _10598_ (
    .A1(io_dmem_s2_xcpt_ae_ld),
    .A2(_03127_),
    .ZN(_03133_)
  );
  AND2_X1 _10599_ (
    .A1(io_dmem_s2_xcpt_ae_st),
    .A2(_03127_),
    .ZN(_03134_)
  );
  OR2_X1 _10600_ (
    .A1(_03133_),
    .A2(_03134_),
    .ZN(_03135_)
  );
  OR2_X1 _10601_ (
    .A1(_03132_),
    .A2(_03135_),
    .ZN(_03136_)
  );
  AND2_X1 _10602_ (
    .A1(io_dmem_s2_xcpt_ma_ld),
    .A2(_03127_),
    .ZN(_03137_)
  );
  AND2_X1 _10603_ (
    .A1(io_dmem_s2_xcpt_ma_st),
    .A2(_03127_),
    .ZN(_03138_)
  );
  OR2_X1 _10604_ (
    .A1(_03137_),
    .A2(_03138_),
    .ZN(_03139_)
  );
  OR2_X1 _10605_ (
    .A1(_03136_),
    .A2(_03139_),
    .ZN(csr_io_exception)
  );
  INV_X1 _10606_ (
    .A(csr_io_exception),
    .ZN(_03140_)
  );
  AND2_X1 _10607_ (
    .A1(_03086_),
    .A2(_03087_),
    .ZN(_03141_)
  );
  OR2_X1 _10608_ (
    .A1(io_dmem_s2_nack),
    .A2(wb_reg_replay),
    .ZN(_03142_)
  );
  AND2_X1 _10609_ (
    .A1(wb_reg_valid),
    .A2(_03141_),
    .ZN(_03143_)
  );
  AND2_X1 _10610_ (
    .A1(_03140_),
    .A2(_03143_),
    .ZN(csr_io_retire)
  );
  AND2_X1 _10611_ (
    .A1(wb_ctrl_wxd),
    .A2(csr_io_retire),
    .ZN(_03144_)
  );
  AND2_X1 _10612_ (
    .A1(_03126_),
    .A2(_03144_),
    .ZN(_03145_)
  );
  AND2_X1 _10613_ (
    .A1(_03029_),
    .A2(_03145_),
    .ZN(_03146_)
  );
  AND2_X1 _10614_ (
    .A1(_03124_),
    .A2(_03146_),
    .ZN(_03147_)
  );
  OR2_X1 _10615_ (
    .A1(_03121_),
    .A2(_03147_),
    .ZN(_03148_)
  );
  AND2_X1 _10616_ (
    .A1(_02979_),
    .A2(_03148_),
    .ZN(_00036_)
  );
  OR2_X1 _10617_ (
    .A1(_03101_),
    .A2(_03102_),
    .ZN(_03149_)
  );
  OR2_X1 _10618_ (
    .A1(_03106_),
    .A2(_03149_),
    .ZN(_03150_)
  );
  OR2_X1 _10619_ (
    .A1(_03119_),
    .A2(_03150_),
    .ZN(_03151_)
  );
  AND2_X1 _10620_ (
    .A1(_r[2]),
    .A2(_03151_),
    .ZN(_03152_)
  );
  AND2_X1 _10621_ (
    .A1(wb_reg_inst[8]),
    .A2(_00029_),
    .ZN(_03153_)
  );
  AND2_X1 _10622_ (
    .A1(_03027_),
    .A2(_03153_),
    .ZN(_03154_)
  );
  AND2_X1 _10623_ (
    .A1(_03028_),
    .A2(_03154_),
    .ZN(_03155_)
  );
  AND2_X1 _10624_ (
    .A1(_03146_),
    .A2(_03155_),
    .ZN(_03156_)
  );
  OR2_X1 _10625_ (
    .A1(_03152_),
    .A2(_03156_),
    .ZN(_03157_)
  );
  AND2_X1 _10626_ (
    .A1(_02979_),
    .A2(_03157_),
    .ZN(_00037_)
  );
  OR2_X1 _10627_ (
    .A1(_03100_),
    .A2(_03102_),
    .ZN(_03158_)
  );
  OR2_X1 _10628_ (
    .A1(_03106_),
    .A2(_03158_),
    .ZN(_03159_)
  );
  OR2_X1 _10629_ (
    .A1(_03119_),
    .A2(_03159_),
    .ZN(_03160_)
  );
  AND2_X1 _10630_ (
    .A1(_r[3]),
    .A2(_03160_),
    .ZN(_03161_)
  );
  AND2_X1 _10631_ (
    .A1(wb_reg_inst[7]),
    .A2(wb_reg_inst[8]),
    .ZN(_03162_)
  );
  AND2_X1 _10632_ (
    .A1(_03027_),
    .A2(_03162_),
    .ZN(_03163_)
  );
  AND2_X1 _10633_ (
    .A1(_03028_),
    .A2(_03163_),
    .ZN(_03164_)
  );
  AND2_X1 _10634_ (
    .A1(_03146_),
    .A2(_03164_),
    .ZN(_03165_)
  );
  OR2_X1 _10635_ (
    .A1(_03161_),
    .A2(_03165_),
    .ZN(_03166_)
  );
  AND2_X1 _10636_ (
    .A1(_02979_),
    .A2(_03166_),
    .ZN(_00038_)
  );
  OR2_X1 _10637_ (
    .A1(_03101_),
    .A2(_03103_),
    .ZN(_03167_)
  );
  OR2_X1 _10638_ (
    .A1(_03105_),
    .A2(_03167_),
    .ZN(_03168_)
  );
  OR2_X1 _10639_ (
    .A1(_03119_),
    .A2(_03168_),
    .ZN(_03169_)
  );
  AND2_X1 _10640_ (
    .A1(_r[4]),
    .A2(_03169_),
    .ZN(_03170_)
  );
  AND2_X1 _10641_ (
    .A1(_03026_),
    .A2(_00029_),
    .ZN(_03171_)
  );
  AND2_X1 _10642_ (
    .A1(wb_reg_inst[9]),
    .A2(_03171_),
    .ZN(_03172_)
  );
  AND2_X1 _10643_ (
    .A1(_03028_),
    .A2(_03172_),
    .ZN(_03173_)
  );
  AND2_X1 _10644_ (
    .A1(_03146_),
    .A2(_03173_),
    .ZN(_03174_)
  );
  OR2_X1 _10645_ (
    .A1(_03170_),
    .A2(_03174_),
    .ZN(_03175_)
  );
  AND2_X1 _10646_ (
    .A1(_02979_),
    .A2(_03175_),
    .ZN(_00039_)
  );
  OR2_X1 _10647_ (
    .A1(_03104_),
    .A2(_03105_),
    .ZN(_03176_)
  );
  OR2_X1 _10648_ (
    .A1(_03119_),
    .A2(_03176_),
    .ZN(_03177_)
  );
  AND2_X1 _10649_ (
    .A1(_r[5]),
    .A2(_03177_),
    .ZN(_03178_)
  );
  AND2_X1 _10650_ (
    .A1(wb_reg_inst[9]),
    .A2(_03122_),
    .ZN(_03179_)
  );
  AND2_X1 _10651_ (
    .A1(_03028_),
    .A2(_03179_),
    .ZN(_03180_)
  );
  AND2_X1 _10652_ (
    .A1(_03146_),
    .A2(_03180_),
    .ZN(_03181_)
  );
  OR2_X1 _10653_ (
    .A1(_03178_),
    .A2(_03181_),
    .ZN(_03182_)
  );
  AND2_X1 _10654_ (
    .A1(_02979_),
    .A2(_03182_),
    .ZN(_00040_)
  );
  OR2_X1 _10655_ (
    .A1(_03105_),
    .A2(_03149_),
    .ZN(_03183_)
  );
  OR2_X1 _10656_ (
    .A1(_03119_),
    .A2(_03183_),
    .ZN(_03184_)
  );
  AND2_X1 _10657_ (
    .A1(_r[6]),
    .A2(_03184_),
    .ZN(_03185_)
  );
  AND2_X1 _10658_ (
    .A1(wb_reg_inst[9]),
    .A2(_03153_),
    .ZN(_03186_)
  );
  AND2_X1 _10659_ (
    .A1(_03028_),
    .A2(_03186_),
    .ZN(_03187_)
  );
  AND2_X1 _10660_ (
    .A1(_03146_),
    .A2(_03187_),
    .ZN(_03188_)
  );
  OR2_X1 _10661_ (
    .A1(_03185_),
    .A2(_03188_),
    .ZN(_03189_)
  );
  AND2_X1 _10662_ (
    .A1(_02979_),
    .A2(_03189_),
    .ZN(_00041_)
  );
  OR2_X1 _10663_ (
    .A1(_03105_),
    .A2(_03158_),
    .ZN(_03190_)
  );
  OR2_X1 _10664_ (
    .A1(_03119_),
    .A2(_03190_),
    .ZN(_03191_)
  );
  AND2_X1 _10665_ (
    .A1(_r[7]),
    .A2(_03191_),
    .ZN(_03192_)
  );
  AND2_X1 _10666_ (
    .A1(wb_reg_inst[9]),
    .A2(_03162_),
    .ZN(_03193_)
  );
  AND2_X1 _10667_ (
    .A1(_03028_),
    .A2(_03193_),
    .ZN(_03194_)
  );
  AND2_X1 _10668_ (
    .A1(_03146_),
    .A2(_03194_),
    .ZN(_03195_)
  );
  OR2_X1 _10669_ (
    .A1(_03192_),
    .A2(_03195_),
    .ZN(_03196_)
  );
  AND2_X1 _10670_ (
    .A1(_02979_),
    .A2(_03196_),
    .ZN(_00042_)
  );
  OR2_X1 _10671_ (
    .A1(_03106_),
    .A2(_03167_),
    .ZN(_03197_)
  );
  OR2_X1 _10672_ (
    .A1(_03108_),
    .A2(_03197_),
    .ZN(_03198_)
  );
  OR2_X1 _10673_ (
    .A1(_03118_),
    .A2(_03198_),
    .ZN(_03199_)
  );
  AND2_X1 _10674_ (
    .A1(_r[8]),
    .A2(_03199_),
    .ZN(_03200_)
  );
  AND2_X1 _10675_ (
    .A1(_03027_),
    .A2(_03171_),
    .ZN(_03201_)
  );
  AND2_X1 _10676_ (
    .A1(wb_reg_inst[10]),
    .A2(_03145_),
    .ZN(_03202_)
  );
  AND2_X1 _10677_ (
    .A1(_03201_),
    .A2(_03202_),
    .ZN(_03203_)
  );
  AND2_X1 _10678_ (
    .A1(_03029_),
    .A2(_03203_),
    .ZN(_03204_)
  );
  OR2_X1 _10679_ (
    .A1(_03200_),
    .A2(_03204_),
    .ZN(_03205_)
  );
  AND2_X1 _10680_ (
    .A1(_02979_),
    .A2(_03205_),
    .ZN(_00043_)
  );
  OR2_X1 _10681_ (
    .A1(_03107_),
    .A2(_03108_),
    .ZN(_03206_)
  );
  OR2_X1 _10682_ (
    .A1(_03118_),
    .A2(_03206_),
    .ZN(_03207_)
  );
  AND2_X1 _10683_ (
    .A1(_r[9]),
    .A2(_03207_),
    .ZN(_03208_)
  );
  AND2_X1 _10684_ (
    .A1(_03123_),
    .A2(_03202_),
    .ZN(_03209_)
  );
  AND2_X1 _10685_ (
    .A1(_03029_),
    .A2(_03209_),
    .ZN(_03210_)
  );
  OR2_X1 _10686_ (
    .A1(_03208_),
    .A2(_03210_),
    .ZN(_03211_)
  );
  AND2_X1 _10687_ (
    .A1(_02979_),
    .A2(_03211_),
    .ZN(_00044_)
  );
  OR2_X1 _10688_ (
    .A1(_03108_),
    .A2(_03150_),
    .ZN(_03212_)
  );
  OR2_X1 _10689_ (
    .A1(_03118_),
    .A2(_03212_),
    .ZN(_03213_)
  );
  AND2_X1 _10690_ (
    .A1(_r[10]),
    .A2(_03213_),
    .ZN(_03214_)
  );
  AND2_X1 _10691_ (
    .A1(_03154_),
    .A2(_03202_),
    .ZN(_03215_)
  );
  AND2_X1 _10692_ (
    .A1(_03029_),
    .A2(_03215_),
    .ZN(_03216_)
  );
  OR2_X1 _10693_ (
    .A1(_03214_),
    .A2(_03216_),
    .ZN(_03217_)
  );
  AND2_X1 _10694_ (
    .A1(_02979_),
    .A2(_03217_),
    .ZN(_00045_)
  );
  OR2_X1 _10695_ (
    .A1(_03108_),
    .A2(_03159_),
    .ZN(_03218_)
  );
  OR2_X1 _10696_ (
    .A1(_03118_),
    .A2(_03218_),
    .ZN(_03219_)
  );
  AND2_X1 _10697_ (
    .A1(_r[11]),
    .A2(_03219_),
    .ZN(_03220_)
  );
  AND2_X1 _10698_ (
    .A1(_03163_),
    .A2(_03202_),
    .ZN(_03221_)
  );
  AND2_X1 _10699_ (
    .A1(_03029_),
    .A2(_03221_),
    .ZN(_03222_)
  );
  OR2_X1 _10700_ (
    .A1(_03220_),
    .A2(_03222_),
    .ZN(_03223_)
  );
  AND2_X1 _10701_ (
    .A1(_02979_),
    .A2(_03223_),
    .ZN(_00046_)
  );
  OR2_X1 _10702_ (
    .A1(_03108_),
    .A2(_03168_),
    .ZN(_03224_)
  );
  OR2_X1 _10703_ (
    .A1(_03118_),
    .A2(_03224_),
    .ZN(_03225_)
  );
  AND2_X1 _10704_ (
    .A1(_r[12]),
    .A2(_03225_),
    .ZN(_03226_)
  );
  AND2_X1 _10705_ (
    .A1(_03172_),
    .A2(_03202_),
    .ZN(_03227_)
  );
  AND2_X1 _10706_ (
    .A1(_03029_),
    .A2(_03227_),
    .ZN(_03228_)
  );
  OR2_X1 _10707_ (
    .A1(_03226_),
    .A2(_03228_),
    .ZN(_03229_)
  );
  AND2_X1 _10708_ (
    .A1(_02979_),
    .A2(_03229_),
    .ZN(_00047_)
  );
  OR2_X1 _10709_ (
    .A1(_03108_),
    .A2(_03176_),
    .ZN(_03230_)
  );
  OR2_X1 _10710_ (
    .A1(_03118_),
    .A2(_03230_),
    .ZN(_03231_)
  );
  AND2_X1 _10711_ (
    .A1(_r[13]),
    .A2(_03231_),
    .ZN(_03232_)
  );
  AND2_X1 _10712_ (
    .A1(_03179_),
    .A2(_03202_),
    .ZN(_03233_)
  );
  AND2_X1 _10713_ (
    .A1(_03029_),
    .A2(_03233_),
    .ZN(_03234_)
  );
  OR2_X1 _10714_ (
    .A1(_03232_),
    .A2(_03234_),
    .ZN(_03235_)
  );
  AND2_X1 _10715_ (
    .A1(_02979_),
    .A2(_03235_),
    .ZN(_00048_)
  );
  OR2_X1 _10716_ (
    .A1(_03108_),
    .A2(_03183_),
    .ZN(_03236_)
  );
  OR2_X1 _10717_ (
    .A1(_03118_),
    .A2(_03236_),
    .ZN(_03237_)
  );
  AND2_X1 _10718_ (
    .A1(_r[14]),
    .A2(_03237_),
    .ZN(_03238_)
  );
  AND2_X1 _10719_ (
    .A1(_03186_),
    .A2(_03202_),
    .ZN(_03239_)
  );
  AND2_X1 _10720_ (
    .A1(_03029_),
    .A2(_03239_),
    .ZN(_03240_)
  );
  OR2_X1 _10721_ (
    .A1(_03238_),
    .A2(_03240_),
    .ZN(_03241_)
  );
  AND2_X1 _10722_ (
    .A1(_02979_),
    .A2(_03241_),
    .ZN(_00049_)
  );
  OR2_X1 _10723_ (
    .A1(_03108_),
    .A2(_03190_),
    .ZN(_03242_)
  );
  OR2_X1 _10724_ (
    .A1(_03118_),
    .A2(_03242_),
    .ZN(_03243_)
  );
  AND2_X1 _10725_ (
    .A1(_r[15]),
    .A2(_03243_),
    .ZN(_03244_)
  );
  AND2_X1 _10726_ (
    .A1(_03193_),
    .A2(_03202_),
    .ZN(_03245_)
  );
  AND2_X1 _10727_ (
    .A1(_03029_),
    .A2(_03245_),
    .ZN(_03246_)
  );
  OR2_X1 _10728_ (
    .A1(_03244_),
    .A2(_03246_),
    .ZN(_03247_)
  );
  AND2_X1 _10729_ (
    .A1(_02979_),
    .A2(_03247_),
    .ZN(_00050_)
  );
  OR2_X1 _10730_ (
    .A1(_03111_),
    .A2(_03116_),
    .ZN(_03248_)
  );
  OR2_X1 _10731_ (
    .A1(_03109_),
    .A2(_03248_),
    .ZN(_03249_)
  );
  OR2_X1 _10732_ (
    .A1(_03197_),
    .A2(_03249_),
    .ZN(_03250_)
  );
  AND2_X1 _10733_ (
    .A1(_r[16]),
    .A2(_03250_),
    .ZN(_03251_)
  );
  AND2_X1 _10734_ (
    .A1(wb_reg_inst[11]),
    .A2(_03145_),
    .ZN(_03252_)
  );
  AND2_X1 _10735_ (
    .A1(_03201_),
    .A2(_03252_),
    .ZN(_03253_)
  );
  AND2_X1 _10736_ (
    .A1(_03028_),
    .A2(_03253_),
    .ZN(_03254_)
  );
  OR2_X1 _10737_ (
    .A1(_03251_),
    .A2(_03254_),
    .ZN(_03255_)
  );
  AND2_X1 _10738_ (
    .A1(_02979_),
    .A2(_03255_),
    .ZN(_00051_)
  );
  OR2_X1 _10739_ (
    .A1(_03107_),
    .A2(_03249_),
    .ZN(_03256_)
  );
  AND2_X1 _10740_ (
    .A1(_r[17]),
    .A2(_03256_),
    .ZN(_03257_)
  );
  AND2_X1 _10741_ (
    .A1(_03124_),
    .A2(_03252_),
    .ZN(_03258_)
  );
  OR2_X1 _10742_ (
    .A1(_03257_),
    .A2(_03258_),
    .ZN(_03259_)
  );
  AND2_X1 _10743_ (
    .A1(_02979_),
    .A2(_03259_),
    .ZN(_00052_)
  );
  OR2_X1 _10744_ (
    .A1(_03150_),
    .A2(_03249_),
    .ZN(_03260_)
  );
  AND2_X1 _10745_ (
    .A1(_r[18]),
    .A2(_03260_),
    .ZN(_03261_)
  );
  AND2_X1 _10746_ (
    .A1(_03155_),
    .A2(_03252_),
    .ZN(_03262_)
  );
  OR2_X1 _10747_ (
    .A1(_03261_),
    .A2(_03262_),
    .ZN(_03263_)
  );
  AND2_X1 _10748_ (
    .A1(_02979_),
    .A2(_03263_),
    .ZN(_00053_)
  );
  OR2_X1 _10749_ (
    .A1(_03159_),
    .A2(_03249_),
    .ZN(_03264_)
  );
  AND2_X1 _10750_ (
    .A1(_r[19]),
    .A2(_03264_),
    .ZN(_03265_)
  );
  AND2_X1 _10751_ (
    .A1(_03164_),
    .A2(_03252_),
    .ZN(_03266_)
  );
  OR2_X1 _10752_ (
    .A1(_03265_),
    .A2(_03266_),
    .ZN(_03267_)
  );
  AND2_X1 _10753_ (
    .A1(_02979_),
    .A2(_03267_),
    .ZN(_00054_)
  );
  OR2_X1 _10754_ (
    .A1(_03168_),
    .A2(_03249_),
    .ZN(_03268_)
  );
  AND2_X1 _10755_ (
    .A1(_r[20]),
    .A2(_03268_),
    .ZN(_03269_)
  );
  AND2_X1 _10756_ (
    .A1(_03173_),
    .A2(_03252_),
    .ZN(_03270_)
  );
  OR2_X1 _10757_ (
    .A1(_03269_),
    .A2(_03270_),
    .ZN(_03271_)
  );
  AND2_X1 _10758_ (
    .A1(_02979_),
    .A2(_03271_),
    .ZN(_00055_)
  );
  OR2_X1 _10759_ (
    .A1(_03176_),
    .A2(_03249_),
    .ZN(_03272_)
  );
  AND2_X1 _10760_ (
    .A1(_r[21]),
    .A2(_03272_),
    .ZN(_03273_)
  );
  AND2_X1 _10761_ (
    .A1(_03180_),
    .A2(_03252_),
    .ZN(_03274_)
  );
  OR2_X1 _10762_ (
    .A1(_03273_),
    .A2(_03274_),
    .ZN(_03275_)
  );
  AND2_X1 _10763_ (
    .A1(_02979_),
    .A2(_03275_),
    .ZN(_00056_)
  );
  OR2_X1 _10764_ (
    .A1(_03183_),
    .A2(_03249_),
    .ZN(_03276_)
  );
  AND2_X1 _10765_ (
    .A1(_r[22]),
    .A2(_03276_),
    .ZN(_03277_)
  );
  AND2_X1 _10766_ (
    .A1(_03187_),
    .A2(_03252_),
    .ZN(_03278_)
  );
  OR2_X1 _10767_ (
    .A1(_03277_),
    .A2(_03278_),
    .ZN(_03279_)
  );
  AND2_X1 _10768_ (
    .A1(_02979_),
    .A2(_03279_),
    .ZN(_00057_)
  );
  OR2_X1 _10769_ (
    .A1(_03190_),
    .A2(_03249_),
    .ZN(_03280_)
  );
  AND2_X1 _10770_ (
    .A1(_r[23]),
    .A2(_03280_),
    .ZN(_03281_)
  );
  AND2_X1 _10771_ (
    .A1(_03194_),
    .A2(_03252_),
    .ZN(_03282_)
  );
  OR2_X1 _10772_ (
    .A1(_03281_),
    .A2(_03282_),
    .ZN(_03283_)
  );
  AND2_X1 _10773_ (
    .A1(_02979_),
    .A2(_03283_),
    .ZN(_00058_)
  );
  OR2_X1 _10774_ (
    .A1(_03198_),
    .A2(_03248_),
    .ZN(_03284_)
  );
  AND2_X1 _10775_ (
    .A1(_r[24]),
    .A2(_03284_),
    .ZN(_03285_)
  );
  AND2_X1 _10776_ (
    .A1(wb_reg_inst[10]),
    .A2(_03253_),
    .ZN(_03286_)
  );
  OR2_X1 _10777_ (
    .A1(_03285_),
    .A2(_03286_),
    .ZN(_03287_)
  );
  AND2_X1 _10778_ (
    .A1(_02979_),
    .A2(_03287_),
    .ZN(_00059_)
  );
  OR2_X1 _10779_ (
    .A1(_03206_),
    .A2(_03248_),
    .ZN(_03288_)
  );
  AND2_X1 _10780_ (
    .A1(_r[25]),
    .A2(_03288_),
    .ZN(_03289_)
  );
  AND2_X1 _10781_ (
    .A1(wb_reg_inst[11]),
    .A2(_03209_),
    .ZN(_03290_)
  );
  OR2_X1 _10782_ (
    .A1(_03289_),
    .A2(_03290_),
    .ZN(_03291_)
  );
  AND2_X1 _10783_ (
    .A1(_02979_),
    .A2(_03291_),
    .ZN(_00060_)
  );
  OR2_X1 _10784_ (
    .A1(_03212_),
    .A2(_03248_),
    .ZN(_03292_)
  );
  AND2_X1 _10785_ (
    .A1(_r[26]),
    .A2(_03292_),
    .ZN(_03293_)
  );
  AND2_X1 _10786_ (
    .A1(wb_reg_inst[11]),
    .A2(_03215_),
    .ZN(_03294_)
  );
  OR2_X1 _10787_ (
    .A1(_03293_),
    .A2(_03294_),
    .ZN(_03295_)
  );
  AND2_X1 _10788_ (
    .A1(_02979_),
    .A2(_03295_),
    .ZN(_00061_)
  );
  OR2_X1 _10789_ (
    .A1(_03218_),
    .A2(_03248_),
    .ZN(_03296_)
  );
  AND2_X1 _10790_ (
    .A1(_r[27]),
    .A2(_03296_),
    .ZN(_03297_)
  );
  AND2_X1 _10791_ (
    .A1(wb_reg_inst[11]),
    .A2(_03221_),
    .ZN(_03298_)
  );
  OR2_X1 _10792_ (
    .A1(_03297_),
    .A2(_03298_),
    .ZN(_03299_)
  );
  AND2_X1 _10793_ (
    .A1(_02979_),
    .A2(_03299_),
    .ZN(_00062_)
  );
  OR2_X1 _10794_ (
    .A1(_03224_),
    .A2(_03248_),
    .ZN(_03300_)
  );
  AND2_X1 _10795_ (
    .A1(_r[28]),
    .A2(_03300_),
    .ZN(_03301_)
  );
  AND2_X1 _10796_ (
    .A1(wb_reg_inst[11]),
    .A2(_03227_),
    .ZN(_03302_)
  );
  OR2_X1 _10797_ (
    .A1(_03301_),
    .A2(_03302_),
    .ZN(_03303_)
  );
  AND2_X1 _10798_ (
    .A1(_02979_),
    .A2(_03303_),
    .ZN(_00063_)
  );
  OR2_X1 _10799_ (
    .A1(_03230_),
    .A2(_03248_),
    .ZN(_03304_)
  );
  AND2_X1 _10800_ (
    .A1(_r[29]),
    .A2(_03304_),
    .ZN(_03305_)
  );
  AND2_X1 _10801_ (
    .A1(wb_reg_inst[11]),
    .A2(_03233_),
    .ZN(_03306_)
  );
  OR2_X1 _10802_ (
    .A1(_03305_),
    .A2(_03306_),
    .ZN(_03307_)
  );
  AND2_X1 _10803_ (
    .A1(_02979_),
    .A2(_03307_),
    .ZN(_00064_)
  );
  OR2_X1 _10804_ (
    .A1(_03236_),
    .A2(_03248_),
    .ZN(_03308_)
  );
  AND2_X1 _10805_ (
    .A1(_r[30]),
    .A2(_03308_),
    .ZN(_03309_)
  );
  AND2_X1 _10806_ (
    .A1(wb_reg_inst[11]),
    .A2(_03239_),
    .ZN(_03310_)
  );
  OR2_X1 _10807_ (
    .A1(_03309_),
    .A2(_03310_),
    .ZN(_03311_)
  );
  AND2_X1 _10808_ (
    .A1(_02979_),
    .A2(_03311_),
    .ZN(_00065_)
  );
  OR2_X1 _10809_ (
    .A1(_03242_),
    .A2(_03248_),
    .ZN(_03312_)
  );
  AND2_X1 _10810_ (
    .A1(_r[31]),
    .A2(_03312_),
    .ZN(_03313_)
  );
  AND2_X1 _10811_ (
    .A1(wb_reg_inst[11]),
    .A2(_03245_),
    .ZN(_03314_)
  );
  OR2_X1 _10812_ (
    .A1(_03313_),
    .A2(_03314_),
    .ZN(_03315_)
  );
  AND2_X1 _10813_ (
    .A1(_02979_),
    .A2(_03315_),
    .ZN(_00066_)
  );
  AND2_X1 _10814_ (
    .A1(csr_io_decode_0_inst[1]),
    .A2(_03037_),
    .ZN(_03316_)
  );
  AND2_X1 _10815_ (
    .A1(_03040_),
    .A2(_03316_),
    .ZN(_03317_)
  );
  AND2_X1 _10816_ (
    .A1(csr_io_decode_0_inst[0]),
    .A2(csr_io_decode_0_inst[1]),
    .ZN(_03318_)
  );
  AND2_X1 _10817_ (
    .A1(csr_io_decode_0_inst[0]),
    .A2(_03317_),
    .ZN(_03319_)
  );
  AND2_X1 _10818_ (
    .A1(_03036_),
    .A2(_03319_),
    .ZN(_03320_)
  );
  AND2_X1 _10819_ (
    .A1(_03038_),
    .A2(_03320_),
    .ZN(_03321_)
  );
  AND2_X1 _10820_ (
    .A1(_03000_),
    .A2(_03001_),
    .ZN(_03322_)
  );
  OR2_X1 _10821_ (
    .A1(csr_io_decode_0_inst[12]),
    .A2(csr_io_decode_0_inst[13]),
    .ZN(_03323_)
  );
  AND2_X1 _10822_ (
    .A1(_03321_),
    .A2(_03322_),
    .ZN(_03324_)
  );
  AND2_X1 _10823_ (
    .A1(_03001_),
    .A2(_03039_),
    .ZN(_03325_)
  );
  OR2_X1 _10824_ (
    .A1(csr_io_decode_0_inst[13]),
    .A2(csr_io_decode_0_inst[4]),
    .ZN(_03326_)
  );
  AND2_X1 _10825_ (
    .A1(_03001_),
    .A2(_03002_),
    .ZN(_03327_)
  );
  OR2_X1 _10826_ (
    .A1(csr_io_decode_0_inst[13]),
    .A2(csr_io_decode_0_inst[14]),
    .ZN(_03328_)
  );
  OR2_X1 _10827_ (
    .A1(csr_io_decode_0_inst[4]),
    .A2(_03328_),
    .ZN(_03329_)
  );
  AND2_X1 _10828_ (
    .A1(_03000_),
    .A2(_03002_),
    .ZN(_03330_)
  );
  OR2_X1 _10829_ (
    .A1(csr_io_decode_0_inst[12]),
    .A2(csr_io_decode_0_inst[14]),
    .ZN(_03331_)
  );
  OR2_X1 _10830_ (
    .A1(csr_io_decode_0_inst[4]),
    .A2(_03331_),
    .ZN(_03332_)
  );
  INV_X1 _10831_ (
    .A(_03332_),
    .ZN(_03333_)
  );
  OR2_X1 _10832_ (
    .A1(csr_io_decode_0_inst[5]),
    .A2(_03326_),
    .ZN(_03334_)
  );
  INV_X1 _10833_ (
    .A(_03334_),
    .ZN(_03335_)
  );
  AND2_X1 _10834_ (
    .A1(_03332_),
    .A2(_03334_),
    .ZN(_03336_)
  );
  AND2_X1 _10835_ (
    .A1(_03329_),
    .A2(_03336_),
    .ZN(_03337_)
  );
  INV_X1 _10836_ (
    .A(_03337_),
    .ZN(_03338_)
  );
  AND2_X1 _10837_ (
    .A1(_03320_),
    .A2(_03338_),
    .ZN(_03339_)
  );
  OR2_X1 _10838_ (
    .A1(_03324_),
    .A2(_03339_),
    .ZN(_03340_)
  );
  AND2_X1 _10839_ (
    .A1(_03040_),
    .A2(_03318_),
    .ZN(_03341_)
  );
  AND2_X1 _10840_ (
    .A1(csr_io_decode_0_inst[6]),
    .A2(csr_io_decode_0_inst[5]),
    .ZN(_03342_)
  );
  AND2_X1 _10841_ (
    .A1(_03325_),
    .A2(_03342_),
    .ZN(_03343_)
  );
  AND2_X1 _10842_ (
    .A1(_03330_),
    .A2(_03343_),
    .ZN(_03344_)
  );
  AND2_X1 _10843_ (
    .A1(_03341_),
    .A2(_03344_),
    .ZN(_03345_)
  );
  AND2_X1 _10844_ (
    .A1(csr_io_decode_0_inst[0]),
    .A2(csr_io_decode_0_inst[4]),
    .ZN(_03346_)
  );
  AND2_X1 _10845_ (
    .A1(_03317_),
    .A2(_03346_),
    .ZN(_03347_)
  );
  AND2_X1 _10846_ (
    .A1(csr_io_decode_0_inst[12]),
    .A2(_03036_),
    .ZN(_03348_)
  );
  AND2_X1 _10847_ (
    .A1(_03347_),
    .A2(_03348_),
    .ZN(_03349_)
  );
  OR2_X1 _10848_ (
    .A1(csr_io_decode_0_inst[25]),
    .A2(csr_io_decode_0_inst[26]),
    .ZN(_03350_)
  );
  INV_X1 _10849_ (
    .A(_03350_),
    .ZN(_03351_)
  );
  AND2_X1 _10850_ (
    .A1(_03005_),
    .A2(_03006_),
    .ZN(_03352_)
  );
  AND2_X1 _10851_ (
    .A1(_03001_),
    .A2(_03004_),
    .ZN(_03353_)
  );
  AND2_X1 _10852_ (
    .A1(_03352_),
    .A2(_03353_),
    .ZN(_03354_)
  );
  OR2_X1 _10853_ (
    .A1(csr_io_decode_0_inst[30]),
    .A2(csr_io_decode_0_inst[31]),
    .ZN(_03355_)
  );
  INV_X1 _10854_ (
    .A(_03355_),
    .ZN(_03356_)
  );
  AND2_X1 _10855_ (
    .A1(_03008_),
    .A2(_03009_),
    .ZN(_03357_)
  );
  AND2_X1 _10856_ (
    .A1(_03008_),
    .A2(_03356_),
    .ZN(_03358_)
  );
  AND2_X1 _10857_ (
    .A1(_03007_),
    .A2(_03357_),
    .ZN(_03359_)
  );
  AND2_X1 _10858_ (
    .A1(_03007_),
    .A2(_03358_),
    .ZN(_03360_)
  );
  AND2_X1 _10859_ (
    .A1(_03354_),
    .A2(_03360_),
    .ZN(_03361_)
  );
  AND2_X1 _10860_ (
    .A1(_03349_),
    .A2(_03361_),
    .ZN(_03362_)
  );
  OR2_X1 _10861_ (
    .A1(_03345_),
    .A2(_03362_),
    .ZN(_03363_)
  );
  OR2_X1 _10862_ (
    .A1(_03340_),
    .A2(_03363_),
    .ZN(_03364_)
  );
  AND2_X1 _10863_ (
    .A1(_03039_),
    .A2(_03319_),
    .ZN(_03365_)
  );
  AND2_X1 _10864_ (
    .A1(_03342_),
    .A2(_03365_),
    .ZN(_03366_)
  );
  AND2_X1 _10865_ (
    .A1(csr_io_decode_0_inst[14]),
    .A2(_03342_),
    .ZN(_03367_)
  );
  AND2_X1 _10866_ (
    .A1(_03365_),
    .A2(_03367_),
    .ZN(_03368_)
  );
  AND2_X1 _10867_ (
    .A1(csr_io_decode_0_inst[14]),
    .A2(_03354_),
    .ZN(_03369_)
  );
  AND2_X1 _10868_ (
    .A1(_03349_),
    .A2(_03369_),
    .ZN(_03370_)
  );
  AND2_X1 _10869_ (
    .A1(_03359_),
    .A2(_03370_),
    .ZN(_03371_)
  );
  AND2_X1 _10870_ (
    .A1(csr_io_decode_0_inst[14]),
    .A2(_03348_),
    .ZN(_03372_)
  );
  AND2_X1 _10871_ (
    .A1(_03354_),
    .A2(_03372_),
    .ZN(_03373_)
  );
  AND2_X1 _10872_ (
    .A1(_03347_),
    .A2(_03373_),
    .ZN(_03374_)
  );
  AND2_X1 _10873_ (
    .A1(_03359_),
    .A2(_03374_),
    .ZN(_03375_)
  );
  OR2_X1 _10874_ (
    .A1(_03368_),
    .A2(_03375_),
    .ZN(_03376_)
  );
  AND2_X1 _10875_ (
    .A1(csr_io_decode_0_inst[13]),
    .A2(_03036_),
    .ZN(_03377_)
  );
  AND2_X1 _10876_ (
    .A1(_03038_),
    .A2(_03347_),
    .ZN(_03378_)
  );
  AND2_X1 _10877_ (
    .A1(_03377_),
    .A2(_03378_),
    .ZN(_03379_)
  );
  AND2_X1 _10878_ (
    .A1(_03006_),
    .A2(_03007_),
    .ZN(_03380_)
  );
  AND2_X1 _10879_ (
    .A1(csr_io_decode_0_inst[5]),
    .A2(_03333_),
    .ZN(_03381_)
  );
  AND2_X1 _10880_ (
    .A1(csr_io_decode_0_inst[2]),
    .A2(csr_io_decode_0_inst[3]),
    .ZN(_03382_)
  );
  AND2_X1 _10881_ (
    .A1(_03318_),
    .A2(_03382_),
    .ZN(_03383_)
  );
  AND2_X1 _10882_ (
    .A1(_03377_),
    .A2(_03383_),
    .ZN(_03384_)
  );
  AND2_X1 _10883_ (
    .A1(_03381_),
    .A2(_03384_),
    .ZN(_03385_)
  );
  AND2_X1 _10884_ (
    .A1(_03380_),
    .A2(_03385_),
    .ZN(_03386_)
  );
  OR2_X1 _10885_ (
    .A1(_03379_),
    .A2(_03386_),
    .ZN(_03387_)
  );
  AND2_X1 _10886_ (
    .A1(csr_io_decode_0_inst[13]),
    .A2(_03002_),
    .ZN(_03388_)
  );
  INV_X1 _10887_ (
    .A(_03388_),
    .ZN(_03389_)
  );
  AND2_X1 _10888_ (
    .A1(csr_io_decode_0_inst[5]),
    .A2(csr_io_decode_0_inst[4]),
    .ZN(_03390_)
  );
  AND2_X1 _10889_ (
    .A1(_03342_),
    .A2(_03346_),
    .ZN(_03391_)
  );
  AND2_X1 _10890_ (
    .A1(_03317_),
    .A2(_03391_),
    .ZN(_03392_)
  );
  AND2_X1 _10891_ (
    .A1(_03388_),
    .A2(_03392_),
    .ZN(_03393_)
  );
  AND2_X1 _10892_ (
    .A1(csr_io_decode_0_inst[12]),
    .A2(_03342_),
    .ZN(_03394_)
  );
  AND2_X1 _10893_ (
    .A1(_03319_),
    .A2(_03327_),
    .ZN(_03395_)
  );
  AND2_X1 _10894_ (
    .A1(_03394_),
    .A2(_03395_),
    .ZN(_03396_)
  );
  OR2_X1 _10895_ (
    .A1(_03393_),
    .A2(_03396_),
    .ZN(_03397_)
  );
  OR2_X1 _10896_ (
    .A1(_03387_),
    .A2(_03397_),
    .ZN(_03398_)
  );
  AND2_X1 _10897_ (
    .A1(csr_io_decode_0_inst[5]),
    .A2(_03039_),
    .ZN(_03399_)
  );
  AND2_X1 _10898_ (
    .A1(_03383_),
    .A2(_03399_),
    .ZN(_03400_)
  );
  AND2_X1 _10899_ (
    .A1(_03000_),
    .A2(_03036_),
    .ZN(_03401_)
  );
  OR2_X1 _10900_ (
    .A1(csr_io_decode_0_inst[12]),
    .A2(csr_io_decode_0_inst[6]),
    .ZN(_03402_)
  );
  AND2_X1 _10901_ (
    .A1(_03388_),
    .A2(_03401_),
    .ZN(_03403_)
  );
  AND2_X1 _10902_ (
    .A1(_03400_),
    .A2(_03403_),
    .ZN(_03404_)
  );
  AND2_X1 _10903_ (
    .A1(_03380_),
    .A2(_03404_),
    .ZN(_03405_)
  );
  OR2_X1 _10904_ (
    .A1(_03376_),
    .A2(_03398_),
    .ZN(_03406_)
  );
  AND2_X1 _10905_ (
    .A1(_03036_),
    .A2(_03038_),
    .ZN(_03407_)
  );
  AND2_X1 _10906_ (
    .A1(_03319_),
    .A2(_03407_),
    .ZN(_03408_)
  );
  AND2_X1 _10907_ (
    .A1(_03325_),
    .A2(_03408_),
    .ZN(_03409_)
  );
  AND2_X1 _10908_ (
    .A1(_03329_),
    .A2(_03332_),
    .ZN(_03410_)
  );
  INV_X1 _10909_ (
    .A(_03410_),
    .ZN(_03411_)
  );
  AND2_X1 _10910_ (
    .A1(_03320_),
    .A2(_03411_),
    .ZN(_03412_)
  );
  OR2_X1 _10911_ (
    .A1(_03364_),
    .A2(_03406_),
    .ZN(_03413_)
  );
  AND2_X1 _10912_ (
    .A1(csr_io_decode_0_inst[28]),
    .A2(_03358_),
    .ZN(_03414_)
  );
  OR2_X1 _10913_ (
    .A1(csr_io_decode_0_inst[24]),
    .A2(csr_io_decode_0_inst[27]),
    .ZN(_03415_)
  );
  INV_X1 _10914_ (
    .A(_03415_),
    .ZN(_03416_)
  );
  OR2_X1 _10915_ (
    .A1(csr_io_decode_0_inst[21]),
    .A2(csr_io_decode_0_inst[23]),
    .ZN(_03417_)
  );
  OR2_X1 _10916_ (
    .A1(csr_io_decode_0_inst[20]),
    .A2(csr_io_decode_0_inst[22]),
    .ZN(_03418_)
  );
  INV_X1 _10917_ (
    .A(_03418_),
    .ZN(_03419_)
  );
  OR2_X1 _10918_ (
    .A1(_03417_),
    .A2(_03418_),
    .ZN(_03420_)
  );
  INV_X1 _10919_ (
    .A(_03420_),
    .ZN(_03421_)
  );
  AND2_X1 _10920_ (
    .A1(_03416_),
    .A2(_03421_),
    .ZN(_03422_)
  );
  AND2_X1 _10921_ (
    .A1(_03414_),
    .A2(_03422_),
    .ZN(_03423_)
  );
  AND2_X1 _10922_ (
    .A1(_03036_),
    .A2(_03400_),
    .ZN(_03424_)
  );
  AND2_X1 _10923_ (
    .A1(_03423_),
    .A2(_03424_),
    .ZN(_03425_)
  );
  AND2_X1 _10924_ (
    .A1(csr_io_decode_0_inst[27]),
    .A2(_03385_),
    .ZN(_03426_)
  );
  AND2_X1 _10925_ (
    .A1(_03358_),
    .A2(_03426_),
    .ZN(_03427_)
  );
  OR2_X1 _10926_ (
    .A1(_03425_),
    .A2(_03427_),
    .ZN(_03428_)
  );
  AND2_X1 _10927_ (
    .A1(_03352_),
    .A2(_03360_),
    .ZN(_03429_)
  );
  AND2_X1 _10928_ (
    .A1(csr_io_decode_0_inst[5]),
    .A2(_03347_),
    .ZN(_03430_)
  );
  AND2_X1 _10929_ (
    .A1(_03036_),
    .A2(_03430_),
    .ZN(_03431_)
  );
  AND2_X1 _10930_ (
    .A1(_03429_),
    .A2(_03431_),
    .ZN(_03432_)
  );
  OR2_X1 _10931_ (
    .A1(csr_io_decode_0_inst[27]),
    .A2(_03402_),
    .ZN(_03433_)
  );
  OR2_X1 _10932_ (
    .A1(_03328_),
    .A2(_03350_),
    .ZN(_03434_)
  );
  OR2_X1 _10933_ (
    .A1(_03433_),
    .A2(_03434_),
    .ZN(_03435_)
  );
  INV_X1 _10934_ (
    .A(_03435_),
    .ZN(_03436_)
  );
  AND2_X1 _10935_ (
    .A1(_03359_),
    .A2(_03436_),
    .ZN(_03437_)
  );
  AND2_X1 _10936_ (
    .A1(_03430_),
    .A2(_03437_),
    .ZN(_03438_)
  );
  OR2_X1 _10937_ (
    .A1(_03432_),
    .A2(_03438_),
    .ZN(_03439_)
  );
  OR2_X1 _10938_ (
    .A1(_03428_),
    .A2(_03439_),
    .ZN(_03440_)
  );
  AND2_X1 _10939_ (
    .A1(_03036_),
    .A2(_03423_),
    .ZN(_03441_)
  );
  AND2_X1 _10940_ (
    .A1(_03400_),
    .A2(_03441_),
    .ZN(_03442_)
  );
  AND2_X1 _10941_ (
    .A1(csr_io_decode_0_inst[27]),
    .A2(_03358_),
    .ZN(_03443_)
  );
  AND2_X1 _10942_ (
    .A1(_03404_),
    .A2(_03443_),
    .ZN(_03444_)
  );
  OR2_X1 _10943_ (
    .A1(_03364_),
    .A2(_03376_),
    .ZN(_03445_)
  );
  AND2_X1 _10944_ (
    .A1(_03039_),
    .A2(_03383_),
    .ZN(_03446_)
  );
  OR2_X1 _10945_ (
    .A1(_03413_),
    .A2(_03440_),
    .ZN(_03447_)
  );
  OR2_X1 _10946_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[3]),
    .ZN(_03448_)
  );
  OR2_X1 _10947_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_03449_)
  );
  OR2_X1 _10948_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_03449_),
    .ZN(_03450_)
  );
  OR2_X1 _10949_ (
    .A1(_03448_),
    .A2(_03450_),
    .ZN(_03451_)
  );
  AND2_X1 _10950_ (
    .A1(ex_ctrl_wxd),
    .A2(ex_reg_valid),
    .ZN(_03452_)
  );
  OR2_X1 _10951_ (
    .A1(_02983_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[0]),
    .ZN(_03453_)
  );
  OR2_X1 _10952_ (
    .A1(_02985_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_03454_)
  );
  AND2_X1 _10953_ (
    .A1(_03453_),
    .A2(_03454_),
    .ZN(_03455_)
  );
  OR2_X1 _10954_ (
    .A1(ex_reg_inst[8]),
    .A2(_03045_),
    .ZN(_03456_)
  );
  OR2_X1 _10955_ (
    .A1(ex_reg_inst[7]),
    .A2(_03044_),
    .ZN(_03457_)
  );
  AND2_X1 _10956_ (
    .A1(_03456_),
    .A2(_03457_),
    .ZN(_03458_)
  );
  AND2_X1 _10957_ (
    .A1(_03455_),
    .A2(_03458_),
    .ZN(_03459_)
  );
  XOR2_X1 _10958_ (
    .A(ex_reg_inst[9]),
    .B(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_03460_)
  );
  XOR2_X1 _10959_ (
    .A(ex_reg_inst[11]),
    .B(ibuf_io_inst_0_bits_inst_rs1[4]),
    .Z(_03461_)
  );
  XOR2_X1 _10960_ (
    .A(ex_reg_inst[10]),
    .B(ibuf_io_inst_0_bits_inst_rs1[3]),
    .Z(_03462_)
  );
  OR2_X1 _10961_ (
    .A1(_03461_),
    .A2(_03462_),
    .ZN(_03463_)
  );
  OR2_X1 _10962_ (
    .A1(_03460_),
    .A2(_03463_),
    .ZN(_03464_)
  );
  INV_X1 _10963_ (
    .A(_03464_),
    .ZN(_03465_)
  );
  AND2_X1 _10964_ (
    .A1(_03459_),
    .A2(_03465_),
    .ZN(_03466_)
  );
  AND2_X1 _10965_ (
    .A1(_03452_),
    .A2(_03466_),
    .ZN(_03467_)
  );
  INV_X1 _10966_ (
    .A(_03467_),
    .ZN(_03468_)
  );
  AND2_X1 _10967_ (
    .A1(_03451_),
    .A2(_03468_),
    .ZN(_03469_)
  );
  INV_X1 _10968_ (
    .A(_03469_),
    .ZN(_03470_)
  );
  AND2_X1 _10969_ (
    .A1(mem_ctrl_wxd),
    .A2(mem_reg_valid),
    .ZN(_03471_)
  );
  INV_X1 _10970_ (
    .A(_03471_),
    .ZN(_03472_)
  );
  AND2_X1 _10971_ (
    .A1(mem_reg_inst[7]),
    .A2(_03044_),
    .ZN(_03473_)
  );
  AND2_X1 _10972_ (
    .A1(mem_reg_inst[8]),
    .A2(_03045_),
    .ZN(_03474_)
  );
  OR2_X1 _10973_ (
    .A1(_03473_),
    .A2(_03474_),
    .ZN(_03475_)
  );
  AND2_X1 _10974_ (
    .A1(_02984_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_03476_)
  );
  AND2_X1 _10975_ (
    .A1(_02982_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[0]),
    .ZN(_03477_)
  );
  OR2_X1 _10976_ (
    .A1(_03476_),
    .A2(_03477_),
    .ZN(_03478_)
  );
  OR2_X1 _10977_ (
    .A1(_03475_),
    .A2(_03478_),
    .ZN(_03479_)
  );
  XOR2_X1 _10978_ (
    .A(mem_reg_inst[9]),
    .B(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_03480_)
  );
  XOR2_X1 _10979_ (
    .A(mem_reg_inst[11]),
    .B(ibuf_io_inst_0_bits_inst_rs1[4]),
    .Z(_03481_)
  );
  XOR2_X1 _10980_ (
    .A(mem_reg_inst[10]),
    .B(ibuf_io_inst_0_bits_inst_rs1[3]),
    .Z(_03482_)
  );
  OR2_X1 _10981_ (
    .A1(_03481_),
    .A2(_03482_),
    .ZN(_03483_)
  );
  OR2_X1 _10982_ (
    .A1(_03480_),
    .A2(_03483_),
    .ZN(_03484_)
  );
  OR2_X1 _10983_ (
    .A1(_03479_),
    .A2(_03484_),
    .ZN(_03485_)
  );
  INV_X1 _10984_ (
    .A(_03485_),
    .ZN(_03486_)
  );
  AND2_X1 _10985_ (
    .A1(_03471_),
    .A2(_03486_),
    .ZN(_03487_)
  );
  OR2_X1 _10986_ (
    .A1(_03470_),
    .A2(_03487_),
    .ZN(_03488_)
  );
  INV_X1 _10987_ (
    .A(_03488_),
    .ZN(_03489_)
  );
  AND2_X1 _10988_ (
    .A1(_03447_),
    .A2(_03489_),
    .ZN(_03490_)
  );
  AND2_X1 _10989_ (
    .A1(_03036_),
    .A2(csr_io_decode_0_inst[4]),
    .ZN(_03491_)
  );
  AND2_X1 _10990_ (
    .A1(csr_io_decode_0_inst[2]),
    .A2(_03491_),
    .ZN(_03492_)
  );
  AND2_X1 _10991_ (
    .A1(_03341_),
    .A2(_03492_),
    .ZN(_03493_)
  );
  OR2_X1 _10992_ (
    .A1(_03439_),
    .A2(_03493_),
    .ZN(_03494_)
  );
  AND2_X1 _10993_ (
    .A1(_03351_),
    .A2(_03416_),
    .ZN(_03495_)
  );
  OR2_X1 _10994_ (
    .A1(_03355_),
    .A2(_03417_),
    .ZN(_03496_)
  );
  INV_X1 _10995_ (
    .A(_03496_),
    .ZN(_03497_)
  );
  AND2_X1 _10996_ (
    .A1(_03391_),
    .A2(_03497_),
    .ZN(_03498_)
  );
  AND2_X1 _10997_ (
    .A1(_03495_),
    .A2(_03498_),
    .ZN(_03499_)
  );
  OR2_X1 _10998_ (
    .A1(csr_io_decode_0_inst[16]),
    .A2(csr_io_decode_0_inst[17]),
    .ZN(_03500_)
  );
  OR2_X1 _10999_ (
    .A1(csr_io_decode_0_inst[15]),
    .A2(csr_io_decode_0_inst[18]),
    .ZN(_03501_)
  );
  OR2_X1 _11000_ (
    .A1(_03500_),
    .A2(_03501_),
    .ZN(_03502_)
  );
  OR2_X1 _11001_ (
    .A1(csr_io_decode_0_inst[10]),
    .A2(csr_io_decode_0_inst[14]),
    .ZN(_03503_)
  );
  OR2_X1 _11002_ (
    .A1(csr_io_decode_0_inst[9]),
    .A2(_03503_),
    .ZN(_03504_)
  );
  OR2_X1 _11003_ (
    .A1(_03502_),
    .A2(_03504_),
    .ZN(_03505_)
  );
  INV_X1 _11004_ (
    .A(_03505_),
    .ZN(_03506_)
  );
  OR2_X1 _11005_ (
    .A1(csr_io_decode_0_inst[7]),
    .A2(csr_io_decode_0_inst[8]),
    .ZN(_03507_)
  );
  OR2_X1 _11006_ (
    .A1(csr_io_decode_0_inst[11]),
    .A2(csr_io_decode_0_inst[19]),
    .ZN(_03508_)
  );
  OR2_X1 _11007_ (
    .A1(_03507_),
    .A2(_03508_),
    .ZN(_03509_)
  );
  OR2_X1 _11008_ (
    .A1(_03323_),
    .A2(_03509_),
    .ZN(_03510_)
  );
  INV_X1 _11009_ (
    .A(_03510_),
    .ZN(_03511_)
  );
  AND2_X1 _11010_ (
    .A1(_03506_),
    .A2(_03511_),
    .ZN(_03512_)
  );
  OR2_X1 _11011_ (
    .A1(csr_io_decode_0_inst[22]),
    .A2(csr_io_decode_0_inst[28]),
    .ZN(_03513_)
  );
  OR2_X1 _11012_ (
    .A1(csr_io_decode_0_inst[29]),
    .A2(_03513_),
    .ZN(_03514_)
  );
  INV_X1 _11013_ (
    .A(_03514_),
    .ZN(_03515_)
  );
  AND2_X1 _11014_ (
    .A1(csr_io_decode_0_inst[20]),
    .A2(csr_io_decode_0_inst[22]),
    .ZN(_03516_)
  );
  AND2_X1 _11015_ (
    .A1(csr_io_decode_0_inst[28]),
    .A2(_03516_),
    .ZN(_03517_)
  );
  OR2_X1 _11016_ (
    .A1(_03515_),
    .A2(_03517_),
    .ZN(_03518_)
  );
  AND2_X1 _11017_ (
    .A1(_03512_),
    .A2(_03518_),
    .ZN(_03519_)
  );
  AND2_X1 _11018_ (
    .A1(_03499_),
    .A2(_03519_),
    .ZN(_03520_)
  );
  AND2_X1 _11019_ (
    .A1(_03317_),
    .A2(_03520_),
    .ZN(_03521_)
  );
  OR2_X1 _11020_ (
    .A1(_03494_),
    .A2(_03521_),
    .ZN(_03522_)
  );
  OR2_X1 _11021_ (
    .A1(_03445_),
    .A2(_03522_),
    .ZN(_03523_)
  );
  AND2_X1 _11022_ (
    .A1(_03001_),
    .A2(_03394_),
    .ZN(_03524_)
  );
  AND2_X1 _11023_ (
    .A1(csr_io_decode_0_inst[28]),
    .A2(csr_io_decode_0_inst[29]),
    .ZN(_03525_)
  );
  AND2_X1 _11024_ (
    .A1(_03009_),
    .A2(csr_io_decode_0_inst[6]),
    .ZN(_03526_)
  );
  AND2_X1 _11025_ (
    .A1(_03525_),
    .A2(_03526_),
    .ZN(_03527_)
  );
  AND2_X1 _11026_ (
    .A1(csr_io_decode_0_inst[21]),
    .A2(_03003_),
    .ZN(_03528_)
  );
  AND2_X1 _11027_ (
    .A1(_03419_),
    .A2(_03528_),
    .ZN(_03529_)
  );
  AND2_X1 _11028_ (
    .A1(_03390_),
    .A2(_03529_),
    .ZN(_03530_)
  );
  AND2_X1 _11029_ (
    .A1(_03527_),
    .A2(_03530_),
    .ZN(_03531_)
  );
  AND2_X1 _11030_ (
    .A1(csr_io_decode_0_inst[25]),
    .A2(csr_io_decode_0_inst[27]),
    .ZN(_03532_)
  );
  AND2_X1 _11031_ (
    .A1(csr_io_decode_0_inst[24]),
    .A2(_03532_),
    .ZN(_03533_)
  );
  AND2_X1 _11032_ (
    .A1(_03005_),
    .A2(_03533_),
    .ZN(_03534_)
  );
  MUX2_X1 _11033_ (
    .A(_03495_),
    .B(_03534_),
    .S(csr_io_decode_0_inst[30]),
    .Z(_03535_)
  );
  AND2_X1 _11034_ (
    .A1(_03512_),
    .A2(_03535_),
    .ZN(_03536_)
  );
  AND2_X1 _11035_ (
    .A1(_03531_),
    .A2(_03536_),
    .ZN(_03537_)
  );
  OR2_X1 _11036_ (
    .A1(_03524_),
    .A2(_03537_),
    .ZN(_03538_)
  );
  AND2_X1 _11037_ (
    .A1(_03319_),
    .A2(_03538_),
    .ZN(_03539_)
  );
  AND2_X1 _11038_ (
    .A1(_03385_),
    .A2(_03423_),
    .ZN(_03540_)
  );
  AND2_X1 _11039_ (
    .A1(csr_io_decode_0_inst[13]),
    .A2(_03392_),
    .ZN(_03541_)
  );
  INV_X1 _11040_ (
    .A(_03541_),
    .ZN(_03542_)
  );
  AND2_X1 _11041_ (
    .A1(csr_io_decode_0_inst[6]),
    .A2(_03400_),
    .ZN(_03543_)
  );
  AND2_X1 _11042_ (
    .A1(_03342_),
    .A2(_03446_),
    .ZN(_03544_)
  );
  OR2_X1 _11043_ (
    .A1(_03541_),
    .A2(_03544_),
    .ZN(_03545_)
  );
  OR2_X1 _11044_ (
    .A1(csr_io_decode_0_inst[14]),
    .A2(csr_io_decode_0_inst[6]),
    .ZN(_03546_)
  );
  INV_X1 _11045_ (
    .A(_03546_),
    .ZN(_03547_)
  );
  AND2_X1 _11046_ (
    .A1(_03383_),
    .A2(_03547_),
    .ZN(_03548_)
  );
  AND2_X1 _11047_ (
    .A1(_03335_),
    .A2(_03548_),
    .ZN(_03549_)
  );
  OR2_X1 _11048_ (
    .A1(_03545_),
    .A2(_03549_),
    .ZN(_03550_)
  );
  OR2_X1 _11049_ (
    .A1(_03540_),
    .A2(_03550_),
    .ZN(_03551_)
  );
  OR2_X1 _11050_ (
    .A1(_03387_),
    .A2(_03427_),
    .ZN(_03552_)
  );
  OR2_X1 _11051_ (
    .A1(_03551_),
    .A2(_03552_),
    .ZN(_03553_)
  );
  OR2_X1 _11052_ (
    .A1(_03539_),
    .A2(_03553_),
    .ZN(_03554_)
  );
  OR2_X1 _11053_ (
    .A1(_03405_),
    .A2(_03444_),
    .ZN(_03555_)
  );
  AND2_X1 _11054_ (
    .A1(_03404_),
    .A2(_03423_),
    .ZN(_03556_)
  );
  AND2_X1 _11055_ (
    .A1(_03327_),
    .A2(_03446_),
    .ZN(_03557_)
  );
  AND2_X1 _11056_ (
    .A1(_03407_),
    .A2(_03557_),
    .ZN(_03558_)
  );
  OR2_X1 _11057_ (
    .A1(_03523_),
    .A2(_03554_),
    .ZN(_03559_)
  );
  INV_X1 _11058_ (
    .A(_03559_),
    .ZN(_03560_)
  );
  AND2_X1 _11059_ (
    .A1(csr_io_decode_0_inst[12]),
    .A2(_03392_),
    .ZN(_03561_)
  );
  AND2_X1 _11060_ (
    .A1(_03323_),
    .A2(_03392_),
    .ZN(_03562_)
  );
  INV_X1 _11061_ (
    .A(_03562_),
    .ZN(_03563_)
  );
  OR2_X1 _11062_ (
    .A1(_03520_),
    .A2(_03562_),
    .ZN(_03564_)
  );
  OR2_X1 _11063_ (
    .A1(_03537_),
    .A2(_03564_),
    .ZN(_03565_)
  );
  AND2_X1 _11064_ (
    .A1(_03563_),
    .A2(_03565_),
    .ZN(_03566_)
  );
  AND2_X1 _11065_ (
    .A1(_03065_),
    .A2(csr_io_decode_0_system_illegal),
    .ZN(_03567_)
  );
  AND2_X1 _11066_ (
    .A1(_03566_),
    .A2(_03567_),
    .ZN(_03568_)
  );
  OR2_X1 _11067_ (
    .A1(_03451_),
    .A2(_03542_),
    .ZN(_03569_)
  );
  AND2_X1 _11068_ (
    .A1(csr_io_decode_0_write_illegal),
    .A2(_03569_),
    .ZN(_03570_)
  );
  OR2_X1 _11069_ (
    .A1(csr_io_decode_0_read_illegal),
    .A2(_03570_),
    .ZN(_03571_)
  );
  AND2_X1 _11070_ (
    .A1(_03562_),
    .A2(_03571_),
    .ZN(_03572_)
  );
  AND2_X1 _11071_ (
    .A1(ibuf_io_inst_0_bits_rvc),
    .A2(_03079_),
    .ZN(_03573_)
  );
  AND2_X1 _11072_ (
    .A1(csr_io_decode_0_inst[25]),
    .A2(_03432_),
    .ZN(_03574_)
  );
  AND2_X1 _11073_ (
    .A1(_03077_),
    .A2(_03574_),
    .ZN(_03575_)
  );
  OR2_X1 _11074_ (
    .A1(_03573_),
    .A2(_03575_),
    .ZN(_03576_)
  );
  OR2_X1 _11075_ (
    .A1(_03572_),
    .A2(_03576_),
    .ZN(_03577_)
  );
  OR2_X1 _11076_ (
    .A1(_03442_),
    .A2(_03555_),
    .ZN(_03578_)
  );
  AND2_X1 _11077_ (
    .A1(_03078_),
    .A2(_03578_),
    .ZN(_03579_)
  );
  OR2_X1 _11078_ (
    .A1(_03577_),
    .A2(_03579_),
    .ZN(_03580_)
  );
  OR2_X1 _11079_ (
    .A1(_03568_),
    .A2(_03580_),
    .ZN(_03581_)
  );
  OR2_X1 _11080_ (
    .A1(_03560_),
    .A2(_03581_),
    .ZN(_03582_)
  );
  INV_X1 _11081_ (
    .A(_03582_),
    .ZN(_03583_)
  );
  OR2_X1 _11082_ (
    .A1(_03490_),
    .A2(_03582_),
    .ZN(_03584_)
  );
  INV_X1 _11083_ (
    .A(_03584_),
    .ZN(_03585_)
  );
  OR2_X1 _11084_ (
    .A1(csr_io_interrupt),
    .A2(ibuf_io_inst_0_bits_replay),
    .ZN(_03586_)
  );
  OR2_X1 _11085_ (
    .A1(_03362_),
    .A2(_03371_),
    .ZN(_03587_)
  );
  OR2_X1 _11086_ (
    .A1(_03493_),
    .A2(_03561_),
    .ZN(_03588_)
  );
  OR2_X1 _11087_ (
    .A1(_03545_),
    .A2(_03588_),
    .ZN(_03589_)
  );
  AND2_X1 _11088_ (
    .A1(csr_io_decode_0_inst[2]),
    .A2(_03345_),
    .ZN(_03590_)
  );
  AND2_X1 _11089_ (
    .A1(csr_io_decode_0_inst[13]),
    .A2(csr_io_decode_0_inst[14]),
    .ZN(_03591_)
  );
  OR2_X1 _11090_ (
    .A1(csr_io_decode_0_inst[12]),
    .A2(_03591_),
    .ZN(_03592_)
  );
  INV_X1 _11091_ (
    .A(_03592_),
    .ZN(_03593_)
  );
  OR2_X1 _11092_ (
    .A1(_03325_),
    .A2(_03593_),
    .ZN(_03594_)
  );
  AND2_X1 _11093_ (
    .A1(_03321_),
    .A2(_03594_),
    .ZN(_03595_)
  );
  OR2_X1 _11094_ (
    .A1(_03590_),
    .A2(_03595_),
    .ZN(_03596_)
  );
  OR2_X1 _11095_ (
    .A1(_03589_),
    .A2(_03596_),
    .ZN(_03597_)
  );
  OR2_X1 _11096_ (
    .A1(_03387_),
    .A2(_03597_),
    .ZN(_03598_)
  );
  OR2_X1 _11097_ (
    .A1(_03362_),
    .A2(_03375_),
    .ZN(_03599_)
  );
  OR2_X1 _11098_ (
    .A1(_03587_),
    .A2(_03598_),
    .ZN(_03600_)
  );
  OR2_X1 _11099_ (
    .A1(_03440_),
    .A2(_03600_),
    .ZN(_03601_)
  );
  OR2_X1 _11100_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[0]),
    .A2(ibuf_io_inst_0_bits_inst_rd[1]),
    .ZN(_03602_)
  );
  OR2_X1 _11101_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[2]),
    .A2(ibuf_io_inst_0_bits_inst_rd[4]),
    .ZN(_03603_)
  );
  OR2_X1 _11102_ (
    .A1(_03602_),
    .A2(_03603_),
    .ZN(_03604_)
  );
  OR2_X1 _11103_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[3]),
    .A2(_03604_),
    .ZN(_03605_)
  );
  AND2_X1 _11104_ (
    .A1(_03601_),
    .A2(_03605_),
    .ZN(_03606_)
  );
  AND2_X1 _11105_ (
    .A1(_03053_),
    .A2(_03103_),
    .ZN(_03607_)
  );
  AND2_X1 _11106_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[1]),
    .A2(_03102_),
    .ZN(_03608_)
  );
  XOR2_X1 _11107_ (
    .A(_03052_),
    .B(_03100_),
    .Z(_03609_)
  );
  OR2_X1 _11108_ (
    .A1(_03607_),
    .A2(_03609_),
    .ZN(_03610_)
  );
  XOR2_X1 _11109_ (
    .A(_03054_),
    .B(_03105_),
    .Z(_03611_)
  );
  XOR2_X1 _11110_ (
    .A(_03055_),
    .B(_03108_),
    .Z(_03612_)
  );
  OR2_X1 _11111_ (
    .A1(_03611_),
    .A2(_03612_),
    .ZN(_03613_)
  );
  XOR2_X1 _11112_ (
    .A(ibuf_io_inst_0_bits_inst_rd[4]),
    .B(_03110_),
    .Z(_03614_)
  );
  OR2_X1 _11113_ (
    .A1(_03116_),
    .A2(_03608_),
    .ZN(_03615_)
  );
  OR2_X1 _11114_ (
    .A1(_03614_),
    .A2(_03615_),
    .ZN(_03616_)
  );
  OR2_X1 _11115_ (
    .A1(_03613_),
    .A2(_03616_),
    .ZN(_03617_)
  );
  OR2_X1 _11116_ (
    .A1(_03610_),
    .A2(_03617_),
    .ZN(_03618_)
  );
  MUX2_X1 _11117_ (
    .A(_r[24]),
    .B(_r[25]),
    .S(ibuf_io_inst_0_bits_inst_rd[0]),
    .Z(_03619_)
  );
  AND2_X1 _11118_ (
    .A1(_03054_),
    .A2(_03619_),
    .ZN(_03620_)
  );
  MUX2_X1 _11119_ (
    .A(_r[28]),
    .B(_r[29]),
    .S(ibuf_io_inst_0_bits_inst_rd[0]),
    .Z(_03621_)
  );
  AND2_X1 _11120_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[2]),
    .A2(_03621_),
    .ZN(_03622_)
  );
  OR2_X1 _11121_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[1]),
    .A2(_03622_),
    .ZN(_03623_)
  );
  OR2_X1 _11122_ (
    .A1(_03620_),
    .A2(_03623_),
    .ZN(_03624_)
  );
  MUX2_X1 _11123_ (
    .A(_r[26]),
    .B(_r[27]),
    .S(ibuf_io_inst_0_bits_inst_rd[0]),
    .Z(_03625_)
  );
  AND2_X1 _11124_ (
    .A1(_03054_),
    .A2(_03625_),
    .ZN(_03626_)
  );
  MUX2_X1 _11125_ (
    .A(_r[30]),
    .B(_r[31]),
    .S(ibuf_io_inst_0_bits_inst_rd[0]),
    .Z(_03627_)
  );
  AND2_X1 _11126_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[2]),
    .A2(_03627_),
    .ZN(_03628_)
  );
  OR2_X1 _11127_ (
    .A1(_03053_),
    .A2(_03628_),
    .ZN(_03629_)
  );
  OR2_X1 _11128_ (
    .A1(_03626_),
    .A2(_03629_),
    .ZN(_03630_)
  );
  AND2_X1 _11129_ (
    .A1(_03624_),
    .A2(_03630_),
    .ZN(_03631_)
  );
  AND2_X1 _11130_ (
    .A1(_r[17]),
    .A2(_03053_),
    .ZN(_03632_)
  );
  AND2_X1 _11131_ (
    .A1(_r[19]),
    .A2(ibuf_io_inst_0_bits_inst_rd[1]),
    .ZN(_03633_)
  );
  OR2_X1 _11132_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[2]),
    .A2(_03633_),
    .ZN(_03634_)
  );
  OR2_X1 _11133_ (
    .A1(_03632_),
    .A2(_03634_),
    .ZN(_03635_)
  );
  AND2_X1 _11134_ (
    .A1(_r[21]),
    .A2(_03053_),
    .ZN(_03636_)
  );
  AND2_X1 _11135_ (
    .A1(_r[23]),
    .A2(ibuf_io_inst_0_bits_inst_rd[1]),
    .ZN(_03637_)
  );
  OR2_X1 _11136_ (
    .A1(_03054_),
    .A2(_03637_),
    .ZN(_03638_)
  );
  OR2_X1 _11137_ (
    .A1(_03636_),
    .A2(_03638_),
    .ZN(_03639_)
  );
  AND2_X1 _11138_ (
    .A1(_03635_),
    .A2(_03639_),
    .ZN(_03640_)
  );
  AND2_X1 _11139_ (
    .A1(_r[16]),
    .A2(_03053_),
    .ZN(_03641_)
  );
  AND2_X1 _11140_ (
    .A1(_r[18]),
    .A2(ibuf_io_inst_0_bits_inst_rd[1]),
    .ZN(_03642_)
  );
  OR2_X1 _11141_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[2]),
    .A2(_03642_),
    .ZN(_03643_)
  );
  OR2_X1 _11142_ (
    .A1(_03641_),
    .A2(_03643_),
    .ZN(_03644_)
  );
  AND2_X1 _11143_ (
    .A1(_r[20]),
    .A2(_03053_),
    .ZN(_03645_)
  );
  AND2_X1 _11144_ (
    .A1(_r[22]),
    .A2(ibuf_io_inst_0_bits_inst_rd[1]),
    .ZN(_03646_)
  );
  OR2_X1 _11145_ (
    .A1(_03054_),
    .A2(_03646_),
    .ZN(_03647_)
  );
  OR2_X1 _11146_ (
    .A1(_03645_),
    .A2(_03647_),
    .ZN(_03648_)
  );
  AND2_X1 _11147_ (
    .A1(_03644_),
    .A2(_03648_),
    .ZN(_03649_)
  );
  MUX2_X1 _11148_ (
    .A(_03640_),
    .B(_03649_),
    .S(_03052_),
    .Z(_03650_)
  );
  MUX2_X1 _11149_ (
    .A(_03631_),
    .B(_03650_),
    .S(_03055_),
    .Z(_03651_)
  );
  MUX2_X1 _11150_ (
    .A(_r[1]),
    .B(_r[5]),
    .S(ibuf_io_inst_0_bits_inst_rd[2]),
    .Z(_03652_)
  );
  OR2_X1 _11151_ (
    .A1(_r[14]),
    .A2(_03054_),
    .ZN(_03653_)
  );
  OR2_X1 _11152_ (
    .A1(_r[10]),
    .A2(ibuf_io_inst_0_bits_inst_rd[2]),
    .ZN(_03654_)
  );
  AND2_X1 _11153_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[1]),
    .A2(_03654_),
    .ZN(_03655_)
  );
  AND2_X1 _11154_ (
    .A1(_03653_),
    .A2(_03655_),
    .ZN(_03656_)
  );
  MUX2_X1 _11155_ (
    .A(_r[8]),
    .B(_r[12]),
    .S(ibuf_io_inst_0_bits_inst_rd[2]),
    .Z(_03657_)
  );
  AND2_X1 _11156_ (
    .A1(_03053_),
    .A2(_03657_),
    .ZN(_03658_)
  );
  OR2_X1 _11157_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[0]),
    .A2(_03658_),
    .ZN(_03659_)
  );
  OR2_X1 _11158_ (
    .A1(_03656_),
    .A2(_03659_),
    .ZN(_03660_)
  );
  MUX2_X1 _11159_ (
    .A(_r[9]),
    .B(_r[13]),
    .S(ibuf_io_inst_0_bits_inst_rd[2]),
    .Z(_03661_)
  );
  AND2_X1 _11160_ (
    .A1(_03053_),
    .A2(_03661_),
    .ZN(_03662_)
  );
  OR2_X1 _11161_ (
    .A1(_r[11]),
    .A2(ibuf_io_inst_0_bits_inst_rd[2]),
    .ZN(_03663_)
  );
  OR2_X1 _11162_ (
    .A1(_r[15]),
    .A2(_03054_),
    .ZN(_03664_)
  );
  AND2_X1 _11163_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[1]),
    .A2(_03664_),
    .ZN(_03665_)
  );
  AND2_X1 _11164_ (
    .A1(_03663_),
    .A2(_03665_),
    .ZN(_03666_)
  );
  OR2_X1 _11165_ (
    .A1(_03052_),
    .A2(_03666_),
    .ZN(_03667_)
  );
  OR2_X1 _11166_ (
    .A1(_03662_),
    .A2(_03667_),
    .ZN(_03668_)
  );
  AND2_X1 _11167_ (
    .A1(_03660_),
    .A2(_03668_),
    .ZN(_03669_)
  );
  OR2_X1 _11168_ (
    .A1(_r[3]),
    .A2(ibuf_io_inst_0_bits_inst_rd[2]),
    .ZN(_03670_)
  );
  OR2_X1 _11169_ (
    .A1(_r[7]),
    .A2(_03054_),
    .ZN(_03671_)
  );
  AND2_X1 _11170_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[1]),
    .A2(_03670_),
    .ZN(_03672_)
  );
  AND2_X1 _11171_ (
    .A1(_03671_),
    .A2(_03672_),
    .ZN(_03673_)
  );
  AND2_X1 _11172_ (
    .A1(_03053_),
    .A2(_03652_),
    .ZN(_03674_)
  );
  OR2_X1 _11173_ (
    .A1(_03052_),
    .A2(_03674_),
    .ZN(_03675_)
  );
  OR2_X1 _11174_ (
    .A1(_03673_),
    .A2(_03675_),
    .ZN(_03676_)
  );
  OR2_X1 _11175_ (
    .A1(_r[6]),
    .A2(_03054_),
    .ZN(_03677_)
  );
  OR2_X1 _11176_ (
    .A1(_r[2]),
    .A2(ibuf_io_inst_0_bits_inst_rd[2]),
    .ZN(_03678_)
  );
  AND2_X1 _11177_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[1]),
    .A2(_03678_),
    .ZN(_03679_)
  );
  AND2_X1 _11178_ (
    .A1(_03677_),
    .A2(_03679_),
    .ZN(_03680_)
  );
  AND2_X1 _11179_ (
    .A1(_r[4]),
    .A2(ibuf_io_inst_0_bits_inst_rd[2]),
    .ZN(_03681_)
  );
  AND2_X1 _11180_ (
    .A1(_03053_),
    .A2(_03681_),
    .ZN(_03682_)
  );
  OR2_X1 _11181_ (
    .A1(ibuf_io_inst_0_bits_inst_rd[0]),
    .A2(_03682_),
    .ZN(_03683_)
  );
  OR2_X1 _11182_ (
    .A1(_03680_),
    .A2(_03683_),
    .ZN(_03684_)
  );
  AND2_X1 _11183_ (
    .A1(_03676_),
    .A2(_03684_),
    .ZN(_03685_)
  );
  MUX2_X1 _11184_ (
    .A(_03669_),
    .B(_03685_),
    .S(_03055_),
    .Z(_03686_)
  );
  MUX2_X1 _11185_ (
    .A(_03686_),
    .B(_03651_),
    .S(ibuf_io_inst_0_bits_inst_rd[4]),
    .Z(_03687_)
  );
  AND2_X1 _11186_ (
    .A1(_03618_),
    .A2(_03687_),
    .ZN(_03688_)
  );
  AND2_X1 _11187_ (
    .A1(_03606_),
    .A2(_03688_),
    .ZN(_03689_)
  );
  AND2_X1 _11188_ (
    .A1(ex_ctrl_mem),
    .A2(ex_reg_valid),
    .ZN(io_dmem_req_valid)
  );
  OR2_X1 _11189_ (
    .A1(_03080_),
    .A2(io_dmem_req_valid),
    .ZN(_03690_)
  );
  AND2_X1 _11190_ (
    .A1(_03084_),
    .A2(_03114_),
    .ZN(_03691_)
  );
  AND2_X1 _11191_ (
    .A1(ex_ctrl_div),
    .A2(ex_reg_valid),
    .ZN(div_io_req_valid)
  );
  OR2_X1 _11192_ (
    .A1(_03691_),
    .A2(div_io_req_valid),
    .ZN(_03692_)
  );
  AND2_X1 _11193_ (
    .A1(_03574_),
    .A2(_03692_),
    .ZN(_03693_)
  );
  OR2_X1 _11194_ (
    .A1(ex_reg_valid),
    .A2(mem_reg_valid),
    .ZN(_03694_)
  );
  OR2_X1 _11195_ (
    .A1(wb_reg_valid),
    .A2(_03694_),
    .ZN(_03695_)
  );
  AND2_X1 _11196_ (
    .A1(csr_io_singleStep),
    .A2(_03695_),
    .ZN(_03696_)
  );
  OR2_X1 _11197_ (
    .A1(id_reg_pause),
    .A2(csr_io_csr_stall),
    .ZN(_03697_)
  );
  OR2_X1 _11198_ (
    .A1(_03696_),
    .A2(_03697_),
    .ZN(_03698_)
  );
  OR2_X1 _11199_ (
    .A1(_03693_),
    .A2(_03698_),
    .ZN(_03699_)
  );
  AND2_X1 _11200_ (
    .A1(_03083_),
    .A2(blocked),
    .ZN(_03700_)
  );
  AND2_X1 _11201_ (
    .A1(id_reg_fence),
    .A2(_03690_),
    .ZN(_03701_)
  );
  OR2_X1 _11202_ (
    .A1(_03700_),
    .A2(_03701_),
    .ZN(_03702_)
  );
  AND2_X1 _11203_ (
    .A1(_03447_),
    .A2(_03451_),
    .ZN(_03703_)
  );
  AND2_X1 _11204_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_03100_),
    .ZN(_03704_)
  );
  AND2_X1 _11205_ (
    .A1(_03044_),
    .A2(_03101_),
    .ZN(_03705_)
  );
  XOR2_X1 _11206_ (
    .A(ibuf_io_inst_0_bits_inst_rs1[4]),
    .B(_03110_),
    .Z(_03706_)
  );
  XOR2_X1 _11207_ (
    .A(_03046_),
    .B(_03105_),
    .Z(_03707_)
  );
  XOR2_X1 _11208_ (
    .A(_03047_),
    .B(_03108_),
    .Z(_03708_)
  );
  XOR2_X1 _11209_ (
    .A(_03045_),
    .B(_03102_),
    .Z(_03709_)
  );
  OR2_X1 _11210_ (
    .A1(_03116_),
    .A2(_03704_),
    .ZN(_03710_)
  );
  OR2_X1 _11211_ (
    .A1(_03705_),
    .A2(_03710_),
    .ZN(_03711_)
  );
  OR2_X1 _11212_ (
    .A1(_03706_),
    .A2(_03709_),
    .ZN(_03712_)
  );
  OR2_X1 _11213_ (
    .A1(_03708_),
    .A2(_03712_),
    .ZN(_03713_)
  );
  OR2_X1 _11214_ (
    .A1(_03707_),
    .A2(_03713_),
    .ZN(_03714_)
  );
  OR2_X1 _11215_ (
    .A1(_03711_),
    .A2(_03714_),
    .ZN(_03715_)
  );
  MUX2_X1 _11216_ (
    .A(_r[26]),
    .B(_r[30]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_03716_)
  );
  AND2_X1 _11217_ (
    .A1(_03044_),
    .A2(_03716_),
    .ZN(_03717_)
  );
  OR2_X1 _11218_ (
    .A1(_r[27]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_03718_)
  );
  OR2_X1 _11219_ (
    .A1(_r[31]),
    .A2(_03046_),
    .ZN(_03719_)
  );
  AND2_X1 _11220_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_03719_),
    .ZN(_03720_)
  );
  AND2_X1 _11221_ (
    .A1(_03718_),
    .A2(_03720_),
    .ZN(_03721_)
  );
  OR2_X1 _11222_ (
    .A1(_03045_),
    .A2(_03721_),
    .ZN(_03722_)
  );
  OR2_X1 _11223_ (
    .A1(_03717_),
    .A2(_03722_),
    .ZN(_03723_)
  );
  OR2_X1 _11224_ (
    .A1(_r[29]),
    .A2(_03046_),
    .ZN(_03724_)
  );
  OR2_X1 _11225_ (
    .A1(_r[25]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_03725_)
  );
  AND2_X1 _11226_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_03725_),
    .ZN(_03726_)
  );
  AND2_X1 _11227_ (
    .A1(_03724_),
    .A2(_03726_),
    .ZN(_03727_)
  );
  MUX2_X1 _11228_ (
    .A(_r[24]),
    .B(_r[28]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_03728_)
  );
  AND2_X1 _11229_ (
    .A1(_03044_),
    .A2(_03728_),
    .ZN(_03729_)
  );
  OR2_X1 _11230_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_03729_),
    .ZN(_03730_)
  );
  OR2_X1 _11231_ (
    .A1(_03727_),
    .A2(_03730_),
    .ZN(_03731_)
  );
  AND2_X1 _11232_ (
    .A1(_03723_),
    .A2(_03731_),
    .ZN(_03732_)
  );
  AND2_X1 _11233_ (
    .A1(_r[17]),
    .A2(_03045_),
    .ZN(_03733_)
  );
  AND2_X1 _11234_ (
    .A1(_r[19]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_03734_)
  );
  OR2_X1 _11235_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_03734_),
    .ZN(_03735_)
  );
  OR2_X1 _11236_ (
    .A1(_03733_),
    .A2(_03735_),
    .ZN(_03736_)
  );
  AND2_X1 _11237_ (
    .A1(_r[21]),
    .A2(_03045_),
    .ZN(_03737_)
  );
  AND2_X1 _11238_ (
    .A1(_r[23]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_03738_)
  );
  OR2_X1 _11239_ (
    .A1(_03046_),
    .A2(_03738_),
    .ZN(_03739_)
  );
  OR2_X1 _11240_ (
    .A1(_03737_),
    .A2(_03739_),
    .ZN(_03740_)
  );
  AND2_X1 _11241_ (
    .A1(_03736_),
    .A2(_03740_),
    .ZN(_03741_)
  );
  AND2_X1 _11242_ (
    .A1(_r[16]),
    .A2(_03045_),
    .ZN(_03742_)
  );
  AND2_X1 _11243_ (
    .A1(_r[18]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_03743_)
  );
  OR2_X1 _11244_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_03743_),
    .ZN(_03744_)
  );
  OR2_X1 _11245_ (
    .A1(_03742_),
    .A2(_03744_),
    .ZN(_03745_)
  );
  AND2_X1 _11246_ (
    .A1(_r[20]),
    .A2(_03045_),
    .ZN(_03746_)
  );
  AND2_X1 _11247_ (
    .A1(_r[22]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_03747_)
  );
  OR2_X1 _11248_ (
    .A1(_03046_),
    .A2(_03747_),
    .ZN(_03748_)
  );
  OR2_X1 _11249_ (
    .A1(_03746_),
    .A2(_03748_),
    .ZN(_03749_)
  );
  AND2_X1 _11250_ (
    .A1(_03745_),
    .A2(_03749_),
    .ZN(_03750_)
  );
  MUX2_X1 _11251_ (
    .A(_03741_),
    .B(_03750_),
    .S(_03044_),
    .Z(_03751_)
  );
  MUX2_X1 _11252_ (
    .A(_03732_),
    .B(_03751_),
    .S(_03047_),
    .Z(_03752_)
  );
  MUX2_X1 _11253_ (
    .A(_r[6]),
    .B(_r[7]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_03753_)
  );
  MUX2_X1 _11254_ (
    .A(_r[2]),
    .B(_r[3]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_03754_)
  );
  MUX2_X1 _11255_ (
    .A(_03753_),
    .B(_03754_),
    .S(_03046_),
    .Z(_03755_)
  );
  OR2_X1 _11256_ (
    .A1(_r[5]),
    .A2(_03046_),
    .ZN(_03756_)
  );
  OR2_X1 _11257_ (
    .A1(_r[1]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_03757_)
  );
  AND2_X1 _11258_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_03757_),
    .ZN(_03758_)
  );
  AND2_X1 _11259_ (
    .A1(_03756_),
    .A2(_03758_),
    .ZN(_03759_)
  );
  AND2_X1 _11260_ (
    .A1(_03044_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_03760_)
  );
  AND2_X1 _11261_ (
    .A1(_r[4]),
    .A2(_03760_),
    .ZN(_03761_)
  );
  OR2_X1 _11262_ (
    .A1(_03759_),
    .A2(_03761_),
    .ZN(_03762_)
  );
  MUX2_X1 _11263_ (
    .A(_03755_),
    .B(_03762_),
    .S(_03045_),
    .Z(_03763_)
  );
  OR2_X1 _11264_ (
    .A1(_r[15]),
    .A2(_03046_),
    .ZN(_03764_)
  );
  OR2_X1 _11265_ (
    .A1(_r[11]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_03765_)
  );
  AND2_X1 _11266_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_03765_),
    .ZN(_03766_)
  );
  AND2_X1 _11267_ (
    .A1(_03764_),
    .A2(_03766_),
    .ZN(_03767_)
  );
  MUX2_X1 _11268_ (
    .A(_r[10]),
    .B(_r[14]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_03768_)
  );
  AND2_X1 _11269_ (
    .A1(_03044_),
    .A2(_03768_),
    .ZN(_03769_)
  );
  OR2_X1 _11270_ (
    .A1(_03045_),
    .A2(_03769_),
    .ZN(_03770_)
  );
  OR2_X1 _11271_ (
    .A1(_03767_),
    .A2(_03770_),
    .ZN(_03771_)
  );
  OR2_X1 _11272_ (
    .A1(_r[13]),
    .A2(_03046_),
    .ZN(_03772_)
  );
  OR2_X1 _11273_ (
    .A1(_r[9]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_03773_)
  );
  AND2_X1 _11274_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_03773_),
    .ZN(_03774_)
  );
  AND2_X1 _11275_ (
    .A1(_03772_),
    .A2(_03774_),
    .ZN(_03775_)
  );
  MUX2_X1 _11276_ (
    .A(_r[8]),
    .B(_r[12]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_03776_)
  );
  AND2_X1 _11277_ (
    .A1(_03044_),
    .A2(_03776_),
    .ZN(_03777_)
  );
  OR2_X1 _11278_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_03777_),
    .ZN(_03778_)
  );
  OR2_X1 _11279_ (
    .A1(_03775_),
    .A2(_03778_),
    .ZN(_03779_)
  );
  AND2_X1 _11280_ (
    .A1(_03771_),
    .A2(_03779_),
    .ZN(_03780_)
  );
  MUX2_X1 _11281_ (
    .A(_03763_),
    .B(_03780_),
    .S(ibuf_io_inst_0_bits_inst_rs1[3]),
    .Z(_03781_)
  );
  MUX2_X1 _11282_ (
    .A(_03752_),
    .B(_03781_),
    .S(_03063_),
    .Z(_03782_)
  );
  AND2_X1 _11283_ (
    .A1(_03715_),
    .A2(_03782_),
    .ZN(_03783_)
  );
  AND2_X1 _11284_ (
    .A1(_03703_),
    .A2(_03783_),
    .ZN(_03784_)
  );
  AND2_X1 _11285_ (
    .A1(_03048_),
    .A2(_03101_),
    .ZN(_03785_)
  );
  XOR2_X1 _11286_ (
    .A(_03050_),
    .B(_03105_),
    .Z(_03786_)
  );
  OR2_X1 _11287_ (
    .A1(_03785_),
    .A2(_03786_),
    .ZN(_03787_)
  );
  AND2_X1 _11288_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03100_),
    .ZN(_03788_)
  );
  XOR2_X1 _11289_ (
    .A(_03051_),
    .B(_03108_),
    .Z(_03789_)
  );
  XOR2_X1 _11290_ (
    .A(_03049_),
    .B(_03102_),
    .Z(_03790_)
  );
  XOR2_X1 _11291_ (
    .A(ibuf_io_inst_0_bits_inst_rs2[4]),
    .B(_03110_),
    .Z(_03791_)
  );
  OR2_X1 _11292_ (
    .A1(_03790_),
    .A2(_03791_),
    .ZN(_03792_)
  );
  OR2_X1 _11293_ (
    .A1(_03789_),
    .A2(_03792_),
    .ZN(_03793_)
  );
  OR2_X1 _11294_ (
    .A1(_03116_),
    .A2(_03788_),
    .ZN(_03794_)
  );
  OR2_X1 _11295_ (
    .A1(_03787_),
    .A2(_03794_),
    .ZN(_03795_)
  );
  OR2_X1 _11296_ (
    .A1(_03793_),
    .A2(_03795_),
    .ZN(_03796_)
  );
  OR2_X1 _11297_ (
    .A1(_03368_),
    .A2(_03386_),
    .ZN(_03797_)
  );
  AND2_X1 _11298_ (
    .A1(_03395_),
    .A2(_03399_),
    .ZN(_03798_)
  );
  AND2_X1 _11299_ (
    .A1(_03320_),
    .A2(_03381_),
    .ZN(_03799_)
  );
  OR2_X1 _11300_ (
    .A1(_03798_),
    .A2(_03799_),
    .ZN(_03800_)
  );
  AND2_X1 _11301_ (
    .A1(_03348_),
    .A2(_03359_),
    .ZN(_03801_)
  );
  AND2_X1 _11302_ (
    .A1(_03430_),
    .A2(_03801_),
    .ZN(_03802_)
  );
  AND2_X1 _11303_ (
    .A1(_03369_),
    .A2(_03802_),
    .ZN(_03803_)
  );
  OR2_X1 _11304_ (
    .A1(_03800_),
    .A2(_03803_),
    .ZN(_03804_)
  );
  OR2_X1 _11305_ (
    .A1(_03797_),
    .A2(_03804_),
    .ZN(_03805_)
  );
  OR2_X1 _11306_ (
    .A1(_03440_),
    .A2(_03805_),
    .ZN(_03806_)
  );
  INV_X1 _11307_ (
    .A(_03806_),
    .ZN(_03807_)
  );
  OR2_X1 _11308_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[3]),
    .ZN(_03808_)
  );
  OR2_X1 _11309_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03809_)
  );
  OR2_X1 _11310_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[4]),
    .A2(_03809_),
    .ZN(_03810_)
  );
  OR2_X1 _11311_ (
    .A1(_03808_),
    .A2(_03810_),
    .ZN(_03811_)
  );
  AND2_X1 _11312_ (
    .A1(_03806_),
    .A2(_03811_),
    .ZN(_03812_)
  );
  OR2_X1 _11313_ (
    .A1(_r[5]),
    .A2(_03050_),
    .ZN(_03813_)
  );
  OR2_X1 _11314_ (
    .A1(_r[1]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03814_)
  );
  AND2_X1 _11315_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03814_),
    .ZN(_03815_)
  );
  AND2_X1 _11316_ (
    .A1(_03813_),
    .A2(_03815_),
    .ZN(_03816_)
  );
  AND2_X1 _11317_ (
    .A1(_03048_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03817_)
  );
  AND2_X1 _11318_ (
    .A1(_r[4]),
    .A2(_03817_),
    .ZN(_03818_)
  );
  OR2_X1 _11319_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03818_),
    .ZN(_03819_)
  );
  OR2_X1 _11320_ (
    .A1(_03816_),
    .A2(_03819_),
    .ZN(_03820_)
  );
  OR2_X1 _11321_ (
    .A1(_r[3]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03821_)
  );
  OR2_X1 _11322_ (
    .A1(_r[7]),
    .A2(_03050_),
    .ZN(_03822_)
  );
  AND2_X1 _11323_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03822_),
    .ZN(_03823_)
  );
  AND2_X1 _11324_ (
    .A1(_03821_),
    .A2(_03823_),
    .ZN(_03824_)
  );
  MUX2_X1 _11325_ (
    .A(_r[2]),
    .B(_r[6]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03825_)
  );
  AND2_X1 _11326_ (
    .A1(_03048_),
    .A2(_03825_),
    .ZN(_03826_)
  );
  OR2_X1 _11327_ (
    .A1(_03049_),
    .A2(_03826_),
    .ZN(_03827_)
  );
  OR2_X1 _11328_ (
    .A1(_03824_),
    .A2(_03827_),
    .ZN(_03828_)
  );
  AND2_X1 _11329_ (
    .A1(_03820_),
    .A2(_03828_),
    .ZN(_03829_)
  );
  MUX2_X1 _11330_ (
    .A(_r[10]),
    .B(_r[14]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03830_)
  );
  AND2_X1 _11331_ (
    .A1(_03048_),
    .A2(_03830_),
    .ZN(_03831_)
  );
  OR2_X1 _11332_ (
    .A1(_r[15]),
    .A2(_03050_),
    .ZN(_03832_)
  );
  OR2_X1 _11333_ (
    .A1(_r[11]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03833_)
  );
  AND2_X1 _11334_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03833_),
    .ZN(_03834_)
  );
  AND2_X1 _11335_ (
    .A1(_03832_),
    .A2(_03834_),
    .ZN(_03835_)
  );
  OR2_X1 _11336_ (
    .A1(_03049_),
    .A2(_03835_),
    .ZN(_03836_)
  );
  OR2_X1 _11337_ (
    .A1(_03831_),
    .A2(_03836_),
    .ZN(_03837_)
  );
  MUX2_X1 _11338_ (
    .A(_r[8]),
    .B(_r[12]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03838_)
  );
  AND2_X1 _11339_ (
    .A1(_03048_),
    .A2(_03838_),
    .ZN(_03839_)
  );
  OR2_X1 _11340_ (
    .A1(_r[13]),
    .A2(_03050_),
    .ZN(_03840_)
  );
  OR2_X1 _11341_ (
    .A1(_r[9]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03841_)
  );
  AND2_X1 _11342_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03841_),
    .ZN(_03842_)
  );
  AND2_X1 _11343_ (
    .A1(_03840_),
    .A2(_03842_),
    .ZN(_03843_)
  );
  OR2_X1 _11344_ (
    .A1(_03839_),
    .A2(_03843_),
    .ZN(_03844_)
  );
  OR2_X1 _11345_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03844_),
    .ZN(_03845_)
  );
  AND2_X1 _11346_ (
    .A1(_03837_),
    .A2(_03845_),
    .ZN(_03846_)
  );
  MUX2_X1 _11347_ (
    .A(_03829_),
    .B(_03846_),
    .S(ibuf_io_inst_0_bits_inst_rs2[3]),
    .Z(_03847_)
  );
  AND2_X1 _11348_ (
    .A1(_03064_),
    .A2(_03847_),
    .ZN(_03848_)
  );
  MUX2_X1 _11349_ (
    .A(_r[17]),
    .B(_r[21]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03849_)
  );
  MUX2_X1 _11350_ (
    .A(_r[16]),
    .B(_r[20]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03850_)
  );
  MUX2_X1 _11351_ (
    .A(_r[19]),
    .B(_r[23]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03851_)
  );
  MUX2_X1 _11352_ (
    .A(_r[18]),
    .B(_r[22]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03852_)
  );
  MUX2_X1 _11353_ (
    .A(_03849_),
    .B(_03850_),
    .S(_03048_),
    .Z(_03853_)
  );
  MUX2_X1 _11354_ (
    .A(_03851_),
    .B(_03852_),
    .S(_03048_),
    .Z(_03854_)
  );
  MUX2_X1 _11355_ (
    .A(_03853_),
    .B(_03854_),
    .S(ibuf_io_inst_0_bits_inst_rs2[1]),
    .Z(_03855_)
  );
  OR2_X1 _11356_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_03855_),
    .ZN(_03856_)
  );
  OR2_X1 _11357_ (
    .A1(_r[29]),
    .A2(_03050_),
    .ZN(_03857_)
  );
  OR2_X1 _11358_ (
    .A1(_r[25]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03858_)
  );
  AND2_X1 _11359_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03858_),
    .ZN(_03859_)
  );
  AND2_X1 _11360_ (
    .A1(_03857_),
    .A2(_03859_),
    .ZN(_03860_)
  );
  MUX2_X1 _11361_ (
    .A(_r[24]),
    .B(_r[28]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03861_)
  );
  AND2_X1 _11362_ (
    .A1(_03048_),
    .A2(_03861_),
    .ZN(_03862_)
  );
  OR2_X1 _11363_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_03862_),
    .ZN(_03863_)
  );
  OR2_X1 _11364_ (
    .A1(_03860_),
    .A2(_03863_),
    .ZN(_03864_)
  );
  OR2_X1 _11365_ (
    .A1(_r[27]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_03865_)
  );
  OR2_X1 _11366_ (
    .A1(_r[31]),
    .A2(_03050_),
    .ZN(_03866_)
  );
  AND2_X1 _11367_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_03866_),
    .ZN(_03867_)
  );
  AND2_X1 _11368_ (
    .A1(_03865_),
    .A2(_03867_),
    .ZN(_03868_)
  );
  MUX2_X1 _11369_ (
    .A(_r[26]),
    .B(_r[30]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03869_)
  );
  AND2_X1 _11370_ (
    .A1(_03048_),
    .A2(_03869_),
    .ZN(_03870_)
  );
  OR2_X1 _11371_ (
    .A1(_03049_),
    .A2(_03870_),
    .ZN(_03871_)
  );
  OR2_X1 _11372_ (
    .A1(_03868_),
    .A2(_03871_),
    .ZN(_03872_)
  );
  AND2_X1 _11373_ (
    .A1(_03864_),
    .A2(_03872_),
    .ZN(_03873_)
  );
  OR2_X1 _11374_ (
    .A1(_03051_),
    .A2(_03873_),
    .ZN(_03874_)
  );
  AND2_X1 _11375_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[4]),
    .A2(_03856_),
    .ZN(_03875_)
  );
  AND2_X1 _11376_ (
    .A1(_03874_),
    .A2(_03875_),
    .ZN(_03876_)
  );
  OR2_X1 _11377_ (
    .A1(_03848_),
    .A2(_03876_),
    .ZN(_03877_)
  );
  AND2_X1 _11378_ (
    .A1(_03796_),
    .A2(_03877_),
    .ZN(_03878_)
  );
  AND2_X1 _11379_ (
    .A1(_03812_),
    .A2(_03878_),
    .ZN(_03879_)
  );
  OR2_X1 _11380_ (
    .A1(_03689_),
    .A2(_03879_),
    .ZN(_03880_)
  );
  AND2_X1 _11381_ (
    .A1(csr_io_decode_0_inst[25]),
    .A2(_03578_),
    .ZN(_03881_)
  );
  AND2_X1 _11382_ (
    .A1(csr_io_decode_0_inst[12]),
    .A2(_03558_),
    .ZN(_03882_)
  );
  OR2_X1 _11383_ (
    .A1(_03881_),
    .A2(_03882_),
    .ZN(_03883_)
  );
  AND2_X1 _11384_ (
    .A1(_03690_),
    .A2(_03883_),
    .ZN(_03884_)
  );
  OR2_X1 _11385_ (
    .A1(_03699_),
    .A2(_03884_),
    .ZN(_03885_)
  );
  OR2_X1 _11386_ (
    .A1(_03409_),
    .A2(_03412_),
    .ZN(_03886_)
  );
  OR2_X1 _11387_ (
    .A1(_03556_),
    .A2(_03886_),
    .ZN(_03887_)
  );
  OR2_X1 _11388_ (
    .A1(_03555_),
    .A2(_03887_),
    .ZN(_03888_)
  );
  AND2_X1 _11389_ (
    .A1(_03702_),
    .A2(_03888_),
    .ZN(_03889_)
  );
  OR2_X1 _11390_ (
    .A1(_03784_),
    .A2(_03889_),
    .ZN(_03890_)
  );
  OR2_X1 _11391_ (
    .A1(_03885_),
    .A2(_03890_),
    .ZN(_03891_)
  );
  OR2_X1 _11392_ (
    .A1(_03880_),
    .A2(_03891_),
    .ZN(_03892_)
  );
  AND2_X1 _11393_ (
    .A1(mem_reg_slow_bypass),
    .A2(mem_ctrl_mem),
    .ZN(_03893_)
  );
  OR2_X1 _11394_ (
    .A1(mem_ctrl_csr[0]),
    .A2(mem_ctrl_csr[1]),
    .ZN(_03894_)
  );
  OR2_X1 _11395_ (
    .A1(mem_ctrl_csr[2]),
    .A2(mem_ctrl_div),
    .ZN(_03895_)
  );
  OR2_X1 _11396_ (
    .A1(_03894_),
    .A2(_03895_),
    .ZN(_03896_)
  );
  OR2_X1 _11397_ (
    .A1(_03893_),
    .A2(_03896_),
    .ZN(_03897_)
  );
  AND2_X1 _11398_ (
    .A1(mem_reg_inst[8]),
    .A2(_03049_),
    .ZN(_03898_)
  );
  AND2_X1 _11399_ (
    .A1(mem_reg_inst[11]),
    .A2(_03064_),
    .ZN(_03899_)
  );
  OR2_X1 _11400_ (
    .A1(_03898_),
    .A2(_03899_),
    .ZN(_03900_)
  );
  AND2_X1 _11401_ (
    .A1(_02984_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_03901_)
  );
  AND2_X1 _11402_ (
    .A1(_02989_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[4]),
    .ZN(_03902_)
  );
  OR2_X1 _11403_ (
    .A1(_03901_),
    .A2(_03902_),
    .ZN(_03903_)
  );
  OR2_X1 _11404_ (
    .A1(_03900_),
    .A2(_03903_),
    .ZN(_03904_)
  );
  XOR2_X1 _11405_ (
    .A(mem_reg_inst[7]),
    .B(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_03905_)
  );
  XOR2_X1 _11406_ (
    .A(mem_reg_inst[9]),
    .B(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03906_)
  );
  XOR2_X1 _11407_ (
    .A(mem_reg_inst[10]),
    .B(ibuf_io_inst_0_bits_inst_rs2[3]),
    .Z(_03907_)
  );
  OR2_X1 _11408_ (
    .A1(_03906_),
    .A2(_03907_),
    .ZN(_03908_)
  );
  OR2_X1 _11409_ (
    .A1(_03905_),
    .A2(_03908_),
    .ZN(_03909_)
  );
  OR2_X1 _11410_ (
    .A1(_03904_),
    .A2(_03909_),
    .ZN(_03910_)
  );
  INV_X1 _11411_ (
    .A(_03910_),
    .ZN(_03911_)
  );
  AND2_X1 _11412_ (
    .A1(_03471_),
    .A2(_03911_),
    .ZN(_03912_)
  );
  AND2_X1 _11413_ (
    .A1(_03812_),
    .A2(_03912_),
    .ZN(_03913_)
  );
  AND2_X1 _11414_ (
    .A1(_03487_),
    .A2(_03703_),
    .ZN(_03914_)
  );
  OR2_X1 _11415_ (
    .A1(_03913_),
    .A2(_03914_),
    .ZN(_03915_)
  );
  OR2_X1 _11416_ (
    .A1(mem_reg_inst[10]),
    .A2(_03055_),
    .ZN(_03916_)
  );
  OR2_X1 _11417_ (
    .A1(_02986_),
    .A2(ibuf_io_inst_0_bits_inst_rd[2]),
    .ZN(_03917_)
  );
  OR2_X1 _11418_ (
    .A1(_02987_),
    .A2(ibuf_io_inst_0_bits_inst_rd[3]),
    .ZN(_03918_)
  );
  OR2_X1 _11419_ (
    .A1(_02984_),
    .A2(ibuf_io_inst_0_bits_inst_rd[1]),
    .ZN(_03919_)
  );
  OR2_X1 _11420_ (
    .A1(mem_reg_inst[9]),
    .A2(_03054_),
    .ZN(_03920_)
  );
  OR2_X1 _11421_ (
    .A1(mem_reg_inst[8]),
    .A2(_03053_),
    .ZN(_03921_)
  );
  XOR2_X1 _11422_ (
    .A(_02989_),
    .B(ibuf_io_inst_0_bits_inst_rd[4]),
    .Z(_03922_)
  );
  AND2_X1 _11423_ (
    .A1(_03916_),
    .A2(_03921_),
    .ZN(_03923_)
  );
  AND2_X1 _11424_ (
    .A1(_03919_),
    .A2(_03923_),
    .ZN(_03924_)
  );
  AND2_X1 _11425_ (
    .A1(_03471_),
    .A2(_03917_),
    .ZN(_03925_)
  );
  XOR2_X1 _11426_ (
    .A(_02982_),
    .B(ibuf_io_inst_0_bits_inst_rd[0]),
    .Z(_03926_)
  );
  AND2_X1 _11427_ (
    .A1(_03925_),
    .A2(_03926_),
    .ZN(_03927_)
  );
  AND2_X1 _11428_ (
    .A1(_03918_),
    .A2(_03920_),
    .ZN(_03928_)
  );
  AND2_X1 _11429_ (
    .A1(_03922_),
    .A2(_03928_),
    .ZN(_03929_)
  );
  AND2_X1 _11430_ (
    .A1(_03927_),
    .A2(_03929_),
    .ZN(_03930_)
  );
  AND2_X1 _11431_ (
    .A1(_03606_),
    .A2(_03930_),
    .ZN(_03931_)
  );
  AND2_X1 _11432_ (
    .A1(_03924_),
    .A2(_03931_),
    .ZN(_03932_)
  );
  OR2_X1 _11433_ (
    .A1(_03915_),
    .A2(_03932_),
    .ZN(_03933_)
  );
  AND2_X1 _11434_ (
    .A1(_03897_),
    .A2(_03933_),
    .ZN(_03934_)
  );
  OR2_X1 _11435_ (
    .A1(_03892_),
    .A2(_03934_),
    .ZN(_03935_)
  );
  INV_X1 _11436_ (
    .A(_03935_),
    .ZN(_03936_)
  );
  AND2_X1 _11437_ (
    .A1(_03112_),
    .A2(_03126_),
    .ZN(_03937_)
  );
  XOR2_X1 _11438_ (
    .A(wb_reg_inst[7]),
    .B(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_03938_)
  );
  XOR2_X1 _11439_ (
    .A(wb_reg_inst[10]),
    .B(ibuf_io_inst_0_bits_inst_rs2[3]),
    .Z(_03939_)
  );
  OR2_X1 _11440_ (
    .A1(_03938_),
    .A2(_03939_),
    .ZN(_03940_)
  );
  XOR2_X1 _11441_ (
    .A(wb_reg_inst[9]),
    .B(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03941_)
  );
  XOR2_X1 _11442_ (
    .A(wb_reg_inst[11]),
    .B(ibuf_io_inst_0_bits_inst_rs2[4]),
    .Z(_03942_)
  );
  XOR2_X1 _11443_ (
    .A(wb_reg_inst[8]),
    .B(ibuf_io_inst_0_bits_inst_rs2[1]),
    .Z(_03943_)
  );
  OR2_X1 _11444_ (
    .A1(_03942_),
    .A2(_03943_),
    .ZN(_03944_)
  );
  OR2_X1 _11445_ (
    .A1(_03941_),
    .A2(_03944_),
    .ZN(_03945_)
  );
  OR2_X1 _11446_ (
    .A1(_03940_),
    .A2(_03945_),
    .ZN(_03946_)
  );
  INV_X1 _11447_ (
    .A(_03946_),
    .ZN(_03947_)
  );
  AND2_X1 _11448_ (
    .A1(_03812_),
    .A2(_03947_),
    .ZN(_03948_)
  );
  AND2_X1 _11449_ (
    .A1(_03028_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[3]),
    .ZN(_03949_)
  );
  AND2_X1 _11450_ (
    .A1(wb_reg_inst[9]),
    .A2(_03046_),
    .ZN(_03950_)
  );
  AND2_X1 _11451_ (
    .A1(_03027_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_03951_)
  );
  XOR2_X1 _11452_ (
    .A(wb_reg_inst[11]),
    .B(ibuf_io_inst_0_bits_inst_rs1[4]),
    .Z(_03952_)
  );
  XOR2_X1 _11453_ (
    .A(wb_reg_inst[7]),
    .B(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_03953_)
  );
  AND2_X1 _11454_ (
    .A1(wb_reg_inst[10]),
    .A2(_03047_),
    .ZN(_03954_)
  );
  OR2_X1 _11455_ (
    .A1(_03950_),
    .A2(_03954_),
    .ZN(_03955_)
  );
  OR2_X1 _11456_ (
    .A1(_03953_),
    .A2(_03955_),
    .ZN(_03956_)
  );
  OR2_X1 _11457_ (
    .A1(_03949_),
    .A2(_03951_),
    .ZN(_03957_)
  );
  XOR2_X1 _11458_ (
    .A(wb_reg_inst[8]),
    .B(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_03958_)
  );
  OR2_X1 _11459_ (
    .A1(_03952_),
    .A2(_03958_),
    .ZN(_03959_)
  );
  OR2_X1 _11460_ (
    .A1(_03957_),
    .A2(_03959_),
    .ZN(_03960_)
  );
  OR2_X1 _11461_ (
    .A1(_03956_),
    .A2(_03960_),
    .ZN(_03961_)
  );
  INV_X1 _11462_ (
    .A(_03961_),
    .ZN(_03962_)
  );
  AND2_X1 _11463_ (
    .A1(_03703_),
    .A2(_03962_),
    .ZN(_03963_)
  );
  OR2_X1 _11464_ (
    .A1(_03948_),
    .A2(_03963_),
    .ZN(_03964_)
  );
  AND2_X1 _11465_ (
    .A1(_03028_),
    .A2(ibuf_io_inst_0_bits_inst_rd[3]),
    .ZN(_03965_)
  );
  AND2_X1 _11466_ (
    .A1(_03026_),
    .A2(ibuf_io_inst_0_bits_inst_rd[1]),
    .ZN(_03966_)
  );
  OR2_X1 _11467_ (
    .A1(_03965_),
    .A2(_03966_),
    .ZN(_03967_)
  );
  XOR2_X1 _11468_ (
    .A(wb_reg_inst[11]),
    .B(ibuf_io_inst_0_bits_inst_rd[4]),
    .Z(_03968_)
  );
  OR2_X1 _11469_ (
    .A1(_03967_),
    .A2(_03968_),
    .ZN(_03969_)
  );
  XOR2_X1 _11470_ (
    .A(wb_reg_inst[9]),
    .B(ibuf_io_inst_0_bits_inst_rd[2]),
    .Z(_03970_)
  );
  XOR2_X1 _11471_ (
    .A(wb_reg_inst[7]),
    .B(ibuf_io_inst_0_bits_inst_rd[0]),
    .Z(_03971_)
  );
  AND2_X1 _11472_ (
    .A1(wb_reg_inst[8]),
    .A2(_03053_),
    .ZN(_03972_)
  );
  AND2_X1 _11473_ (
    .A1(wb_reg_inst[10]),
    .A2(_03055_),
    .ZN(_03973_)
  );
  OR2_X1 _11474_ (
    .A1(_03972_),
    .A2(_03973_),
    .ZN(_03974_)
  );
  OR2_X1 _11475_ (
    .A1(_03971_),
    .A2(_03974_),
    .ZN(_03975_)
  );
  OR2_X1 _11476_ (
    .A1(_03970_),
    .A2(_03975_),
    .ZN(_03976_)
  );
  OR2_X1 _11477_ (
    .A1(_03969_),
    .A2(_03976_),
    .ZN(_03977_)
  );
  INV_X1 _11478_ (
    .A(_03977_),
    .ZN(_03978_)
  );
  AND2_X1 _11479_ (
    .A1(_03606_),
    .A2(_03978_),
    .ZN(_03979_)
  );
  OR2_X1 _11480_ (
    .A1(_03964_),
    .A2(_03979_),
    .ZN(_03980_)
  );
  AND2_X1 _11481_ (
    .A1(_03937_),
    .A2(_03980_),
    .ZN(_03981_)
  );
  OR2_X1 _11482_ (
    .A1(ex_ctrl_csr[0]),
    .A2(ex_ctrl_csr[1]),
    .ZN(_03982_)
  );
  OR2_X1 _11483_ (
    .A1(ex_ctrl_csr[2]),
    .A2(ex_ctrl_jalr),
    .ZN(_03983_)
  );
  OR2_X1 _11484_ (
    .A1(ex_ctrl_div),
    .A2(ex_ctrl_mem),
    .ZN(_03984_)
  );
  OR2_X1 _11485_ (
    .A1(_03982_),
    .A2(_03984_),
    .ZN(_03985_)
  );
  OR2_X1 _11486_ (
    .A1(_03983_),
    .A2(_03985_),
    .ZN(_03986_)
  );
  AND2_X1 _11487_ (
    .A1(_03452_),
    .A2(_03986_),
    .ZN(_03987_)
  );
  AND2_X1 _11488_ (
    .A1(_03466_),
    .A2(_03703_),
    .ZN(_03988_)
  );
  OR2_X1 _11489_ (
    .A1(_02985_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_03989_)
  );
  OR2_X1 _11490_ (
    .A1(_02990_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[4]),
    .ZN(_03990_)
  );
  AND2_X1 _11491_ (
    .A1(_03989_),
    .A2(_03990_),
    .ZN(_03991_)
  );
  OR2_X1 _11492_ (
    .A1(ex_reg_inst[8]),
    .A2(_03049_),
    .ZN(_03992_)
  );
  OR2_X1 _11493_ (
    .A1(ex_reg_inst[11]),
    .A2(_03064_),
    .ZN(_03993_)
  );
  AND2_X1 _11494_ (
    .A1(_03992_),
    .A2(_03993_),
    .ZN(_03994_)
  );
  AND2_X1 _11495_ (
    .A1(_03991_),
    .A2(_03994_),
    .ZN(_03995_)
  );
  XOR2_X1 _11496_ (
    .A(ex_reg_inst[7]),
    .B(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_03996_)
  );
  XOR2_X1 _11497_ (
    .A(ex_reg_inst[9]),
    .B(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_03997_)
  );
  XOR2_X1 _11498_ (
    .A(ex_reg_inst[10]),
    .B(ibuf_io_inst_0_bits_inst_rs2[3]),
    .Z(_03998_)
  );
  OR2_X1 _11499_ (
    .A1(_03997_),
    .A2(_03998_),
    .ZN(_03999_)
  );
  OR2_X1 _11500_ (
    .A1(_03996_),
    .A2(_03999_),
    .ZN(_04000_)
  );
  INV_X1 _11501_ (
    .A(_04000_),
    .ZN(_04001_)
  );
  AND2_X1 _11502_ (
    .A1(_03995_),
    .A2(_04001_),
    .ZN(_04002_)
  );
  AND2_X1 _11503_ (
    .A1(_03812_),
    .A2(_04002_),
    .ZN(_04003_)
  );
  XOR2_X1 _11504_ (
    .A(ex_reg_inst[11]),
    .B(ibuf_io_inst_0_bits_inst_rd[4]),
    .Z(_04004_)
  );
  AND2_X1 _11505_ (
    .A1(_02988_),
    .A2(ibuf_io_inst_0_bits_inst_rd[3]),
    .ZN(_04005_)
  );
  AND2_X1 _11506_ (
    .A1(_02983_),
    .A2(ibuf_io_inst_0_bits_inst_rd[0]),
    .ZN(_04006_)
  );
  OR2_X1 _11507_ (
    .A1(_04005_),
    .A2(_04006_),
    .ZN(_04007_)
  );
  OR2_X1 _11508_ (
    .A1(_04004_),
    .A2(_04007_),
    .ZN(_04008_)
  );
  XOR2_X1 _11509_ (
    .A(ex_reg_inst[9]),
    .B(ibuf_io_inst_0_bits_inst_rd[2]),
    .Z(_04009_)
  );
  XOR2_X1 _11510_ (
    .A(ex_reg_inst[8]),
    .B(ibuf_io_inst_0_bits_inst_rd[1]),
    .Z(_04010_)
  );
  AND2_X1 _11511_ (
    .A1(ex_reg_inst[10]),
    .A2(_03055_),
    .ZN(_04011_)
  );
  AND2_X1 _11512_ (
    .A1(ex_reg_inst[7]),
    .A2(_03052_),
    .ZN(_04012_)
  );
  OR2_X1 _11513_ (
    .A1(_04011_),
    .A2(_04012_),
    .ZN(_04013_)
  );
  OR2_X1 _11514_ (
    .A1(_04010_),
    .A2(_04013_),
    .ZN(_04014_)
  );
  OR2_X1 _11515_ (
    .A1(_04009_),
    .A2(_04014_),
    .ZN(_04015_)
  );
  OR2_X1 _11516_ (
    .A1(_04008_),
    .A2(_04015_),
    .ZN(_04016_)
  );
  INV_X1 _11517_ (
    .A(_04016_),
    .ZN(_04017_)
  );
  AND2_X1 _11518_ (
    .A1(_03606_),
    .A2(_04017_),
    .ZN(_04018_)
  );
  OR2_X1 _11519_ (
    .A1(_04003_),
    .A2(_04018_),
    .ZN(_04019_)
  );
  OR2_X1 _11520_ (
    .A1(_03988_),
    .A2(_04019_),
    .ZN(_04020_)
  );
  AND2_X1 _11521_ (
    .A1(_03987_),
    .A2(_04020_),
    .ZN(_04021_)
  );
  OR2_X1 _11522_ (
    .A1(_03981_),
    .A2(_04021_),
    .ZN(_04022_)
  );
  INV_X1 _11523_ (
    .A(_04022_),
    .ZN(_04023_)
  );
  AND2_X1 _11524_ (
    .A1(_03936_),
    .A2(_04023_),
    .ZN(ibuf_io_inst_0_ready)
  );
  INV_X1 _11525_ (
    .A(ibuf_io_inst_0_ready),
    .ZN(_04024_)
  );
  AND2_X1 _11526_ (
    .A1(_03090_),
    .A2(_03140_),
    .ZN(_04025_)
  );
  OR2_X1 _11527_ (
    .A1(csr_io_eret),
    .A2(csr_io_exception),
    .ZN(_04026_)
  );
  OR2_X1 _11528_ (
    .A1(wb_reg_flush_pipe),
    .A2(_03142_),
    .ZN(_04027_)
  );
  INV_X1 _11529_ (
    .A(_04027_),
    .ZN(_04028_)
  );
  AND2_X1 _11530_ (
    .A1(_04025_),
    .A2(_04028_),
    .ZN(io_imem_req_bits_speculative)
  );
  INV_X1 _11531_ (
    .A(io_imem_req_bits_speculative),
    .ZN(_04029_)
  );
  AND2_X1 _11532_ (
    .A1(mem_br_taken),
    .A2(mem_ctrl_branch),
    .ZN(_04030_)
  );
  OR2_X1 _11533_ (
    .A1(mem_ctrl_jal),
    .A2(_04030_),
    .ZN(_04031_)
  );
  OR2_X1 _11534_ (
    .A1(mem_ctrl_jalr),
    .A2(_04031_),
    .ZN(_04032_)
  );
  AND2_X1 _11535_ (
    .A1(mem_reg_valid),
    .A2(_take_pc_mem_T),
    .ZN(_04033_)
  );
  AND2_X1 _11536_ (
    .A1(_04032_),
    .A2(_04033_),
    .ZN(_04034_)
  );
  INV_X1 _11537_ (
    .A(_04034_),
    .ZN(_04035_)
  );
  AND2_X1 _11538_ (
    .A1(io_imem_req_bits_speculative),
    .A2(_04035_),
    .ZN(_04036_)
  );
  INV_X1 _11539_ (
    .A(_04036_),
    .ZN(ibuf_io_kill)
  );
  AND2_X1 _11540_ (
    .A1(ibuf_io_inst_0_valid),
    .A2(_04036_),
    .ZN(_04037_)
  );
  INV_X1 _11541_ (
    .A(_04037_),
    .ZN(_04038_)
  );
  AND2_X1 _11542_ (
    .A1(ibuf_io_inst_0_ready),
    .A2(_04037_),
    .ZN(_04039_)
  );
  INV_X1 _11543_ (
    .A(_04039_),
    .ZN(_04040_)
  );
  OR2_X1 _11544_ (
    .A1(_03586_),
    .A2(_04040_),
    .ZN(_04041_)
  );
  INV_X1 _11545_ (
    .A(_04041_),
    .ZN(_ex_reg_valid_T)
  );
  AND2_X1 _11546_ (
    .A1(_03584_),
    .A2(_ex_reg_valid_T),
    .ZN(_04042_)
  );
  AND2_X1 _11547_ (
    .A1(ibuf_io_inst_0_bits_raw[2]),
    .A2(_03582_),
    .ZN(_04043_)
  );
  AND2_X1 _11548_ (
    .A1(_03490_),
    .A2(_03583_),
    .ZN(_04044_)
  );
  INV_X1 _11549_ (
    .A(_04044_),
    .ZN(_04045_)
  );
  OR2_X1 _11550_ (
    .A1(_03117_),
    .A2(_03144_),
    .ZN(_04046_)
  );
  MUX2_X1 _11551_ (
    .A(wb_reg_inst[8]),
    .B(_03103_),
    .S(_03117_),
    .Z(_04047_)
  );
  INV_X1 _11552_ (
    .A(_04047_),
    .ZN(_04048_)
  );
  MUX2_X1 _11553_ (
    .A(wb_reg_inst[7]),
    .B(_03101_),
    .S(_03117_),
    .Z(_04049_)
  );
  INV_X1 _11554_ (
    .A(_04049_),
    .ZN(_04050_)
  );
  OR2_X1 _11555_ (
    .A1(_04047_),
    .A2(_04049_),
    .ZN(_04051_)
  );
  MUX2_X1 _11556_ (
    .A(_03027_),
    .B(_03105_),
    .S(_03117_),
    .Z(_04052_)
  );
  MUX2_X1 _11557_ (
    .A(wb_reg_inst[9]),
    .B(_03106_),
    .S(_03117_),
    .Z(_04053_)
  );
  MUX2_X1 _11558_ (
    .A(wb_reg_inst[11]),
    .B(_03110_),
    .S(_03117_),
    .Z(_04054_)
  );
  INV_X1 _11559_ (
    .A(_04054_),
    .ZN(_04055_)
  );
  MUX2_X1 _11560_ (
    .A(wb_reg_inst[10]),
    .B(_03109_),
    .S(_03117_),
    .Z(_04056_)
  );
  INV_X1 _11561_ (
    .A(_04056_),
    .ZN(_04057_)
  );
  AND2_X1 _11562_ (
    .A1(_04055_),
    .A2(_04057_),
    .ZN(_04058_)
  );
  AND2_X1 _11563_ (
    .A1(_04052_),
    .A2(_04058_),
    .ZN(_04059_)
  );
  INV_X1 _11564_ (
    .A(_04059_),
    .ZN(_04060_)
  );
  OR2_X1 _11565_ (
    .A1(_04051_),
    .A2(_04060_),
    .ZN(_04061_)
  );
  AND2_X1 _11566_ (
    .A1(_04046_),
    .A2(_04061_),
    .ZN(_04062_)
  );
  INV_X1 _11567_ (
    .A(_04062_),
    .ZN(_04063_)
  );
  XOR2_X1 _11568_ (
    .A(ibuf_io_inst_0_bits_inst_rs1[4]),
    .B(_04054_),
    .Z(_04064_)
  );
  XOR2_X1 _11569_ (
    .A(_03046_),
    .B(_04052_),
    .Z(_04065_)
  );
  OR2_X1 _11570_ (
    .A1(_04064_),
    .A2(_04065_),
    .ZN(_04066_)
  );
  XOR2_X1 _11571_ (
    .A(ibuf_io_inst_0_bits_inst_rs1[1]),
    .B(_04047_),
    .Z(_04067_)
  );
  XOR2_X1 _11572_ (
    .A(ibuf_io_inst_0_bits_inst_rs1[3]),
    .B(_04056_),
    .Z(_04068_)
  );
  XOR2_X1 _11573_ (
    .A(ibuf_io_inst_0_bits_inst_rs1[0]),
    .B(_04049_),
    .Z(_04069_)
  );
  OR2_X1 _11574_ (
    .A1(_04068_),
    .A2(_04069_),
    .ZN(_04070_)
  );
  OR2_X1 _11575_ (
    .A1(_04067_),
    .A2(_04070_),
    .ZN(_04071_)
  );
  OR2_X1 _11576_ (
    .A1(_04066_),
    .A2(_04071_),
    .ZN(_04072_)
  );
  INV_X1 _11577_ (
    .A(_04072_),
    .ZN(_04073_)
  );
  AND2_X1 _11578_ (
    .A1(_04062_),
    .A2(_04073_),
    .ZN(_04074_)
  );
  OR2_X1 _11579_ (
    .A1(_04063_),
    .A2(_04072_),
    .ZN(_04075_)
  );
  OR2_X1 _11580_ (
    .A1(wb_ctrl_csr[0]),
    .A2(wb_ctrl_csr[1]),
    .ZN(_04076_)
  );
  OR2_X1 _11581_ (
    .A1(wb_ctrl_csr[2]),
    .A2(_04076_),
    .ZN(_04077_)
  );
  MUX2_X1 _11582_ (
    .A(wb_reg_wdata[2]),
    .B(csr_io_rw_rdata[2]),
    .S(_04077_),
    .Z(_04078_)
  );
  MUX2_X1 _11583_ (
    .A(div_io_resp_bits_data[2]),
    .B(_04078_),
    .S(_03114_),
    .Z(_04079_)
  );
  MUX2_X1 _11584_ (
    .A(_04079_),
    .B(io_dmem_resp_bits_data[2]),
    .S(_03097_),
    .Z(_04080_)
  );
  OR2_X1 _11585_ (
    .A1(\rf[26] [2]),
    .A2(_03046_),
    .ZN(_04081_)
  );
  OR2_X1 _11586_ (
    .A1(\rf[30] [2]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04082_)
  );
  AND2_X1 _11587_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04082_),
    .ZN(_04083_)
  );
  AND2_X1 _11588_ (
    .A1(_04081_),
    .A2(_04083_),
    .ZN(_04084_)
  );
  AND2_X1 _11589_ (
    .A1(\rf[27] [2]),
    .A2(_03760_),
    .ZN(_04085_)
  );
  OR2_X1 _11590_ (
    .A1(_04084_),
    .A2(_04085_),
    .ZN(_04086_)
  );
  MUX2_X1 _11591_ (
    .A(\rf[23] [2]),
    .B(\rf[19] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04087_)
  );
  AND2_X1 _11592_ (
    .A1(_03044_),
    .A2(_04087_),
    .ZN(_04088_)
  );
  OR2_X1 _11593_ (
    .A1(\rf[22] [2]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04089_)
  );
  OR2_X1 _11594_ (
    .A1(\rf[18] [2]),
    .A2(_03046_),
    .ZN(_04090_)
  );
  AND2_X1 _11595_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04090_),
    .ZN(_04091_)
  );
  AND2_X1 _11596_ (
    .A1(_04089_),
    .A2(_04091_),
    .ZN(_04092_)
  );
  OR2_X1 _11597_ (
    .A1(_03047_),
    .A2(_04092_),
    .ZN(_04093_)
  );
  OR2_X1 _11598_ (
    .A1(_04088_),
    .A2(_04093_),
    .ZN(_04094_)
  );
  OR2_X1 _11599_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_04086_),
    .ZN(_04095_)
  );
  AND2_X1 _11600_ (
    .A1(_03045_),
    .A2(_04095_),
    .ZN(_04096_)
  );
  AND2_X1 _11601_ (
    .A1(_04094_),
    .A2(_04096_),
    .ZN(_04097_)
  );
  MUX2_X1 _11602_ (
    .A(\rf[21] [2]),
    .B(\rf[17] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04098_)
  );
  AND2_X1 _11603_ (
    .A1(_03044_),
    .A2(_04098_),
    .ZN(_04099_)
  );
  OR2_X1 _11604_ (
    .A1(\rf[20] [2]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04100_)
  );
  OR2_X1 _11605_ (
    .A1(\rf[16] [2]),
    .A2(_03046_),
    .ZN(_04101_)
  );
  AND2_X1 _11606_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04100_),
    .ZN(_04102_)
  );
  AND2_X1 _11607_ (
    .A1(_04101_),
    .A2(_04102_),
    .ZN(_04103_)
  );
  OR2_X1 _11608_ (
    .A1(_03047_),
    .A2(_04099_),
    .ZN(_04104_)
  );
  OR2_X1 _11609_ (
    .A1(_04103_),
    .A2(_04104_),
    .ZN(_04105_)
  );
  OR2_X1 _11610_ (
    .A1(\rf[24] [2]),
    .A2(_03046_),
    .ZN(_04106_)
  );
  OR2_X1 _11611_ (
    .A1(\rf[28] [2]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04107_)
  );
  AND2_X1 _11612_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04107_),
    .ZN(_04108_)
  );
  AND2_X1 _11613_ (
    .A1(_04106_),
    .A2(_04108_),
    .ZN(_04109_)
  );
  MUX2_X1 _11614_ (
    .A(\rf[29] [2]),
    .B(\rf[25] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04110_)
  );
  AND2_X1 _11615_ (
    .A1(_03044_),
    .A2(_04110_),
    .ZN(_04111_)
  );
  OR2_X1 _11616_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_04111_),
    .ZN(_04112_)
  );
  OR2_X1 _11617_ (
    .A1(_04109_),
    .A2(_04112_),
    .ZN(_04113_)
  );
  AND2_X1 _11618_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04113_),
    .ZN(_04114_)
  );
  AND2_X1 _11619_ (
    .A1(_04105_),
    .A2(_04114_),
    .ZN(_04115_)
  );
  OR2_X1 _11620_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_04115_),
    .ZN(_04116_)
  );
  OR2_X1 _11621_ (
    .A1(_04097_),
    .A2(_04116_),
    .ZN(_04117_)
  );
  MUX2_X1 _11622_ (
    .A(\rf[1] [2]),
    .B(\rf[0] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_04118_)
  );
  MUX2_X1 _11623_ (
    .A(\rf[5] [2]),
    .B(\rf[4] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_04119_)
  );
  MUX2_X1 _11624_ (
    .A(_04118_),
    .B(_04119_),
    .S(_03046_),
    .Z(_04120_)
  );
  OR2_X1 _11625_ (
    .A1(_03047_),
    .A2(_04120_),
    .ZN(_04121_)
  );
  MUX2_X1 _11626_ (
    .A(\rf[13] [2]),
    .B(\rf[9] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04122_)
  );
  OR2_X1 _11627_ (
    .A1(_03448_),
    .A2(_04122_),
    .ZN(_04123_)
  );
  OR2_X1 _11628_ (
    .A1(_03044_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[3]),
    .ZN(_04124_)
  );
  MUX2_X1 _11629_ (
    .A(\rf[12] [2]),
    .B(\rf[8] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04125_)
  );
  OR2_X1 _11630_ (
    .A1(_04124_),
    .A2(_04125_),
    .ZN(_04126_)
  );
  AND2_X1 _11631_ (
    .A1(_04123_),
    .A2(_04126_),
    .ZN(_04127_)
  );
  AND2_X1 _11632_ (
    .A1(_04121_),
    .A2(_04127_),
    .ZN(_04128_)
  );
  MUX2_X1 _11633_ (
    .A(\rf[3] [2]),
    .B(\rf[2] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_04129_)
  );
  MUX2_X1 _11634_ (
    .A(\rf[7] [2]),
    .B(\rf[6] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_04130_)
  );
  MUX2_X1 _11635_ (
    .A(_04129_),
    .B(_04130_),
    .S(_03046_),
    .Z(_04131_)
  );
  OR2_X1 _11636_ (
    .A1(_03047_),
    .A2(_04131_),
    .ZN(_04132_)
  );
  MUX2_X1 _11637_ (
    .A(\rf[14] [2]),
    .B(\rf[10] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04133_)
  );
  OR2_X1 _11638_ (
    .A1(_04124_),
    .A2(_04133_),
    .ZN(_04134_)
  );
  MUX2_X1 _11639_ (
    .A(\rf[15] [2]),
    .B(\rf[11] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04135_)
  );
  OR2_X1 _11640_ (
    .A1(_03448_),
    .A2(_04135_),
    .ZN(_04136_)
  );
  AND2_X1 _11641_ (
    .A1(_04134_),
    .A2(_04136_),
    .ZN(_04137_)
  );
  AND2_X1 _11642_ (
    .A1(_04132_),
    .A2(_04137_),
    .ZN(_04138_)
  );
  MUX2_X1 _11643_ (
    .A(_04128_),
    .B(_04138_),
    .S(_03045_),
    .Z(_04139_)
  );
  OR2_X1 _11644_ (
    .A1(_03063_),
    .A2(_04139_),
    .ZN(_04140_)
  );
  AND2_X1 _11645_ (
    .A1(_04117_),
    .A2(_04140_),
    .ZN(_04141_)
  );
  MUX2_X1 _11646_ (
    .A(_04141_),
    .B(_04080_),
    .S(_04074_),
    .Z(_04142_)
  );
  AND2_X1 _11647_ (
    .A1(_04044_),
    .A2(_04142_),
    .ZN(_04143_)
  );
  OR2_X1 _11648_ (
    .A1(_04043_),
    .A2(_04143_),
    .ZN(_04144_)
  );
  OR2_X1 _11649_ (
    .A1(_03586_),
    .A2(_04038_),
    .ZN(_04145_)
  );
  OR2_X1 _11650_ (
    .A1(_04024_),
    .A2(_04145_),
    .ZN(_04146_)
  );
  MUX2_X1 _11651_ (
    .A(ex_reg_rs_msb_0[0]),
    .B(_04144_),
    .S(_04042_),
    .Z(_00067_)
  );
  AND2_X1 _11652_ (
    .A1(ibuf_io_inst_0_bits_raw[3]),
    .A2(_03582_),
    .ZN(_04147_)
  );
  MUX2_X1 _11653_ (
    .A(wb_reg_wdata[3]),
    .B(csr_io_rw_rdata[3]),
    .S(_04077_),
    .Z(_04148_)
  );
  MUX2_X1 _11654_ (
    .A(div_io_resp_bits_data[3]),
    .B(_04148_),
    .S(_03114_),
    .Z(_04149_)
  );
  MUX2_X1 _11655_ (
    .A(_04149_),
    .B(io_dmem_resp_bits_data[3]),
    .S(_03097_),
    .Z(_04150_)
  );
  MUX2_X1 _11656_ (
    .A(\rf[15] [3]),
    .B(\rf[11] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04151_)
  );
  OR2_X1 _11657_ (
    .A1(\rf[14] [3]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04152_)
  );
  OR2_X1 _11658_ (
    .A1(\rf[10] [3]),
    .A2(_03046_),
    .ZN(_04153_)
  );
  MUX2_X1 _11659_ (
    .A(\rf[13] [3]),
    .B(\rf[9] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04154_)
  );
  OR2_X1 _11660_ (
    .A1(\rf[8] [3]),
    .A2(_03046_),
    .ZN(_04155_)
  );
  OR2_X1 _11661_ (
    .A1(\rf[12] [3]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04156_)
  );
  AND2_X1 _11662_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04152_),
    .ZN(_04157_)
  );
  AND2_X1 _11663_ (
    .A1(_04153_),
    .A2(_04157_),
    .ZN(_04158_)
  );
  AND2_X1 _11664_ (
    .A1(_03044_),
    .A2(_04151_),
    .ZN(_04159_)
  );
  OR2_X1 _11665_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04159_),
    .ZN(_04160_)
  );
  OR2_X1 _11666_ (
    .A1(_04158_),
    .A2(_04160_),
    .ZN(_04161_)
  );
  AND2_X1 _11667_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04156_),
    .ZN(_04162_)
  );
  AND2_X1 _11668_ (
    .A1(_04155_),
    .A2(_04162_),
    .ZN(_04163_)
  );
  AND2_X1 _11669_ (
    .A1(_03044_),
    .A2(_04154_),
    .ZN(_04164_)
  );
  OR2_X1 _11670_ (
    .A1(_03045_),
    .A2(_04164_),
    .ZN(_04165_)
  );
  OR2_X1 _11671_ (
    .A1(_04163_),
    .A2(_04165_),
    .ZN(_04166_)
  );
  AND2_X1 _11672_ (
    .A1(_03047_),
    .A2(_04166_),
    .ZN(_04167_)
  );
  AND2_X1 _11673_ (
    .A1(_04161_),
    .A2(_04167_),
    .ZN(_04168_)
  );
  OR2_X1 _11674_ (
    .A1(\rf[0] [3]),
    .A2(_03046_),
    .ZN(_04169_)
  );
  OR2_X1 _11675_ (
    .A1(\rf[4] [3]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04170_)
  );
  AND2_X1 _11676_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04170_),
    .ZN(_04171_)
  );
  AND2_X1 _11677_ (
    .A1(_04169_),
    .A2(_04171_),
    .ZN(_04172_)
  );
  MUX2_X1 _11678_ (
    .A(\rf[5] [3]),
    .B(\rf[1] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04173_)
  );
  AND2_X1 _11679_ (
    .A1(_03044_),
    .A2(_04173_),
    .ZN(_04174_)
  );
  OR2_X1 _11680_ (
    .A1(_03045_),
    .A2(_04174_),
    .ZN(_04175_)
  );
  OR2_X1 _11681_ (
    .A1(_04172_),
    .A2(_04175_),
    .ZN(_04176_)
  );
  MUX2_X1 _11682_ (
    .A(\rf[7] [3]),
    .B(\rf[3] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04177_)
  );
  AND2_X1 _11683_ (
    .A1(_03044_),
    .A2(_04177_),
    .ZN(_04178_)
  );
  OR2_X1 _11684_ (
    .A1(\rf[2] [3]),
    .A2(_03046_),
    .ZN(_04179_)
  );
  OR2_X1 _11685_ (
    .A1(\rf[6] [3]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04180_)
  );
  AND2_X1 _11686_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04180_),
    .ZN(_04181_)
  );
  AND2_X1 _11687_ (
    .A1(_04179_),
    .A2(_04181_),
    .ZN(_04182_)
  );
  OR2_X1 _11688_ (
    .A1(_04178_),
    .A2(_04182_),
    .ZN(_04183_)
  );
  OR2_X1 _11689_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04183_),
    .ZN(_04184_)
  );
  AND2_X1 _11690_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_04176_),
    .ZN(_04185_)
  );
  AND2_X1 _11691_ (
    .A1(_04184_),
    .A2(_04185_),
    .ZN(_04186_)
  );
  OR2_X1 _11692_ (
    .A1(_03063_),
    .A2(_04168_),
    .ZN(_04187_)
  );
  OR2_X1 _11693_ (
    .A1(_04186_),
    .A2(_04187_),
    .ZN(_04188_)
  );
  OR2_X1 _11694_ (
    .A1(\rf[26] [3]),
    .A2(_03046_),
    .ZN(_04189_)
  );
  OR2_X1 _11695_ (
    .A1(\rf[30] [3]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04190_)
  );
  AND2_X1 _11696_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04190_),
    .ZN(_04191_)
  );
  AND2_X1 _11697_ (
    .A1(_04189_),
    .A2(_04191_),
    .ZN(_04192_)
  );
  AND2_X1 _11698_ (
    .A1(\rf[27] [3]),
    .A2(_03760_),
    .ZN(_04193_)
  );
  OR2_X1 _11699_ (
    .A1(_04192_),
    .A2(_04193_),
    .ZN(_04194_)
  );
  MUX2_X1 _11700_ (
    .A(\rf[29] [3]),
    .B(\rf[25] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04195_)
  );
  AND2_X1 _11701_ (
    .A1(_03044_),
    .A2(_04195_),
    .ZN(_04196_)
  );
  OR2_X1 _11702_ (
    .A1(\rf[28] [3]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04197_)
  );
  OR2_X1 _11703_ (
    .A1(\rf[24] [3]),
    .A2(_03046_),
    .ZN(_04198_)
  );
  AND2_X1 _11704_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04198_),
    .ZN(_04199_)
  );
  AND2_X1 _11705_ (
    .A1(_04197_),
    .A2(_04199_),
    .ZN(_04200_)
  );
  OR2_X1 _11706_ (
    .A1(_03045_),
    .A2(_04200_),
    .ZN(_04201_)
  );
  OR2_X1 _11707_ (
    .A1(_04196_),
    .A2(_04201_),
    .ZN(_04202_)
  );
  OR2_X1 _11708_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04194_),
    .ZN(_04203_)
  );
  AND2_X1 _11709_ (
    .A1(_03047_),
    .A2(_04203_),
    .ZN(_04204_)
  );
  AND2_X1 _11710_ (
    .A1(_04202_),
    .A2(_04204_),
    .ZN(_04205_)
  );
  MUX2_X1 _11711_ (
    .A(\rf[21] [3]),
    .B(\rf[17] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04206_)
  );
  AND2_X1 _11712_ (
    .A1(_03044_),
    .A2(_04206_),
    .ZN(_04207_)
  );
  OR2_X1 _11713_ (
    .A1(\rf[20] [3]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04208_)
  );
  OR2_X1 _11714_ (
    .A1(\rf[16] [3]),
    .A2(_03046_),
    .ZN(_04209_)
  );
  AND2_X1 _11715_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04208_),
    .ZN(_04210_)
  );
  AND2_X1 _11716_ (
    .A1(_04209_),
    .A2(_04210_),
    .ZN(_04211_)
  );
  OR2_X1 _11717_ (
    .A1(_03045_),
    .A2(_04207_),
    .ZN(_04212_)
  );
  OR2_X1 _11718_ (
    .A1(_04211_),
    .A2(_04212_),
    .ZN(_04213_)
  );
  OR2_X1 _11719_ (
    .A1(\rf[18] [3]),
    .A2(_03046_),
    .ZN(_04214_)
  );
  OR2_X1 _11720_ (
    .A1(\rf[22] [3]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04215_)
  );
  AND2_X1 _11721_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04215_),
    .ZN(_04216_)
  );
  AND2_X1 _11722_ (
    .A1(_04214_),
    .A2(_04216_),
    .ZN(_04217_)
  );
  MUX2_X1 _11723_ (
    .A(\rf[23] [3]),
    .B(\rf[19] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04218_)
  );
  AND2_X1 _11724_ (
    .A1(_03044_),
    .A2(_04218_),
    .ZN(_04219_)
  );
  OR2_X1 _11725_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04219_),
    .ZN(_04220_)
  );
  OR2_X1 _11726_ (
    .A1(_04217_),
    .A2(_04220_),
    .ZN(_04221_)
  );
  AND2_X1 _11727_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_04221_),
    .ZN(_04222_)
  );
  AND2_X1 _11728_ (
    .A1(_04213_),
    .A2(_04222_),
    .ZN(_04223_)
  );
  OR2_X1 _11729_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_04223_),
    .ZN(_04224_)
  );
  OR2_X1 _11730_ (
    .A1(_04205_),
    .A2(_04224_),
    .ZN(_04225_)
  );
  AND2_X1 _11731_ (
    .A1(_04188_),
    .A2(_04225_),
    .ZN(_04226_)
  );
  MUX2_X1 _11732_ (
    .A(_04226_),
    .B(_04150_),
    .S(_04074_),
    .Z(_04227_)
  );
  AND2_X1 _11733_ (
    .A1(_04044_),
    .A2(_04227_),
    .ZN(_04228_)
  );
  OR2_X1 _11734_ (
    .A1(_04147_),
    .A2(_04228_),
    .ZN(_04229_)
  );
  MUX2_X1 _11735_ (
    .A(ex_reg_rs_msb_0[1]),
    .B(_04229_),
    .S(_04042_),
    .Z(_00068_)
  );
  AND2_X1 _11736_ (
    .A1(ibuf_io_inst_0_bits_raw[4]),
    .A2(_03582_),
    .ZN(_04230_)
  );
  MUX2_X1 _11737_ (
    .A(wb_reg_wdata[4]),
    .B(csr_io_rw_rdata[4]),
    .S(_04077_),
    .Z(_04231_)
  );
  MUX2_X1 _11738_ (
    .A(div_io_resp_bits_data[4]),
    .B(_04231_),
    .S(_03114_),
    .Z(_04232_)
  );
  MUX2_X1 _11739_ (
    .A(_04232_),
    .B(io_dmem_resp_bits_data[4]),
    .S(_03097_),
    .Z(_04233_)
  );
  MUX2_X1 _11740_ (
    .A(\rf[3] [4]),
    .B(\rf[1] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_04234_)
  );
  MUX2_X1 _11741_ (
    .A(\rf[7] [4]),
    .B(\rf[5] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_04235_)
  );
  MUX2_X1 _11742_ (
    .A(_04234_),
    .B(_04235_),
    .S(_03046_),
    .Z(_04236_)
  );
  AND2_X1 _11743_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_04236_),
    .ZN(_04237_)
  );
  MUX2_X1 _11744_ (
    .A(\rf[13] [4]),
    .B(\rf[9] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04238_)
  );
  OR2_X1 _11745_ (
    .A1(_03045_),
    .A2(_04238_),
    .ZN(_04239_)
  );
  MUX2_X1 _11746_ (
    .A(\rf[15] [4]),
    .B(\rf[11] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04240_)
  );
  OR2_X1 _11747_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04240_),
    .ZN(_04241_)
  );
  AND2_X1 _11748_ (
    .A1(_03047_),
    .A2(_04241_),
    .ZN(_04242_)
  );
  AND2_X1 _11749_ (
    .A1(_04239_),
    .A2(_04242_),
    .ZN(_04243_)
  );
  OR2_X1 _11750_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04243_),
    .ZN(_04244_)
  );
  OR2_X1 _11751_ (
    .A1(_04237_),
    .A2(_04244_),
    .ZN(_04245_)
  );
  MUX2_X1 _11752_ (
    .A(\rf[2] [4]),
    .B(\rf[0] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_04246_)
  );
  MUX2_X1 _11753_ (
    .A(\rf[6] [4]),
    .B(\rf[4] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_04247_)
  );
  MUX2_X1 _11754_ (
    .A(_04246_),
    .B(_04247_),
    .S(_03046_),
    .Z(_04248_)
  );
  AND2_X1 _11755_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_04248_),
    .ZN(_04249_)
  );
  MUX2_X1 _11756_ (
    .A(\rf[12] [4]),
    .B(\rf[8] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04250_)
  );
  OR2_X1 _11757_ (
    .A1(_03045_),
    .A2(_04250_),
    .ZN(_04251_)
  );
  MUX2_X1 _11758_ (
    .A(\rf[14] [4]),
    .B(\rf[10] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04252_)
  );
  OR2_X1 _11759_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04252_),
    .ZN(_04253_)
  );
  AND2_X1 _11760_ (
    .A1(_03047_),
    .A2(_04253_),
    .ZN(_04254_)
  );
  AND2_X1 _11761_ (
    .A1(_04251_),
    .A2(_04254_),
    .ZN(_04255_)
  );
  OR2_X1 _11762_ (
    .A1(_03044_),
    .A2(_04255_),
    .ZN(_04256_)
  );
  OR2_X1 _11763_ (
    .A1(_04249_),
    .A2(_04256_),
    .ZN(_04257_)
  );
  AND2_X1 _11764_ (
    .A1(_04245_),
    .A2(_04257_),
    .ZN(_04258_)
  );
  AND2_X1 _11765_ (
    .A1(\rf[21] [4]),
    .A2(_03046_),
    .ZN(_04259_)
  );
  AND2_X1 _11766_ (
    .A1(\rf[17] [4]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04260_)
  );
  OR2_X1 _11767_ (
    .A1(_03045_),
    .A2(_04260_),
    .ZN(_04261_)
  );
  OR2_X1 _11768_ (
    .A1(_04259_),
    .A2(_04261_),
    .ZN(_04262_)
  );
  AND2_X1 _11769_ (
    .A1(\rf[19] [4]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04263_)
  );
  AND2_X1 _11770_ (
    .A1(\rf[23] [4]),
    .A2(_03046_),
    .ZN(_04264_)
  );
  OR2_X1 _11771_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04264_),
    .ZN(_04265_)
  );
  OR2_X1 _11772_ (
    .A1(_04263_),
    .A2(_04265_),
    .ZN(_04266_)
  );
  AND2_X1 _11773_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_04266_),
    .ZN(_04267_)
  );
  AND2_X1 _11774_ (
    .A1(_04262_),
    .A2(_04267_),
    .ZN(_04268_)
  );
  OR2_X1 _11775_ (
    .A1(\rf[25] [4]),
    .A2(_03046_),
    .ZN(_04269_)
  );
  OR2_X1 _11776_ (
    .A1(\rf[29] [4]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04270_)
  );
  AND2_X1 _11777_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04270_),
    .ZN(_04271_)
  );
  AND2_X1 _11778_ (
    .A1(_04269_),
    .A2(_04271_),
    .ZN(_04272_)
  );
  AND2_X1 _11779_ (
    .A1(_03045_),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04273_)
  );
  AND2_X1 _11780_ (
    .A1(\rf[27] [4]),
    .A2(_04273_),
    .ZN(_04274_)
  );
  OR2_X1 _11781_ (
    .A1(_04272_),
    .A2(_04274_),
    .ZN(_04275_)
  );
  AND2_X1 _11782_ (
    .A1(_03047_),
    .A2(_04275_),
    .ZN(_04276_)
  );
  OR2_X1 _11783_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04276_),
    .ZN(_04277_)
  );
  OR2_X1 _11784_ (
    .A1(_04268_),
    .A2(_04277_),
    .ZN(_04278_)
  );
  MUX2_X1 _11785_ (
    .A(\rf[30] [4]),
    .B(\rf[26] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04279_)
  );
  OR2_X1 _11786_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04279_),
    .ZN(_04280_)
  );
  MUX2_X1 _11787_ (
    .A(\rf[28] [4]),
    .B(\rf[24] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04281_)
  );
  OR2_X1 _11788_ (
    .A1(_03045_),
    .A2(_04281_),
    .ZN(_04282_)
  );
  AND2_X1 _11789_ (
    .A1(_03047_),
    .A2(_04282_),
    .ZN(_04283_)
  );
  AND2_X1 _11790_ (
    .A1(_04280_),
    .A2(_04283_),
    .ZN(_04284_)
  );
  AND2_X1 _11791_ (
    .A1(\rf[16] [4]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04285_)
  );
  AND2_X1 _11792_ (
    .A1(\rf[20] [4]),
    .A2(_03046_),
    .ZN(_04286_)
  );
  OR2_X1 _11793_ (
    .A1(_03045_),
    .A2(_04286_),
    .ZN(_04287_)
  );
  OR2_X1 _11794_ (
    .A1(_04285_),
    .A2(_04287_),
    .ZN(_04288_)
  );
  AND2_X1 _11795_ (
    .A1(\rf[18] [4]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04289_)
  );
  AND2_X1 _11796_ (
    .A1(\rf[22] [4]),
    .A2(_03046_),
    .ZN(_04290_)
  );
  OR2_X1 _11797_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04290_),
    .ZN(_04291_)
  );
  OR2_X1 _11798_ (
    .A1(_04289_),
    .A2(_04291_),
    .ZN(_04292_)
  );
  AND2_X1 _11799_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_04292_),
    .ZN(_04293_)
  );
  AND2_X1 _11800_ (
    .A1(_04288_),
    .A2(_04293_),
    .ZN(_04294_)
  );
  OR2_X1 _11801_ (
    .A1(_03044_),
    .A2(_04294_),
    .ZN(_04295_)
  );
  OR2_X1 _11802_ (
    .A1(_04284_),
    .A2(_04295_),
    .ZN(_04296_)
  );
  AND2_X1 _11803_ (
    .A1(_04278_),
    .A2(_04296_),
    .ZN(_04297_)
  );
  MUX2_X1 _11804_ (
    .A(_04258_),
    .B(_04297_),
    .S(_03063_),
    .Z(_04298_)
  );
  MUX2_X1 _11805_ (
    .A(_04298_),
    .B(_04233_),
    .S(_04074_),
    .Z(_04299_)
  );
  AND2_X1 _11806_ (
    .A1(_04044_),
    .A2(_04299_),
    .ZN(_04300_)
  );
  OR2_X1 _11807_ (
    .A1(_04230_),
    .A2(_04300_),
    .ZN(_04301_)
  );
  MUX2_X1 _11808_ (
    .A(ex_reg_rs_msb_0[2]),
    .B(_04301_),
    .S(_04042_),
    .Z(_00069_)
  );
  AND2_X1 _11809_ (
    .A1(ibuf_io_inst_0_bits_raw[5]),
    .A2(_03582_),
    .ZN(_04302_)
  );
  MUX2_X1 _11810_ (
    .A(wb_reg_wdata[5]),
    .B(csr_io_rw_rdata[5]),
    .S(_04077_),
    .Z(_04303_)
  );
  MUX2_X1 _11811_ (
    .A(div_io_resp_bits_data[5]),
    .B(_04303_),
    .S(_03114_),
    .Z(_04304_)
  );
  MUX2_X1 _11812_ (
    .A(_04304_),
    .B(io_dmem_resp_bits_data[5]),
    .S(_03097_),
    .Z(_04305_)
  );
  MUX2_X1 _11813_ (
    .A(\rf[5] [5]),
    .B(\rf[1] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04306_)
  );
  MUX2_X1 _11814_ (
    .A(\rf[7] [5]),
    .B(\rf[3] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04307_)
  );
  MUX2_X1 _11815_ (
    .A(_04306_),
    .B(_04307_),
    .S(_03045_),
    .Z(_04308_)
  );
  AND2_X1 _11816_ (
    .A1(_03044_),
    .A2(_04308_),
    .ZN(_04309_)
  );
  MUX2_X1 _11817_ (
    .A(\rf[4] [5]),
    .B(\rf[0] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04310_)
  );
  MUX2_X1 _11818_ (
    .A(\rf[6] [5]),
    .B(\rf[2] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04311_)
  );
  MUX2_X1 _11819_ (
    .A(_04310_),
    .B(_04311_),
    .S(_03045_),
    .Z(_04312_)
  );
  AND2_X1 _11820_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04312_),
    .ZN(_04313_)
  );
  OR2_X1 _11821_ (
    .A1(_03063_),
    .A2(_04313_),
    .ZN(_04314_)
  );
  OR2_X1 _11822_ (
    .A1(_04309_),
    .A2(_04314_),
    .ZN(_04315_)
  );
  OR2_X1 _11823_ (
    .A1(\rf[20] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04316_)
  );
  OR2_X1 _11824_ (
    .A1(\rf[16] [5]),
    .A2(_03046_),
    .ZN(_04317_)
  );
  AND2_X1 _11825_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04317_),
    .ZN(_04318_)
  );
  AND2_X1 _11826_ (
    .A1(_04316_),
    .A2(_04318_),
    .ZN(_04319_)
  );
  MUX2_X1 _11827_ (
    .A(\rf[22] [5]),
    .B(\rf[18] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04320_)
  );
  AND2_X1 _11828_ (
    .A1(_03045_),
    .A2(_04320_),
    .ZN(_04321_)
  );
  OR2_X1 _11829_ (
    .A1(_03044_),
    .A2(_04321_),
    .ZN(_04322_)
  );
  OR2_X1 _11830_ (
    .A1(_04319_),
    .A2(_04322_),
    .ZN(_04323_)
  );
  OR2_X1 _11831_ (
    .A1(\rf[17] [5]),
    .A2(_03046_),
    .ZN(_04324_)
  );
  OR2_X1 _11832_ (
    .A1(\rf[21] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04325_)
  );
  AND2_X1 _11833_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04325_),
    .ZN(_04326_)
  );
  AND2_X1 _11834_ (
    .A1(_04324_),
    .A2(_04326_),
    .ZN(_04327_)
  );
  MUX2_X1 _11835_ (
    .A(\rf[23] [5]),
    .B(\rf[19] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04328_)
  );
  AND2_X1 _11836_ (
    .A1(_03045_),
    .A2(_04328_),
    .ZN(_04329_)
  );
  OR2_X1 _11837_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04329_),
    .ZN(_04330_)
  );
  OR2_X1 _11838_ (
    .A1(_04327_),
    .A2(_04330_),
    .ZN(_04331_)
  );
  AND2_X1 _11839_ (
    .A1(_04323_),
    .A2(_04331_),
    .ZN(_04332_)
  );
  OR2_X1 _11840_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_04332_),
    .ZN(_04333_)
  );
  AND2_X1 _11841_ (
    .A1(_04315_),
    .A2(_04333_),
    .ZN(_04334_)
  );
  AND2_X1 _11842_ (
    .A1(\rf[10] [5]),
    .A2(_03045_),
    .ZN(_04335_)
  );
  AND2_X1 _11843_ (
    .A1(\rf[8] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_04336_)
  );
  OR2_X1 _11844_ (
    .A1(_03046_),
    .A2(_04336_),
    .ZN(_04337_)
  );
  OR2_X1 _11845_ (
    .A1(_04335_),
    .A2(_04337_),
    .ZN(_04338_)
  );
  AND2_X1 _11846_ (
    .A1(\rf[14] [5]),
    .A2(_03045_),
    .ZN(_04339_)
  );
  AND2_X1 _11847_ (
    .A1(\rf[12] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_04340_)
  );
  OR2_X1 _11848_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_04340_),
    .ZN(_04341_)
  );
  OR2_X1 _11849_ (
    .A1(_04339_),
    .A2(_04341_),
    .ZN(_04342_)
  );
  AND2_X1 _11850_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04342_),
    .ZN(_04343_)
  );
  AND2_X1 _11851_ (
    .A1(_04338_),
    .A2(_04343_),
    .ZN(_04344_)
  );
  AND2_X1 _11852_ (
    .A1(\rf[11] [5]),
    .A2(_03045_),
    .ZN(_04345_)
  );
  AND2_X1 _11853_ (
    .A1(\rf[9] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_04346_)
  );
  OR2_X1 _11854_ (
    .A1(_03046_),
    .A2(_04346_),
    .ZN(_04347_)
  );
  OR2_X1 _11855_ (
    .A1(_04345_),
    .A2(_04347_),
    .ZN(_04348_)
  );
  AND2_X1 _11856_ (
    .A1(\rf[15] [5]),
    .A2(_03045_),
    .ZN(_04349_)
  );
  AND2_X1 _11857_ (
    .A1(\rf[13] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_04350_)
  );
  OR2_X1 _11858_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_04350_),
    .ZN(_04351_)
  );
  OR2_X1 _11859_ (
    .A1(_04349_),
    .A2(_04351_),
    .ZN(_04352_)
  );
  AND2_X1 _11860_ (
    .A1(_03044_),
    .A2(_04352_),
    .ZN(_04353_)
  );
  AND2_X1 _11861_ (
    .A1(_04348_),
    .A2(_04353_),
    .ZN(_04354_)
  );
  OR2_X1 _11862_ (
    .A1(_03063_),
    .A2(_04354_),
    .ZN(_04355_)
  );
  OR2_X1 _11863_ (
    .A1(_04344_),
    .A2(_04355_),
    .ZN(_04356_)
  );
  OR2_X1 _11864_ (
    .A1(\rf[28] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04357_)
  );
  OR2_X1 _11865_ (
    .A1(\rf[24] [5]),
    .A2(_03046_),
    .ZN(_04358_)
  );
  AND2_X1 _11866_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04357_),
    .ZN(_04359_)
  );
  AND2_X1 _11867_ (
    .A1(_04358_),
    .A2(_04359_),
    .ZN(_04360_)
  );
  MUX2_X1 _11868_ (
    .A(\rf[30] [5]),
    .B(\rf[26] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04361_)
  );
  AND2_X1 _11869_ (
    .A1(_03045_),
    .A2(_04361_),
    .ZN(_04362_)
  );
  OR2_X1 _11870_ (
    .A1(_03044_),
    .A2(_04362_),
    .ZN(_04363_)
  );
  OR2_X1 _11871_ (
    .A1(_04360_),
    .A2(_04363_),
    .ZN(_04364_)
  );
  MUX2_X1 _11872_ (
    .A(\rf[29] [5]),
    .B(\rf[25] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04365_)
  );
  AND2_X1 _11873_ (
    .A1(\rf[27] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04366_)
  );
  MUX2_X1 _11874_ (
    .A(_04365_),
    .B(_04366_),
    .S(_03045_),
    .Z(_04367_)
  );
  OR2_X1 _11875_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04367_),
    .ZN(_04368_)
  );
  AND2_X1 _11876_ (
    .A1(_04364_),
    .A2(_04368_),
    .ZN(_04369_)
  );
  OR2_X1 _11877_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_04369_),
    .ZN(_04370_)
  );
  AND2_X1 _11878_ (
    .A1(_04356_),
    .A2(_04370_),
    .ZN(_04371_)
  );
  MUX2_X1 _11879_ (
    .A(_04334_),
    .B(_04371_),
    .S(_03047_),
    .Z(_04372_)
  );
  MUX2_X1 _11880_ (
    .A(_04372_),
    .B(_04305_),
    .S(_04074_),
    .Z(_04373_)
  );
  AND2_X1 _11881_ (
    .A1(_04044_),
    .A2(_04373_),
    .ZN(_04374_)
  );
  OR2_X1 _11882_ (
    .A1(_04302_),
    .A2(_04374_),
    .ZN(_04375_)
  );
  MUX2_X1 _11883_ (
    .A(ex_reg_rs_msb_0[3]),
    .B(_04375_),
    .S(_04042_),
    .Z(_00070_)
  );
  AND2_X1 _11884_ (
    .A1(ibuf_io_inst_0_bits_raw[6]),
    .A2(_03582_),
    .ZN(_04376_)
  );
  MUX2_X1 _11885_ (
    .A(wb_reg_wdata[6]),
    .B(csr_io_rw_rdata[6]),
    .S(_04077_),
    .Z(_04377_)
  );
  MUX2_X1 _11886_ (
    .A(div_io_resp_bits_data[6]),
    .B(_04377_),
    .S(_03114_),
    .Z(_04378_)
  );
  MUX2_X1 _11887_ (
    .A(_04378_),
    .B(io_dmem_resp_bits_data[6]),
    .S(_03097_),
    .Z(_04379_)
  );
  MUX2_X1 _11888_ (
    .A(\rf[3] [6]),
    .B(\rf[1] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_04380_)
  );
  MUX2_X1 _11889_ (
    .A(\rf[7] [6]),
    .B(\rf[5] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_04381_)
  );
  MUX2_X1 _11890_ (
    .A(_04380_),
    .B(_04381_),
    .S(_03046_),
    .Z(_04382_)
  );
  AND2_X1 _11891_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_04382_),
    .ZN(_04383_)
  );
  MUX2_X1 _11892_ (
    .A(\rf[13] [6]),
    .B(\rf[9] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04384_)
  );
  OR2_X1 _11893_ (
    .A1(_03045_),
    .A2(_04384_),
    .ZN(_04385_)
  );
  MUX2_X1 _11894_ (
    .A(\rf[15] [6]),
    .B(\rf[11] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04386_)
  );
  OR2_X1 _11895_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04386_),
    .ZN(_04387_)
  );
  AND2_X1 _11896_ (
    .A1(_03047_),
    .A2(_04387_),
    .ZN(_04388_)
  );
  AND2_X1 _11897_ (
    .A1(_04385_),
    .A2(_04388_),
    .ZN(_04389_)
  );
  OR2_X1 _11898_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04389_),
    .ZN(_04390_)
  );
  OR2_X1 _11899_ (
    .A1(_04383_),
    .A2(_04390_),
    .ZN(_04391_)
  );
  MUX2_X1 _11900_ (
    .A(\rf[2] [6]),
    .B(\rf[0] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_04392_)
  );
  MUX2_X1 _11901_ (
    .A(\rf[6] [6]),
    .B(\rf[4] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_04393_)
  );
  MUX2_X1 _11902_ (
    .A(_04392_),
    .B(_04393_),
    .S(_03046_),
    .Z(_04394_)
  );
  AND2_X1 _11903_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_04394_),
    .ZN(_04395_)
  );
  MUX2_X1 _11904_ (
    .A(\rf[12] [6]),
    .B(\rf[8] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04396_)
  );
  OR2_X1 _11905_ (
    .A1(_03045_),
    .A2(_04396_),
    .ZN(_04397_)
  );
  MUX2_X1 _11906_ (
    .A(\rf[14] [6]),
    .B(\rf[10] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04398_)
  );
  OR2_X1 _11907_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04398_),
    .ZN(_04399_)
  );
  AND2_X1 _11908_ (
    .A1(_03047_),
    .A2(_04399_),
    .ZN(_04400_)
  );
  AND2_X1 _11909_ (
    .A1(_04397_),
    .A2(_04400_),
    .ZN(_04401_)
  );
  OR2_X1 _11910_ (
    .A1(_03044_),
    .A2(_04401_),
    .ZN(_04402_)
  );
  OR2_X1 _11911_ (
    .A1(_04395_),
    .A2(_04402_),
    .ZN(_04403_)
  );
  AND2_X1 _11912_ (
    .A1(_04391_),
    .A2(_04403_),
    .ZN(_04404_)
  );
  OR2_X1 _11913_ (
    .A1(_03063_),
    .A2(_04404_),
    .ZN(_04405_)
  );
  OR2_X1 _11914_ (
    .A1(\rf[25] [6]),
    .A2(_03046_),
    .ZN(_04406_)
  );
  OR2_X1 _11915_ (
    .A1(\rf[29] [6]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04407_)
  );
  AND2_X1 _11916_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04407_),
    .ZN(_04408_)
  );
  AND2_X1 _11917_ (
    .A1(_04406_),
    .A2(_04408_),
    .ZN(_04409_)
  );
  AND2_X1 _11918_ (
    .A1(\rf[27] [6]),
    .A2(_04273_),
    .ZN(_04410_)
  );
  OR2_X1 _11919_ (
    .A1(_04409_),
    .A2(_04410_),
    .ZN(_04411_)
  );
  MUX2_X1 _11920_ (
    .A(\rf[30] [6]),
    .B(\rf[26] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04412_)
  );
  OR2_X1 _11921_ (
    .A1(\rf[24] [6]),
    .A2(_03046_),
    .ZN(_04413_)
  );
  OR2_X1 _11922_ (
    .A1(\rf[28] [6]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04414_)
  );
  AND2_X1 _11923_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04414_),
    .ZN(_04415_)
  );
  AND2_X1 _11924_ (
    .A1(_04413_),
    .A2(_04415_),
    .ZN(_04416_)
  );
  AND2_X1 _11925_ (
    .A1(_03045_),
    .A2(_04412_),
    .ZN(_04417_)
  );
  OR2_X1 _11926_ (
    .A1(_03044_),
    .A2(_04417_),
    .ZN(_04418_)
  );
  OR2_X1 _11927_ (
    .A1(_04416_),
    .A2(_04418_),
    .ZN(_04419_)
  );
  OR2_X1 _11928_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04411_),
    .ZN(_04420_)
  );
  AND2_X1 _11929_ (
    .A1(_04419_),
    .A2(_04420_),
    .ZN(_04421_)
  );
  AND2_X1 _11930_ (
    .A1(_03047_),
    .A2(_04421_),
    .ZN(_04422_)
  );
  OR2_X1 _11931_ (
    .A1(\rf[20] [6]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04423_)
  );
  OR2_X1 _11932_ (
    .A1(\rf[16] [6]),
    .A2(_03046_),
    .ZN(_04424_)
  );
  AND2_X1 _11933_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04424_),
    .ZN(_04425_)
  );
  AND2_X1 _11934_ (
    .A1(_04423_),
    .A2(_04425_),
    .ZN(_04426_)
  );
  MUX2_X1 _11935_ (
    .A(\rf[22] [6]),
    .B(\rf[18] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04427_)
  );
  AND2_X1 _11936_ (
    .A1(_03045_),
    .A2(_04427_),
    .ZN(_04428_)
  );
  OR2_X1 _11937_ (
    .A1(_03044_),
    .A2(_04428_),
    .ZN(_04429_)
  );
  OR2_X1 _11938_ (
    .A1(_04426_),
    .A2(_04429_),
    .ZN(_04430_)
  );
  OR2_X1 _11939_ (
    .A1(\rf[17] [6]),
    .A2(_03046_),
    .ZN(_04431_)
  );
  OR2_X1 _11940_ (
    .A1(\rf[21] [6]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04432_)
  );
  AND2_X1 _11941_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04432_),
    .ZN(_04433_)
  );
  AND2_X1 _11942_ (
    .A1(_04431_),
    .A2(_04433_),
    .ZN(_04434_)
  );
  MUX2_X1 _11943_ (
    .A(\rf[23] [6]),
    .B(\rf[19] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04435_)
  );
  AND2_X1 _11944_ (
    .A1(_03045_),
    .A2(_04435_),
    .ZN(_04436_)
  );
  OR2_X1 _11945_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04436_),
    .ZN(_04437_)
  );
  OR2_X1 _11946_ (
    .A1(_04434_),
    .A2(_04437_),
    .ZN(_04438_)
  );
  AND2_X1 _11947_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_04438_),
    .ZN(_04439_)
  );
  AND2_X1 _11948_ (
    .A1(_04430_),
    .A2(_04439_),
    .ZN(_04440_)
  );
  OR2_X1 _11949_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_04440_),
    .ZN(_04441_)
  );
  OR2_X1 _11950_ (
    .A1(_04422_),
    .A2(_04441_),
    .ZN(_04442_)
  );
  AND2_X1 _11951_ (
    .A1(_04405_),
    .A2(_04442_),
    .ZN(_04443_)
  );
  MUX2_X1 _11952_ (
    .A(_04443_),
    .B(_04379_),
    .S(_04074_),
    .Z(_04444_)
  );
  AND2_X1 _11953_ (
    .A1(_04044_),
    .A2(_04444_),
    .ZN(_04445_)
  );
  OR2_X1 _11954_ (
    .A1(_04376_),
    .A2(_04445_),
    .ZN(_04446_)
  );
  MUX2_X1 _11955_ (
    .A(ex_reg_rs_msb_0[4]),
    .B(_04446_),
    .S(_04042_),
    .Z(_00071_)
  );
  AND2_X1 _11956_ (
    .A1(ibuf_io_inst_0_bits_raw[7]),
    .A2(_03582_),
    .ZN(_04447_)
  );
  MUX2_X1 _11957_ (
    .A(wb_reg_wdata[7]),
    .B(csr_io_rw_rdata[7]),
    .S(_04077_),
    .Z(_04448_)
  );
  MUX2_X1 _11958_ (
    .A(div_io_resp_bits_data[7]),
    .B(_04448_),
    .S(_03114_),
    .Z(_04449_)
  );
  MUX2_X1 _11959_ (
    .A(_04449_),
    .B(io_dmem_resp_bits_data[7]),
    .S(_03097_),
    .Z(_04450_)
  );
  MUX2_X1 _11960_ (
    .A(\rf[3] [7]),
    .B(\rf[1] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_04451_)
  );
  MUX2_X1 _11961_ (
    .A(\rf[7] [7]),
    .B(\rf[5] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_04452_)
  );
  MUX2_X1 _11962_ (
    .A(_04451_),
    .B(_04452_),
    .S(_03046_),
    .Z(_04453_)
  );
  AND2_X1 _11963_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_04453_),
    .ZN(_04454_)
  );
  MUX2_X1 _11964_ (
    .A(\rf[13] [7]),
    .B(\rf[9] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04455_)
  );
  OR2_X1 _11965_ (
    .A1(_03045_),
    .A2(_04455_),
    .ZN(_04456_)
  );
  MUX2_X1 _11966_ (
    .A(\rf[15] [7]),
    .B(\rf[11] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04457_)
  );
  OR2_X1 _11967_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04457_),
    .ZN(_04458_)
  );
  AND2_X1 _11968_ (
    .A1(_03047_),
    .A2(_04458_),
    .ZN(_04459_)
  );
  AND2_X1 _11969_ (
    .A1(_04456_),
    .A2(_04459_),
    .ZN(_04460_)
  );
  OR2_X1 _11970_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04460_),
    .ZN(_04461_)
  );
  OR2_X1 _11971_ (
    .A1(_04454_),
    .A2(_04461_),
    .ZN(_04462_)
  );
  MUX2_X1 _11972_ (
    .A(\rf[2] [7]),
    .B(\rf[0] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_04463_)
  );
  MUX2_X1 _11973_ (
    .A(\rf[6] [7]),
    .B(\rf[4] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_04464_)
  );
  MUX2_X1 _11974_ (
    .A(_04463_),
    .B(_04464_),
    .S(_03046_),
    .Z(_04465_)
  );
  AND2_X1 _11975_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_04465_),
    .ZN(_04466_)
  );
  MUX2_X1 _11976_ (
    .A(\rf[12] [7]),
    .B(\rf[8] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04467_)
  );
  OR2_X1 _11977_ (
    .A1(_03045_),
    .A2(_04467_),
    .ZN(_04468_)
  );
  MUX2_X1 _11978_ (
    .A(\rf[14] [7]),
    .B(\rf[10] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04469_)
  );
  OR2_X1 _11979_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04469_),
    .ZN(_04470_)
  );
  AND2_X1 _11980_ (
    .A1(_03047_),
    .A2(_04470_),
    .ZN(_04471_)
  );
  AND2_X1 _11981_ (
    .A1(_04468_),
    .A2(_04471_),
    .ZN(_04472_)
  );
  OR2_X1 _11982_ (
    .A1(_03044_),
    .A2(_04472_),
    .ZN(_04473_)
  );
  OR2_X1 _11983_ (
    .A1(_04466_),
    .A2(_04473_),
    .ZN(_04474_)
  );
  AND2_X1 _11984_ (
    .A1(_04462_),
    .A2(_04474_),
    .ZN(_04475_)
  );
  OR2_X1 _11985_ (
    .A1(_03063_),
    .A2(_04475_),
    .ZN(_04476_)
  );
  OR2_X1 _11986_ (
    .A1(\rf[25] [7]),
    .A2(_03046_),
    .ZN(_04477_)
  );
  OR2_X1 _11987_ (
    .A1(\rf[29] [7]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04478_)
  );
  AND2_X1 _11988_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04478_),
    .ZN(_04479_)
  );
  AND2_X1 _11989_ (
    .A1(_04477_),
    .A2(_04479_),
    .ZN(_04480_)
  );
  AND2_X1 _11990_ (
    .A1(\rf[27] [7]),
    .A2(_04273_),
    .ZN(_04481_)
  );
  OR2_X1 _11991_ (
    .A1(_04480_),
    .A2(_04481_),
    .ZN(_04482_)
  );
  MUX2_X1 _11992_ (
    .A(\rf[30] [7]),
    .B(\rf[26] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04483_)
  );
  OR2_X1 _11993_ (
    .A1(\rf[24] [7]),
    .A2(_03046_),
    .ZN(_04484_)
  );
  OR2_X1 _11994_ (
    .A1(\rf[28] [7]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04485_)
  );
  AND2_X1 _11995_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04485_),
    .ZN(_04486_)
  );
  AND2_X1 _11996_ (
    .A1(_04484_),
    .A2(_04486_),
    .ZN(_04487_)
  );
  AND2_X1 _11997_ (
    .A1(_03045_),
    .A2(_04483_),
    .ZN(_04488_)
  );
  OR2_X1 _11998_ (
    .A1(_03044_),
    .A2(_04488_),
    .ZN(_04489_)
  );
  OR2_X1 _11999_ (
    .A1(_04487_),
    .A2(_04489_),
    .ZN(_04490_)
  );
  OR2_X1 _12000_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04482_),
    .ZN(_04491_)
  );
  AND2_X1 _12001_ (
    .A1(_04490_),
    .A2(_04491_),
    .ZN(_04492_)
  );
  AND2_X1 _12002_ (
    .A1(_03047_),
    .A2(_04492_),
    .ZN(_04493_)
  );
  OR2_X1 _12003_ (
    .A1(\rf[20] [7]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04494_)
  );
  OR2_X1 _12004_ (
    .A1(\rf[16] [7]),
    .A2(_03046_),
    .ZN(_04495_)
  );
  AND2_X1 _12005_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04495_),
    .ZN(_04496_)
  );
  AND2_X1 _12006_ (
    .A1(_04494_),
    .A2(_04496_),
    .ZN(_04497_)
  );
  MUX2_X1 _12007_ (
    .A(\rf[22] [7]),
    .B(\rf[18] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04498_)
  );
  AND2_X1 _12008_ (
    .A1(_03045_),
    .A2(_04498_),
    .ZN(_04499_)
  );
  OR2_X1 _12009_ (
    .A1(_03044_),
    .A2(_04499_),
    .ZN(_04500_)
  );
  OR2_X1 _12010_ (
    .A1(_04497_),
    .A2(_04500_),
    .ZN(_04501_)
  );
  OR2_X1 _12011_ (
    .A1(\rf[17] [7]),
    .A2(_03046_),
    .ZN(_04502_)
  );
  OR2_X1 _12012_ (
    .A1(\rf[21] [7]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04503_)
  );
  AND2_X1 _12013_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04503_),
    .ZN(_04504_)
  );
  AND2_X1 _12014_ (
    .A1(_04502_),
    .A2(_04504_),
    .ZN(_04505_)
  );
  MUX2_X1 _12015_ (
    .A(\rf[23] [7]),
    .B(\rf[19] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04506_)
  );
  AND2_X1 _12016_ (
    .A1(_03045_),
    .A2(_04506_),
    .ZN(_04507_)
  );
  OR2_X1 _12017_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04507_),
    .ZN(_04508_)
  );
  OR2_X1 _12018_ (
    .A1(_04505_),
    .A2(_04508_),
    .ZN(_04509_)
  );
  AND2_X1 _12019_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_04509_),
    .ZN(_04510_)
  );
  AND2_X1 _12020_ (
    .A1(_04501_),
    .A2(_04510_),
    .ZN(_04511_)
  );
  OR2_X1 _12021_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_04511_),
    .ZN(_04512_)
  );
  OR2_X1 _12022_ (
    .A1(_04493_),
    .A2(_04512_),
    .ZN(_04513_)
  );
  AND2_X1 _12023_ (
    .A1(_04476_),
    .A2(_04513_),
    .ZN(_04514_)
  );
  MUX2_X1 _12024_ (
    .A(_04514_),
    .B(_04450_),
    .S(_04074_),
    .Z(_04515_)
  );
  AND2_X1 _12025_ (
    .A1(_04044_),
    .A2(_04515_),
    .ZN(_04516_)
  );
  OR2_X1 _12026_ (
    .A1(_04447_),
    .A2(_04516_),
    .ZN(_04517_)
  );
  MUX2_X1 _12027_ (
    .A(ex_reg_rs_msb_0[5]),
    .B(_04517_),
    .S(_04042_),
    .Z(_00072_)
  );
  AND2_X1 _12028_ (
    .A1(ibuf_io_inst_0_bits_raw[8]),
    .A2(_03582_),
    .ZN(_04518_)
  );
  MUX2_X1 _12029_ (
    .A(wb_reg_wdata[8]),
    .B(csr_io_rw_rdata[8]),
    .S(_04077_),
    .Z(_04519_)
  );
  MUX2_X1 _12030_ (
    .A(div_io_resp_bits_data[8]),
    .B(_04519_),
    .S(_03114_),
    .Z(_04520_)
  );
  MUX2_X1 _12031_ (
    .A(_04520_),
    .B(io_dmem_resp_bits_data[8]),
    .S(_03097_),
    .Z(_04521_)
  );
  OR2_X1 _12032_ (
    .A1(\rf[25] [8]),
    .A2(_03046_),
    .ZN(_04522_)
  );
  OR2_X1 _12033_ (
    .A1(\rf[29] [8]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04523_)
  );
  AND2_X1 _12034_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04523_),
    .ZN(_04524_)
  );
  AND2_X1 _12035_ (
    .A1(_04522_),
    .A2(_04524_),
    .ZN(_04525_)
  );
  AND2_X1 _12036_ (
    .A1(\rf[27] [8]),
    .A2(_04273_),
    .ZN(_04526_)
  );
  OR2_X1 _12037_ (
    .A1(_04525_),
    .A2(_04526_),
    .ZN(_04527_)
  );
  MUX2_X1 _12038_ (
    .A(\rf[30] [8]),
    .B(\rf[26] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04528_)
  );
  OR2_X1 _12039_ (
    .A1(\rf[24] [8]),
    .A2(_03046_),
    .ZN(_04529_)
  );
  OR2_X1 _12040_ (
    .A1(\rf[28] [8]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04530_)
  );
  AND2_X1 _12041_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04530_),
    .ZN(_04531_)
  );
  AND2_X1 _12042_ (
    .A1(_04529_),
    .A2(_04531_),
    .ZN(_04532_)
  );
  AND2_X1 _12043_ (
    .A1(_03045_),
    .A2(_04528_),
    .ZN(_04533_)
  );
  OR2_X1 _12044_ (
    .A1(_03044_),
    .A2(_04533_),
    .ZN(_04534_)
  );
  OR2_X1 _12045_ (
    .A1(_04532_),
    .A2(_04534_),
    .ZN(_04535_)
  );
  OR2_X1 _12046_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04527_),
    .ZN(_04536_)
  );
  AND2_X1 _12047_ (
    .A1(_04535_),
    .A2(_04536_),
    .ZN(_04537_)
  );
  AND2_X1 _12048_ (
    .A1(_03047_),
    .A2(_04537_),
    .ZN(_04538_)
  );
  OR2_X1 _12049_ (
    .A1(\rf[20] [8]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04539_)
  );
  OR2_X1 _12050_ (
    .A1(\rf[16] [8]),
    .A2(_03046_),
    .ZN(_04540_)
  );
  AND2_X1 _12051_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04540_),
    .ZN(_04541_)
  );
  AND2_X1 _12052_ (
    .A1(_04539_),
    .A2(_04541_),
    .ZN(_04542_)
  );
  MUX2_X1 _12053_ (
    .A(\rf[22] [8]),
    .B(\rf[18] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04543_)
  );
  AND2_X1 _12054_ (
    .A1(_03045_),
    .A2(_04543_),
    .ZN(_04544_)
  );
  OR2_X1 _12055_ (
    .A1(_03044_),
    .A2(_04544_),
    .ZN(_04545_)
  );
  OR2_X1 _12056_ (
    .A1(_04542_),
    .A2(_04545_),
    .ZN(_04546_)
  );
  OR2_X1 _12057_ (
    .A1(\rf[17] [8]),
    .A2(_03046_),
    .ZN(_04547_)
  );
  OR2_X1 _12058_ (
    .A1(\rf[21] [8]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04548_)
  );
  AND2_X1 _12059_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04548_),
    .ZN(_04549_)
  );
  AND2_X1 _12060_ (
    .A1(_04547_),
    .A2(_04549_),
    .ZN(_04550_)
  );
  MUX2_X1 _12061_ (
    .A(\rf[23] [8]),
    .B(\rf[19] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04551_)
  );
  AND2_X1 _12062_ (
    .A1(_03045_),
    .A2(_04551_),
    .ZN(_04552_)
  );
  OR2_X1 _12063_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04552_),
    .ZN(_04553_)
  );
  OR2_X1 _12064_ (
    .A1(_04550_),
    .A2(_04553_),
    .ZN(_04554_)
  );
  AND2_X1 _12065_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_04554_),
    .ZN(_04555_)
  );
  AND2_X1 _12066_ (
    .A1(_04546_),
    .A2(_04555_),
    .ZN(_04556_)
  );
  OR2_X1 _12067_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_04556_),
    .ZN(_04557_)
  );
  OR2_X1 _12068_ (
    .A1(_04538_),
    .A2(_04557_),
    .ZN(_04558_)
  );
  MUX2_X1 _12069_ (
    .A(\rf[1] [8]),
    .B(\rf[0] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_04559_)
  );
  MUX2_X1 _12070_ (
    .A(\rf[5] [8]),
    .B(\rf[4] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_04560_)
  );
  MUX2_X1 _12071_ (
    .A(_04559_),
    .B(_04560_),
    .S(_03046_),
    .Z(_04561_)
  );
  OR2_X1 _12072_ (
    .A1(_03047_),
    .A2(_04561_),
    .ZN(_04562_)
  );
  MUX2_X1 _12073_ (
    .A(\rf[12] [8]),
    .B(\rf[8] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04563_)
  );
  OR2_X1 _12074_ (
    .A1(_04124_),
    .A2(_04563_),
    .ZN(_04564_)
  );
  MUX2_X1 _12075_ (
    .A(\rf[13] [8]),
    .B(\rf[9] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04565_)
  );
  OR2_X1 _12076_ (
    .A1(_03448_),
    .A2(_04565_),
    .ZN(_04566_)
  );
  AND2_X1 _12077_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04566_),
    .ZN(_04567_)
  );
  AND2_X1 _12078_ (
    .A1(_04564_),
    .A2(_04567_),
    .ZN(_04568_)
  );
  AND2_X1 _12079_ (
    .A1(_04562_),
    .A2(_04568_),
    .ZN(_04569_)
  );
  MUX2_X1 _12080_ (
    .A(\rf[3] [8]),
    .B(\rf[2] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_04570_)
  );
  MUX2_X1 _12081_ (
    .A(\rf[7] [8]),
    .B(\rf[6] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_04571_)
  );
  MUX2_X1 _12082_ (
    .A(_04570_),
    .B(_04571_),
    .S(_03046_),
    .Z(_04572_)
  );
  OR2_X1 _12083_ (
    .A1(_03047_),
    .A2(_04572_),
    .ZN(_04573_)
  );
  MUX2_X1 _12084_ (
    .A(\rf[15] [8]),
    .B(\rf[11] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04574_)
  );
  OR2_X1 _12085_ (
    .A1(_03448_),
    .A2(_04574_),
    .ZN(_04575_)
  );
  MUX2_X1 _12086_ (
    .A(\rf[14] [8]),
    .B(\rf[10] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04576_)
  );
  OR2_X1 _12087_ (
    .A1(_04124_),
    .A2(_04576_),
    .ZN(_04577_)
  );
  AND2_X1 _12088_ (
    .A1(_04575_),
    .A2(_04577_),
    .ZN(_04578_)
  );
  AND2_X1 _12089_ (
    .A1(_04573_),
    .A2(_04578_),
    .ZN(_04579_)
  );
  AND2_X1 _12090_ (
    .A1(_03045_),
    .A2(_04579_),
    .ZN(_04580_)
  );
  OR2_X1 _12091_ (
    .A1(_03063_),
    .A2(_04569_),
    .ZN(_04581_)
  );
  OR2_X1 _12092_ (
    .A1(_04580_),
    .A2(_04581_),
    .ZN(_04582_)
  );
  AND2_X1 _12093_ (
    .A1(_04558_),
    .A2(_04582_),
    .ZN(_04583_)
  );
  MUX2_X1 _12094_ (
    .A(_04583_),
    .B(_04521_),
    .S(_04074_),
    .Z(_04584_)
  );
  AND2_X1 _12095_ (
    .A1(_04044_),
    .A2(_04584_),
    .ZN(_04585_)
  );
  OR2_X1 _12096_ (
    .A1(_04518_),
    .A2(_04585_),
    .ZN(_04586_)
  );
  MUX2_X1 _12097_ (
    .A(ex_reg_rs_msb_0[6]),
    .B(_04586_),
    .S(_04042_),
    .Z(_00073_)
  );
  AND2_X1 _12098_ (
    .A1(ibuf_io_inst_0_bits_raw[9]),
    .A2(_03582_),
    .ZN(_04587_)
  );
  MUX2_X1 _12099_ (
    .A(wb_reg_wdata[9]),
    .B(csr_io_rw_rdata[9]),
    .S(_04077_),
    .Z(_04588_)
  );
  MUX2_X1 _12100_ (
    .A(div_io_resp_bits_data[9]),
    .B(_04588_),
    .S(_03114_),
    .Z(_04589_)
  );
  MUX2_X1 _12101_ (
    .A(_04589_),
    .B(io_dmem_resp_bits_data[9]),
    .S(_03097_),
    .Z(_04590_)
  );
  OR2_X1 _12102_ (
    .A1(\rf[25] [9]),
    .A2(_03046_),
    .ZN(_04591_)
  );
  OR2_X1 _12103_ (
    .A1(\rf[29] [9]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04592_)
  );
  AND2_X1 _12104_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04592_),
    .ZN(_04593_)
  );
  AND2_X1 _12105_ (
    .A1(_04591_),
    .A2(_04593_),
    .ZN(_04594_)
  );
  AND2_X1 _12106_ (
    .A1(\rf[27] [9]),
    .A2(_04273_),
    .ZN(_04595_)
  );
  OR2_X1 _12107_ (
    .A1(_04594_),
    .A2(_04595_),
    .ZN(_04596_)
  );
  MUX2_X1 _12108_ (
    .A(\rf[30] [9]),
    .B(\rf[26] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04597_)
  );
  OR2_X1 _12109_ (
    .A1(\rf[24] [9]),
    .A2(_03046_),
    .ZN(_04598_)
  );
  OR2_X1 _12110_ (
    .A1(\rf[28] [9]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04599_)
  );
  AND2_X1 _12111_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04599_),
    .ZN(_04600_)
  );
  AND2_X1 _12112_ (
    .A1(_04598_),
    .A2(_04600_),
    .ZN(_04601_)
  );
  AND2_X1 _12113_ (
    .A1(_03045_),
    .A2(_04597_),
    .ZN(_04602_)
  );
  OR2_X1 _12114_ (
    .A1(_03044_),
    .A2(_04602_),
    .ZN(_04603_)
  );
  OR2_X1 _12115_ (
    .A1(_04601_),
    .A2(_04603_),
    .ZN(_04604_)
  );
  OR2_X1 _12116_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04596_),
    .ZN(_04605_)
  );
  AND2_X1 _12117_ (
    .A1(_04604_),
    .A2(_04605_),
    .ZN(_04606_)
  );
  AND2_X1 _12118_ (
    .A1(_03047_),
    .A2(_04606_),
    .ZN(_04607_)
  );
  OR2_X1 _12119_ (
    .A1(\rf[20] [9]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04608_)
  );
  OR2_X1 _12120_ (
    .A1(\rf[16] [9]),
    .A2(_03046_),
    .ZN(_04609_)
  );
  AND2_X1 _12121_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04609_),
    .ZN(_04610_)
  );
  AND2_X1 _12122_ (
    .A1(_04608_),
    .A2(_04610_),
    .ZN(_04611_)
  );
  MUX2_X1 _12123_ (
    .A(\rf[22] [9]),
    .B(\rf[18] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04612_)
  );
  AND2_X1 _12124_ (
    .A1(_03045_),
    .A2(_04612_),
    .ZN(_04613_)
  );
  OR2_X1 _12125_ (
    .A1(_03044_),
    .A2(_04613_),
    .ZN(_04614_)
  );
  OR2_X1 _12126_ (
    .A1(_04611_),
    .A2(_04614_),
    .ZN(_04615_)
  );
  OR2_X1 _12127_ (
    .A1(\rf[17] [9]),
    .A2(_03046_),
    .ZN(_04616_)
  );
  OR2_X1 _12128_ (
    .A1(\rf[21] [9]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04617_)
  );
  AND2_X1 _12129_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04617_),
    .ZN(_04618_)
  );
  AND2_X1 _12130_ (
    .A1(_04616_),
    .A2(_04618_),
    .ZN(_04619_)
  );
  MUX2_X1 _12131_ (
    .A(\rf[23] [9]),
    .B(\rf[19] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04620_)
  );
  AND2_X1 _12132_ (
    .A1(_03045_),
    .A2(_04620_),
    .ZN(_04621_)
  );
  OR2_X1 _12133_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04621_),
    .ZN(_04622_)
  );
  OR2_X1 _12134_ (
    .A1(_04619_),
    .A2(_04622_),
    .ZN(_04623_)
  );
  AND2_X1 _12135_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_04623_),
    .ZN(_04624_)
  );
  AND2_X1 _12136_ (
    .A1(_04615_),
    .A2(_04624_),
    .ZN(_04625_)
  );
  OR2_X1 _12137_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_04625_),
    .ZN(_04626_)
  );
  OR2_X1 _12138_ (
    .A1(_04607_),
    .A2(_04626_),
    .ZN(_04627_)
  );
  MUX2_X1 _12139_ (
    .A(\rf[1] [9]),
    .B(\rf[0] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_04628_)
  );
  MUX2_X1 _12140_ (
    .A(\rf[5] [9]),
    .B(\rf[4] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_04629_)
  );
  MUX2_X1 _12141_ (
    .A(_04628_),
    .B(_04629_),
    .S(_03046_),
    .Z(_04630_)
  );
  OR2_X1 _12142_ (
    .A1(_03047_),
    .A2(_04630_),
    .ZN(_04631_)
  );
  MUX2_X1 _12143_ (
    .A(\rf[12] [9]),
    .B(\rf[8] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04632_)
  );
  OR2_X1 _12144_ (
    .A1(_04124_),
    .A2(_04632_),
    .ZN(_04633_)
  );
  MUX2_X1 _12145_ (
    .A(\rf[13] [9]),
    .B(\rf[9] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04634_)
  );
  OR2_X1 _12146_ (
    .A1(_03448_),
    .A2(_04634_),
    .ZN(_04635_)
  );
  AND2_X1 _12147_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04635_),
    .ZN(_04636_)
  );
  AND2_X1 _12148_ (
    .A1(_04633_),
    .A2(_04636_),
    .ZN(_04637_)
  );
  AND2_X1 _12149_ (
    .A1(_04631_),
    .A2(_04637_),
    .ZN(_04638_)
  );
  MUX2_X1 _12150_ (
    .A(\rf[3] [9]),
    .B(\rf[2] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_04639_)
  );
  MUX2_X1 _12151_ (
    .A(\rf[7] [9]),
    .B(\rf[6] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_04640_)
  );
  MUX2_X1 _12152_ (
    .A(_04639_),
    .B(_04640_),
    .S(_03046_),
    .Z(_04641_)
  );
  OR2_X1 _12153_ (
    .A1(_03047_),
    .A2(_04641_),
    .ZN(_04642_)
  );
  MUX2_X1 _12154_ (
    .A(\rf[14] [9]),
    .B(\rf[10] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04643_)
  );
  OR2_X1 _12155_ (
    .A1(_04124_),
    .A2(_04643_),
    .ZN(_04644_)
  );
  MUX2_X1 _12156_ (
    .A(\rf[15] [9]),
    .B(\rf[11] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04645_)
  );
  OR2_X1 _12157_ (
    .A1(_03448_),
    .A2(_04645_),
    .ZN(_04646_)
  );
  AND2_X1 _12158_ (
    .A1(_03045_),
    .A2(_04646_),
    .ZN(_04647_)
  );
  AND2_X1 _12159_ (
    .A1(_04644_),
    .A2(_04647_),
    .ZN(_04648_)
  );
  AND2_X1 _12160_ (
    .A1(_04642_),
    .A2(_04648_),
    .ZN(_04649_)
  );
  OR2_X1 _12161_ (
    .A1(_03063_),
    .A2(_04638_),
    .ZN(_04650_)
  );
  OR2_X1 _12162_ (
    .A1(_04649_),
    .A2(_04650_),
    .ZN(_04651_)
  );
  AND2_X1 _12163_ (
    .A1(_04627_),
    .A2(_04651_),
    .ZN(_04652_)
  );
  MUX2_X1 _12164_ (
    .A(_04652_),
    .B(_04590_),
    .S(_04074_),
    .Z(_04653_)
  );
  AND2_X1 _12165_ (
    .A1(_04044_),
    .A2(_04653_),
    .ZN(_04654_)
  );
  OR2_X1 _12166_ (
    .A1(_04587_),
    .A2(_04654_),
    .ZN(_04655_)
  );
  MUX2_X1 _12167_ (
    .A(ex_reg_rs_msb_0[7]),
    .B(_04655_),
    .S(_04042_),
    .Z(_00074_)
  );
  AND2_X1 _12168_ (
    .A1(ibuf_io_inst_0_bits_raw[10]),
    .A2(_03582_),
    .ZN(_04656_)
  );
  MUX2_X1 _12169_ (
    .A(wb_reg_wdata[10]),
    .B(csr_io_rw_rdata[10]),
    .S(_04077_),
    .Z(_04657_)
  );
  MUX2_X1 _12170_ (
    .A(div_io_resp_bits_data[10]),
    .B(_04657_),
    .S(_03114_),
    .Z(_04658_)
  );
  MUX2_X1 _12171_ (
    .A(_04658_),
    .B(io_dmem_resp_bits_data[10]),
    .S(_03097_),
    .Z(_04659_)
  );
  MUX2_X1 _12172_ (
    .A(\rf[15] [10]),
    .B(\rf[11] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04660_)
  );
  OR2_X1 _12173_ (
    .A1(\rf[14] [10]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04661_)
  );
  OR2_X1 _12174_ (
    .A1(\rf[10] [10]),
    .A2(_03046_),
    .ZN(_04662_)
  );
  MUX2_X1 _12175_ (
    .A(\rf[13] [10]),
    .B(\rf[9] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04663_)
  );
  OR2_X1 _12176_ (
    .A1(\rf[8] [10]),
    .A2(_03046_),
    .ZN(_04664_)
  );
  OR2_X1 _12177_ (
    .A1(\rf[12] [10]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04665_)
  );
  AND2_X1 _12178_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04661_),
    .ZN(_04666_)
  );
  AND2_X1 _12179_ (
    .A1(_04662_),
    .A2(_04666_),
    .ZN(_04667_)
  );
  AND2_X1 _12180_ (
    .A1(_03044_),
    .A2(_04660_),
    .ZN(_04668_)
  );
  OR2_X1 _12181_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04668_),
    .ZN(_04669_)
  );
  OR2_X1 _12182_ (
    .A1(_04667_),
    .A2(_04669_),
    .ZN(_04670_)
  );
  AND2_X1 _12183_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04665_),
    .ZN(_04671_)
  );
  AND2_X1 _12184_ (
    .A1(_04664_),
    .A2(_04671_),
    .ZN(_04672_)
  );
  AND2_X1 _12185_ (
    .A1(_03044_),
    .A2(_04663_),
    .ZN(_04673_)
  );
  OR2_X1 _12186_ (
    .A1(_03045_),
    .A2(_04673_),
    .ZN(_04674_)
  );
  OR2_X1 _12187_ (
    .A1(_04672_),
    .A2(_04674_),
    .ZN(_04675_)
  );
  AND2_X1 _12188_ (
    .A1(_03047_),
    .A2(_04675_),
    .ZN(_04676_)
  );
  AND2_X1 _12189_ (
    .A1(_04670_),
    .A2(_04676_),
    .ZN(_04677_)
  );
  OR2_X1 _12190_ (
    .A1(\rf[0] [10]),
    .A2(_03046_),
    .ZN(_04678_)
  );
  OR2_X1 _12191_ (
    .A1(\rf[4] [10]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04679_)
  );
  AND2_X1 _12192_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04679_),
    .ZN(_04680_)
  );
  AND2_X1 _12193_ (
    .A1(_04678_),
    .A2(_04680_),
    .ZN(_04681_)
  );
  MUX2_X1 _12194_ (
    .A(\rf[5] [10]),
    .B(\rf[1] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04682_)
  );
  AND2_X1 _12195_ (
    .A1(_03044_),
    .A2(_04682_),
    .ZN(_04683_)
  );
  OR2_X1 _12196_ (
    .A1(_03045_),
    .A2(_04683_),
    .ZN(_04684_)
  );
  OR2_X1 _12197_ (
    .A1(_04681_),
    .A2(_04684_),
    .ZN(_04685_)
  );
  MUX2_X1 _12198_ (
    .A(\rf[7] [10]),
    .B(\rf[3] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04686_)
  );
  AND2_X1 _12199_ (
    .A1(_03044_),
    .A2(_04686_),
    .ZN(_04687_)
  );
  OR2_X1 _12200_ (
    .A1(\rf[2] [10]),
    .A2(_03046_),
    .ZN(_04688_)
  );
  OR2_X1 _12201_ (
    .A1(\rf[6] [10]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04689_)
  );
  AND2_X1 _12202_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04689_),
    .ZN(_04690_)
  );
  AND2_X1 _12203_ (
    .A1(_04688_),
    .A2(_04690_),
    .ZN(_04691_)
  );
  OR2_X1 _12204_ (
    .A1(_04687_),
    .A2(_04691_),
    .ZN(_04692_)
  );
  OR2_X1 _12205_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04692_),
    .ZN(_04693_)
  );
  AND2_X1 _12206_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_04685_),
    .ZN(_04694_)
  );
  AND2_X1 _12207_ (
    .A1(_04693_),
    .A2(_04694_),
    .ZN(_04695_)
  );
  OR2_X1 _12208_ (
    .A1(_03063_),
    .A2(_04677_),
    .ZN(_04696_)
  );
  OR2_X1 _12209_ (
    .A1(_04695_),
    .A2(_04696_),
    .ZN(_04697_)
  );
  OR2_X1 _12210_ (
    .A1(\rf[26] [10]),
    .A2(_03046_),
    .ZN(_04698_)
  );
  OR2_X1 _12211_ (
    .A1(\rf[30] [10]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04699_)
  );
  AND2_X1 _12212_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04699_),
    .ZN(_04700_)
  );
  AND2_X1 _12213_ (
    .A1(_04698_),
    .A2(_04700_),
    .ZN(_04701_)
  );
  AND2_X1 _12214_ (
    .A1(\rf[27] [10]),
    .A2(_03760_),
    .ZN(_04702_)
  );
  OR2_X1 _12215_ (
    .A1(_04701_),
    .A2(_04702_),
    .ZN(_04703_)
  );
  MUX2_X1 _12216_ (
    .A(\rf[29] [10]),
    .B(\rf[25] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04704_)
  );
  AND2_X1 _12217_ (
    .A1(_03044_),
    .A2(_04704_),
    .ZN(_04705_)
  );
  OR2_X1 _12218_ (
    .A1(\rf[28] [10]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04706_)
  );
  OR2_X1 _12219_ (
    .A1(\rf[24] [10]),
    .A2(_03046_),
    .ZN(_04707_)
  );
  AND2_X1 _12220_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04707_),
    .ZN(_04708_)
  );
  AND2_X1 _12221_ (
    .A1(_04706_),
    .A2(_04708_),
    .ZN(_04709_)
  );
  OR2_X1 _12222_ (
    .A1(_03045_),
    .A2(_04709_),
    .ZN(_04710_)
  );
  OR2_X1 _12223_ (
    .A1(_04705_),
    .A2(_04710_),
    .ZN(_04711_)
  );
  OR2_X1 _12224_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04703_),
    .ZN(_04712_)
  );
  AND2_X1 _12225_ (
    .A1(_03047_),
    .A2(_04712_),
    .ZN(_04713_)
  );
  AND2_X1 _12226_ (
    .A1(_04711_),
    .A2(_04713_),
    .ZN(_04714_)
  );
  MUX2_X1 _12227_ (
    .A(\rf[21] [10]),
    .B(\rf[17] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04715_)
  );
  AND2_X1 _12228_ (
    .A1(_03044_),
    .A2(_04715_),
    .ZN(_04716_)
  );
  OR2_X1 _12229_ (
    .A1(\rf[20] [10]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04717_)
  );
  OR2_X1 _12230_ (
    .A1(\rf[16] [10]),
    .A2(_03046_),
    .ZN(_04718_)
  );
  AND2_X1 _12231_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04717_),
    .ZN(_04719_)
  );
  AND2_X1 _12232_ (
    .A1(_04718_),
    .A2(_04719_),
    .ZN(_04720_)
  );
  OR2_X1 _12233_ (
    .A1(_03045_),
    .A2(_04716_),
    .ZN(_04721_)
  );
  OR2_X1 _12234_ (
    .A1(_04720_),
    .A2(_04721_),
    .ZN(_04722_)
  );
  OR2_X1 _12235_ (
    .A1(\rf[18] [10]),
    .A2(_03046_),
    .ZN(_04723_)
  );
  OR2_X1 _12236_ (
    .A1(\rf[22] [10]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04724_)
  );
  AND2_X1 _12237_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04724_),
    .ZN(_04725_)
  );
  AND2_X1 _12238_ (
    .A1(_04723_),
    .A2(_04725_),
    .ZN(_04726_)
  );
  MUX2_X1 _12239_ (
    .A(\rf[23] [10]),
    .B(\rf[19] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04727_)
  );
  AND2_X1 _12240_ (
    .A1(_03044_),
    .A2(_04727_),
    .ZN(_04728_)
  );
  OR2_X1 _12241_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04728_),
    .ZN(_04729_)
  );
  OR2_X1 _12242_ (
    .A1(_04726_),
    .A2(_04729_),
    .ZN(_04730_)
  );
  AND2_X1 _12243_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_04730_),
    .ZN(_04731_)
  );
  AND2_X1 _12244_ (
    .A1(_04722_),
    .A2(_04731_),
    .ZN(_04732_)
  );
  OR2_X1 _12245_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_04732_),
    .ZN(_04733_)
  );
  OR2_X1 _12246_ (
    .A1(_04714_),
    .A2(_04733_),
    .ZN(_04734_)
  );
  AND2_X1 _12247_ (
    .A1(_04697_),
    .A2(_04734_),
    .ZN(_04735_)
  );
  MUX2_X1 _12248_ (
    .A(_04735_),
    .B(_04659_),
    .S(_04074_),
    .Z(_04736_)
  );
  AND2_X1 _12249_ (
    .A1(_04044_),
    .A2(_04736_),
    .ZN(_04737_)
  );
  OR2_X1 _12250_ (
    .A1(_04656_),
    .A2(_04737_),
    .ZN(_04738_)
  );
  MUX2_X1 _12251_ (
    .A(ex_reg_rs_msb_0[8]),
    .B(_04738_),
    .S(_04042_),
    .Z(_00075_)
  );
  AND2_X1 _12252_ (
    .A1(ibuf_io_inst_0_bits_raw[11]),
    .A2(_03582_),
    .ZN(_04739_)
  );
  MUX2_X1 _12253_ (
    .A(wb_reg_wdata[11]),
    .B(csr_io_rw_rdata[11]),
    .S(_04077_),
    .Z(_04740_)
  );
  MUX2_X1 _12254_ (
    .A(div_io_resp_bits_data[11]),
    .B(_04740_),
    .S(_03114_),
    .Z(_04741_)
  );
  MUX2_X1 _12255_ (
    .A(_04741_),
    .B(io_dmem_resp_bits_data[11]),
    .S(_03097_),
    .Z(_04742_)
  );
  OR2_X1 _12256_ (
    .A1(\rf[25] [11]),
    .A2(_03046_),
    .ZN(_04743_)
  );
  OR2_X1 _12257_ (
    .A1(\rf[29] [11]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04744_)
  );
  AND2_X1 _12258_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04744_),
    .ZN(_04745_)
  );
  AND2_X1 _12259_ (
    .A1(_04743_),
    .A2(_04745_),
    .ZN(_04746_)
  );
  AND2_X1 _12260_ (
    .A1(\rf[27] [11]),
    .A2(_04273_),
    .ZN(_04747_)
  );
  OR2_X1 _12261_ (
    .A1(_04746_),
    .A2(_04747_),
    .ZN(_04748_)
  );
  MUX2_X1 _12262_ (
    .A(\rf[30] [11]),
    .B(\rf[26] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04749_)
  );
  OR2_X1 _12263_ (
    .A1(\rf[24] [11]),
    .A2(_03046_),
    .ZN(_04750_)
  );
  OR2_X1 _12264_ (
    .A1(\rf[28] [11]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04751_)
  );
  AND2_X1 _12265_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04751_),
    .ZN(_04752_)
  );
  AND2_X1 _12266_ (
    .A1(_04750_),
    .A2(_04752_),
    .ZN(_04753_)
  );
  AND2_X1 _12267_ (
    .A1(_03045_),
    .A2(_04749_),
    .ZN(_04754_)
  );
  OR2_X1 _12268_ (
    .A1(_03044_),
    .A2(_04754_),
    .ZN(_04755_)
  );
  OR2_X1 _12269_ (
    .A1(_04753_),
    .A2(_04755_),
    .ZN(_04756_)
  );
  OR2_X1 _12270_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04748_),
    .ZN(_04757_)
  );
  AND2_X1 _12271_ (
    .A1(_04756_),
    .A2(_04757_),
    .ZN(_04758_)
  );
  AND2_X1 _12272_ (
    .A1(_03047_),
    .A2(_04758_),
    .ZN(_04759_)
  );
  OR2_X1 _12273_ (
    .A1(\rf[20] [11]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04760_)
  );
  OR2_X1 _12274_ (
    .A1(\rf[16] [11]),
    .A2(_03046_),
    .ZN(_04761_)
  );
  AND2_X1 _12275_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04761_),
    .ZN(_04762_)
  );
  AND2_X1 _12276_ (
    .A1(_04760_),
    .A2(_04762_),
    .ZN(_04763_)
  );
  MUX2_X1 _12277_ (
    .A(\rf[22] [11]),
    .B(\rf[18] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04764_)
  );
  AND2_X1 _12278_ (
    .A1(_03045_),
    .A2(_04764_),
    .ZN(_04765_)
  );
  OR2_X1 _12279_ (
    .A1(_03044_),
    .A2(_04765_),
    .ZN(_04766_)
  );
  OR2_X1 _12280_ (
    .A1(_04763_),
    .A2(_04766_),
    .ZN(_04767_)
  );
  OR2_X1 _12281_ (
    .A1(\rf[17] [11]),
    .A2(_03046_),
    .ZN(_04768_)
  );
  OR2_X1 _12282_ (
    .A1(\rf[21] [11]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04769_)
  );
  AND2_X1 _12283_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04769_),
    .ZN(_04770_)
  );
  AND2_X1 _12284_ (
    .A1(_04768_),
    .A2(_04770_),
    .ZN(_04771_)
  );
  MUX2_X1 _12285_ (
    .A(\rf[23] [11]),
    .B(\rf[19] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04772_)
  );
  AND2_X1 _12286_ (
    .A1(_03045_),
    .A2(_04772_),
    .ZN(_04773_)
  );
  OR2_X1 _12287_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04773_),
    .ZN(_04774_)
  );
  OR2_X1 _12288_ (
    .A1(_04771_),
    .A2(_04774_),
    .ZN(_04775_)
  );
  AND2_X1 _12289_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_04775_),
    .ZN(_04776_)
  );
  AND2_X1 _12290_ (
    .A1(_04767_),
    .A2(_04776_),
    .ZN(_04777_)
  );
  OR2_X1 _12291_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_04777_),
    .ZN(_04778_)
  );
  OR2_X1 _12292_ (
    .A1(_04759_),
    .A2(_04778_),
    .ZN(_04779_)
  );
  MUX2_X1 _12293_ (
    .A(\rf[1] [11]),
    .B(\rf[0] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_04780_)
  );
  MUX2_X1 _12294_ (
    .A(\rf[5] [11]),
    .B(\rf[4] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_04781_)
  );
  MUX2_X1 _12295_ (
    .A(_04780_),
    .B(_04781_),
    .S(_03046_),
    .Z(_04782_)
  );
  OR2_X1 _12296_ (
    .A1(_03047_),
    .A2(_04782_),
    .ZN(_04783_)
  );
  MUX2_X1 _12297_ (
    .A(\rf[12] [11]),
    .B(\rf[8] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04784_)
  );
  OR2_X1 _12298_ (
    .A1(_04124_),
    .A2(_04784_),
    .ZN(_04785_)
  );
  MUX2_X1 _12299_ (
    .A(\rf[13] [11]),
    .B(\rf[9] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04786_)
  );
  OR2_X1 _12300_ (
    .A1(_03448_),
    .A2(_04786_),
    .ZN(_04787_)
  );
  AND2_X1 _12301_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04787_),
    .ZN(_04788_)
  );
  AND2_X1 _12302_ (
    .A1(_04785_),
    .A2(_04788_),
    .ZN(_04789_)
  );
  AND2_X1 _12303_ (
    .A1(_04783_),
    .A2(_04789_),
    .ZN(_04790_)
  );
  MUX2_X1 _12304_ (
    .A(\rf[3] [11]),
    .B(\rf[2] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_04791_)
  );
  MUX2_X1 _12305_ (
    .A(\rf[7] [11]),
    .B(\rf[6] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_04792_)
  );
  MUX2_X1 _12306_ (
    .A(_04791_),
    .B(_04792_),
    .S(_03046_),
    .Z(_04793_)
  );
  OR2_X1 _12307_ (
    .A1(_03047_),
    .A2(_04793_),
    .ZN(_04794_)
  );
  MUX2_X1 _12308_ (
    .A(\rf[14] [11]),
    .B(\rf[10] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04795_)
  );
  OR2_X1 _12309_ (
    .A1(_04124_),
    .A2(_04795_),
    .ZN(_04796_)
  );
  MUX2_X1 _12310_ (
    .A(\rf[15] [11]),
    .B(\rf[11] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04797_)
  );
  OR2_X1 _12311_ (
    .A1(_03448_),
    .A2(_04797_),
    .ZN(_04798_)
  );
  AND2_X1 _12312_ (
    .A1(_03045_),
    .A2(_04798_),
    .ZN(_04799_)
  );
  AND2_X1 _12313_ (
    .A1(_04796_),
    .A2(_04799_),
    .ZN(_04800_)
  );
  AND2_X1 _12314_ (
    .A1(_04794_),
    .A2(_04800_),
    .ZN(_04801_)
  );
  OR2_X1 _12315_ (
    .A1(_03063_),
    .A2(_04790_),
    .ZN(_04802_)
  );
  OR2_X1 _12316_ (
    .A1(_04801_),
    .A2(_04802_),
    .ZN(_04803_)
  );
  AND2_X1 _12317_ (
    .A1(_04779_),
    .A2(_04803_),
    .ZN(_04804_)
  );
  MUX2_X1 _12318_ (
    .A(_04804_),
    .B(_04742_),
    .S(_04074_),
    .Z(_04805_)
  );
  AND2_X1 _12319_ (
    .A1(_04044_),
    .A2(_04805_),
    .ZN(_04806_)
  );
  OR2_X1 _12320_ (
    .A1(_04739_),
    .A2(_04806_),
    .ZN(_04807_)
  );
  MUX2_X1 _12321_ (
    .A(ex_reg_rs_msb_0[9]),
    .B(_04807_),
    .S(_04042_),
    .Z(_00076_)
  );
  AND2_X1 _12322_ (
    .A1(ibuf_io_inst_0_bits_raw[12]),
    .A2(_03582_),
    .ZN(_04808_)
  );
  MUX2_X1 _12323_ (
    .A(wb_reg_wdata[12]),
    .B(csr_io_rw_rdata[12]),
    .S(_04077_),
    .Z(_04809_)
  );
  MUX2_X1 _12324_ (
    .A(div_io_resp_bits_data[12]),
    .B(_04809_),
    .S(_03114_),
    .Z(_04810_)
  );
  MUX2_X1 _12325_ (
    .A(_04810_),
    .B(io_dmem_resp_bits_data[12]),
    .S(_03097_),
    .Z(_04811_)
  );
  MUX2_X1 _12326_ (
    .A(\rf[3] [12]),
    .B(\rf[1] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_04812_)
  );
  MUX2_X1 _12327_ (
    .A(\rf[7] [12]),
    .B(\rf[5] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_04813_)
  );
  MUX2_X1 _12328_ (
    .A(_04812_),
    .B(_04813_),
    .S(_03046_),
    .Z(_04814_)
  );
  AND2_X1 _12329_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_04814_),
    .ZN(_04815_)
  );
  MUX2_X1 _12330_ (
    .A(\rf[13] [12]),
    .B(\rf[9] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04816_)
  );
  OR2_X1 _12331_ (
    .A1(_03045_),
    .A2(_04816_),
    .ZN(_04817_)
  );
  MUX2_X1 _12332_ (
    .A(\rf[15] [12]),
    .B(\rf[11] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04818_)
  );
  OR2_X1 _12333_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04818_),
    .ZN(_04819_)
  );
  AND2_X1 _12334_ (
    .A1(_03047_),
    .A2(_04819_),
    .ZN(_04820_)
  );
  AND2_X1 _12335_ (
    .A1(_04817_),
    .A2(_04820_),
    .ZN(_04821_)
  );
  OR2_X1 _12336_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04821_),
    .ZN(_04822_)
  );
  OR2_X1 _12337_ (
    .A1(_04815_),
    .A2(_04822_),
    .ZN(_04823_)
  );
  MUX2_X1 _12338_ (
    .A(\rf[2] [12]),
    .B(\rf[0] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_04824_)
  );
  MUX2_X1 _12339_ (
    .A(\rf[6] [12]),
    .B(\rf[4] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_04825_)
  );
  MUX2_X1 _12340_ (
    .A(_04824_),
    .B(_04825_),
    .S(_03046_),
    .Z(_04826_)
  );
  AND2_X1 _12341_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_04826_),
    .ZN(_04827_)
  );
  MUX2_X1 _12342_ (
    .A(\rf[12] [12]),
    .B(\rf[8] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04828_)
  );
  OR2_X1 _12343_ (
    .A1(_03045_),
    .A2(_04828_),
    .ZN(_04829_)
  );
  MUX2_X1 _12344_ (
    .A(\rf[14] [12]),
    .B(\rf[10] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04830_)
  );
  OR2_X1 _12345_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04830_),
    .ZN(_04831_)
  );
  AND2_X1 _12346_ (
    .A1(_03047_),
    .A2(_04831_),
    .ZN(_04832_)
  );
  AND2_X1 _12347_ (
    .A1(_04829_),
    .A2(_04832_),
    .ZN(_04833_)
  );
  OR2_X1 _12348_ (
    .A1(_03044_),
    .A2(_04833_),
    .ZN(_04834_)
  );
  OR2_X1 _12349_ (
    .A1(_04827_),
    .A2(_04834_),
    .ZN(_04835_)
  );
  AND2_X1 _12350_ (
    .A1(_04823_),
    .A2(_04835_),
    .ZN(_04836_)
  );
  OR2_X1 _12351_ (
    .A1(_03063_),
    .A2(_04836_),
    .ZN(_04837_)
  );
  OR2_X1 _12352_ (
    .A1(\rf[25] [12]),
    .A2(_03046_),
    .ZN(_04838_)
  );
  OR2_X1 _12353_ (
    .A1(\rf[29] [12]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04839_)
  );
  AND2_X1 _12354_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04839_),
    .ZN(_04840_)
  );
  AND2_X1 _12355_ (
    .A1(_04838_),
    .A2(_04840_),
    .ZN(_04841_)
  );
  AND2_X1 _12356_ (
    .A1(\rf[27] [12]),
    .A2(_04273_),
    .ZN(_04842_)
  );
  OR2_X1 _12357_ (
    .A1(_04841_),
    .A2(_04842_),
    .ZN(_04843_)
  );
  MUX2_X1 _12358_ (
    .A(\rf[30] [12]),
    .B(\rf[26] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04844_)
  );
  OR2_X1 _12359_ (
    .A1(\rf[24] [12]),
    .A2(_03046_),
    .ZN(_04845_)
  );
  OR2_X1 _12360_ (
    .A1(\rf[28] [12]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04846_)
  );
  AND2_X1 _12361_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04846_),
    .ZN(_04847_)
  );
  AND2_X1 _12362_ (
    .A1(_04845_),
    .A2(_04847_),
    .ZN(_04848_)
  );
  AND2_X1 _12363_ (
    .A1(_03045_),
    .A2(_04844_),
    .ZN(_04849_)
  );
  OR2_X1 _12364_ (
    .A1(_03044_),
    .A2(_04849_),
    .ZN(_04850_)
  );
  OR2_X1 _12365_ (
    .A1(_04848_),
    .A2(_04850_),
    .ZN(_04851_)
  );
  OR2_X1 _12366_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04843_),
    .ZN(_04852_)
  );
  AND2_X1 _12367_ (
    .A1(_04851_),
    .A2(_04852_),
    .ZN(_04853_)
  );
  AND2_X1 _12368_ (
    .A1(_03047_),
    .A2(_04853_),
    .ZN(_04854_)
  );
  OR2_X1 _12369_ (
    .A1(\rf[20] [12]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04855_)
  );
  OR2_X1 _12370_ (
    .A1(\rf[16] [12]),
    .A2(_03046_),
    .ZN(_04856_)
  );
  AND2_X1 _12371_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04856_),
    .ZN(_04857_)
  );
  AND2_X1 _12372_ (
    .A1(_04855_),
    .A2(_04857_),
    .ZN(_04858_)
  );
  MUX2_X1 _12373_ (
    .A(\rf[22] [12]),
    .B(\rf[18] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04859_)
  );
  AND2_X1 _12374_ (
    .A1(_03045_),
    .A2(_04859_),
    .ZN(_04860_)
  );
  OR2_X1 _12375_ (
    .A1(_03044_),
    .A2(_04860_),
    .ZN(_04861_)
  );
  OR2_X1 _12376_ (
    .A1(_04858_),
    .A2(_04861_),
    .ZN(_04862_)
  );
  OR2_X1 _12377_ (
    .A1(\rf[17] [12]),
    .A2(_03046_),
    .ZN(_04863_)
  );
  OR2_X1 _12378_ (
    .A1(\rf[21] [12]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04864_)
  );
  AND2_X1 _12379_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04864_),
    .ZN(_04865_)
  );
  AND2_X1 _12380_ (
    .A1(_04863_),
    .A2(_04865_),
    .ZN(_04866_)
  );
  MUX2_X1 _12381_ (
    .A(\rf[23] [12]),
    .B(\rf[19] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04867_)
  );
  AND2_X1 _12382_ (
    .A1(_03045_),
    .A2(_04867_),
    .ZN(_04868_)
  );
  OR2_X1 _12383_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04868_),
    .ZN(_04869_)
  );
  OR2_X1 _12384_ (
    .A1(_04866_),
    .A2(_04869_),
    .ZN(_04870_)
  );
  AND2_X1 _12385_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_04870_),
    .ZN(_04871_)
  );
  AND2_X1 _12386_ (
    .A1(_04862_),
    .A2(_04871_),
    .ZN(_04872_)
  );
  OR2_X1 _12387_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_04872_),
    .ZN(_04873_)
  );
  OR2_X1 _12388_ (
    .A1(_04854_),
    .A2(_04873_),
    .ZN(_04874_)
  );
  AND2_X1 _12389_ (
    .A1(_04837_),
    .A2(_04874_),
    .ZN(_04875_)
  );
  MUX2_X1 _12390_ (
    .A(_04875_),
    .B(_04811_),
    .S(_04074_),
    .Z(_04876_)
  );
  AND2_X1 _12391_ (
    .A1(_04044_),
    .A2(_04876_),
    .ZN(_04877_)
  );
  OR2_X1 _12392_ (
    .A1(_04808_),
    .A2(_04877_),
    .ZN(_04878_)
  );
  MUX2_X1 _12393_ (
    .A(ex_reg_rs_msb_0[10]),
    .B(_04878_),
    .S(_04042_),
    .Z(_00077_)
  );
  AND2_X1 _12394_ (
    .A1(ibuf_io_inst_0_bits_raw[13]),
    .A2(_03582_),
    .ZN(_04879_)
  );
  MUX2_X1 _12395_ (
    .A(wb_reg_wdata[13]),
    .B(csr_io_rw_rdata[13]),
    .S(_04077_),
    .Z(_04880_)
  );
  MUX2_X1 _12396_ (
    .A(div_io_resp_bits_data[13]),
    .B(_04880_),
    .S(_03114_),
    .Z(_04881_)
  );
  MUX2_X1 _12397_ (
    .A(_04881_),
    .B(io_dmem_resp_bits_data[13]),
    .S(_03097_),
    .Z(_04882_)
  );
  MUX2_X1 _12398_ (
    .A(\rf[3] [13]),
    .B(\rf[1] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_04883_)
  );
  MUX2_X1 _12399_ (
    .A(\rf[7] [13]),
    .B(\rf[5] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_04884_)
  );
  MUX2_X1 _12400_ (
    .A(_04883_),
    .B(_04884_),
    .S(_03046_),
    .Z(_04885_)
  );
  AND2_X1 _12401_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_04885_),
    .ZN(_04886_)
  );
  MUX2_X1 _12402_ (
    .A(\rf[13] [13]),
    .B(\rf[9] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04887_)
  );
  OR2_X1 _12403_ (
    .A1(_03045_),
    .A2(_04887_),
    .ZN(_04888_)
  );
  MUX2_X1 _12404_ (
    .A(\rf[15] [13]),
    .B(\rf[11] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04889_)
  );
  OR2_X1 _12405_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04889_),
    .ZN(_04890_)
  );
  AND2_X1 _12406_ (
    .A1(_03047_),
    .A2(_04890_),
    .ZN(_04891_)
  );
  AND2_X1 _12407_ (
    .A1(_04888_),
    .A2(_04891_),
    .ZN(_04892_)
  );
  OR2_X1 _12408_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04892_),
    .ZN(_04893_)
  );
  OR2_X1 _12409_ (
    .A1(_04886_),
    .A2(_04893_),
    .ZN(_04894_)
  );
  MUX2_X1 _12410_ (
    .A(\rf[2] [13]),
    .B(\rf[0] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_04895_)
  );
  MUX2_X1 _12411_ (
    .A(\rf[6] [13]),
    .B(\rf[4] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs1[1]),
    .Z(_04896_)
  );
  MUX2_X1 _12412_ (
    .A(_04895_),
    .B(_04896_),
    .S(_03046_),
    .Z(_04897_)
  );
  AND2_X1 _12413_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_04897_),
    .ZN(_04898_)
  );
  MUX2_X1 _12414_ (
    .A(\rf[12] [13]),
    .B(\rf[8] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04899_)
  );
  OR2_X1 _12415_ (
    .A1(_03045_),
    .A2(_04899_),
    .ZN(_04900_)
  );
  MUX2_X1 _12416_ (
    .A(\rf[14] [13]),
    .B(\rf[10] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04901_)
  );
  OR2_X1 _12417_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04901_),
    .ZN(_04902_)
  );
  AND2_X1 _12418_ (
    .A1(_03047_),
    .A2(_04902_),
    .ZN(_04903_)
  );
  AND2_X1 _12419_ (
    .A1(_04900_),
    .A2(_04903_),
    .ZN(_04904_)
  );
  OR2_X1 _12420_ (
    .A1(_03044_),
    .A2(_04904_),
    .ZN(_04905_)
  );
  OR2_X1 _12421_ (
    .A1(_04898_),
    .A2(_04905_),
    .ZN(_04906_)
  );
  AND2_X1 _12422_ (
    .A1(_04894_),
    .A2(_04906_),
    .ZN(_04907_)
  );
  OR2_X1 _12423_ (
    .A1(_03063_),
    .A2(_04907_),
    .ZN(_04908_)
  );
  OR2_X1 _12424_ (
    .A1(\rf[25] [13]),
    .A2(_03046_),
    .ZN(_04909_)
  );
  OR2_X1 _12425_ (
    .A1(\rf[29] [13]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04910_)
  );
  AND2_X1 _12426_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04910_),
    .ZN(_04911_)
  );
  AND2_X1 _12427_ (
    .A1(_04909_),
    .A2(_04911_),
    .ZN(_04912_)
  );
  AND2_X1 _12428_ (
    .A1(\rf[27] [13]),
    .A2(_04273_),
    .ZN(_04913_)
  );
  OR2_X1 _12429_ (
    .A1(_04912_),
    .A2(_04913_),
    .ZN(_04914_)
  );
  MUX2_X1 _12430_ (
    .A(\rf[30] [13]),
    .B(\rf[26] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04915_)
  );
  OR2_X1 _12431_ (
    .A1(\rf[24] [13]),
    .A2(_03046_),
    .ZN(_04916_)
  );
  OR2_X1 _12432_ (
    .A1(\rf[28] [13]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04917_)
  );
  AND2_X1 _12433_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04917_),
    .ZN(_04918_)
  );
  AND2_X1 _12434_ (
    .A1(_04916_),
    .A2(_04918_),
    .ZN(_04919_)
  );
  AND2_X1 _12435_ (
    .A1(_03045_),
    .A2(_04915_),
    .ZN(_04920_)
  );
  OR2_X1 _12436_ (
    .A1(_03044_),
    .A2(_04920_),
    .ZN(_04921_)
  );
  OR2_X1 _12437_ (
    .A1(_04919_),
    .A2(_04921_),
    .ZN(_04922_)
  );
  OR2_X1 _12438_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04914_),
    .ZN(_04923_)
  );
  AND2_X1 _12439_ (
    .A1(_04922_),
    .A2(_04923_),
    .ZN(_04924_)
  );
  AND2_X1 _12440_ (
    .A1(_03047_),
    .A2(_04924_),
    .ZN(_04925_)
  );
  OR2_X1 _12441_ (
    .A1(\rf[20] [13]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04926_)
  );
  OR2_X1 _12442_ (
    .A1(\rf[16] [13]),
    .A2(_03046_),
    .ZN(_04927_)
  );
  AND2_X1 _12443_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04927_),
    .ZN(_04928_)
  );
  AND2_X1 _12444_ (
    .A1(_04926_),
    .A2(_04928_),
    .ZN(_04929_)
  );
  MUX2_X1 _12445_ (
    .A(\rf[22] [13]),
    .B(\rf[18] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04930_)
  );
  AND2_X1 _12446_ (
    .A1(_03045_),
    .A2(_04930_),
    .ZN(_04931_)
  );
  OR2_X1 _12447_ (
    .A1(_03044_),
    .A2(_04931_),
    .ZN(_04932_)
  );
  OR2_X1 _12448_ (
    .A1(_04929_),
    .A2(_04932_),
    .ZN(_04933_)
  );
  OR2_X1 _12449_ (
    .A1(\rf[17] [13]),
    .A2(_03046_),
    .ZN(_04934_)
  );
  OR2_X1 _12450_ (
    .A1(\rf[21] [13]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04935_)
  );
  AND2_X1 _12451_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04935_),
    .ZN(_04936_)
  );
  AND2_X1 _12452_ (
    .A1(_04934_),
    .A2(_04936_),
    .ZN(_04937_)
  );
  MUX2_X1 _12453_ (
    .A(\rf[23] [13]),
    .B(\rf[19] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04938_)
  );
  AND2_X1 _12454_ (
    .A1(_03045_),
    .A2(_04938_),
    .ZN(_04939_)
  );
  OR2_X1 _12455_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04939_),
    .ZN(_04940_)
  );
  OR2_X1 _12456_ (
    .A1(_04937_),
    .A2(_04940_),
    .ZN(_04941_)
  );
  AND2_X1 _12457_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_04941_),
    .ZN(_04942_)
  );
  AND2_X1 _12458_ (
    .A1(_04933_),
    .A2(_04942_),
    .ZN(_04943_)
  );
  OR2_X1 _12459_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_04943_),
    .ZN(_04944_)
  );
  OR2_X1 _12460_ (
    .A1(_04925_),
    .A2(_04944_),
    .ZN(_04945_)
  );
  AND2_X1 _12461_ (
    .A1(_04908_),
    .A2(_04945_),
    .ZN(_04946_)
  );
  MUX2_X1 _12462_ (
    .A(_04946_),
    .B(_04882_),
    .S(_04074_),
    .Z(_04947_)
  );
  AND2_X1 _12463_ (
    .A1(_04044_),
    .A2(_04947_),
    .ZN(_04948_)
  );
  OR2_X1 _12464_ (
    .A1(_04879_),
    .A2(_04948_),
    .ZN(_04949_)
  );
  MUX2_X1 _12465_ (
    .A(ex_reg_rs_msb_0[11]),
    .B(_04949_),
    .S(_04042_),
    .Z(_00078_)
  );
  AND2_X1 _12466_ (
    .A1(ibuf_io_inst_0_bits_raw[14]),
    .A2(_03582_),
    .ZN(_04950_)
  );
  MUX2_X1 _12467_ (
    .A(wb_reg_wdata[14]),
    .B(csr_io_rw_rdata[14]),
    .S(_04077_),
    .Z(_04951_)
  );
  MUX2_X1 _12468_ (
    .A(div_io_resp_bits_data[14]),
    .B(_04951_),
    .S(_03114_),
    .Z(_04952_)
  );
  MUX2_X1 _12469_ (
    .A(_04952_),
    .B(io_dmem_resp_bits_data[14]),
    .S(_03097_),
    .Z(_04953_)
  );
  MUX2_X1 _12470_ (
    .A(\rf[5] [14]),
    .B(\rf[1] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04954_)
  );
  MUX2_X1 _12471_ (
    .A(\rf[7] [14]),
    .B(\rf[3] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04955_)
  );
  MUX2_X1 _12472_ (
    .A(_04954_),
    .B(_04955_),
    .S(_03045_),
    .Z(_04956_)
  );
  AND2_X1 _12473_ (
    .A1(_03044_),
    .A2(_04956_),
    .ZN(_04957_)
  );
  MUX2_X1 _12474_ (
    .A(\rf[4] [14]),
    .B(\rf[0] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04958_)
  );
  MUX2_X1 _12475_ (
    .A(\rf[6] [14]),
    .B(\rf[2] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04959_)
  );
  MUX2_X1 _12476_ (
    .A(_04958_),
    .B(_04959_),
    .S(_03045_),
    .Z(_04960_)
  );
  AND2_X1 _12477_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04960_),
    .ZN(_04961_)
  );
  OR2_X1 _12478_ (
    .A1(_03063_),
    .A2(_04961_),
    .ZN(_04962_)
  );
  OR2_X1 _12479_ (
    .A1(_04957_),
    .A2(_04962_),
    .ZN(_04963_)
  );
  OR2_X1 _12480_ (
    .A1(\rf[20] [14]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04964_)
  );
  OR2_X1 _12481_ (
    .A1(\rf[16] [14]),
    .A2(_03046_),
    .ZN(_04965_)
  );
  AND2_X1 _12482_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04965_),
    .ZN(_04966_)
  );
  AND2_X1 _12483_ (
    .A1(_04964_),
    .A2(_04966_),
    .ZN(_04967_)
  );
  MUX2_X1 _12484_ (
    .A(\rf[22] [14]),
    .B(\rf[18] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04968_)
  );
  AND2_X1 _12485_ (
    .A1(_03045_),
    .A2(_04968_),
    .ZN(_04969_)
  );
  OR2_X1 _12486_ (
    .A1(_03044_),
    .A2(_04969_),
    .ZN(_04970_)
  );
  OR2_X1 _12487_ (
    .A1(_04967_),
    .A2(_04970_),
    .ZN(_04971_)
  );
  OR2_X1 _12488_ (
    .A1(\rf[17] [14]),
    .A2(_03046_),
    .ZN(_04972_)
  );
  OR2_X1 _12489_ (
    .A1(\rf[21] [14]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_04973_)
  );
  AND2_X1 _12490_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_04973_),
    .ZN(_04974_)
  );
  AND2_X1 _12491_ (
    .A1(_04972_),
    .A2(_04974_),
    .ZN(_04975_)
  );
  MUX2_X1 _12492_ (
    .A(\rf[23] [14]),
    .B(\rf[19] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_04976_)
  );
  AND2_X1 _12493_ (
    .A1(_03045_),
    .A2(_04976_),
    .ZN(_04977_)
  );
  OR2_X1 _12494_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04977_),
    .ZN(_04978_)
  );
  OR2_X1 _12495_ (
    .A1(_04975_),
    .A2(_04978_),
    .ZN(_04979_)
  );
  AND2_X1 _12496_ (
    .A1(_04971_),
    .A2(_04979_),
    .ZN(_04980_)
  );
  OR2_X1 _12497_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_04980_),
    .ZN(_04981_)
  );
  AND2_X1 _12498_ (
    .A1(_04963_),
    .A2(_04981_),
    .ZN(_04982_)
  );
  AND2_X1 _12499_ (
    .A1(\rf[10] [14]),
    .A2(_03045_),
    .ZN(_04983_)
  );
  AND2_X1 _12500_ (
    .A1(\rf[8] [14]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_04984_)
  );
  OR2_X1 _12501_ (
    .A1(_03046_),
    .A2(_04984_),
    .ZN(_04985_)
  );
  OR2_X1 _12502_ (
    .A1(_04983_),
    .A2(_04985_),
    .ZN(_04986_)
  );
  AND2_X1 _12503_ (
    .A1(\rf[14] [14]),
    .A2(_03045_),
    .ZN(_04987_)
  );
  AND2_X1 _12504_ (
    .A1(\rf[12] [14]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_04988_)
  );
  OR2_X1 _12505_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_04988_),
    .ZN(_04989_)
  );
  OR2_X1 _12506_ (
    .A1(_04987_),
    .A2(_04989_),
    .ZN(_04990_)
  );
  AND2_X1 _12507_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_04990_),
    .ZN(_04991_)
  );
  AND2_X1 _12508_ (
    .A1(_04986_),
    .A2(_04991_),
    .ZN(_04992_)
  );
  AND2_X1 _12509_ (
    .A1(\rf[11] [14]),
    .A2(_03045_),
    .ZN(_04993_)
  );
  AND2_X1 _12510_ (
    .A1(\rf[9] [14]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_04994_)
  );
  OR2_X1 _12511_ (
    .A1(_03046_),
    .A2(_04994_),
    .ZN(_04995_)
  );
  OR2_X1 _12512_ (
    .A1(_04993_),
    .A2(_04995_),
    .ZN(_04996_)
  );
  AND2_X1 _12513_ (
    .A1(\rf[15] [14]),
    .A2(_03045_),
    .ZN(_04997_)
  );
  AND2_X1 _12514_ (
    .A1(\rf[13] [14]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_04998_)
  );
  OR2_X1 _12515_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_04998_),
    .ZN(_04999_)
  );
  OR2_X1 _12516_ (
    .A1(_04997_),
    .A2(_04999_),
    .ZN(_05000_)
  );
  AND2_X1 _12517_ (
    .A1(_03044_),
    .A2(_05000_),
    .ZN(_05001_)
  );
  AND2_X1 _12518_ (
    .A1(_04996_),
    .A2(_05001_),
    .ZN(_05002_)
  );
  OR2_X1 _12519_ (
    .A1(_03063_),
    .A2(_05002_),
    .ZN(_05003_)
  );
  OR2_X1 _12520_ (
    .A1(_04992_),
    .A2(_05003_),
    .ZN(_05004_)
  );
  OR2_X1 _12521_ (
    .A1(\rf[28] [14]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05005_)
  );
  OR2_X1 _12522_ (
    .A1(\rf[24] [14]),
    .A2(_03046_),
    .ZN(_05006_)
  );
  AND2_X1 _12523_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05005_),
    .ZN(_05007_)
  );
  AND2_X1 _12524_ (
    .A1(_05006_),
    .A2(_05007_),
    .ZN(_05008_)
  );
  MUX2_X1 _12525_ (
    .A(\rf[30] [14]),
    .B(\rf[26] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05009_)
  );
  AND2_X1 _12526_ (
    .A1(_03045_),
    .A2(_05009_),
    .ZN(_05010_)
  );
  OR2_X1 _12527_ (
    .A1(_03044_),
    .A2(_05010_),
    .ZN(_05011_)
  );
  OR2_X1 _12528_ (
    .A1(_05008_),
    .A2(_05011_),
    .ZN(_05012_)
  );
  MUX2_X1 _12529_ (
    .A(\rf[29] [14]),
    .B(\rf[25] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05013_)
  );
  AND2_X1 _12530_ (
    .A1(\rf[27] [14]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05014_)
  );
  MUX2_X1 _12531_ (
    .A(_05013_),
    .B(_05014_),
    .S(_03045_),
    .Z(_05015_)
  );
  OR2_X1 _12532_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05015_),
    .ZN(_05016_)
  );
  AND2_X1 _12533_ (
    .A1(_05012_),
    .A2(_05016_),
    .ZN(_05017_)
  );
  OR2_X1 _12534_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_05017_),
    .ZN(_05018_)
  );
  AND2_X1 _12535_ (
    .A1(_05004_),
    .A2(_05018_),
    .ZN(_05019_)
  );
  MUX2_X1 _12536_ (
    .A(_04982_),
    .B(_05019_),
    .S(_03047_),
    .Z(_05020_)
  );
  MUX2_X1 _12537_ (
    .A(_05020_),
    .B(_04953_),
    .S(_04074_),
    .Z(_05021_)
  );
  AND2_X1 _12538_ (
    .A1(_04044_),
    .A2(_05021_),
    .ZN(_05022_)
  );
  OR2_X1 _12539_ (
    .A1(_04950_),
    .A2(_05022_),
    .ZN(_05023_)
  );
  MUX2_X1 _12540_ (
    .A(ex_reg_rs_msb_0[12]),
    .B(_05023_),
    .S(_04042_),
    .Z(_00079_)
  );
  AND2_X1 _12541_ (
    .A1(ibuf_io_inst_0_bits_raw[15]),
    .A2(_03582_),
    .ZN(_05024_)
  );
  MUX2_X1 _12542_ (
    .A(wb_reg_wdata[15]),
    .B(csr_io_rw_rdata[15]),
    .S(_04077_),
    .Z(_05025_)
  );
  MUX2_X1 _12543_ (
    .A(div_io_resp_bits_data[15]),
    .B(_05025_),
    .S(_03114_),
    .Z(_05026_)
  );
  MUX2_X1 _12544_ (
    .A(_05026_),
    .B(io_dmem_resp_bits_data[15]),
    .S(_03097_),
    .Z(_05027_)
  );
  OR2_X1 _12545_ (
    .A1(\rf[26] [15]),
    .A2(_03046_),
    .ZN(_05028_)
  );
  OR2_X1 _12546_ (
    .A1(\rf[30] [15]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05029_)
  );
  AND2_X1 _12547_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05029_),
    .ZN(_05030_)
  );
  AND2_X1 _12548_ (
    .A1(_05028_),
    .A2(_05030_),
    .ZN(_05031_)
  );
  AND2_X1 _12549_ (
    .A1(\rf[27] [15]),
    .A2(_03760_),
    .ZN(_05032_)
  );
  OR2_X1 _12550_ (
    .A1(_05031_),
    .A2(_05032_),
    .ZN(_05033_)
  );
  MUX2_X1 _12551_ (
    .A(\rf[23] [15]),
    .B(\rf[19] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05034_)
  );
  AND2_X1 _12552_ (
    .A1(_03044_),
    .A2(_05034_),
    .ZN(_05035_)
  );
  OR2_X1 _12553_ (
    .A1(\rf[22] [15]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05036_)
  );
  OR2_X1 _12554_ (
    .A1(\rf[18] [15]),
    .A2(_03046_),
    .ZN(_05037_)
  );
  AND2_X1 _12555_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05037_),
    .ZN(_05038_)
  );
  AND2_X1 _12556_ (
    .A1(_05036_),
    .A2(_05038_),
    .ZN(_05039_)
  );
  OR2_X1 _12557_ (
    .A1(_03047_),
    .A2(_05039_),
    .ZN(_05040_)
  );
  OR2_X1 _12558_ (
    .A1(_05035_),
    .A2(_05040_),
    .ZN(_05041_)
  );
  OR2_X1 _12559_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_05033_),
    .ZN(_05042_)
  );
  AND2_X1 _12560_ (
    .A1(_03045_),
    .A2(_05042_),
    .ZN(_05043_)
  );
  AND2_X1 _12561_ (
    .A1(_05041_),
    .A2(_05043_),
    .ZN(_05044_)
  );
  MUX2_X1 _12562_ (
    .A(\rf[21] [15]),
    .B(\rf[17] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05045_)
  );
  AND2_X1 _12563_ (
    .A1(_03044_),
    .A2(_05045_),
    .ZN(_05046_)
  );
  OR2_X1 _12564_ (
    .A1(\rf[20] [15]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05047_)
  );
  OR2_X1 _12565_ (
    .A1(\rf[16] [15]),
    .A2(_03046_),
    .ZN(_05048_)
  );
  AND2_X1 _12566_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05047_),
    .ZN(_05049_)
  );
  AND2_X1 _12567_ (
    .A1(_05048_),
    .A2(_05049_),
    .ZN(_05050_)
  );
  OR2_X1 _12568_ (
    .A1(_03047_),
    .A2(_05046_),
    .ZN(_05051_)
  );
  OR2_X1 _12569_ (
    .A1(_05050_),
    .A2(_05051_),
    .ZN(_05052_)
  );
  OR2_X1 _12570_ (
    .A1(\rf[24] [15]),
    .A2(_03046_),
    .ZN(_05053_)
  );
  OR2_X1 _12571_ (
    .A1(\rf[28] [15]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05054_)
  );
  AND2_X1 _12572_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05054_),
    .ZN(_05055_)
  );
  AND2_X1 _12573_ (
    .A1(_05053_),
    .A2(_05055_),
    .ZN(_05056_)
  );
  MUX2_X1 _12574_ (
    .A(\rf[29] [15]),
    .B(\rf[25] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05057_)
  );
  AND2_X1 _12575_ (
    .A1(_03044_),
    .A2(_05057_),
    .ZN(_05058_)
  );
  OR2_X1 _12576_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_05058_),
    .ZN(_05059_)
  );
  OR2_X1 _12577_ (
    .A1(_05056_),
    .A2(_05059_),
    .ZN(_05060_)
  );
  AND2_X1 _12578_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05060_),
    .ZN(_05061_)
  );
  AND2_X1 _12579_ (
    .A1(_05052_),
    .A2(_05061_),
    .ZN(_05062_)
  );
  OR2_X1 _12580_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_05062_),
    .ZN(_05063_)
  );
  OR2_X1 _12581_ (
    .A1(_05044_),
    .A2(_05063_),
    .ZN(_05064_)
  );
  MUX2_X1 _12582_ (
    .A(\rf[1] [15]),
    .B(\rf[0] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_05065_)
  );
  MUX2_X1 _12583_ (
    .A(\rf[5] [15]),
    .B(\rf[4] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_05066_)
  );
  MUX2_X1 _12584_ (
    .A(_05065_),
    .B(_05066_),
    .S(_03046_),
    .Z(_05067_)
  );
  OR2_X1 _12585_ (
    .A1(_03047_),
    .A2(_05067_),
    .ZN(_05068_)
  );
  MUX2_X1 _12586_ (
    .A(\rf[12] [15]),
    .B(\rf[8] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05069_)
  );
  OR2_X1 _12587_ (
    .A1(_04124_),
    .A2(_05069_),
    .ZN(_05070_)
  );
  MUX2_X1 _12588_ (
    .A(\rf[13] [15]),
    .B(\rf[9] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05071_)
  );
  OR2_X1 _12589_ (
    .A1(_03448_),
    .A2(_05071_),
    .ZN(_05072_)
  );
  AND2_X1 _12590_ (
    .A1(_05070_),
    .A2(_05072_),
    .ZN(_05073_)
  );
  AND2_X1 _12591_ (
    .A1(_05068_),
    .A2(_05073_),
    .ZN(_05074_)
  );
  MUX2_X1 _12592_ (
    .A(\rf[3] [15]),
    .B(\rf[2] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_05075_)
  );
  MUX2_X1 _12593_ (
    .A(\rf[7] [15]),
    .B(\rf[6] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_05076_)
  );
  MUX2_X1 _12594_ (
    .A(_05075_),
    .B(_05076_),
    .S(_03046_),
    .Z(_05077_)
  );
  OR2_X1 _12595_ (
    .A1(_03047_),
    .A2(_05077_),
    .ZN(_05078_)
  );
  MUX2_X1 _12596_ (
    .A(\rf[14] [15]),
    .B(\rf[10] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05079_)
  );
  OR2_X1 _12597_ (
    .A1(_04124_),
    .A2(_05079_),
    .ZN(_05080_)
  );
  MUX2_X1 _12598_ (
    .A(\rf[15] [15]),
    .B(\rf[11] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05081_)
  );
  OR2_X1 _12599_ (
    .A1(_03448_),
    .A2(_05081_),
    .ZN(_05082_)
  );
  AND2_X1 _12600_ (
    .A1(_05080_),
    .A2(_05082_),
    .ZN(_05083_)
  );
  AND2_X1 _12601_ (
    .A1(_05078_),
    .A2(_05083_),
    .ZN(_05084_)
  );
  MUX2_X1 _12602_ (
    .A(_05074_),
    .B(_05084_),
    .S(_03045_),
    .Z(_05085_)
  );
  OR2_X1 _12603_ (
    .A1(_03063_),
    .A2(_05085_),
    .ZN(_05086_)
  );
  AND2_X1 _12604_ (
    .A1(_05064_),
    .A2(_05086_),
    .ZN(_05087_)
  );
  MUX2_X1 _12605_ (
    .A(_05087_),
    .B(_05027_),
    .S(_04074_),
    .Z(_05088_)
  );
  AND2_X1 _12606_ (
    .A1(_04044_),
    .A2(_05088_),
    .ZN(_05089_)
  );
  OR2_X1 _12607_ (
    .A1(_05024_),
    .A2(_05089_),
    .ZN(_05090_)
  );
  MUX2_X1 _12608_ (
    .A(ex_reg_rs_msb_0[13]),
    .B(_05090_),
    .S(_04042_),
    .Z(_00080_)
  );
  AND2_X1 _12609_ (
    .A1(_03065_),
    .A2(ibuf_io_inst_0_bits_raw[16]),
    .ZN(_05091_)
  );
  AND2_X1 _12610_ (
    .A1(_03582_),
    .A2(_05091_),
    .ZN(_05092_)
  );
  MUX2_X1 _12611_ (
    .A(wb_reg_wdata[16]),
    .B(csr_io_rw_rdata[16]),
    .S(_04077_),
    .Z(_05093_)
  );
  MUX2_X1 _12612_ (
    .A(div_io_resp_bits_data[16]),
    .B(_05093_),
    .S(_03114_),
    .Z(_05094_)
  );
  MUX2_X1 _12613_ (
    .A(_05094_),
    .B(io_dmem_resp_bits_data[16]),
    .S(_03097_),
    .Z(_05095_)
  );
  MUX2_X1 _12614_ (
    .A(\rf[5] [16]),
    .B(\rf[1] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05096_)
  );
  MUX2_X1 _12615_ (
    .A(\rf[7] [16]),
    .B(\rf[3] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05097_)
  );
  MUX2_X1 _12616_ (
    .A(_05096_),
    .B(_05097_),
    .S(_03045_),
    .Z(_05098_)
  );
  AND2_X1 _12617_ (
    .A1(_03044_),
    .A2(_05098_),
    .ZN(_05099_)
  );
  MUX2_X1 _12618_ (
    .A(\rf[4] [16]),
    .B(\rf[0] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05100_)
  );
  MUX2_X1 _12619_ (
    .A(\rf[6] [16]),
    .B(\rf[2] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05101_)
  );
  MUX2_X1 _12620_ (
    .A(_05100_),
    .B(_05101_),
    .S(_03045_),
    .Z(_05102_)
  );
  AND2_X1 _12621_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05102_),
    .ZN(_05103_)
  );
  OR2_X1 _12622_ (
    .A1(_03063_),
    .A2(_05103_),
    .ZN(_05104_)
  );
  OR2_X1 _12623_ (
    .A1(_05099_),
    .A2(_05104_),
    .ZN(_05105_)
  );
  OR2_X1 _12624_ (
    .A1(\rf[20] [16]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05106_)
  );
  OR2_X1 _12625_ (
    .A1(\rf[16] [16]),
    .A2(_03046_),
    .ZN(_05107_)
  );
  AND2_X1 _12626_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05107_),
    .ZN(_05108_)
  );
  AND2_X1 _12627_ (
    .A1(_05106_),
    .A2(_05108_),
    .ZN(_05109_)
  );
  MUX2_X1 _12628_ (
    .A(\rf[22] [16]),
    .B(\rf[18] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05110_)
  );
  AND2_X1 _12629_ (
    .A1(_03045_),
    .A2(_05110_),
    .ZN(_05111_)
  );
  OR2_X1 _12630_ (
    .A1(_03044_),
    .A2(_05111_),
    .ZN(_05112_)
  );
  OR2_X1 _12631_ (
    .A1(_05109_),
    .A2(_05112_),
    .ZN(_05113_)
  );
  OR2_X1 _12632_ (
    .A1(\rf[17] [16]),
    .A2(_03046_),
    .ZN(_05114_)
  );
  OR2_X1 _12633_ (
    .A1(\rf[21] [16]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05115_)
  );
  AND2_X1 _12634_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05115_),
    .ZN(_05116_)
  );
  AND2_X1 _12635_ (
    .A1(_05114_),
    .A2(_05116_),
    .ZN(_05117_)
  );
  MUX2_X1 _12636_ (
    .A(\rf[23] [16]),
    .B(\rf[19] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05118_)
  );
  AND2_X1 _12637_ (
    .A1(_03045_),
    .A2(_05118_),
    .ZN(_05119_)
  );
  OR2_X1 _12638_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05119_),
    .ZN(_05120_)
  );
  OR2_X1 _12639_ (
    .A1(_05117_),
    .A2(_05120_),
    .ZN(_05121_)
  );
  AND2_X1 _12640_ (
    .A1(_05113_),
    .A2(_05121_),
    .ZN(_05122_)
  );
  OR2_X1 _12641_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_05122_),
    .ZN(_05123_)
  );
  AND2_X1 _12642_ (
    .A1(_05105_),
    .A2(_05123_),
    .ZN(_05124_)
  );
  AND2_X1 _12643_ (
    .A1(\rf[10] [16]),
    .A2(_03045_),
    .ZN(_05125_)
  );
  AND2_X1 _12644_ (
    .A1(\rf[8] [16]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05126_)
  );
  OR2_X1 _12645_ (
    .A1(_03046_),
    .A2(_05126_),
    .ZN(_05127_)
  );
  OR2_X1 _12646_ (
    .A1(_05125_),
    .A2(_05127_),
    .ZN(_05128_)
  );
  AND2_X1 _12647_ (
    .A1(\rf[14] [16]),
    .A2(_03045_),
    .ZN(_05129_)
  );
  AND2_X1 _12648_ (
    .A1(\rf[12] [16]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05130_)
  );
  OR2_X1 _12649_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_05130_),
    .ZN(_05131_)
  );
  OR2_X1 _12650_ (
    .A1(_05129_),
    .A2(_05131_),
    .ZN(_05132_)
  );
  AND2_X1 _12651_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05132_),
    .ZN(_05133_)
  );
  AND2_X1 _12652_ (
    .A1(_05128_),
    .A2(_05133_),
    .ZN(_05134_)
  );
  AND2_X1 _12653_ (
    .A1(\rf[11] [16]),
    .A2(_03045_),
    .ZN(_05135_)
  );
  AND2_X1 _12654_ (
    .A1(\rf[9] [16]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05136_)
  );
  OR2_X1 _12655_ (
    .A1(_03046_),
    .A2(_05136_),
    .ZN(_05137_)
  );
  OR2_X1 _12656_ (
    .A1(_05135_),
    .A2(_05137_),
    .ZN(_05138_)
  );
  AND2_X1 _12657_ (
    .A1(\rf[15] [16]),
    .A2(_03045_),
    .ZN(_05139_)
  );
  AND2_X1 _12658_ (
    .A1(\rf[13] [16]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05140_)
  );
  OR2_X1 _12659_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_05140_),
    .ZN(_05141_)
  );
  OR2_X1 _12660_ (
    .A1(_05139_),
    .A2(_05141_),
    .ZN(_05142_)
  );
  AND2_X1 _12661_ (
    .A1(_03044_),
    .A2(_05142_),
    .ZN(_05143_)
  );
  AND2_X1 _12662_ (
    .A1(_05138_),
    .A2(_05143_),
    .ZN(_05144_)
  );
  OR2_X1 _12663_ (
    .A1(_03063_),
    .A2(_05144_),
    .ZN(_05145_)
  );
  OR2_X1 _12664_ (
    .A1(_05134_),
    .A2(_05145_),
    .ZN(_05146_)
  );
  OR2_X1 _12665_ (
    .A1(\rf[28] [16]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05147_)
  );
  OR2_X1 _12666_ (
    .A1(\rf[24] [16]),
    .A2(_03046_),
    .ZN(_05148_)
  );
  AND2_X1 _12667_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05147_),
    .ZN(_05149_)
  );
  AND2_X1 _12668_ (
    .A1(_05148_),
    .A2(_05149_),
    .ZN(_05150_)
  );
  MUX2_X1 _12669_ (
    .A(\rf[30] [16]),
    .B(\rf[26] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05151_)
  );
  AND2_X1 _12670_ (
    .A1(_03045_),
    .A2(_05151_),
    .ZN(_05152_)
  );
  OR2_X1 _12671_ (
    .A1(_03044_),
    .A2(_05152_),
    .ZN(_05153_)
  );
  OR2_X1 _12672_ (
    .A1(_05150_),
    .A2(_05153_),
    .ZN(_05154_)
  );
  MUX2_X1 _12673_ (
    .A(\rf[29] [16]),
    .B(\rf[25] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05155_)
  );
  AND2_X1 _12674_ (
    .A1(\rf[27] [16]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05156_)
  );
  MUX2_X1 _12675_ (
    .A(_05155_),
    .B(_05156_),
    .S(_03045_),
    .Z(_05157_)
  );
  OR2_X1 _12676_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05157_),
    .ZN(_05158_)
  );
  AND2_X1 _12677_ (
    .A1(_05154_),
    .A2(_05158_),
    .ZN(_05159_)
  );
  OR2_X1 _12678_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_05159_),
    .ZN(_05160_)
  );
  AND2_X1 _12679_ (
    .A1(_05146_),
    .A2(_05160_),
    .ZN(_05161_)
  );
  MUX2_X1 _12680_ (
    .A(_05124_),
    .B(_05161_),
    .S(_03047_),
    .Z(_05162_)
  );
  MUX2_X1 _12681_ (
    .A(_05162_),
    .B(_05095_),
    .S(_04074_),
    .Z(_05163_)
  );
  AND2_X1 _12682_ (
    .A1(_04044_),
    .A2(_05163_),
    .ZN(_05164_)
  );
  OR2_X1 _12683_ (
    .A1(_05092_),
    .A2(_05164_),
    .ZN(_05165_)
  );
  MUX2_X1 _12684_ (
    .A(ex_reg_rs_msb_0[14]),
    .B(_05165_),
    .S(_04042_),
    .Z(_00081_)
  );
  AND2_X1 _12685_ (
    .A1(_03065_),
    .A2(ibuf_io_inst_0_bits_raw[17]),
    .ZN(_05166_)
  );
  AND2_X1 _12686_ (
    .A1(_03582_),
    .A2(_05166_),
    .ZN(_05167_)
  );
  MUX2_X1 _12687_ (
    .A(wb_reg_wdata[17]),
    .B(csr_io_rw_rdata[17]),
    .S(_04077_),
    .Z(_05168_)
  );
  MUX2_X1 _12688_ (
    .A(div_io_resp_bits_data[17]),
    .B(_05168_),
    .S(_03114_),
    .Z(_05169_)
  );
  MUX2_X1 _12689_ (
    .A(_05169_),
    .B(io_dmem_resp_bits_data[17]),
    .S(_03097_),
    .Z(_05170_)
  );
  MUX2_X1 _12690_ (
    .A(\rf[5] [17]),
    .B(\rf[1] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05171_)
  );
  MUX2_X1 _12691_ (
    .A(\rf[7] [17]),
    .B(\rf[3] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05172_)
  );
  MUX2_X1 _12692_ (
    .A(_05171_),
    .B(_05172_),
    .S(_03045_),
    .Z(_05173_)
  );
  AND2_X1 _12693_ (
    .A1(_03044_),
    .A2(_05173_),
    .ZN(_05174_)
  );
  MUX2_X1 _12694_ (
    .A(\rf[4] [17]),
    .B(\rf[0] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05175_)
  );
  MUX2_X1 _12695_ (
    .A(\rf[6] [17]),
    .B(\rf[2] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05176_)
  );
  MUX2_X1 _12696_ (
    .A(_05175_),
    .B(_05176_),
    .S(_03045_),
    .Z(_05177_)
  );
  AND2_X1 _12697_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05177_),
    .ZN(_05178_)
  );
  OR2_X1 _12698_ (
    .A1(_03063_),
    .A2(_05178_),
    .ZN(_05179_)
  );
  OR2_X1 _12699_ (
    .A1(_05174_),
    .A2(_05179_),
    .ZN(_05180_)
  );
  OR2_X1 _12700_ (
    .A1(\rf[20] [17]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05181_)
  );
  OR2_X1 _12701_ (
    .A1(\rf[16] [17]),
    .A2(_03046_),
    .ZN(_05182_)
  );
  AND2_X1 _12702_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05182_),
    .ZN(_05183_)
  );
  AND2_X1 _12703_ (
    .A1(_05181_),
    .A2(_05183_),
    .ZN(_05184_)
  );
  MUX2_X1 _12704_ (
    .A(\rf[22] [17]),
    .B(\rf[18] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05185_)
  );
  AND2_X1 _12705_ (
    .A1(_03045_),
    .A2(_05185_),
    .ZN(_05186_)
  );
  OR2_X1 _12706_ (
    .A1(_03044_),
    .A2(_05186_),
    .ZN(_05187_)
  );
  OR2_X1 _12707_ (
    .A1(_05184_),
    .A2(_05187_),
    .ZN(_05188_)
  );
  OR2_X1 _12708_ (
    .A1(\rf[17] [17]),
    .A2(_03046_),
    .ZN(_05189_)
  );
  OR2_X1 _12709_ (
    .A1(\rf[21] [17]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05190_)
  );
  AND2_X1 _12710_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05190_),
    .ZN(_05191_)
  );
  AND2_X1 _12711_ (
    .A1(_05189_),
    .A2(_05191_),
    .ZN(_05192_)
  );
  MUX2_X1 _12712_ (
    .A(\rf[23] [17]),
    .B(\rf[19] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05193_)
  );
  AND2_X1 _12713_ (
    .A1(_03045_),
    .A2(_05193_),
    .ZN(_05194_)
  );
  OR2_X1 _12714_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05194_),
    .ZN(_05195_)
  );
  OR2_X1 _12715_ (
    .A1(_05192_),
    .A2(_05195_),
    .ZN(_05196_)
  );
  AND2_X1 _12716_ (
    .A1(_05188_),
    .A2(_05196_),
    .ZN(_05197_)
  );
  OR2_X1 _12717_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_05197_),
    .ZN(_05198_)
  );
  AND2_X1 _12718_ (
    .A1(_05180_),
    .A2(_05198_),
    .ZN(_05199_)
  );
  AND2_X1 _12719_ (
    .A1(\rf[10] [17]),
    .A2(_03045_),
    .ZN(_05200_)
  );
  AND2_X1 _12720_ (
    .A1(\rf[8] [17]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05201_)
  );
  OR2_X1 _12721_ (
    .A1(_03046_),
    .A2(_05201_),
    .ZN(_05202_)
  );
  OR2_X1 _12722_ (
    .A1(_05200_),
    .A2(_05202_),
    .ZN(_05203_)
  );
  AND2_X1 _12723_ (
    .A1(\rf[14] [17]),
    .A2(_03045_),
    .ZN(_05204_)
  );
  AND2_X1 _12724_ (
    .A1(\rf[12] [17]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05205_)
  );
  OR2_X1 _12725_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_05205_),
    .ZN(_05206_)
  );
  OR2_X1 _12726_ (
    .A1(_05204_),
    .A2(_05206_),
    .ZN(_05207_)
  );
  AND2_X1 _12727_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05207_),
    .ZN(_05208_)
  );
  AND2_X1 _12728_ (
    .A1(_05203_),
    .A2(_05208_),
    .ZN(_05209_)
  );
  AND2_X1 _12729_ (
    .A1(\rf[11] [17]),
    .A2(_03045_),
    .ZN(_05210_)
  );
  AND2_X1 _12730_ (
    .A1(\rf[9] [17]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05211_)
  );
  OR2_X1 _12731_ (
    .A1(_03046_),
    .A2(_05211_),
    .ZN(_05212_)
  );
  OR2_X1 _12732_ (
    .A1(_05210_),
    .A2(_05212_),
    .ZN(_05213_)
  );
  AND2_X1 _12733_ (
    .A1(\rf[15] [17]),
    .A2(_03045_),
    .ZN(_05214_)
  );
  AND2_X1 _12734_ (
    .A1(\rf[13] [17]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05215_)
  );
  OR2_X1 _12735_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_05215_),
    .ZN(_05216_)
  );
  OR2_X1 _12736_ (
    .A1(_05214_),
    .A2(_05216_),
    .ZN(_05217_)
  );
  AND2_X1 _12737_ (
    .A1(_03044_),
    .A2(_05217_),
    .ZN(_05218_)
  );
  AND2_X1 _12738_ (
    .A1(_05213_),
    .A2(_05218_),
    .ZN(_05219_)
  );
  OR2_X1 _12739_ (
    .A1(_03063_),
    .A2(_05219_),
    .ZN(_05220_)
  );
  OR2_X1 _12740_ (
    .A1(_05209_),
    .A2(_05220_),
    .ZN(_05221_)
  );
  OR2_X1 _12741_ (
    .A1(\rf[28] [17]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05222_)
  );
  OR2_X1 _12742_ (
    .A1(\rf[24] [17]),
    .A2(_03046_),
    .ZN(_05223_)
  );
  AND2_X1 _12743_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05222_),
    .ZN(_05224_)
  );
  AND2_X1 _12744_ (
    .A1(_05223_),
    .A2(_05224_),
    .ZN(_05225_)
  );
  MUX2_X1 _12745_ (
    .A(\rf[30] [17]),
    .B(\rf[26] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05226_)
  );
  AND2_X1 _12746_ (
    .A1(_03045_),
    .A2(_05226_),
    .ZN(_05227_)
  );
  OR2_X1 _12747_ (
    .A1(_03044_),
    .A2(_05227_),
    .ZN(_05228_)
  );
  OR2_X1 _12748_ (
    .A1(_05225_),
    .A2(_05228_),
    .ZN(_05229_)
  );
  MUX2_X1 _12749_ (
    .A(\rf[29] [17]),
    .B(\rf[25] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05230_)
  );
  AND2_X1 _12750_ (
    .A1(\rf[27] [17]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05231_)
  );
  MUX2_X1 _12751_ (
    .A(_05230_),
    .B(_05231_),
    .S(_03045_),
    .Z(_05232_)
  );
  OR2_X1 _12752_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05232_),
    .ZN(_05233_)
  );
  AND2_X1 _12753_ (
    .A1(_05229_),
    .A2(_05233_),
    .ZN(_05234_)
  );
  OR2_X1 _12754_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_05234_),
    .ZN(_05235_)
  );
  AND2_X1 _12755_ (
    .A1(_05221_),
    .A2(_05235_),
    .ZN(_05236_)
  );
  MUX2_X1 _12756_ (
    .A(_05199_),
    .B(_05236_),
    .S(_03047_),
    .Z(_05237_)
  );
  MUX2_X1 _12757_ (
    .A(_05237_),
    .B(_05170_),
    .S(_04074_),
    .Z(_05238_)
  );
  AND2_X1 _12758_ (
    .A1(_04044_),
    .A2(_05238_),
    .ZN(_05239_)
  );
  OR2_X1 _12759_ (
    .A1(_05167_),
    .A2(_05239_),
    .ZN(_05240_)
  );
  MUX2_X1 _12760_ (
    .A(ex_reg_rs_msb_0[15]),
    .B(_05240_),
    .S(_04042_),
    .Z(_00082_)
  );
  AND2_X1 _12761_ (
    .A1(_03065_),
    .A2(ibuf_io_inst_0_bits_raw[18]),
    .ZN(_05241_)
  );
  AND2_X1 _12762_ (
    .A1(_03582_),
    .A2(_05241_),
    .ZN(_05242_)
  );
  MUX2_X1 _12763_ (
    .A(\rf[3] [18]),
    .B(\rf[2] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_05243_)
  );
  MUX2_X1 _12764_ (
    .A(\rf[7] [18]),
    .B(\rf[6] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_05244_)
  );
  MUX2_X1 _12765_ (
    .A(_05243_),
    .B(_05244_),
    .S(_03046_),
    .Z(_05245_)
  );
  OR2_X1 _12766_ (
    .A1(_03047_),
    .A2(_05245_),
    .ZN(_05246_)
  );
  MUX2_X1 _12767_ (
    .A(\rf[14] [18]),
    .B(\rf[10] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05247_)
  );
  OR2_X1 _12768_ (
    .A1(_04124_),
    .A2(_05247_),
    .ZN(_05248_)
  );
  MUX2_X1 _12769_ (
    .A(\rf[15] [18]),
    .B(\rf[11] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05249_)
  );
  OR2_X1 _12770_ (
    .A1(_03448_),
    .A2(_05249_),
    .ZN(_05250_)
  );
  AND2_X1 _12771_ (
    .A1(_03045_),
    .A2(_05250_),
    .ZN(_05251_)
  );
  AND2_X1 _12772_ (
    .A1(_05248_),
    .A2(_05251_),
    .ZN(_05252_)
  );
  AND2_X1 _12773_ (
    .A1(_05246_),
    .A2(_05252_),
    .ZN(_05253_)
  );
  MUX2_X1 _12774_ (
    .A(\rf[1] [18]),
    .B(\rf[0] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_05254_)
  );
  MUX2_X1 _12775_ (
    .A(\rf[5] [18]),
    .B(\rf[4] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_05255_)
  );
  MUX2_X1 _12776_ (
    .A(_05254_),
    .B(_05255_),
    .S(_03046_),
    .Z(_05256_)
  );
  OR2_X1 _12777_ (
    .A1(_03047_),
    .A2(_05256_),
    .ZN(_05257_)
  );
  MUX2_X1 _12778_ (
    .A(\rf[13] [18]),
    .B(\rf[9] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05258_)
  );
  OR2_X1 _12779_ (
    .A1(_03448_),
    .A2(_05258_),
    .ZN(_05259_)
  );
  MUX2_X1 _12780_ (
    .A(\rf[12] [18]),
    .B(\rf[8] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05260_)
  );
  OR2_X1 _12781_ (
    .A1(_04124_),
    .A2(_05260_),
    .ZN(_05261_)
  );
  AND2_X1 _12782_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05259_),
    .ZN(_05262_)
  );
  AND2_X1 _12783_ (
    .A1(_05261_),
    .A2(_05262_),
    .ZN(_05263_)
  );
  AND2_X1 _12784_ (
    .A1(_05257_),
    .A2(_05263_),
    .ZN(_05264_)
  );
  OR2_X1 _12785_ (
    .A1(_03063_),
    .A2(_05264_),
    .ZN(_05265_)
  );
  OR2_X1 _12786_ (
    .A1(_05253_),
    .A2(_05265_),
    .ZN(_05266_)
  );
  OR2_X1 _12787_ (
    .A1(\rf[28] [18]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05267_)
  );
  OR2_X1 _12788_ (
    .A1(\rf[24] [18]),
    .A2(_03046_),
    .ZN(_05268_)
  );
  AND2_X1 _12789_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05267_),
    .ZN(_05269_)
  );
  AND2_X1 _12790_ (
    .A1(_05268_),
    .A2(_05269_),
    .ZN(_05270_)
  );
  MUX2_X1 _12791_ (
    .A(\rf[30] [18]),
    .B(\rf[26] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05271_)
  );
  AND2_X1 _12792_ (
    .A1(_03045_),
    .A2(_05271_),
    .ZN(_05272_)
  );
  OR2_X1 _12793_ (
    .A1(_03044_),
    .A2(_05272_),
    .ZN(_05273_)
  );
  OR2_X1 _12794_ (
    .A1(_05270_),
    .A2(_05273_),
    .ZN(_05274_)
  );
  MUX2_X1 _12795_ (
    .A(\rf[29] [18]),
    .B(\rf[25] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05275_)
  );
  AND2_X1 _12796_ (
    .A1(\rf[27] [18]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05276_)
  );
  MUX2_X1 _12797_ (
    .A(_05275_),
    .B(_05276_),
    .S(_03045_),
    .Z(_05277_)
  );
  OR2_X1 _12798_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05277_),
    .ZN(_05278_)
  );
  AND2_X1 _12799_ (
    .A1(_05274_),
    .A2(_05278_),
    .ZN(_05279_)
  );
  OR2_X1 _12800_ (
    .A1(\rf[20] [18]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05280_)
  );
  OR2_X1 _12801_ (
    .A1(\rf[16] [18]),
    .A2(_03046_),
    .ZN(_05281_)
  );
  AND2_X1 _12802_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05281_),
    .ZN(_05282_)
  );
  AND2_X1 _12803_ (
    .A1(_05280_),
    .A2(_05282_),
    .ZN(_05283_)
  );
  MUX2_X1 _12804_ (
    .A(\rf[22] [18]),
    .B(\rf[18] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05284_)
  );
  AND2_X1 _12805_ (
    .A1(_03045_),
    .A2(_05284_),
    .ZN(_05285_)
  );
  OR2_X1 _12806_ (
    .A1(_03044_),
    .A2(_05285_),
    .ZN(_05286_)
  );
  OR2_X1 _12807_ (
    .A1(_05283_),
    .A2(_05286_),
    .ZN(_05287_)
  );
  OR2_X1 _12808_ (
    .A1(\rf[17] [18]),
    .A2(_03046_),
    .ZN(_05288_)
  );
  OR2_X1 _12809_ (
    .A1(\rf[21] [18]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05289_)
  );
  AND2_X1 _12810_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05289_),
    .ZN(_05290_)
  );
  AND2_X1 _12811_ (
    .A1(_05288_),
    .A2(_05290_),
    .ZN(_05291_)
  );
  MUX2_X1 _12812_ (
    .A(\rf[23] [18]),
    .B(\rf[19] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05292_)
  );
  AND2_X1 _12813_ (
    .A1(_03045_),
    .A2(_05292_),
    .ZN(_05293_)
  );
  OR2_X1 _12814_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05293_),
    .ZN(_05294_)
  );
  OR2_X1 _12815_ (
    .A1(_05291_),
    .A2(_05294_),
    .ZN(_05295_)
  );
  AND2_X1 _12816_ (
    .A1(_05287_),
    .A2(_05295_),
    .ZN(_05296_)
  );
  MUX2_X1 _12817_ (
    .A(_05279_),
    .B(_05296_),
    .S(ibuf_io_inst_0_bits_inst_rs1[3]),
    .Z(_05297_)
  );
  OR2_X1 _12818_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_05297_),
    .ZN(_05298_)
  );
  AND2_X1 _12819_ (
    .A1(_05266_),
    .A2(_05298_),
    .ZN(_05299_)
  );
  MUX2_X1 _12820_ (
    .A(wb_reg_wdata[18]),
    .B(csr_io_rw_rdata[18]),
    .S(_04077_),
    .Z(_05300_)
  );
  MUX2_X1 _12821_ (
    .A(div_io_resp_bits_data[18]),
    .B(_05300_),
    .S(_03114_),
    .Z(_05301_)
  );
  MUX2_X1 _12822_ (
    .A(_05301_),
    .B(io_dmem_resp_bits_data[18]),
    .S(_03097_),
    .Z(_05302_)
  );
  MUX2_X1 _12823_ (
    .A(_05299_),
    .B(_05302_),
    .S(_04074_),
    .Z(_05303_)
  );
  AND2_X1 _12824_ (
    .A1(_04044_),
    .A2(_05303_),
    .ZN(_05304_)
  );
  OR2_X1 _12825_ (
    .A1(_05242_),
    .A2(_05304_),
    .ZN(_05305_)
  );
  MUX2_X1 _12826_ (
    .A(ex_reg_rs_msb_0[16]),
    .B(_05305_),
    .S(_04042_),
    .Z(_00083_)
  );
  AND2_X1 _12827_ (
    .A1(_03065_),
    .A2(ibuf_io_inst_0_bits_raw[19]),
    .ZN(_05306_)
  );
  AND2_X1 _12828_ (
    .A1(_03582_),
    .A2(_05306_),
    .ZN(_05307_)
  );
  MUX2_X1 _12829_ (
    .A(wb_reg_wdata[19]),
    .B(csr_io_rw_rdata[19]),
    .S(_04077_),
    .Z(_05308_)
  );
  MUX2_X1 _12830_ (
    .A(div_io_resp_bits_data[19]),
    .B(_05308_),
    .S(_03114_),
    .Z(_05309_)
  );
  MUX2_X1 _12831_ (
    .A(_05309_),
    .B(io_dmem_resp_bits_data[19]),
    .S(_03097_),
    .Z(_05310_)
  );
  MUX2_X1 _12832_ (
    .A(\rf[1] [19]),
    .B(\rf[0] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_05311_)
  );
  MUX2_X1 _12833_ (
    .A(\rf[5] [19]),
    .B(\rf[4] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_05312_)
  );
  MUX2_X1 _12834_ (
    .A(_05311_),
    .B(_05312_),
    .S(_03046_),
    .Z(_05313_)
  );
  OR2_X1 _12835_ (
    .A1(_03047_),
    .A2(_05313_),
    .ZN(_05314_)
  );
  MUX2_X1 _12836_ (
    .A(\rf[12] [19]),
    .B(\rf[8] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05315_)
  );
  OR2_X1 _12837_ (
    .A1(_04124_),
    .A2(_05315_),
    .ZN(_05316_)
  );
  MUX2_X1 _12838_ (
    .A(\rf[13] [19]),
    .B(\rf[9] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05317_)
  );
  OR2_X1 _12839_ (
    .A1(_03448_),
    .A2(_05317_),
    .ZN(_05318_)
  );
  AND2_X1 _12840_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05318_),
    .ZN(_05319_)
  );
  AND2_X1 _12841_ (
    .A1(_05316_),
    .A2(_05319_),
    .ZN(_05320_)
  );
  AND2_X1 _12842_ (
    .A1(_05314_),
    .A2(_05320_),
    .ZN(_05321_)
  );
  MUX2_X1 _12843_ (
    .A(\rf[3] [19]),
    .B(\rf[2] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_05322_)
  );
  MUX2_X1 _12844_ (
    .A(\rf[7] [19]),
    .B(\rf[6] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_05323_)
  );
  MUX2_X1 _12845_ (
    .A(_05322_),
    .B(_05323_),
    .S(_03046_),
    .Z(_05324_)
  );
  OR2_X1 _12846_ (
    .A1(_03047_),
    .A2(_05324_),
    .ZN(_05325_)
  );
  MUX2_X1 _12847_ (
    .A(\rf[14] [19]),
    .B(\rf[10] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05326_)
  );
  OR2_X1 _12848_ (
    .A1(_04124_),
    .A2(_05326_),
    .ZN(_05327_)
  );
  MUX2_X1 _12849_ (
    .A(\rf[15] [19]),
    .B(\rf[11] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05328_)
  );
  OR2_X1 _12850_ (
    .A1(_03448_),
    .A2(_05328_),
    .ZN(_05329_)
  );
  AND2_X1 _12851_ (
    .A1(_03045_),
    .A2(_05329_),
    .ZN(_05330_)
  );
  AND2_X1 _12852_ (
    .A1(_05327_),
    .A2(_05330_),
    .ZN(_05331_)
  );
  AND2_X1 _12853_ (
    .A1(_05325_),
    .A2(_05331_),
    .ZN(_05332_)
  );
  OR2_X1 _12854_ (
    .A1(\rf[28] [19]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05333_)
  );
  OR2_X1 _12855_ (
    .A1(\rf[24] [19]),
    .A2(_03046_),
    .ZN(_05334_)
  );
  AND2_X1 _12856_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05333_),
    .ZN(_05335_)
  );
  AND2_X1 _12857_ (
    .A1(_05334_),
    .A2(_05335_),
    .ZN(_05336_)
  );
  MUX2_X1 _12858_ (
    .A(\rf[30] [19]),
    .B(\rf[26] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05337_)
  );
  AND2_X1 _12859_ (
    .A1(_03045_),
    .A2(_05337_),
    .ZN(_05338_)
  );
  OR2_X1 _12860_ (
    .A1(_03044_),
    .A2(_05338_),
    .ZN(_05339_)
  );
  OR2_X1 _12861_ (
    .A1(_05336_),
    .A2(_05339_),
    .ZN(_05340_)
  );
  MUX2_X1 _12862_ (
    .A(\rf[29] [19]),
    .B(\rf[25] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05341_)
  );
  AND2_X1 _12863_ (
    .A1(\rf[27] [19]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05342_)
  );
  MUX2_X1 _12864_ (
    .A(_05341_),
    .B(_05342_),
    .S(_03045_),
    .Z(_05343_)
  );
  OR2_X1 _12865_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05343_),
    .ZN(_05344_)
  );
  AND2_X1 _12866_ (
    .A1(_05340_),
    .A2(_05344_),
    .ZN(_05345_)
  );
  OR2_X1 _12867_ (
    .A1(\rf[20] [19]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05346_)
  );
  OR2_X1 _12868_ (
    .A1(\rf[16] [19]),
    .A2(_03046_),
    .ZN(_05347_)
  );
  AND2_X1 _12869_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05347_),
    .ZN(_05348_)
  );
  AND2_X1 _12870_ (
    .A1(_05346_),
    .A2(_05348_),
    .ZN(_05349_)
  );
  MUX2_X1 _12871_ (
    .A(\rf[22] [19]),
    .B(\rf[18] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05350_)
  );
  AND2_X1 _12872_ (
    .A1(_03045_),
    .A2(_05350_),
    .ZN(_05351_)
  );
  OR2_X1 _12873_ (
    .A1(_03044_),
    .A2(_05351_),
    .ZN(_05352_)
  );
  OR2_X1 _12874_ (
    .A1(_05349_),
    .A2(_05352_),
    .ZN(_05353_)
  );
  OR2_X1 _12875_ (
    .A1(\rf[17] [19]),
    .A2(_03046_),
    .ZN(_05354_)
  );
  OR2_X1 _12876_ (
    .A1(\rf[21] [19]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05355_)
  );
  AND2_X1 _12877_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05355_),
    .ZN(_05356_)
  );
  AND2_X1 _12878_ (
    .A1(_05354_),
    .A2(_05356_),
    .ZN(_05357_)
  );
  MUX2_X1 _12879_ (
    .A(\rf[23] [19]),
    .B(\rf[19] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05358_)
  );
  AND2_X1 _12880_ (
    .A1(_03045_),
    .A2(_05358_),
    .ZN(_05359_)
  );
  OR2_X1 _12881_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05359_),
    .ZN(_05360_)
  );
  OR2_X1 _12882_ (
    .A1(_05357_),
    .A2(_05360_),
    .ZN(_05361_)
  );
  AND2_X1 _12883_ (
    .A1(_05353_),
    .A2(_05361_),
    .ZN(_05362_)
  );
  MUX2_X1 _12884_ (
    .A(_05345_),
    .B(_05362_),
    .S(ibuf_io_inst_0_bits_inst_rs1[3]),
    .Z(_05363_)
  );
  OR2_X1 _12885_ (
    .A1(_05321_),
    .A2(_05332_),
    .ZN(_05364_)
  );
  MUX2_X1 _12886_ (
    .A(_05363_),
    .B(_05364_),
    .S(ibuf_io_inst_0_bits_inst_rs1[4]),
    .Z(_05365_)
  );
  MUX2_X1 _12887_ (
    .A(_05365_),
    .B(_05310_),
    .S(_04074_),
    .Z(_05366_)
  );
  AND2_X1 _12888_ (
    .A1(_04044_),
    .A2(_05366_),
    .ZN(_05367_)
  );
  OR2_X1 _12889_ (
    .A1(_05307_),
    .A2(_05367_),
    .ZN(_05368_)
  );
  MUX2_X1 _12890_ (
    .A(ex_reg_rs_msb_0[17]),
    .B(_05368_),
    .S(_04042_),
    .Z(_00084_)
  );
  AND2_X1 _12891_ (
    .A1(_03065_),
    .A2(ibuf_io_inst_0_bits_raw[20]),
    .ZN(_05369_)
  );
  AND2_X1 _12892_ (
    .A1(_03582_),
    .A2(_05369_),
    .ZN(_05370_)
  );
  OR2_X1 _12893_ (
    .A1(\rf[10] [20]),
    .A2(_03046_),
    .ZN(_05371_)
  );
  OR2_X1 _12894_ (
    .A1(\rf[14] [20]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05372_)
  );
  AND2_X1 _12895_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05372_),
    .ZN(_05373_)
  );
  AND2_X1 _12896_ (
    .A1(_05371_),
    .A2(_05373_),
    .ZN(_05374_)
  );
  MUX2_X1 _12897_ (
    .A(\rf[15] [20]),
    .B(\rf[11] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05375_)
  );
  AND2_X1 _12898_ (
    .A1(_03044_),
    .A2(_05375_),
    .ZN(_05376_)
  );
  OR2_X1 _12899_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05376_),
    .ZN(_05377_)
  );
  OR2_X1 _12900_ (
    .A1(_05374_),
    .A2(_05377_),
    .ZN(_05378_)
  );
  OR2_X1 _12901_ (
    .A1(\rf[12] [20]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05379_)
  );
  OR2_X1 _12902_ (
    .A1(\rf[8] [20]),
    .A2(_03046_),
    .ZN(_05380_)
  );
  AND2_X1 _12903_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05379_),
    .ZN(_05381_)
  );
  AND2_X1 _12904_ (
    .A1(_05380_),
    .A2(_05381_),
    .ZN(_05382_)
  );
  MUX2_X1 _12905_ (
    .A(\rf[13] [20]),
    .B(\rf[9] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05383_)
  );
  AND2_X1 _12906_ (
    .A1(_03044_),
    .A2(_05383_),
    .ZN(_05384_)
  );
  OR2_X1 _12907_ (
    .A1(_03045_),
    .A2(_05384_),
    .ZN(_05385_)
  );
  OR2_X1 _12908_ (
    .A1(_05382_),
    .A2(_05385_),
    .ZN(_05386_)
  );
  AND2_X1 _12909_ (
    .A1(_03047_),
    .A2(_05386_),
    .ZN(_05387_)
  );
  AND2_X1 _12910_ (
    .A1(_05378_),
    .A2(_05387_),
    .ZN(_05388_)
  );
  OR2_X1 _12911_ (
    .A1(\rf[0] [20]),
    .A2(_03046_),
    .ZN(_05389_)
  );
  OR2_X1 _12912_ (
    .A1(\rf[4] [20]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05390_)
  );
  AND2_X1 _12913_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05390_),
    .ZN(_05391_)
  );
  AND2_X1 _12914_ (
    .A1(_05389_),
    .A2(_05391_),
    .ZN(_05392_)
  );
  MUX2_X1 _12915_ (
    .A(\rf[5] [20]),
    .B(\rf[1] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05393_)
  );
  AND2_X1 _12916_ (
    .A1(_03044_),
    .A2(_05393_),
    .ZN(_05394_)
  );
  OR2_X1 _12917_ (
    .A1(_03045_),
    .A2(_05394_),
    .ZN(_05395_)
  );
  OR2_X1 _12918_ (
    .A1(_05392_),
    .A2(_05395_),
    .ZN(_05396_)
  );
  MUX2_X1 _12919_ (
    .A(\rf[7] [20]),
    .B(\rf[3] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05397_)
  );
  AND2_X1 _12920_ (
    .A1(_03044_),
    .A2(_05397_),
    .ZN(_05398_)
  );
  OR2_X1 _12921_ (
    .A1(\rf[2] [20]),
    .A2(_03046_),
    .ZN(_05399_)
  );
  OR2_X1 _12922_ (
    .A1(\rf[6] [20]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05400_)
  );
  AND2_X1 _12923_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05400_),
    .ZN(_05401_)
  );
  AND2_X1 _12924_ (
    .A1(_05399_),
    .A2(_05401_),
    .ZN(_05402_)
  );
  OR2_X1 _12925_ (
    .A1(_05398_),
    .A2(_05402_),
    .ZN(_05403_)
  );
  OR2_X1 _12926_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05403_),
    .ZN(_05404_)
  );
  AND2_X1 _12927_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_05396_),
    .ZN(_05405_)
  );
  AND2_X1 _12928_ (
    .A1(_05404_),
    .A2(_05405_),
    .ZN(_05406_)
  );
  OR2_X1 _12929_ (
    .A1(_05388_),
    .A2(_05406_),
    .ZN(_05407_)
  );
  MUX2_X1 _12930_ (
    .A(\rf[30] [20]),
    .B(\rf[26] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05408_)
  );
  AND2_X1 _12931_ (
    .A1(\rf[27] [20]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05409_)
  );
  MUX2_X1 _12932_ (
    .A(_05408_),
    .B(_05409_),
    .S(_03044_),
    .Z(_05410_)
  );
  MUX2_X1 _12933_ (
    .A(\rf[29] [20]),
    .B(\rf[25] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05411_)
  );
  AND2_X1 _12934_ (
    .A1(_03044_),
    .A2(_05411_),
    .ZN(_05412_)
  );
  MUX2_X1 _12935_ (
    .A(\rf[28] [20]),
    .B(\rf[24] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05413_)
  );
  AND2_X1 _12936_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05413_),
    .ZN(_05414_)
  );
  OR2_X1 _12937_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05410_),
    .ZN(_05415_)
  );
  OR2_X1 _12938_ (
    .A1(_03045_),
    .A2(_05414_),
    .ZN(_05416_)
  );
  OR2_X1 _12939_ (
    .A1(_05412_),
    .A2(_05416_),
    .ZN(_05417_)
  );
  AND2_X1 _12940_ (
    .A1(_03047_),
    .A2(_05415_),
    .ZN(_05418_)
  );
  AND2_X1 _12941_ (
    .A1(_05417_),
    .A2(_05418_),
    .ZN(_05419_)
  );
  OR2_X1 _12942_ (
    .A1(\rf[18] [20]),
    .A2(_03046_),
    .ZN(_05420_)
  );
  OR2_X1 _12943_ (
    .A1(\rf[22] [20]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05421_)
  );
  AND2_X1 _12944_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05421_),
    .ZN(_05422_)
  );
  AND2_X1 _12945_ (
    .A1(_05420_),
    .A2(_05422_),
    .ZN(_05423_)
  );
  MUX2_X1 _12946_ (
    .A(\rf[23] [20]),
    .B(\rf[19] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05424_)
  );
  AND2_X1 _12947_ (
    .A1(_03044_),
    .A2(_05424_),
    .ZN(_05425_)
  );
  OR2_X1 _12948_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05425_),
    .ZN(_05426_)
  );
  OR2_X1 _12949_ (
    .A1(_05423_),
    .A2(_05426_),
    .ZN(_05427_)
  );
  MUX2_X1 _12950_ (
    .A(\rf[21] [20]),
    .B(\rf[17] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05428_)
  );
  AND2_X1 _12951_ (
    .A1(_03044_),
    .A2(_05428_),
    .ZN(_05429_)
  );
  OR2_X1 _12952_ (
    .A1(\rf[20] [20]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05430_)
  );
  OR2_X1 _12953_ (
    .A1(\rf[16] [20]),
    .A2(_03046_),
    .ZN(_05431_)
  );
  AND2_X1 _12954_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05430_),
    .ZN(_05432_)
  );
  AND2_X1 _12955_ (
    .A1(_05431_),
    .A2(_05432_),
    .ZN(_05433_)
  );
  OR2_X1 _12956_ (
    .A1(_03045_),
    .A2(_05429_),
    .ZN(_05434_)
  );
  OR2_X1 _12957_ (
    .A1(_05433_),
    .A2(_05434_),
    .ZN(_05435_)
  );
  AND2_X1 _12958_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_05427_),
    .ZN(_05436_)
  );
  AND2_X1 _12959_ (
    .A1(_05435_),
    .A2(_05436_),
    .ZN(_05437_)
  );
  OR2_X1 _12960_ (
    .A1(_05419_),
    .A2(_05437_),
    .ZN(_05438_)
  );
  MUX2_X1 _12961_ (
    .A(_05407_),
    .B(_05438_),
    .S(_03063_),
    .Z(_05439_)
  );
  MUX2_X1 _12962_ (
    .A(wb_reg_wdata[20]),
    .B(csr_io_rw_rdata[20]),
    .S(_04077_),
    .Z(_05440_)
  );
  MUX2_X1 _12963_ (
    .A(div_io_resp_bits_data[20]),
    .B(_05440_),
    .S(_03114_),
    .Z(_05441_)
  );
  MUX2_X1 _12964_ (
    .A(_05441_),
    .B(io_dmem_resp_bits_data[20]),
    .S(_03097_),
    .Z(_05442_)
  );
  MUX2_X1 _12965_ (
    .A(_05439_),
    .B(_05442_),
    .S(_04074_),
    .Z(_05443_)
  );
  AND2_X1 _12966_ (
    .A1(_04044_),
    .A2(_05443_),
    .ZN(_05444_)
  );
  OR2_X1 _12967_ (
    .A1(_05370_),
    .A2(_05444_),
    .ZN(_05445_)
  );
  MUX2_X1 _12968_ (
    .A(ex_reg_rs_msb_0[18]),
    .B(_05445_),
    .S(_04042_),
    .Z(_00085_)
  );
  AND2_X1 _12969_ (
    .A1(_03065_),
    .A2(ibuf_io_inst_0_bits_raw[21]),
    .ZN(_05446_)
  );
  AND2_X1 _12970_ (
    .A1(_03582_),
    .A2(_05446_),
    .ZN(_05447_)
  );
  MUX2_X1 _12971_ (
    .A(wb_reg_wdata[21]),
    .B(csr_io_rw_rdata[21]),
    .S(_04077_),
    .Z(_05448_)
  );
  MUX2_X1 _12972_ (
    .A(div_io_resp_bits_data[21]),
    .B(_05448_),
    .S(_03114_),
    .Z(_05449_)
  );
  MUX2_X1 _12973_ (
    .A(_05449_),
    .B(io_dmem_resp_bits_data[21]),
    .S(_03097_),
    .Z(_05450_)
  );
  MUX2_X1 _12974_ (
    .A(\rf[5] [21]),
    .B(\rf[1] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05451_)
  );
  MUX2_X1 _12975_ (
    .A(\rf[7] [21]),
    .B(\rf[3] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05452_)
  );
  MUX2_X1 _12976_ (
    .A(_05451_),
    .B(_05452_),
    .S(_03045_),
    .Z(_05453_)
  );
  AND2_X1 _12977_ (
    .A1(_03044_),
    .A2(_05453_),
    .ZN(_05454_)
  );
  MUX2_X1 _12978_ (
    .A(\rf[4] [21]),
    .B(\rf[0] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05455_)
  );
  MUX2_X1 _12979_ (
    .A(\rf[6] [21]),
    .B(\rf[2] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05456_)
  );
  MUX2_X1 _12980_ (
    .A(_05455_),
    .B(_05456_),
    .S(_03045_),
    .Z(_05457_)
  );
  AND2_X1 _12981_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05457_),
    .ZN(_05458_)
  );
  OR2_X1 _12982_ (
    .A1(_03063_),
    .A2(_05458_),
    .ZN(_05459_)
  );
  OR2_X1 _12983_ (
    .A1(_05454_),
    .A2(_05459_),
    .ZN(_05460_)
  );
  OR2_X1 _12984_ (
    .A1(\rf[20] [21]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05461_)
  );
  OR2_X1 _12985_ (
    .A1(\rf[16] [21]),
    .A2(_03046_),
    .ZN(_05462_)
  );
  AND2_X1 _12986_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05462_),
    .ZN(_05463_)
  );
  AND2_X1 _12987_ (
    .A1(_05461_),
    .A2(_05463_),
    .ZN(_05464_)
  );
  MUX2_X1 _12988_ (
    .A(\rf[22] [21]),
    .B(\rf[18] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05465_)
  );
  AND2_X1 _12989_ (
    .A1(_03045_),
    .A2(_05465_),
    .ZN(_05466_)
  );
  OR2_X1 _12990_ (
    .A1(_03044_),
    .A2(_05466_),
    .ZN(_05467_)
  );
  OR2_X1 _12991_ (
    .A1(_05464_),
    .A2(_05467_),
    .ZN(_05468_)
  );
  OR2_X1 _12992_ (
    .A1(\rf[17] [21]),
    .A2(_03046_),
    .ZN(_05469_)
  );
  OR2_X1 _12993_ (
    .A1(\rf[21] [21]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05470_)
  );
  AND2_X1 _12994_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05470_),
    .ZN(_05471_)
  );
  AND2_X1 _12995_ (
    .A1(_05469_),
    .A2(_05471_),
    .ZN(_05472_)
  );
  MUX2_X1 _12996_ (
    .A(\rf[23] [21]),
    .B(\rf[19] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05473_)
  );
  AND2_X1 _12997_ (
    .A1(_03045_),
    .A2(_05473_),
    .ZN(_05474_)
  );
  OR2_X1 _12998_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05474_),
    .ZN(_05475_)
  );
  OR2_X1 _12999_ (
    .A1(_05472_),
    .A2(_05475_),
    .ZN(_05476_)
  );
  AND2_X1 _13000_ (
    .A1(_05468_),
    .A2(_05476_),
    .ZN(_05477_)
  );
  OR2_X1 _13001_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_05477_),
    .ZN(_05478_)
  );
  AND2_X1 _13002_ (
    .A1(_05460_),
    .A2(_05478_),
    .ZN(_05479_)
  );
  AND2_X1 _13003_ (
    .A1(\rf[10] [21]),
    .A2(_03045_),
    .ZN(_05480_)
  );
  AND2_X1 _13004_ (
    .A1(\rf[8] [21]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05481_)
  );
  OR2_X1 _13005_ (
    .A1(_03046_),
    .A2(_05481_),
    .ZN(_05482_)
  );
  OR2_X1 _13006_ (
    .A1(_05480_),
    .A2(_05482_),
    .ZN(_05483_)
  );
  AND2_X1 _13007_ (
    .A1(\rf[14] [21]),
    .A2(_03045_),
    .ZN(_05484_)
  );
  AND2_X1 _13008_ (
    .A1(\rf[12] [21]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05485_)
  );
  OR2_X1 _13009_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_05485_),
    .ZN(_05486_)
  );
  OR2_X1 _13010_ (
    .A1(_05484_),
    .A2(_05486_),
    .ZN(_05487_)
  );
  AND2_X1 _13011_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05487_),
    .ZN(_05488_)
  );
  AND2_X1 _13012_ (
    .A1(_05483_),
    .A2(_05488_),
    .ZN(_05489_)
  );
  AND2_X1 _13013_ (
    .A1(\rf[11] [21]),
    .A2(_03045_),
    .ZN(_05490_)
  );
  AND2_X1 _13014_ (
    .A1(\rf[9] [21]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05491_)
  );
  OR2_X1 _13015_ (
    .A1(_03046_),
    .A2(_05491_),
    .ZN(_05492_)
  );
  OR2_X1 _13016_ (
    .A1(_05490_),
    .A2(_05492_),
    .ZN(_05493_)
  );
  AND2_X1 _13017_ (
    .A1(\rf[15] [21]),
    .A2(_03045_),
    .ZN(_05494_)
  );
  AND2_X1 _13018_ (
    .A1(\rf[13] [21]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05495_)
  );
  OR2_X1 _13019_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_05495_),
    .ZN(_05496_)
  );
  OR2_X1 _13020_ (
    .A1(_05494_),
    .A2(_05496_),
    .ZN(_05497_)
  );
  AND2_X1 _13021_ (
    .A1(_03044_),
    .A2(_05497_),
    .ZN(_05498_)
  );
  AND2_X1 _13022_ (
    .A1(_05493_),
    .A2(_05498_),
    .ZN(_05499_)
  );
  OR2_X1 _13023_ (
    .A1(_03063_),
    .A2(_05499_),
    .ZN(_05500_)
  );
  OR2_X1 _13024_ (
    .A1(_05489_),
    .A2(_05500_),
    .ZN(_05501_)
  );
  OR2_X1 _13025_ (
    .A1(\rf[28] [21]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05502_)
  );
  OR2_X1 _13026_ (
    .A1(\rf[24] [21]),
    .A2(_03046_),
    .ZN(_05503_)
  );
  AND2_X1 _13027_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05502_),
    .ZN(_05504_)
  );
  AND2_X1 _13028_ (
    .A1(_05503_),
    .A2(_05504_),
    .ZN(_05505_)
  );
  MUX2_X1 _13029_ (
    .A(\rf[30] [21]),
    .B(\rf[26] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05506_)
  );
  AND2_X1 _13030_ (
    .A1(_03045_),
    .A2(_05506_),
    .ZN(_05507_)
  );
  OR2_X1 _13031_ (
    .A1(_03044_),
    .A2(_05507_),
    .ZN(_05508_)
  );
  OR2_X1 _13032_ (
    .A1(_05505_),
    .A2(_05508_),
    .ZN(_05509_)
  );
  MUX2_X1 _13033_ (
    .A(\rf[29] [21]),
    .B(\rf[25] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05510_)
  );
  AND2_X1 _13034_ (
    .A1(\rf[27] [21]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05511_)
  );
  MUX2_X1 _13035_ (
    .A(_05510_),
    .B(_05511_),
    .S(_03045_),
    .Z(_05512_)
  );
  OR2_X1 _13036_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05512_),
    .ZN(_05513_)
  );
  AND2_X1 _13037_ (
    .A1(_05509_),
    .A2(_05513_),
    .ZN(_05514_)
  );
  OR2_X1 _13038_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_05514_),
    .ZN(_05515_)
  );
  AND2_X1 _13039_ (
    .A1(_05501_),
    .A2(_05515_),
    .ZN(_05516_)
  );
  MUX2_X1 _13040_ (
    .A(_05479_),
    .B(_05516_),
    .S(_03047_),
    .Z(_05517_)
  );
  MUX2_X1 _13041_ (
    .A(_05517_),
    .B(_05450_),
    .S(_04074_),
    .Z(_05518_)
  );
  AND2_X1 _13042_ (
    .A1(_04044_),
    .A2(_05518_),
    .ZN(_05519_)
  );
  OR2_X1 _13043_ (
    .A1(_05447_),
    .A2(_05519_),
    .ZN(_05520_)
  );
  MUX2_X1 _13044_ (
    .A(ex_reg_rs_msb_0[19]),
    .B(_05520_),
    .S(_04042_),
    .Z(_00086_)
  );
  AND2_X1 _13045_ (
    .A1(_03065_),
    .A2(ibuf_io_inst_0_bits_raw[22]),
    .ZN(_05521_)
  );
  AND2_X1 _13046_ (
    .A1(_03582_),
    .A2(_05521_),
    .ZN(_05522_)
  );
  MUX2_X1 _13047_ (
    .A(\rf[5] [22]),
    .B(\rf[1] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05523_)
  );
  MUX2_X1 _13048_ (
    .A(\rf[7] [22]),
    .B(\rf[3] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05524_)
  );
  MUX2_X1 _13049_ (
    .A(_05523_),
    .B(_05524_),
    .S(_03045_),
    .Z(_05525_)
  );
  AND2_X1 _13050_ (
    .A1(_03044_),
    .A2(_05525_),
    .ZN(_05526_)
  );
  MUX2_X1 _13051_ (
    .A(\rf[4] [22]),
    .B(\rf[0] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05527_)
  );
  MUX2_X1 _13052_ (
    .A(\rf[6] [22]),
    .B(\rf[2] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05528_)
  );
  MUX2_X1 _13053_ (
    .A(_05527_),
    .B(_05528_),
    .S(_03045_),
    .Z(_05529_)
  );
  AND2_X1 _13054_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05529_),
    .ZN(_05530_)
  );
  OR2_X1 _13055_ (
    .A1(_03063_),
    .A2(_05530_),
    .ZN(_05531_)
  );
  OR2_X1 _13056_ (
    .A1(_05526_),
    .A2(_05531_),
    .ZN(_05532_)
  );
  OR2_X1 _13057_ (
    .A1(\rf[20] [22]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05533_)
  );
  OR2_X1 _13058_ (
    .A1(\rf[16] [22]),
    .A2(_03046_),
    .ZN(_05534_)
  );
  AND2_X1 _13059_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05534_),
    .ZN(_05535_)
  );
  AND2_X1 _13060_ (
    .A1(_05533_),
    .A2(_05535_),
    .ZN(_05536_)
  );
  MUX2_X1 _13061_ (
    .A(\rf[22] [22]),
    .B(\rf[18] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05537_)
  );
  AND2_X1 _13062_ (
    .A1(_03045_),
    .A2(_05537_),
    .ZN(_05538_)
  );
  OR2_X1 _13063_ (
    .A1(_03044_),
    .A2(_05538_),
    .ZN(_05539_)
  );
  OR2_X1 _13064_ (
    .A1(_05536_),
    .A2(_05539_),
    .ZN(_05540_)
  );
  OR2_X1 _13065_ (
    .A1(\rf[17] [22]),
    .A2(_03046_),
    .ZN(_05541_)
  );
  OR2_X1 _13066_ (
    .A1(\rf[21] [22]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05542_)
  );
  AND2_X1 _13067_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05542_),
    .ZN(_05543_)
  );
  AND2_X1 _13068_ (
    .A1(_05541_),
    .A2(_05543_),
    .ZN(_05544_)
  );
  MUX2_X1 _13069_ (
    .A(\rf[23] [22]),
    .B(\rf[19] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05545_)
  );
  AND2_X1 _13070_ (
    .A1(_03045_),
    .A2(_05545_),
    .ZN(_05546_)
  );
  OR2_X1 _13071_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05546_),
    .ZN(_05547_)
  );
  OR2_X1 _13072_ (
    .A1(_05544_),
    .A2(_05547_),
    .ZN(_05548_)
  );
  AND2_X1 _13073_ (
    .A1(_05540_),
    .A2(_05548_),
    .ZN(_05549_)
  );
  OR2_X1 _13074_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_05549_),
    .ZN(_05550_)
  );
  AND2_X1 _13075_ (
    .A1(_05532_),
    .A2(_05550_),
    .ZN(_05551_)
  );
  AND2_X1 _13076_ (
    .A1(\rf[10] [22]),
    .A2(_03045_),
    .ZN(_05552_)
  );
  AND2_X1 _13077_ (
    .A1(\rf[8] [22]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05553_)
  );
  OR2_X1 _13078_ (
    .A1(_03046_),
    .A2(_05553_),
    .ZN(_05554_)
  );
  OR2_X1 _13079_ (
    .A1(_05552_),
    .A2(_05554_),
    .ZN(_05555_)
  );
  AND2_X1 _13080_ (
    .A1(\rf[14] [22]),
    .A2(_03045_),
    .ZN(_05556_)
  );
  AND2_X1 _13081_ (
    .A1(\rf[12] [22]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05557_)
  );
  OR2_X1 _13082_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_05557_),
    .ZN(_05558_)
  );
  OR2_X1 _13083_ (
    .A1(_05556_),
    .A2(_05558_),
    .ZN(_05559_)
  );
  AND2_X1 _13084_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05559_),
    .ZN(_05560_)
  );
  AND2_X1 _13085_ (
    .A1(_05555_),
    .A2(_05560_),
    .ZN(_05561_)
  );
  AND2_X1 _13086_ (
    .A1(\rf[11] [22]),
    .A2(_03045_),
    .ZN(_05562_)
  );
  AND2_X1 _13087_ (
    .A1(\rf[9] [22]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05563_)
  );
  OR2_X1 _13088_ (
    .A1(_03046_),
    .A2(_05563_),
    .ZN(_05564_)
  );
  OR2_X1 _13089_ (
    .A1(_05562_),
    .A2(_05564_),
    .ZN(_05565_)
  );
  AND2_X1 _13090_ (
    .A1(\rf[15] [22]),
    .A2(_03045_),
    .ZN(_05566_)
  );
  AND2_X1 _13091_ (
    .A1(\rf[13] [22]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05567_)
  );
  OR2_X1 _13092_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_05567_),
    .ZN(_05568_)
  );
  OR2_X1 _13093_ (
    .A1(_05566_),
    .A2(_05568_),
    .ZN(_05569_)
  );
  AND2_X1 _13094_ (
    .A1(_03044_),
    .A2(_05569_),
    .ZN(_05570_)
  );
  AND2_X1 _13095_ (
    .A1(_05565_),
    .A2(_05570_),
    .ZN(_05571_)
  );
  OR2_X1 _13096_ (
    .A1(_03063_),
    .A2(_05571_),
    .ZN(_05572_)
  );
  OR2_X1 _13097_ (
    .A1(_05561_),
    .A2(_05572_),
    .ZN(_05573_)
  );
  OR2_X1 _13098_ (
    .A1(\rf[28] [22]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05574_)
  );
  OR2_X1 _13099_ (
    .A1(\rf[24] [22]),
    .A2(_03046_),
    .ZN(_05575_)
  );
  AND2_X1 _13100_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05574_),
    .ZN(_05576_)
  );
  AND2_X1 _13101_ (
    .A1(_05575_),
    .A2(_05576_),
    .ZN(_05577_)
  );
  MUX2_X1 _13102_ (
    .A(\rf[30] [22]),
    .B(\rf[26] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05578_)
  );
  AND2_X1 _13103_ (
    .A1(_03045_),
    .A2(_05578_),
    .ZN(_05579_)
  );
  OR2_X1 _13104_ (
    .A1(_03044_),
    .A2(_05579_),
    .ZN(_05580_)
  );
  OR2_X1 _13105_ (
    .A1(_05577_),
    .A2(_05580_),
    .ZN(_05581_)
  );
  MUX2_X1 _13106_ (
    .A(\rf[29] [22]),
    .B(\rf[25] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05582_)
  );
  AND2_X1 _13107_ (
    .A1(\rf[27] [22]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05583_)
  );
  MUX2_X1 _13108_ (
    .A(_05582_),
    .B(_05583_),
    .S(_03045_),
    .Z(_05584_)
  );
  OR2_X1 _13109_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05584_),
    .ZN(_05585_)
  );
  AND2_X1 _13110_ (
    .A1(_05581_),
    .A2(_05585_),
    .ZN(_05586_)
  );
  OR2_X1 _13111_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_05586_),
    .ZN(_05587_)
  );
  AND2_X1 _13112_ (
    .A1(_05573_),
    .A2(_05587_),
    .ZN(_05588_)
  );
  MUX2_X1 _13113_ (
    .A(_05551_),
    .B(_05588_),
    .S(_03047_),
    .Z(_05589_)
  );
  MUX2_X1 _13114_ (
    .A(wb_reg_wdata[22]),
    .B(csr_io_rw_rdata[22]),
    .S(_04077_),
    .Z(_05590_)
  );
  MUX2_X1 _13115_ (
    .A(div_io_resp_bits_data[22]),
    .B(_05590_),
    .S(_03114_),
    .Z(_05591_)
  );
  MUX2_X1 _13116_ (
    .A(_05591_),
    .B(io_dmem_resp_bits_data[22]),
    .S(_03097_),
    .Z(_05592_)
  );
  MUX2_X1 _13117_ (
    .A(_05589_),
    .B(_05592_),
    .S(_04074_),
    .Z(_05593_)
  );
  AND2_X1 _13118_ (
    .A1(_04044_),
    .A2(_05593_),
    .ZN(_05594_)
  );
  OR2_X1 _13119_ (
    .A1(_05522_),
    .A2(_05594_),
    .ZN(_05595_)
  );
  MUX2_X1 _13120_ (
    .A(ex_reg_rs_msb_0[20]),
    .B(_05595_),
    .S(_04042_),
    .Z(_00087_)
  );
  AND2_X1 _13121_ (
    .A1(_03065_),
    .A2(ibuf_io_inst_0_bits_raw[23]),
    .ZN(_05596_)
  );
  AND2_X1 _13122_ (
    .A1(_03582_),
    .A2(_05596_),
    .ZN(_05597_)
  );
  MUX2_X1 _13123_ (
    .A(\rf[3] [23]),
    .B(\rf[2] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_05598_)
  );
  MUX2_X1 _13124_ (
    .A(\rf[7] [23]),
    .B(\rf[6] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_05599_)
  );
  MUX2_X1 _13125_ (
    .A(_05598_),
    .B(_05599_),
    .S(_03046_),
    .Z(_05600_)
  );
  OR2_X1 _13126_ (
    .A1(_03047_),
    .A2(_05600_),
    .ZN(_05601_)
  );
  MUX2_X1 _13127_ (
    .A(\rf[15] [23]),
    .B(\rf[11] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05602_)
  );
  OR2_X1 _13128_ (
    .A1(_03448_),
    .A2(_05602_),
    .ZN(_05603_)
  );
  MUX2_X1 _13129_ (
    .A(\rf[14] [23]),
    .B(\rf[10] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05604_)
  );
  OR2_X1 _13130_ (
    .A1(_04124_),
    .A2(_05604_),
    .ZN(_05605_)
  );
  AND2_X1 _13131_ (
    .A1(_05603_),
    .A2(_05605_),
    .ZN(_05606_)
  );
  AND2_X1 _13132_ (
    .A1(_05601_),
    .A2(_05606_),
    .ZN(_05607_)
  );
  AND2_X1 _13133_ (
    .A1(_03045_),
    .A2(_05607_),
    .ZN(_05608_)
  );
  MUX2_X1 _13134_ (
    .A(\rf[1] [23]),
    .B(\rf[0] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_05609_)
  );
  MUX2_X1 _13135_ (
    .A(\rf[5] [23]),
    .B(\rf[4] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs1[0]),
    .Z(_05610_)
  );
  MUX2_X1 _13136_ (
    .A(_05609_),
    .B(_05610_),
    .S(_03046_),
    .Z(_05611_)
  );
  OR2_X1 _13137_ (
    .A1(_03047_),
    .A2(_05611_),
    .ZN(_05612_)
  );
  MUX2_X1 _13138_ (
    .A(\rf[13] [23]),
    .B(\rf[9] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05613_)
  );
  OR2_X1 _13139_ (
    .A1(_03448_),
    .A2(_05613_),
    .ZN(_05614_)
  );
  MUX2_X1 _13140_ (
    .A(\rf[12] [23]),
    .B(\rf[8] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05615_)
  );
  OR2_X1 _13141_ (
    .A1(_04124_),
    .A2(_05615_),
    .ZN(_05616_)
  );
  AND2_X1 _13142_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05614_),
    .ZN(_05617_)
  );
  AND2_X1 _13143_ (
    .A1(_05616_),
    .A2(_05617_),
    .ZN(_05618_)
  );
  AND2_X1 _13144_ (
    .A1(_05612_),
    .A2(_05618_),
    .ZN(_05619_)
  );
  OR2_X1 _13145_ (
    .A1(_03063_),
    .A2(_05619_),
    .ZN(_05620_)
  );
  OR2_X1 _13146_ (
    .A1(_05608_),
    .A2(_05620_),
    .ZN(_05621_)
  );
  OR2_X1 _13147_ (
    .A1(\rf[28] [23]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05622_)
  );
  OR2_X1 _13148_ (
    .A1(\rf[24] [23]),
    .A2(_03046_),
    .ZN(_05623_)
  );
  AND2_X1 _13149_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05622_),
    .ZN(_05624_)
  );
  AND2_X1 _13150_ (
    .A1(_05623_),
    .A2(_05624_),
    .ZN(_05625_)
  );
  MUX2_X1 _13151_ (
    .A(\rf[30] [23]),
    .B(\rf[26] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05626_)
  );
  AND2_X1 _13152_ (
    .A1(_03045_),
    .A2(_05626_),
    .ZN(_05627_)
  );
  OR2_X1 _13153_ (
    .A1(_03044_),
    .A2(_05627_),
    .ZN(_05628_)
  );
  OR2_X1 _13154_ (
    .A1(_05625_),
    .A2(_05628_),
    .ZN(_05629_)
  );
  MUX2_X1 _13155_ (
    .A(\rf[29] [23]),
    .B(\rf[25] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05630_)
  );
  AND2_X1 _13156_ (
    .A1(\rf[27] [23]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05631_)
  );
  MUX2_X1 _13157_ (
    .A(_05630_),
    .B(_05631_),
    .S(_03045_),
    .Z(_05632_)
  );
  OR2_X1 _13158_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05632_),
    .ZN(_05633_)
  );
  AND2_X1 _13159_ (
    .A1(_05629_),
    .A2(_05633_),
    .ZN(_05634_)
  );
  OR2_X1 _13160_ (
    .A1(\rf[20] [23]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05635_)
  );
  OR2_X1 _13161_ (
    .A1(\rf[16] [23]),
    .A2(_03046_),
    .ZN(_05636_)
  );
  AND2_X1 _13162_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05636_),
    .ZN(_05637_)
  );
  AND2_X1 _13163_ (
    .A1(_05635_),
    .A2(_05637_),
    .ZN(_05638_)
  );
  MUX2_X1 _13164_ (
    .A(\rf[22] [23]),
    .B(\rf[18] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05639_)
  );
  AND2_X1 _13165_ (
    .A1(_03045_),
    .A2(_05639_),
    .ZN(_05640_)
  );
  OR2_X1 _13166_ (
    .A1(_03044_),
    .A2(_05640_),
    .ZN(_05641_)
  );
  OR2_X1 _13167_ (
    .A1(_05638_),
    .A2(_05641_),
    .ZN(_05642_)
  );
  OR2_X1 _13168_ (
    .A1(\rf[17] [23]),
    .A2(_03046_),
    .ZN(_05643_)
  );
  OR2_X1 _13169_ (
    .A1(\rf[21] [23]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05644_)
  );
  AND2_X1 _13170_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05644_),
    .ZN(_05645_)
  );
  AND2_X1 _13171_ (
    .A1(_05643_),
    .A2(_05645_),
    .ZN(_05646_)
  );
  MUX2_X1 _13172_ (
    .A(\rf[23] [23]),
    .B(\rf[19] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05647_)
  );
  AND2_X1 _13173_ (
    .A1(_03045_),
    .A2(_05647_),
    .ZN(_05648_)
  );
  OR2_X1 _13174_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05648_),
    .ZN(_05649_)
  );
  OR2_X1 _13175_ (
    .A1(_05646_),
    .A2(_05649_),
    .ZN(_05650_)
  );
  AND2_X1 _13176_ (
    .A1(_05642_),
    .A2(_05650_),
    .ZN(_05651_)
  );
  MUX2_X1 _13177_ (
    .A(_05634_),
    .B(_05651_),
    .S(ibuf_io_inst_0_bits_inst_rs1[3]),
    .Z(_05652_)
  );
  OR2_X1 _13178_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_05652_),
    .ZN(_05653_)
  );
  AND2_X1 _13179_ (
    .A1(_05621_),
    .A2(_05653_),
    .ZN(_05654_)
  );
  MUX2_X1 _13180_ (
    .A(wb_reg_wdata[23]),
    .B(csr_io_rw_rdata[23]),
    .S(_04077_),
    .Z(_05655_)
  );
  MUX2_X1 _13181_ (
    .A(div_io_resp_bits_data[23]),
    .B(_05655_),
    .S(_03114_),
    .Z(_05656_)
  );
  MUX2_X1 _13182_ (
    .A(_05656_),
    .B(io_dmem_resp_bits_data[23]),
    .S(_03097_),
    .Z(_05657_)
  );
  MUX2_X1 _13183_ (
    .A(_05654_),
    .B(_05657_),
    .S(_04074_),
    .Z(_05658_)
  );
  AND2_X1 _13184_ (
    .A1(_04044_),
    .A2(_05658_),
    .ZN(_05659_)
  );
  OR2_X1 _13185_ (
    .A1(_05597_),
    .A2(_05659_),
    .ZN(_05660_)
  );
  MUX2_X1 _13186_ (
    .A(ex_reg_rs_msb_0[21]),
    .B(_05660_),
    .S(_04042_),
    .Z(_00088_)
  );
  AND2_X1 _13187_ (
    .A1(_03065_),
    .A2(ibuf_io_inst_0_bits_raw[24]),
    .ZN(_05661_)
  );
  AND2_X1 _13188_ (
    .A1(_03582_),
    .A2(_05661_),
    .ZN(_05662_)
  );
  MUX2_X1 _13189_ (
    .A(wb_reg_wdata[24]),
    .B(csr_io_rw_rdata[24]),
    .S(_04077_),
    .Z(_05663_)
  );
  MUX2_X1 _13190_ (
    .A(div_io_resp_bits_data[24]),
    .B(_05663_),
    .S(_03114_),
    .Z(_05664_)
  );
  MUX2_X1 _13191_ (
    .A(_05664_),
    .B(io_dmem_resp_bits_data[24]),
    .S(_03097_),
    .Z(_05665_)
  );
  MUX2_X1 _13192_ (
    .A(\rf[5] [24]),
    .B(\rf[1] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05666_)
  );
  MUX2_X1 _13193_ (
    .A(\rf[7] [24]),
    .B(\rf[3] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05667_)
  );
  MUX2_X1 _13194_ (
    .A(_05666_),
    .B(_05667_),
    .S(_03045_),
    .Z(_05668_)
  );
  AND2_X1 _13195_ (
    .A1(_03044_),
    .A2(_05668_),
    .ZN(_05669_)
  );
  MUX2_X1 _13196_ (
    .A(\rf[4] [24]),
    .B(\rf[0] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05670_)
  );
  MUX2_X1 _13197_ (
    .A(\rf[6] [24]),
    .B(\rf[2] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05671_)
  );
  MUX2_X1 _13198_ (
    .A(_05670_),
    .B(_05671_),
    .S(_03045_),
    .Z(_05672_)
  );
  AND2_X1 _13199_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05672_),
    .ZN(_05673_)
  );
  OR2_X1 _13200_ (
    .A1(_03063_),
    .A2(_05673_),
    .ZN(_05674_)
  );
  OR2_X1 _13201_ (
    .A1(_05669_),
    .A2(_05674_),
    .ZN(_05675_)
  );
  OR2_X1 _13202_ (
    .A1(\rf[20] [24]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05676_)
  );
  OR2_X1 _13203_ (
    .A1(\rf[16] [24]),
    .A2(_03046_),
    .ZN(_05677_)
  );
  AND2_X1 _13204_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05677_),
    .ZN(_05678_)
  );
  AND2_X1 _13205_ (
    .A1(_05676_),
    .A2(_05678_),
    .ZN(_05679_)
  );
  MUX2_X1 _13206_ (
    .A(\rf[22] [24]),
    .B(\rf[18] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05680_)
  );
  AND2_X1 _13207_ (
    .A1(_03045_),
    .A2(_05680_),
    .ZN(_05681_)
  );
  OR2_X1 _13208_ (
    .A1(_03044_),
    .A2(_05681_),
    .ZN(_05682_)
  );
  OR2_X1 _13209_ (
    .A1(_05679_),
    .A2(_05682_),
    .ZN(_05683_)
  );
  OR2_X1 _13210_ (
    .A1(\rf[17] [24]),
    .A2(_03046_),
    .ZN(_05684_)
  );
  OR2_X1 _13211_ (
    .A1(\rf[21] [24]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05685_)
  );
  AND2_X1 _13212_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05685_),
    .ZN(_05686_)
  );
  AND2_X1 _13213_ (
    .A1(_05684_),
    .A2(_05686_),
    .ZN(_05687_)
  );
  MUX2_X1 _13214_ (
    .A(\rf[23] [24]),
    .B(\rf[19] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05688_)
  );
  AND2_X1 _13215_ (
    .A1(_03045_),
    .A2(_05688_),
    .ZN(_05689_)
  );
  OR2_X1 _13216_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05689_),
    .ZN(_05690_)
  );
  OR2_X1 _13217_ (
    .A1(_05687_),
    .A2(_05690_),
    .ZN(_05691_)
  );
  AND2_X1 _13218_ (
    .A1(_05683_),
    .A2(_05691_),
    .ZN(_05692_)
  );
  OR2_X1 _13219_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_05692_),
    .ZN(_05693_)
  );
  AND2_X1 _13220_ (
    .A1(_05675_),
    .A2(_05693_),
    .ZN(_05694_)
  );
  AND2_X1 _13221_ (
    .A1(\rf[10] [24]),
    .A2(_03045_),
    .ZN(_05695_)
  );
  AND2_X1 _13222_ (
    .A1(\rf[8] [24]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05696_)
  );
  OR2_X1 _13223_ (
    .A1(_03046_),
    .A2(_05696_),
    .ZN(_05697_)
  );
  OR2_X1 _13224_ (
    .A1(_05695_),
    .A2(_05697_),
    .ZN(_05698_)
  );
  AND2_X1 _13225_ (
    .A1(\rf[14] [24]),
    .A2(_03045_),
    .ZN(_05699_)
  );
  AND2_X1 _13226_ (
    .A1(\rf[12] [24]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05700_)
  );
  OR2_X1 _13227_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_05700_),
    .ZN(_05701_)
  );
  OR2_X1 _13228_ (
    .A1(_05699_),
    .A2(_05701_),
    .ZN(_05702_)
  );
  AND2_X1 _13229_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05702_),
    .ZN(_05703_)
  );
  AND2_X1 _13230_ (
    .A1(_05698_),
    .A2(_05703_),
    .ZN(_05704_)
  );
  AND2_X1 _13231_ (
    .A1(\rf[11] [24]),
    .A2(_03045_),
    .ZN(_05705_)
  );
  AND2_X1 _13232_ (
    .A1(\rf[9] [24]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05706_)
  );
  OR2_X1 _13233_ (
    .A1(_03046_),
    .A2(_05706_),
    .ZN(_05707_)
  );
  OR2_X1 _13234_ (
    .A1(_05705_),
    .A2(_05707_),
    .ZN(_05708_)
  );
  AND2_X1 _13235_ (
    .A1(\rf[15] [24]),
    .A2(_03045_),
    .ZN(_05709_)
  );
  AND2_X1 _13236_ (
    .A1(\rf[13] [24]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05710_)
  );
  OR2_X1 _13237_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_05710_),
    .ZN(_05711_)
  );
  OR2_X1 _13238_ (
    .A1(_05709_),
    .A2(_05711_),
    .ZN(_05712_)
  );
  AND2_X1 _13239_ (
    .A1(_03044_),
    .A2(_05712_),
    .ZN(_05713_)
  );
  AND2_X1 _13240_ (
    .A1(_05708_),
    .A2(_05713_),
    .ZN(_05714_)
  );
  OR2_X1 _13241_ (
    .A1(_03063_),
    .A2(_05714_),
    .ZN(_05715_)
  );
  OR2_X1 _13242_ (
    .A1(_05704_),
    .A2(_05715_),
    .ZN(_05716_)
  );
  OR2_X1 _13243_ (
    .A1(\rf[28] [24]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05717_)
  );
  OR2_X1 _13244_ (
    .A1(\rf[24] [24]),
    .A2(_03046_),
    .ZN(_05718_)
  );
  AND2_X1 _13245_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05717_),
    .ZN(_05719_)
  );
  AND2_X1 _13246_ (
    .A1(_05718_),
    .A2(_05719_),
    .ZN(_05720_)
  );
  MUX2_X1 _13247_ (
    .A(\rf[30] [24]),
    .B(\rf[26] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05721_)
  );
  AND2_X1 _13248_ (
    .A1(_03045_),
    .A2(_05721_),
    .ZN(_05722_)
  );
  OR2_X1 _13249_ (
    .A1(_03044_),
    .A2(_05722_),
    .ZN(_05723_)
  );
  OR2_X1 _13250_ (
    .A1(_05720_),
    .A2(_05723_),
    .ZN(_05724_)
  );
  MUX2_X1 _13251_ (
    .A(\rf[29] [24]),
    .B(\rf[25] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05725_)
  );
  AND2_X1 _13252_ (
    .A1(\rf[27] [24]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05726_)
  );
  MUX2_X1 _13253_ (
    .A(_05725_),
    .B(_05726_),
    .S(_03045_),
    .Z(_05727_)
  );
  OR2_X1 _13254_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05727_),
    .ZN(_05728_)
  );
  AND2_X1 _13255_ (
    .A1(_05724_),
    .A2(_05728_),
    .ZN(_05729_)
  );
  OR2_X1 _13256_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_05729_),
    .ZN(_05730_)
  );
  AND2_X1 _13257_ (
    .A1(_05716_),
    .A2(_05730_),
    .ZN(_05731_)
  );
  MUX2_X1 _13258_ (
    .A(_05694_),
    .B(_05731_),
    .S(_03047_),
    .Z(_05732_)
  );
  MUX2_X1 _13259_ (
    .A(_05732_),
    .B(_05665_),
    .S(_04074_),
    .Z(_05733_)
  );
  AND2_X1 _13260_ (
    .A1(_04044_),
    .A2(_05733_),
    .ZN(_05734_)
  );
  OR2_X1 _13261_ (
    .A1(_05662_),
    .A2(_05734_),
    .ZN(_05735_)
  );
  MUX2_X1 _13262_ (
    .A(ex_reg_rs_msb_0[22]),
    .B(_05735_),
    .S(_04042_),
    .Z(_00089_)
  );
  AND2_X1 _13263_ (
    .A1(_03065_),
    .A2(ibuf_io_inst_0_bits_raw[25]),
    .ZN(_05736_)
  );
  AND2_X1 _13264_ (
    .A1(_03582_),
    .A2(_05736_),
    .ZN(_05737_)
  );
  MUX2_X1 _13265_ (
    .A(wb_reg_wdata[25]),
    .B(csr_io_rw_rdata[25]),
    .S(_04077_),
    .Z(_05738_)
  );
  MUX2_X1 _13266_ (
    .A(div_io_resp_bits_data[25]),
    .B(_05738_),
    .S(_03114_),
    .Z(_05739_)
  );
  MUX2_X1 _13267_ (
    .A(_05739_),
    .B(io_dmem_resp_bits_data[25]),
    .S(_03097_),
    .Z(_05740_)
  );
  MUX2_X1 _13268_ (
    .A(\rf[5] [25]),
    .B(\rf[1] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05741_)
  );
  MUX2_X1 _13269_ (
    .A(\rf[7] [25]),
    .B(\rf[3] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05742_)
  );
  MUX2_X1 _13270_ (
    .A(_05741_),
    .B(_05742_),
    .S(_03045_),
    .Z(_05743_)
  );
  AND2_X1 _13271_ (
    .A1(_03044_),
    .A2(_05743_),
    .ZN(_05744_)
  );
  MUX2_X1 _13272_ (
    .A(\rf[4] [25]),
    .B(\rf[0] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05745_)
  );
  MUX2_X1 _13273_ (
    .A(\rf[6] [25]),
    .B(\rf[2] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05746_)
  );
  MUX2_X1 _13274_ (
    .A(_05745_),
    .B(_05746_),
    .S(_03045_),
    .Z(_05747_)
  );
  AND2_X1 _13275_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05747_),
    .ZN(_05748_)
  );
  OR2_X1 _13276_ (
    .A1(_03063_),
    .A2(_05748_),
    .ZN(_05749_)
  );
  OR2_X1 _13277_ (
    .A1(_05744_),
    .A2(_05749_),
    .ZN(_05750_)
  );
  OR2_X1 _13278_ (
    .A1(\rf[20] [25]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05751_)
  );
  OR2_X1 _13279_ (
    .A1(\rf[16] [25]),
    .A2(_03046_),
    .ZN(_05752_)
  );
  AND2_X1 _13280_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05752_),
    .ZN(_05753_)
  );
  AND2_X1 _13281_ (
    .A1(_05751_),
    .A2(_05753_),
    .ZN(_05754_)
  );
  MUX2_X1 _13282_ (
    .A(\rf[22] [25]),
    .B(\rf[18] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05755_)
  );
  AND2_X1 _13283_ (
    .A1(_03045_),
    .A2(_05755_),
    .ZN(_05756_)
  );
  OR2_X1 _13284_ (
    .A1(_03044_),
    .A2(_05756_),
    .ZN(_05757_)
  );
  OR2_X1 _13285_ (
    .A1(_05754_),
    .A2(_05757_),
    .ZN(_05758_)
  );
  OR2_X1 _13286_ (
    .A1(\rf[17] [25]),
    .A2(_03046_),
    .ZN(_05759_)
  );
  OR2_X1 _13287_ (
    .A1(\rf[21] [25]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05760_)
  );
  AND2_X1 _13288_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05760_),
    .ZN(_05761_)
  );
  AND2_X1 _13289_ (
    .A1(_05759_),
    .A2(_05761_),
    .ZN(_05762_)
  );
  MUX2_X1 _13290_ (
    .A(\rf[23] [25]),
    .B(\rf[19] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05763_)
  );
  AND2_X1 _13291_ (
    .A1(_03045_),
    .A2(_05763_),
    .ZN(_05764_)
  );
  OR2_X1 _13292_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05764_),
    .ZN(_05765_)
  );
  OR2_X1 _13293_ (
    .A1(_05762_),
    .A2(_05765_),
    .ZN(_05766_)
  );
  AND2_X1 _13294_ (
    .A1(_05758_),
    .A2(_05766_),
    .ZN(_05767_)
  );
  OR2_X1 _13295_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_05767_),
    .ZN(_05768_)
  );
  AND2_X1 _13296_ (
    .A1(_05750_),
    .A2(_05768_),
    .ZN(_05769_)
  );
  AND2_X1 _13297_ (
    .A1(\rf[10] [25]),
    .A2(_03045_),
    .ZN(_05770_)
  );
  AND2_X1 _13298_ (
    .A1(\rf[8] [25]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05771_)
  );
  OR2_X1 _13299_ (
    .A1(_03046_),
    .A2(_05771_),
    .ZN(_05772_)
  );
  OR2_X1 _13300_ (
    .A1(_05770_),
    .A2(_05772_),
    .ZN(_05773_)
  );
  AND2_X1 _13301_ (
    .A1(\rf[14] [25]),
    .A2(_03045_),
    .ZN(_05774_)
  );
  AND2_X1 _13302_ (
    .A1(\rf[12] [25]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05775_)
  );
  OR2_X1 _13303_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_05775_),
    .ZN(_05776_)
  );
  OR2_X1 _13304_ (
    .A1(_05774_),
    .A2(_05776_),
    .ZN(_05777_)
  );
  AND2_X1 _13305_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05777_),
    .ZN(_05778_)
  );
  AND2_X1 _13306_ (
    .A1(_05773_),
    .A2(_05778_),
    .ZN(_05779_)
  );
  AND2_X1 _13307_ (
    .A1(\rf[11] [25]),
    .A2(_03045_),
    .ZN(_05780_)
  );
  AND2_X1 _13308_ (
    .A1(\rf[9] [25]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05781_)
  );
  OR2_X1 _13309_ (
    .A1(_03046_),
    .A2(_05781_),
    .ZN(_05782_)
  );
  OR2_X1 _13310_ (
    .A1(_05780_),
    .A2(_05782_),
    .ZN(_05783_)
  );
  AND2_X1 _13311_ (
    .A1(\rf[15] [25]),
    .A2(_03045_),
    .ZN(_05784_)
  );
  AND2_X1 _13312_ (
    .A1(\rf[13] [25]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05785_)
  );
  OR2_X1 _13313_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_05785_),
    .ZN(_05786_)
  );
  OR2_X1 _13314_ (
    .A1(_05784_),
    .A2(_05786_),
    .ZN(_05787_)
  );
  AND2_X1 _13315_ (
    .A1(_03044_),
    .A2(_05787_),
    .ZN(_05788_)
  );
  AND2_X1 _13316_ (
    .A1(_05783_),
    .A2(_05788_),
    .ZN(_05789_)
  );
  OR2_X1 _13317_ (
    .A1(_03063_),
    .A2(_05789_),
    .ZN(_05790_)
  );
  OR2_X1 _13318_ (
    .A1(_05779_),
    .A2(_05790_),
    .ZN(_05791_)
  );
  OR2_X1 _13319_ (
    .A1(\rf[28] [25]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05792_)
  );
  OR2_X1 _13320_ (
    .A1(\rf[24] [25]),
    .A2(_03046_),
    .ZN(_05793_)
  );
  AND2_X1 _13321_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05792_),
    .ZN(_05794_)
  );
  AND2_X1 _13322_ (
    .A1(_05793_),
    .A2(_05794_),
    .ZN(_05795_)
  );
  MUX2_X1 _13323_ (
    .A(\rf[30] [25]),
    .B(\rf[26] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05796_)
  );
  AND2_X1 _13324_ (
    .A1(_03045_),
    .A2(_05796_),
    .ZN(_05797_)
  );
  OR2_X1 _13325_ (
    .A1(_03044_),
    .A2(_05797_),
    .ZN(_05798_)
  );
  OR2_X1 _13326_ (
    .A1(_05795_),
    .A2(_05798_),
    .ZN(_05799_)
  );
  MUX2_X1 _13327_ (
    .A(\rf[29] [25]),
    .B(\rf[25] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05800_)
  );
  AND2_X1 _13328_ (
    .A1(\rf[27] [25]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05801_)
  );
  MUX2_X1 _13329_ (
    .A(_05800_),
    .B(_05801_),
    .S(_03045_),
    .Z(_05802_)
  );
  OR2_X1 _13330_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05802_),
    .ZN(_05803_)
  );
  AND2_X1 _13331_ (
    .A1(_05799_),
    .A2(_05803_),
    .ZN(_05804_)
  );
  OR2_X1 _13332_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_05804_),
    .ZN(_05805_)
  );
  AND2_X1 _13333_ (
    .A1(_05791_),
    .A2(_05805_),
    .ZN(_05806_)
  );
  MUX2_X1 _13334_ (
    .A(_05769_),
    .B(_05806_),
    .S(_03047_),
    .Z(_05807_)
  );
  MUX2_X1 _13335_ (
    .A(_05807_),
    .B(_05740_),
    .S(_04074_),
    .Z(_05808_)
  );
  AND2_X1 _13336_ (
    .A1(_04044_),
    .A2(_05808_),
    .ZN(_05809_)
  );
  OR2_X1 _13337_ (
    .A1(_05737_),
    .A2(_05809_),
    .ZN(_05810_)
  );
  MUX2_X1 _13338_ (
    .A(ex_reg_rs_msb_0[23]),
    .B(_05810_),
    .S(_04042_),
    .Z(_00090_)
  );
  AND2_X1 _13339_ (
    .A1(_03065_),
    .A2(ibuf_io_inst_0_bits_raw[26]),
    .ZN(_05811_)
  );
  AND2_X1 _13340_ (
    .A1(_03582_),
    .A2(_05811_),
    .ZN(_05812_)
  );
  MUX2_X1 _13341_ (
    .A(\rf[5] [26]),
    .B(\rf[1] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05813_)
  );
  MUX2_X1 _13342_ (
    .A(\rf[7] [26]),
    .B(\rf[3] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05814_)
  );
  MUX2_X1 _13343_ (
    .A(_05813_),
    .B(_05814_),
    .S(_03045_),
    .Z(_05815_)
  );
  AND2_X1 _13344_ (
    .A1(_03044_),
    .A2(_05815_),
    .ZN(_05816_)
  );
  MUX2_X1 _13345_ (
    .A(\rf[4] [26]),
    .B(\rf[0] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05817_)
  );
  MUX2_X1 _13346_ (
    .A(\rf[6] [26]),
    .B(\rf[2] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05818_)
  );
  MUX2_X1 _13347_ (
    .A(_05817_),
    .B(_05818_),
    .S(_03045_),
    .Z(_05819_)
  );
  AND2_X1 _13348_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05819_),
    .ZN(_05820_)
  );
  OR2_X1 _13349_ (
    .A1(_03063_),
    .A2(_05820_),
    .ZN(_05821_)
  );
  OR2_X1 _13350_ (
    .A1(_05816_),
    .A2(_05821_),
    .ZN(_05822_)
  );
  OR2_X1 _13351_ (
    .A1(\rf[20] [26]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05823_)
  );
  OR2_X1 _13352_ (
    .A1(\rf[16] [26]),
    .A2(_03046_),
    .ZN(_05824_)
  );
  AND2_X1 _13353_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05824_),
    .ZN(_05825_)
  );
  AND2_X1 _13354_ (
    .A1(_05823_),
    .A2(_05825_),
    .ZN(_05826_)
  );
  MUX2_X1 _13355_ (
    .A(\rf[22] [26]),
    .B(\rf[18] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05827_)
  );
  AND2_X1 _13356_ (
    .A1(_03045_),
    .A2(_05827_),
    .ZN(_05828_)
  );
  OR2_X1 _13357_ (
    .A1(_03044_),
    .A2(_05828_),
    .ZN(_05829_)
  );
  OR2_X1 _13358_ (
    .A1(_05826_),
    .A2(_05829_),
    .ZN(_05830_)
  );
  OR2_X1 _13359_ (
    .A1(\rf[17] [26]),
    .A2(_03046_),
    .ZN(_05831_)
  );
  OR2_X1 _13360_ (
    .A1(\rf[21] [26]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05832_)
  );
  AND2_X1 _13361_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05832_),
    .ZN(_05833_)
  );
  AND2_X1 _13362_ (
    .A1(_05831_),
    .A2(_05833_),
    .ZN(_05834_)
  );
  MUX2_X1 _13363_ (
    .A(\rf[23] [26]),
    .B(\rf[19] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05835_)
  );
  AND2_X1 _13364_ (
    .A1(_03045_),
    .A2(_05835_),
    .ZN(_05836_)
  );
  OR2_X1 _13365_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05836_),
    .ZN(_05837_)
  );
  OR2_X1 _13366_ (
    .A1(_05834_),
    .A2(_05837_),
    .ZN(_05838_)
  );
  AND2_X1 _13367_ (
    .A1(_05830_),
    .A2(_05838_),
    .ZN(_05839_)
  );
  OR2_X1 _13368_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_05839_),
    .ZN(_05840_)
  );
  AND2_X1 _13369_ (
    .A1(_05822_),
    .A2(_05840_),
    .ZN(_05841_)
  );
  AND2_X1 _13370_ (
    .A1(\rf[10] [26]),
    .A2(_03045_),
    .ZN(_05842_)
  );
  AND2_X1 _13371_ (
    .A1(\rf[8] [26]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05843_)
  );
  OR2_X1 _13372_ (
    .A1(_03046_),
    .A2(_05843_),
    .ZN(_05844_)
  );
  OR2_X1 _13373_ (
    .A1(_05842_),
    .A2(_05844_),
    .ZN(_05845_)
  );
  AND2_X1 _13374_ (
    .A1(\rf[14] [26]),
    .A2(_03045_),
    .ZN(_05846_)
  );
  AND2_X1 _13375_ (
    .A1(\rf[12] [26]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05847_)
  );
  OR2_X1 _13376_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_05847_),
    .ZN(_05848_)
  );
  OR2_X1 _13377_ (
    .A1(_05846_),
    .A2(_05848_),
    .ZN(_05849_)
  );
  AND2_X1 _13378_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05849_),
    .ZN(_05850_)
  );
  AND2_X1 _13379_ (
    .A1(_05845_),
    .A2(_05850_),
    .ZN(_05851_)
  );
  AND2_X1 _13380_ (
    .A1(\rf[11] [26]),
    .A2(_03045_),
    .ZN(_05852_)
  );
  AND2_X1 _13381_ (
    .A1(\rf[9] [26]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05853_)
  );
  OR2_X1 _13382_ (
    .A1(_03046_),
    .A2(_05853_),
    .ZN(_05854_)
  );
  OR2_X1 _13383_ (
    .A1(_05852_),
    .A2(_05854_),
    .ZN(_05855_)
  );
  AND2_X1 _13384_ (
    .A1(\rf[15] [26]),
    .A2(_03045_),
    .ZN(_05856_)
  );
  AND2_X1 _13385_ (
    .A1(\rf[13] [26]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05857_)
  );
  OR2_X1 _13386_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_05857_),
    .ZN(_05858_)
  );
  OR2_X1 _13387_ (
    .A1(_05856_),
    .A2(_05858_),
    .ZN(_05859_)
  );
  AND2_X1 _13388_ (
    .A1(_03044_),
    .A2(_05859_),
    .ZN(_05860_)
  );
  AND2_X1 _13389_ (
    .A1(_05855_),
    .A2(_05860_),
    .ZN(_05861_)
  );
  OR2_X1 _13390_ (
    .A1(_03063_),
    .A2(_05861_),
    .ZN(_05862_)
  );
  OR2_X1 _13391_ (
    .A1(_05851_),
    .A2(_05862_),
    .ZN(_05863_)
  );
  OR2_X1 _13392_ (
    .A1(\rf[28] [26]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05864_)
  );
  OR2_X1 _13393_ (
    .A1(\rf[24] [26]),
    .A2(_03046_),
    .ZN(_05865_)
  );
  AND2_X1 _13394_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05864_),
    .ZN(_05866_)
  );
  AND2_X1 _13395_ (
    .A1(_05865_),
    .A2(_05866_),
    .ZN(_05867_)
  );
  MUX2_X1 _13396_ (
    .A(\rf[30] [26]),
    .B(\rf[26] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05868_)
  );
  AND2_X1 _13397_ (
    .A1(_03045_),
    .A2(_05868_),
    .ZN(_05869_)
  );
  OR2_X1 _13398_ (
    .A1(_03044_),
    .A2(_05869_),
    .ZN(_05870_)
  );
  OR2_X1 _13399_ (
    .A1(_05867_),
    .A2(_05870_),
    .ZN(_05871_)
  );
  MUX2_X1 _13400_ (
    .A(\rf[29] [26]),
    .B(\rf[25] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05872_)
  );
  AND2_X1 _13401_ (
    .A1(\rf[27] [26]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05873_)
  );
  MUX2_X1 _13402_ (
    .A(_05872_),
    .B(_05873_),
    .S(_03045_),
    .Z(_05874_)
  );
  OR2_X1 _13403_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05874_),
    .ZN(_05875_)
  );
  AND2_X1 _13404_ (
    .A1(_05871_),
    .A2(_05875_),
    .ZN(_05876_)
  );
  OR2_X1 _13405_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_05876_),
    .ZN(_05877_)
  );
  AND2_X1 _13406_ (
    .A1(_05863_),
    .A2(_05877_),
    .ZN(_05878_)
  );
  MUX2_X1 _13407_ (
    .A(_05841_),
    .B(_05878_),
    .S(_03047_),
    .Z(_05879_)
  );
  MUX2_X1 _13408_ (
    .A(wb_reg_wdata[26]),
    .B(csr_io_rw_rdata[26]),
    .S(_04077_),
    .Z(_05880_)
  );
  MUX2_X1 _13409_ (
    .A(div_io_resp_bits_data[26]),
    .B(_05880_),
    .S(_03114_),
    .Z(_05881_)
  );
  MUX2_X1 _13410_ (
    .A(_05881_),
    .B(io_dmem_resp_bits_data[26]),
    .S(_03097_),
    .Z(_05882_)
  );
  MUX2_X1 _13411_ (
    .A(_05879_),
    .B(_05882_),
    .S(_04074_),
    .Z(_05883_)
  );
  AND2_X1 _13412_ (
    .A1(_04044_),
    .A2(_05883_),
    .ZN(_05884_)
  );
  OR2_X1 _13413_ (
    .A1(_05812_),
    .A2(_05884_),
    .ZN(_05885_)
  );
  MUX2_X1 _13414_ (
    .A(ex_reg_rs_msb_0[24]),
    .B(_05885_),
    .S(_04042_),
    .Z(_00091_)
  );
  AND2_X1 _13415_ (
    .A1(_03065_),
    .A2(ibuf_io_inst_0_bits_raw[27]),
    .ZN(_05886_)
  );
  AND2_X1 _13416_ (
    .A1(_03582_),
    .A2(_05886_),
    .ZN(_05887_)
  );
  MUX2_X1 _13417_ (
    .A(\rf[5] [27]),
    .B(\rf[1] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05888_)
  );
  MUX2_X1 _13418_ (
    .A(\rf[7] [27]),
    .B(\rf[3] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05889_)
  );
  MUX2_X1 _13419_ (
    .A(_05888_),
    .B(_05889_),
    .S(_03045_),
    .Z(_05890_)
  );
  AND2_X1 _13420_ (
    .A1(_03044_),
    .A2(_05890_),
    .ZN(_05891_)
  );
  MUX2_X1 _13421_ (
    .A(\rf[4] [27]),
    .B(\rf[0] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05892_)
  );
  MUX2_X1 _13422_ (
    .A(\rf[6] [27]),
    .B(\rf[2] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05893_)
  );
  MUX2_X1 _13423_ (
    .A(_05892_),
    .B(_05893_),
    .S(_03045_),
    .Z(_05894_)
  );
  AND2_X1 _13424_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05894_),
    .ZN(_05895_)
  );
  OR2_X1 _13425_ (
    .A1(_03063_),
    .A2(_05895_),
    .ZN(_05896_)
  );
  OR2_X1 _13426_ (
    .A1(_05891_),
    .A2(_05896_),
    .ZN(_05897_)
  );
  OR2_X1 _13427_ (
    .A1(\rf[20] [27]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05898_)
  );
  OR2_X1 _13428_ (
    .A1(\rf[16] [27]),
    .A2(_03046_),
    .ZN(_05899_)
  );
  AND2_X1 _13429_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05899_),
    .ZN(_05900_)
  );
  AND2_X1 _13430_ (
    .A1(_05898_),
    .A2(_05900_),
    .ZN(_05901_)
  );
  MUX2_X1 _13431_ (
    .A(\rf[22] [27]),
    .B(\rf[18] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05902_)
  );
  AND2_X1 _13432_ (
    .A1(_03045_),
    .A2(_05902_),
    .ZN(_05903_)
  );
  OR2_X1 _13433_ (
    .A1(_03044_),
    .A2(_05903_),
    .ZN(_05904_)
  );
  OR2_X1 _13434_ (
    .A1(_05901_),
    .A2(_05904_),
    .ZN(_05905_)
  );
  OR2_X1 _13435_ (
    .A1(\rf[17] [27]),
    .A2(_03046_),
    .ZN(_05906_)
  );
  OR2_X1 _13436_ (
    .A1(\rf[21] [27]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05907_)
  );
  AND2_X1 _13437_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05907_),
    .ZN(_05908_)
  );
  AND2_X1 _13438_ (
    .A1(_05906_),
    .A2(_05908_),
    .ZN(_05909_)
  );
  MUX2_X1 _13439_ (
    .A(\rf[23] [27]),
    .B(\rf[19] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05910_)
  );
  AND2_X1 _13440_ (
    .A1(_03045_),
    .A2(_05910_),
    .ZN(_05911_)
  );
  OR2_X1 _13441_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05911_),
    .ZN(_05912_)
  );
  OR2_X1 _13442_ (
    .A1(_05909_),
    .A2(_05912_),
    .ZN(_05913_)
  );
  AND2_X1 _13443_ (
    .A1(_05905_),
    .A2(_05913_),
    .ZN(_05914_)
  );
  OR2_X1 _13444_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_05914_),
    .ZN(_05915_)
  );
  AND2_X1 _13445_ (
    .A1(_05897_),
    .A2(_05915_),
    .ZN(_05916_)
  );
  AND2_X1 _13446_ (
    .A1(\rf[10] [27]),
    .A2(_03045_),
    .ZN(_05917_)
  );
  AND2_X1 _13447_ (
    .A1(\rf[8] [27]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05918_)
  );
  OR2_X1 _13448_ (
    .A1(_03046_),
    .A2(_05918_),
    .ZN(_05919_)
  );
  OR2_X1 _13449_ (
    .A1(_05917_),
    .A2(_05919_),
    .ZN(_05920_)
  );
  AND2_X1 _13450_ (
    .A1(\rf[14] [27]),
    .A2(_03045_),
    .ZN(_05921_)
  );
  AND2_X1 _13451_ (
    .A1(\rf[12] [27]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05922_)
  );
  OR2_X1 _13452_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_05922_),
    .ZN(_05923_)
  );
  OR2_X1 _13453_ (
    .A1(_05921_),
    .A2(_05923_),
    .ZN(_05924_)
  );
  AND2_X1 _13454_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05924_),
    .ZN(_05925_)
  );
  AND2_X1 _13455_ (
    .A1(_05920_),
    .A2(_05925_),
    .ZN(_05926_)
  );
  AND2_X1 _13456_ (
    .A1(\rf[11] [27]),
    .A2(_03045_),
    .ZN(_05927_)
  );
  AND2_X1 _13457_ (
    .A1(\rf[9] [27]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05928_)
  );
  OR2_X1 _13458_ (
    .A1(_03046_),
    .A2(_05928_),
    .ZN(_05929_)
  );
  OR2_X1 _13459_ (
    .A1(_05927_),
    .A2(_05929_),
    .ZN(_05930_)
  );
  AND2_X1 _13460_ (
    .A1(\rf[15] [27]),
    .A2(_03045_),
    .ZN(_05931_)
  );
  AND2_X1 _13461_ (
    .A1(\rf[13] [27]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05932_)
  );
  OR2_X1 _13462_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_05932_),
    .ZN(_05933_)
  );
  OR2_X1 _13463_ (
    .A1(_05931_),
    .A2(_05933_),
    .ZN(_05934_)
  );
  AND2_X1 _13464_ (
    .A1(_03044_),
    .A2(_05934_),
    .ZN(_05935_)
  );
  AND2_X1 _13465_ (
    .A1(_05930_),
    .A2(_05935_),
    .ZN(_05936_)
  );
  OR2_X1 _13466_ (
    .A1(_03063_),
    .A2(_05936_),
    .ZN(_05937_)
  );
  OR2_X1 _13467_ (
    .A1(_05926_),
    .A2(_05937_),
    .ZN(_05938_)
  );
  OR2_X1 _13468_ (
    .A1(\rf[28] [27]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05939_)
  );
  OR2_X1 _13469_ (
    .A1(\rf[24] [27]),
    .A2(_03046_),
    .ZN(_05940_)
  );
  AND2_X1 _13470_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05939_),
    .ZN(_05941_)
  );
  AND2_X1 _13471_ (
    .A1(_05940_),
    .A2(_05941_),
    .ZN(_05942_)
  );
  MUX2_X1 _13472_ (
    .A(\rf[30] [27]),
    .B(\rf[26] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05943_)
  );
  AND2_X1 _13473_ (
    .A1(_03045_),
    .A2(_05943_),
    .ZN(_05944_)
  );
  OR2_X1 _13474_ (
    .A1(_03044_),
    .A2(_05944_),
    .ZN(_05945_)
  );
  OR2_X1 _13475_ (
    .A1(_05942_),
    .A2(_05945_),
    .ZN(_05946_)
  );
  MUX2_X1 _13476_ (
    .A(\rf[29] [27]),
    .B(\rf[25] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05947_)
  );
  AND2_X1 _13477_ (
    .A1(\rf[27] [27]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05948_)
  );
  MUX2_X1 _13478_ (
    .A(_05947_),
    .B(_05948_),
    .S(_03045_),
    .Z(_05949_)
  );
  OR2_X1 _13479_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05949_),
    .ZN(_05950_)
  );
  AND2_X1 _13480_ (
    .A1(_05946_),
    .A2(_05950_),
    .ZN(_05951_)
  );
  OR2_X1 _13481_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_05951_),
    .ZN(_05952_)
  );
  AND2_X1 _13482_ (
    .A1(_05938_),
    .A2(_05952_),
    .ZN(_05953_)
  );
  MUX2_X1 _13483_ (
    .A(_05916_),
    .B(_05953_),
    .S(_03047_),
    .Z(_05954_)
  );
  MUX2_X1 _13484_ (
    .A(wb_reg_wdata[27]),
    .B(csr_io_rw_rdata[27]),
    .S(_04077_),
    .Z(_05955_)
  );
  MUX2_X1 _13485_ (
    .A(div_io_resp_bits_data[27]),
    .B(_05955_),
    .S(_03114_),
    .Z(_05956_)
  );
  MUX2_X1 _13486_ (
    .A(_05956_),
    .B(io_dmem_resp_bits_data[27]),
    .S(_03097_),
    .Z(_05957_)
  );
  MUX2_X1 _13487_ (
    .A(_05954_),
    .B(_05957_),
    .S(_04074_),
    .Z(_05958_)
  );
  AND2_X1 _13488_ (
    .A1(_04044_),
    .A2(_05958_),
    .ZN(_05959_)
  );
  OR2_X1 _13489_ (
    .A1(_05887_),
    .A2(_05959_),
    .ZN(_05960_)
  );
  MUX2_X1 _13490_ (
    .A(ex_reg_rs_msb_0[25]),
    .B(_05960_),
    .S(_04042_),
    .Z(_00092_)
  );
  AND2_X1 _13491_ (
    .A1(_03065_),
    .A2(ibuf_io_inst_0_bits_raw[28]),
    .ZN(_05961_)
  );
  AND2_X1 _13492_ (
    .A1(_03582_),
    .A2(_05961_),
    .ZN(_05962_)
  );
  MUX2_X1 _13493_ (
    .A(\rf[5] [28]),
    .B(\rf[1] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05963_)
  );
  MUX2_X1 _13494_ (
    .A(\rf[7] [28]),
    .B(\rf[3] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05964_)
  );
  MUX2_X1 _13495_ (
    .A(_05963_),
    .B(_05964_),
    .S(_03045_),
    .Z(_05965_)
  );
  AND2_X1 _13496_ (
    .A1(_03044_),
    .A2(_05965_),
    .ZN(_05966_)
  );
  MUX2_X1 _13497_ (
    .A(\rf[4] [28]),
    .B(\rf[0] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05967_)
  );
  MUX2_X1 _13498_ (
    .A(\rf[6] [28]),
    .B(\rf[2] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05968_)
  );
  MUX2_X1 _13499_ (
    .A(_05967_),
    .B(_05968_),
    .S(_03045_),
    .Z(_05969_)
  );
  AND2_X1 _13500_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05969_),
    .ZN(_05970_)
  );
  OR2_X1 _13501_ (
    .A1(_03063_),
    .A2(_05970_),
    .ZN(_05971_)
  );
  OR2_X1 _13502_ (
    .A1(_05966_),
    .A2(_05971_),
    .ZN(_05972_)
  );
  OR2_X1 _13503_ (
    .A1(\rf[20] [28]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05973_)
  );
  OR2_X1 _13504_ (
    .A1(\rf[16] [28]),
    .A2(_03046_),
    .ZN(_05974_)
  );
  AND2_X1 _13505_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05974_),
    .ZN(_05975_)
  );
  AND2_X1 _13506_ (
    .A1(_05973_),
    .A2(_05975_),
    .ZN(_05976_)
  );
  MUX2_X1 _13507_ (
    .A(\rf[22] [28]),
    .B(\rf[18] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05977_)
  );
  AND2_X1 _13508_ (
    .A1(_03045_),
    .A2(_05977_),
    .ZN(_05978_)
  );
  OR2_X1 _13509_ (
    .A1(_03044_),
    .A2(_05978_),
    .ZN(_05979_)
  );
  OR2_X1 _13510_ (
    .A1(_05976_),
    .A2(_05979_),
    .ZN(_05980_)
  );
  OR2_X1 _13511_ (
    .A1(\rf[17] [28]),
    .A2(_03046_),
    .ZN(_05981_)
  );
  OR2_X1 _13512_ (
    .A1(\rf[21] [28]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_05982_)
  );
  AND2_X1 _13513_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_05982_),
    .ZN(_05983_)
  );
  AND2_X1 _13514_ (
    .A1(_05981_),
    .A2(_05983_),
    .ZN(_05984_)
  );
  MUX2_X1 _13515_ (
    .A(\rf[23] [28]),
    .B(\rf[19] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_05985_)
  );
  AND2_X1 _13516_ (
    .A1(_03045_),
    .A2(_05985_),
    .ZN(_05986_)
  );
  OR2_X1 _13517_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05986_),
    .ZN(_05987_)
  );
  OR2_X1 _13518_ (
    .A1(_05984_),
    .A2(_05987_),
    .ZN(_05988_)
  );
  AND2_X1 _13519_ (
    .A1(_05980_),
    .A2(_05988_),
    .ZN(_05989_)
  );
  OR2_X1 _13520_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_05989_),
    .ZN(_05990_)
  );
  AND2_X1 _13521_ (
    .A1(_05972_),
    .A2(_05990_),
    .ZN(_05991_)
  );
  AND2_X1 _13522_ (
    .A1(\rf[10] [28]),
    .A2(_03045_),
    .ZN(_05992_)
  );
  AND2_X1 _13523_ (
    .A1(\rf[8] [28]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05993_)
  );
  OR2_X1 _13524_ (
    .A1(_03046_),
    .A2(_05993_),
    .ZN(_05994_)
  );
  OR2_X1 _13525_ (
    .A1(_05992_),
    .A2(_05994_),
    .ZN(_05995_)
  );
  AND2_X1 _13526_ (
    .A1(\rf[14] [28]),
    .A2(_03045_),
    .ZN(_05996_)
  );
  AND2_X1 _13527_ (
    .A1(\rf[12] [28]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_05997_)
  );
  OR2_X1 _13528_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_05997_),
    .ZN(_05998_)
  );
  OR2_X1 _13529_ (
    .A1(_05996_),
    .A2(_05998_),
    .ZN(_05999_)
  );
  AND2_X1 _13530_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_05999_),
    .ZN(_06000_)
  );
  AND2_X1 _13531_ (
    .A1(_05995_),
    .A2(_06000_),
    .ZN(_06001_)
  );
  AND2_X1 _13532_ (
    .A1(\rf[11] [28]),
    .A2(_03045_),
    .ZN(_06002_)
  );
  AND2_X1 _13533_ (
    .A1(\rf[9] [28]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_06003_)
  );
  OR2_X1 _13534_ (
    .A1(_03046_),
    .A2(_06003_),
    .ZN(_06004_)
  );
  OR2_X1 _13535_ (
    .A1(_06002_),
    .A2(_06004_),
    .ZN(_06005_)
  );
  AND2_X1 _13536_ (
    .A1(\rf[15] [28]),
    .A2(_03045_),
    .ZN(_06006_)
  );
  AND2_X1 _13537_ (
    .A1(\rf[13] [28]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_06007_)
  );
  OR2_X1 _13538_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_06007_),
    .ZN(_06008_)
  );
  OR2_X1 _13539_ (
    .A1(_06006_),
    .A2(_06008_),
    .ZN(_06009_)
  );
  AND2_X1 _13540_ (
    .A1(_03044_),
    .A2(_06009_),
    .ZN(_06010_)
  );
  AND2_X1 _13541_ (
    .A1(_06005_),
    .A2(_06010_),
    .ZN(_06011_)
  );
  OR2_X1 _13542_ (
    .A1(_03063_),
    .A2(_06011_),
    .ZN(_06012_)
  );
  OR2_X1 _13543_ (
    .A1(_06001_),
    .A2(_06012_),
    .ZN(_06013_)
  );
  OR2_X1 _13544_ (
    .A1(\rf[28] [28]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06014_)
  );
  OR2_X1 _13545_ (
    .A1(\rf[24] [28]),
    .A2(_03046_),
    .ZN(_06015_)
  );
  AND2_X1 _13546_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_06014_),
    .ZN(_06016_)
  );
  AND2_X1 _13547_ (
    .A1(_06015_),
    .A2(_06016_),
    .ZN(_06017_)
  );
  MUX2_X1 _13548_ (
    .A(\rf[30] [28]),
    .B(\rf[26] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06018_)
  );
  AND2_X1 _13549_ (
    .A1(_03045_),
    .A2(_06018_),
    .ZN(_06019_)
  );
  OR2_X1 _13550_ (
    .A1(_03044_),
    .A2(_06019_),
    .ZN(_06020_)
  );
  OR2_X1 _13551_ (
    .A1(_06017_),
    .A2(_06020_),
    .ZN(_06021_)
  );
  MUX2_X1 _13552_ (
    .A(\rf[29] [28]),
    .B(\rf[25] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06022_)
  );
  AND2_X1 _13553_ (
    .A1(\rf[27] [28]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06023_)
  );
  MUX2_X1 _13554_ (
    .A(_06022_),
    .B(_06023_),
    .S(_03045_),
    .Z(_06024_)
  );
  OR2_X1 _13555_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_06024_),
    .ZN(_06025_)
  );
  AND2_X1 _13556_ (
    .A1(_06021_),
    .A2(_06025_),
    .ZN(_06026_)
  );
  OR2_X1 _13557_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_06026_),
    .ZN(_06027_)
  );
  AND2_X1 _13558_ (
    .A1(_06013_),
    .A2(_06027_),
    .ZN(_06028_)
  );
  MUX2_X1 _13559_ (
    .A(_05991_),
    .B(_06028_),
    .S(_03047_),
    .Z(_06029_)
  );
  MUX2_X1 _13560_ (
    .A(wb_reg_wdata[28]),
    .B(csr_io_rw_rdata[28]),
    .S(_04077_),
    .Z(_06030_)
  );
  MUX2_X1 _13561_ (
    .A(div_io_resp_bits_data[28]),
    .B(_06030_),
    .S(_03114_),
    .Z(_06031_)
  );
  MUX2_X1 _13562_ (
    .A(_06031_),
    .B(io_dmem_resp_bits_data[28]),
    .S(_03097_),
    .Z(_06032_)
  );
  MUX2_X1 _13563_ (
    .A(_06029_),
    .B(_06032_),
    .S(_04074_),
    .Z(_06033_)
  );
  AND2_X1 _13564_ (
    .A1(_04044_),
    .A2(_06033_),
    .ZN(_06034_)
  );
  OR2_X1 _13565_ (
    .A1(_05962_),
    .A2(_06034_),
    .ZN(_06035_)
  );
  MUX2_X1 _13566_ (
    .A(ex_reg_rs_msb_0[26]),
    .B(_06035_),
    .S(_04042_),
    .Z(_00093_)
  );
  AND2_X1 _13567_ (
    .A1(_03065_),
    .A2(ibuf_io_inst_0_bits_raw[29]),
    .ZN(_06036_)
  );
  AND2_X1 _13568_ (
    .A1(_03582_),
    .A2(_06036_),
    .ZN(_06037_)
  );
  OR2_X1 _13569_ (
    .A1(\rf[10] [29]),
    .A2(_03046_),
    .ZN(_06038_)
  );
  OR2_X1 _13570_ (
    .A1(\rf[14] [29]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06039_)
  );
  AND2_X1 _13571_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_06039_),
    .ZN(_06040_)
  );
  AND2_X1 _13572_ (
    .A1(_06038_),
    .A2(_06040_),
    .ZN(_06041_)
  );
  MUX2_X1 _13573_ (
    .A(\rf[15] [29]),
    .B(\rf[11] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06042_)
  );
  AND2_X1 _13574_ (
    .A1(_03044_),
    .A2(_06042_),
    .ZN(_06043_)
  );
  OR2_X1 _13575_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_06043_),
    .ZN(_06044_)
  );
  OR2_X1 _13576_ (
    .A1(_06041_),
    .A2(_06044_),
    .ZN(_06045_)
  );
  OR2_X1 _13577_ (
    .A1(\rf[12] [29]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06046_)
  );
  OR2_X1 _13578_ (
    .A1(\rf[8] [29]),
    .A2(_03046_),
    .ZN(_06047_)
  );
  AND2_X1 _13579_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_06046_),
    .ZN(_06048_)
  );
  AND2_X1 _13580_ (
    .A1(_06047_),
    .A2(_06048_),
    .ZN(_06049_)
  );
  MUX2_X1 _13581_ (
    .A(\rf[13] [29]),
    .B(\rf[9] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06050_)
  );
  AND2_X1 _13582_ (
    .A1(_03044_),
    .A2(_06050_),
    .ZN(_06051_)
  );
  OR2_X1 _13583_ (
    .A1(_03045_),
    .A2(_06051_),
    .ZN(_06052_)
  );
  OR2_X1 _13584_ (
    .A1(_06049_),
    .A2(_06052_),
    .ZN(_06053_)
  );
  AND2_X1 _13585_ (
    .A1(_03047_),
    .A2(_06053_),
    .ZN(_06054_)
  );
  AND2_X1 _13586_ (
    .A1(_06045_),
    .A2(_06054_),
    .ZN(_06055_)
  );
  OR2_X1 _13587_ (
    .A1(\rf[0] [29]),
    .A2(_03046_),
    .ZN(_06056_)
  );
  OR2_X1 _13588_ (
    .A1(\rf[4] [29]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06057_)
  );
  AND2_X1 _13589_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_06057_),
    .ZN(_06058_)
  );
  AND2_X1 _13590_ (
    .A1(_06056_),
    .A2(_06058_),
    .ZN(_06059_)
  );
  MUX2_X1 _13591_ (
    .A(\rf[5] [29]),
    .B(\rf[1] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06060_)
  );
  AND2_X1 _13592_ (
    .A1(_03044_),
    .A2(_06060_),
    .ZN(_06061_)
  );
  OR2_X1 _13593_ (
    .A1(_03045_),
    .A2(_06061_),
    .ZN(_06062_)
  );
  OR2_X1 _13594_ (
    .A1(_06059_),
    .A2(_06062_),
    .ZN(_06063_)
  );
  MUX2_X1 _13595_ (
    .A(\rf[7] [29]),
    .B(\rf[3] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06064_)
  );
  AND2_X1 _13596_ (
    .A1(_03044_),
    .A2(_06064_),
    .ZN(_06065_)
  );
  OR2_X1 _13597_ (
    .A1(\rf[2] [29]),
    .A2(_03046_),
    .ZN(_06066_)
  );
  OR2_X1 _13598_ (
    .A1(\rf[6] [29]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06067_)
  );
  AND2_X1 _13599_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_06067_),
    .ZN(_06068_)
  );
  AND2_X1 _13600_ (
    .A1(_06066_),
    .A2(_06068_),
    .ZN(_06069_)
  );
  OR2_X1 _13601_ (
    .A1(_06065_),
    .A2(_06069_),
    .ZN(_06070_)
  );
  OR2_X1 _13602_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_06070_),
    .ZN(_06071_)
  );
  AND2_X1 _13603_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_06063_),
    .ZN(_06072_)
  );
  AND2_X1 _13604_ (
    .A1(_06071_),
    .A2(_06072_),
    .ZN(_06073_)
  );
  OR2_X1 _13605_ (
    .A1(_06055_),
    .A2(_06073_),
    .ZN(_06074_)
  );
  MUX2_X1 _13606_ (
    .A(\rf[30] [29]),
    .B(\rf[26] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06075_)
  );
  AND2_X1 _13607_ (
    .A1(\rf[27] [29]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06076_)
  );
  MUX2_X1 _13608_ (
    .A(_06075_),
    .B(_06076_),
    .S(_03044_),
    .Z(_06077_)
  );
  MUX2_X1 _13609_ (
    .A(\rf[29] [29]),
    .B(\rf[25] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06078_)
  );
  AND2_X1 _13610_ (
    .A1(_03044_),
    .A2(_06078_),
    .ZN(_06079_)
  );
  MUX2_X1 _13611_ (
    .A(\rf[28] [29]),
    .B(\rf[24] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06080_)
  );
  AND2_X1 _13612_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_06080_),
    .ZN(_06081_)
  );
  OR2_X1 _13613_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_06077_),
    .ZN(_06082_)
  );
  OR2_X1 _13614_ (
    .A1(_03045_),
    .A2(_06081_),
    .ZN(_06083_)
  );
  OR2_X1 _13615_ (
    .A1(_06079_),
    .A2(_06083_),
    .ZN(_06084_)
  );
  AND2_X1 _13616_ (
    .A1(_03047_),
    .A2(_06082_),
    .ZN(_06085_)
  );
  AND2_X1 _13617_ (
    .A1(_06084_),
    .A2(_06085_),
    .ZN(_06086_)
  );
  OR2_X1 _13618_ (
    .A1(\rf[18] [29]),
    .A2(_03046_),
    .ZN(_06087_)
  );
  OR2_X1 _13619_ (
    .A1(\rf[22] [29]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06088_)
  );
  AND2_X1 _13620_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_06088_),
    .ZN(_06089_)
  );
  AND2_X1 _13621_ (
    .A1(_06087_),
    .A2(_06089_),
    .ZN(_06090_)
  );
  MUX2_X1 _13622_ (
    .A(\rf[23] [29]),
    .B(\rf[19] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06091_)
  );
  AND2_X1 _13623_ (
    .A1(_03044_),
    .A2(_06091_),
    .ZN(_06092_)
  );
  OR2_X1 _13624_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_06092_),
    .ZN(_06093_)
  );
  OR2_X1 _13625_ (
    .A1(_06090_),
    .A2(_06093_),
    .ZN(_06094_)
  );
  MUX2_X1 _13626_ (
    .A(\rf[21] [29]),
    .B(\rf[17] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06095_)
  );
  AND2_X1 _13627_ (
    .A1(_03044_),
    .A2(_06095_),
    .ZN(_06096_)
  );
  OR2_X1 _13628_ (
    .A1(\rf[20] [29]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06097_)
  );
  OR2_X1 _13629_ (
    .A1(\rf[16] [29]),
    .A2(_03046_),
    .ZN(_06098_)
  );
  AND2_X1 _13630_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_06097_),
    .ZN(_06099_)
  );
  AND2_X1 _13631_ (
    .A1(_06098_),
    .A2(_06099_),
    .ZN(_06100_)
  );
  OR2_X1 _13632_ (
    .A1(_03045_),
    .A2(_06096_),
    .ZN(_06101_)
  );
  OR2_X1 _13633_ (
    .A1(_06100_),
    .A2(_06101_),
    .ZN(_06102_)
  );
  AND2_X1 _13634_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_06094_),
    .ZN(_06103_)
  );
  AND2_X1 _13635_ (
    .A1(_06102_),
    .A2(_06103_),
    .ZN(_06104_)
  );
  OR2_X1 _13636_ (
    .A1(_06086_),
    .A2(_06104_),
    .ZN(_06105_)
  );
  MUX2_X1 _13637_ (
    .A(_06074_),
    .B(_06105_),
    .S(_03063_),
    .Z(_06106_)
  );
  MUX2_X1 _13638_ (
    .A(wb_reg_wdata[29]),
    .B(csr_io_rw_rdata[29]),
    .S(_04077_),
    .Z(_06107_)
  );
  MUX2_X1 _13639_ (
    .A(div_io_resp_bits_data[29]),
    .B(_06107_),
    .S(_03114_),
    .Z(_06108_)
  );
  MUX2_X1 _13640_ (
    .A(_06108_),
    .B(io_dmem_resp_bits_data[29]),
    .S(_03097_),
    .Z(_06109_)
  );
  MUX2_X1 _13641_ (
    .A(_06106_),
    .B(_06109_),
    .S(_04074_),
    .Z(_06110_)
  );
  AND2_X1 _13642_ (
    .A1(_04044_),
    .A2(_06110_),
    .ZN(_06111_)
  );
  OR2_X1 _13643_ (
    .A1(_06037_),
    .A2(_06111_),
    .ZN(_06112_)
  );
  MUX2_X1 _13644_ (
    .A(ex_reg_rs_msb_0[27]),
    .B(_06112_),
    .S(_04042_),
    .Z(_00094_)
  );
  AND2_X1 _13645_ (
    .A1(_03065_),
    .A2(ibuf_io_inst_0_bits_raw[30]),
    .ZN(_06113_)
  );
  AND2_X1 _13646_ (
    .A1(_03582_),
    .A2(_06113_),
    .ZN(_06114_)
  );
  MUX2_X1 _13647_ (
    .A(wb_reg_wdata[30]),
    .B(csr_io_rw_rdata[30]),
    .S(_04077_),
    .Z(_06115_)
  );
  MUX2_X1 _13648_ (
    .A(div_io_resp_bits_data[30]),
    .B(_06115_),
    .S(_03114_),
    .Z(_06116_)
  );
  MUX2_X1 _13649_ (
    .A(_06116_),
    .B(io_dmem_resp_bits_data[30]),
    .S(_03097_),
    .Z(_06117_)
  );
  MUX2_X1 _13650_ (
    .A(\rf[5] [30]),
    .B(\rf[1] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06118_)
  );
  MUX2_X1 _13651_ (
    .A(\rf[7] [30]),
    .B(\rf[3] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06119_)
  );
  MUX2_X1 _13652_ (
    .A(_06118_),
    .B(_06119_),
    .S(_03045_),
    .Z(_06120_)
  );
  AND2_X1 _13653_ (
    .A1(_03044_),
    .A2(_06120_),
    .ZN(_06121_)
  );
  MUX2_X1 _13654_ (
    .A(\rf[4] [30]),
    .B(\rf[0] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06122_)
  );
  MUX2_X1 _13655_ (
    .A(\rf[6] [30]),
    .B(\rf[2] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06123_)
  );
  MUX2_X1 _13656_ (
    .A(_06122_),
    .B(_06123_),
    .S(_03045_),
    .Z(_06124_)
  );
  AND2_X1 _13657_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_06124_),
    .ZN(_06125_)
  );
  OR2_X1 _13658_ (
    .A1(_03063_),
    .A2(_06125_),
    .ZN(_06126_)
  );
  OR2_X1 _13659_ (
    .A1(_06121_),
    .A2(_06126_),
    .ZN(_06127_)
  );
  OR2_X1 _13660_ (
    .A1(\rf[20] [30]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06128_)
  );
  OR2_X1 _13661_ (
    .A1(\rf[16] [30]),
    .A2(_03046_),
    .ZN(_06129_)
  );
  AND2_X1 _13662_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_06129_),
    .ZN(_06130_)
  );
  AND2_X1 _13663_ (
    .A1(_06128_),
    .A2(_06130_),
    .ZN(_06131_)
  );
  MUX2_X1 _13664_ (
    .A(\rf[22] [30]),
    .B(\rf[18] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06132_)
  );
  AND2_X1 _13665_ (
    .A1(_03045_),
    .A2(_06132_),
    .ZN(_06133_)
  );
  OR2_X1 _13666_ (
    .A1(_03044_),
    .A2(_06133_),
    .ZN(_06134_)
  );
  OR2_X1 _13667_ (
    .A1(_06131_),
    .A2(_06134_),
    .ZN(_06135_)
  );
  OR2_X1 _13668_ (
    .A1(\rf[17] [30]),
    .A2(_03046_),
    .ZN(_06136_)
  );
  OR2_X1 _13669_ (
    .A1(\rf[21] [30]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06137_)
  );
  AND2_X1 _13670_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_06137_),
    .ZN(_06138_)
  );
  AND2_X1 _13671_ (
    .A1(_06136_),
    .A2(_06138_),
    .ZN(_06139_)
  );
  MUX2_X1 _13672_ (
    .A(\rf[23] [30]),
    .B(\rf[19] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06140_)
  );
  AND2_X1 _13673_ (
    .A1(_03045_),
    .A2(_06140_),
    .ZN(_06141_)
  );
  OR2_X1 _13674_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_06141_),
    .ZN(_06142_)
  );
  OR2_X1 _13675_ (
    .A1(_06139_),
    .A2(_06142_),
    .ZN(_06143_)
  );
  AND2_X1 _13676_ (
    .A1(_06135_),
    .A2(_06143_),
    .ZN(_06144_)
  );
  OR2_X1 _13677_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_06144_),
    .ZN(_06145_)
  );
  AND2_X1 _13678_ (
    .A1(_06127_),
    .A2(_06145_),
    .ZN(_06146_)
  );
  AND2_X1 _13679_ (
    .A1(\rf[10] [30]),
    .A2(_03045_),
    .ZN(_06147_)
  );
  AND2_X1 _13680_ (
    .A1(\rf[8] [30]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_06148_)
  );
  OR2_X1 _13681_ (
    .A1(_03046_),
    .A2(_06148_),
    .ZN(_06149_)
  );
  OR2_X1 _13682_ (
    .A1(_06147_),
    .A2(_06149_),
    .ZN(_06150_)
  );
  AND2_X1 _13683_ (
    .A1(\rf[14] [30]),
    .A2(_03045_),
    .ZN(_06151_)
  );
  AND2_X1 _13684_ (
    .A1(\rf[12] [30]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_06152_)
  );
  OR2_X1 _13685_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_06152_),
    .ZN(_06153_)
  );
  OR2_X1 _13686_ (
    .A1(_06151_),
    .A2(_06153_),
    .ZN(_06154_)
  );
  AND2_X1 _13687_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_06154_),
    .ZN(_06155_)
  );
  AND2_X1 _13688_ (
    .A1(_06150_),
    .A2(_06155_),
    .ZN(_06156_)
  );
  AND2_X1 _13689_ (
    .A1(\rf[11] [30]),
    .A2(_03045_),
    .ZN(_06157_)
  );
  AND2_X1 _13690_ (
    .A1(\rf[9] [30]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_06158_)
  );
  OR2_X1 _13691_ (
    .A1(_03046_),
    .A2(_06158_),
    .ZN(_06159_)
  );
  OR2_X1 _13692_ (
    .A1(_06157_),
    .A2(_06159_),
    .ZN(_06160_)
  );
  AND2_X1 _13693_ (
    .A1(\rf[15] [30]),
    .A2(_03045_),
    .ZN(_06161_)
  );
  AND2_X1 _13694_ (
    .A1(\rf[13] [30]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_06162_)
  );
  OR2_X1 _13695_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_06162_),
    .ZN(_06163_)
  );
  OR2_X1 _13696_ (
    .A1(_06161_),
    .A2(_06163_),
    .ZN(_06164_)
  );
  AND2_X1 _13697_ (
    .A1(_03044_),
    .A2(_06164_),
    .ZN(_06165_)
  );
  AND2_X1 _13698_ (
    .A1(_06160_),
    .A2(_06165_),
    .ZN(_06166_)
  );
  OR2_X1 _13699_ (
    .A1(_03063_),
    .A2(_06166_),
    .ZN(_06167_)
  );
  OR2_X1 _13700_ (
    .A1(_06156_),
    .A2(_06167_),
    .ZN(_06168_)
  );
  OR2_X1 _13701_ (
    .A1(\rf[28] [30]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06169_)
  );
  OR2_X1 _13702_ (
    .A1(\rf[24] [30]),
    .A2(_03046_),
    .ZN(_06170_)
  );
  AND2_X1 _13703_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_06169_),
    .ZN(_06171_)
  );
  AND2_X1 _13704_ (
    .A1(_06170_),
    .A2(_06171_),
    .ZN(_06172_)
  );
  MUX2_X1 _13705_ (
    .A(\rf[30] [30]),
    .B(\rf[26] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06173_)
  );
  AND2_X1 _13706_ (
    .A1(_03045_),
    .A2(_06173_),
    .ZN(_06174_)
  );
  OR2_X1 _13707_ (
    .A1(_03044_),
    .A2(_06174_),
    .ZN(_06175_)
  );
  OR2_X1 _13708_ (
    .A1(_06172_),
    .A2(_06175_),
    .ZN(_06176_)
  );
  MUX2_X1 _13709_ (
    .A(\rf[29] [30]),
    .B(\rf[25] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06177_)
  );
  AND2_X1 _13710_ (
    .A1(\rf[27] [30]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06178_)
  );
  MUX2_X1 _13711_ (
    .A(_06177_),
    .B(_06178_),
    .S(_03045_),
    .Z(_06179_)
  );
  OR2_X1 _13712_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_06179_),
    .ZN(_06180_)
  );
  AND2_X1 _13713_ (
    .A1(_06176_),
    .A2(_06180_),
    .ZN(_06181_)
  );
  OR2_X1 _13714_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_06181_),
    .ZN(_06182_)
  );
  AND2_X1 _13715_ (
    .A1(_06168_),
    .A2(_06182_),
    .ZN(_06183_)
  );
  MUX2_X1 _13716_ (
    .A(_06146_),
    .B(_06183_),
    .S(_03047_),
    .Z(_06184_)
  );
  MUX2_X1 _13717_ (
    .A(_06184_),
    .B(_06117_),
    .S(_04074_),
    .Z(_06185_)
  );
  AND2_X1 _13718_ (
    .A1(_04044_),
    .A2(_06185_),
    .ZN(_06186_)
  );
  OR2_X1 _13719_ (
    .A1(_06114_),
    .A2(_06186_),
    .ZN(_06187_)
  );
  MUX2_X1 _13720_ (
    .A(ex_reg_rs_msb_0[28]),
    .B(_06187_),
    .S(_04042_),
    .Z(_00095_)
  );
  AND2_X1 _13721_ (
    .A1(_03065_),
    .A2(ibuf_io_inst_0_bits_raw[31]),
    .ZN(_06188_)
  );
  AND2_X1 _13722_ (
    .A1(_03582_),
    .A2(_06188_),
    .ZN(_06189_)
  );
  MUX2_X1 _13723_ (
    .A(wb_reg_wdata[31]),
    .B(csr_io_rw_rdata[31]),
    .S(_04077_),
    .Z(_06190_)
  );
  MUX2_X1 _13724_ (
    .A(div_io_resp_bits_data[31]),
    .B(_06190_),
    .S(_03114_),
    .Z(_06191_)
  );
  MUX2_X1 _13725_ (
    .A(_06191_),
    .B(io_dmem_resp_bits_data[31]),
    .S(_03097_),
    .Z(_06192_)
  );
  MUX2_X1 _13726_ (
    .A(\rf[5] [31]),
    .B(\rf[1] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06193_)
  );
  MUX2_X1 _13727_ (
    .A(\rf[7] [31]),
    .B(\rf[3] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06194_)
  );
  MUX2_X1 _13728_ (
    .A(_06193_),
    .B(_06194_),
    .S(_03045_),
    .Z(_06195_)
  );
  AND2_X1 _13729_ (
    .A1(_03044_),
    .A2(_06195_),
    .ZN(_06196_)
  );
  MUX2_X1 _13730_ (
    .A(\rf[4] [31]),
    .B(\rf[0] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06197_)
  );
  MUX2_X1 _13731_ (
    .A(\rf[6] [31]),
    .B(\rf[2] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06198_)
  );
  MUX2_X1 _13732_ (
    .A(_06197_),
    .B(_06198_),
    .S(_03045_),
    .Z(_06199_)
  );
  AND2_X1 _13733_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_06199_),
    .ZN(_06200_)
  );
  OR2_X1 _13734_ (
    .A1(_03063_),
    .A2(_06200_),
    .ZN(_06201_)
  );
  OR2_X1 _13735_ (
    .A1(_06196_),
    .A2(_06201_),
    .ZN(_06202_)
  );
  OR2_X1 _13736_ (
    .A1(\rf[20] [31]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06203_)
  );
  OR2_X1 _13737_ (
    .A1(\rf[16] [31]),
    .A2(_03046_),
    .ZN(_06204_)
  );
  AND2_X1 _13738_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_06204_),
    .ZN(_06205_)
  );
  AND2_X1 _13739_ (
    .A1(_06203_),
    .A2(_06205_),
    .ZN(_06206_)
  );
  MUX2_X1 _13740_ (
    .A(\rf[22] [31]),
    .B(\rf[18] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06207_)
  );
  AND2_X1 _13741_ (
    .A1(_03045_),
    .A2(_06207_),
    .ZN(_06208_)
  );
  OR2_X1 _13742_ (
    .A1(_03044_),
    .A2(_06208_),
    .ZN(_06209_)
  );
  OR2_X1 _13743_ (
    .A1(_06206_),
    .A2(_06209_),
    .ZN(_06210_)
  );
  OR2_X1 _13744_ (
    .A1(\rf[17] [31]),
    .A2(_03046_),
    .ZN(_06211_)
  );
  OR2_X1 _13745_ (
    .A1(\rf[21] [31]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06212_)
  );
  AND2_X1 _13746_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_06212_),
    .ZN(_06213_)
  );
  AND2_X1 _13747_ (
    .A1(_06211_),
    .A2(_06213_),
    .ZN(_06214_)
  );
  MUX2_X1 _13748_ (
    .A(\rf[23] [31]),
    .B(\rf[19] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06215_)
  );
  AND2_X1 _13749_ (
    .A1(_03045_),
    .A2(_06215_),
    .ZN(_06216_)
  );
  OR2_X1 _13750_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_06216_),
    .ZN(_06217_)
  );
  OR2_X1 _13751_ (
    .A1(_06214_),
    .A2(_06217_),
    .ZN(_06218_)
  );
  AND2_X1 _13752_ (
    .A1(_06210_),
    .A2(_06218_),
    .ZN(_06219_)
  );
  OR2_X1 _13753_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_06219_),
    .ZN(_06220_)
  );
  AND2_X1 _13754_ (
    .A1(_06202_),
    .A2(_06220_),
    .ZN(_06221_)
  );
  AND2_X1 _13755_ (
    .A1(\rf[10] [31]),
    .A2(_03045_),
    .ZN(_06222_)
  );
  AND2_X1 _13756_ (
    .A1(\rf[8] [31]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_06223_)
  );
  OR2_X1 _13757_ (
    .A1(_03046_),
    .A2(_06223_),
    .ZN(_06224_)
  );
  OR2_X1 _13758_ (
    .A1(_06222_),
    .A2(_06224_),
    .ZN(_06225_)
  );
  AND2_X1 _13759_ (
    .A1(\rf[14] [31]),
    .A2(_03045_),
    .ZN(_06226_)
  );
  AND2_X1 _13760_ (
    .A1(\rf[12] [31]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_06227_)
  );
  OR2_X1 _13761_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_06227_),
    .ZN(_06228_)
  );
  OR2_X1 _13762_ (
    .A1(_06226_),
    .A2(_06228_),
    .ZN(_06229_)
  );
  AND2_X1 _13763_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_06229_),
    .ZN(_06230_)
  );
  AND2_X1 _13764_ (
    .A1(_06225_),
    .A2(_06230_),
    .ZN(_06231_)
  );
  AND2_X1 _13765_ (
    .A1(\rf[11] [31]),
    .A2(_03045_),
    .ZN(_06232_)
  );
  AND2_X1 _13766_ (
    .A1(\rf[9] [31]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_06233_)
  );
  OR2_X1 _13767_ (
    .A1(_03046_),
    .A2(_06233_),
    .ZN(_06234_)
  );
  OR2_X1 _13768_ (
    .A1(_06232_),
    .A2(_06234_),
    .ZN(_06235_)
  );
  AND2_X1 _13769_ (
    .A1(\rf[15] [31]),
    .A2(_03045_),
    .ZN(_06236_)
  );
  AND2_X1 _13770_ (
    .A1(\rf[13] [31]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[1]),
    .ZN(_06237_)
  );
  OR2_X1 _13771_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[2]),
    .A2(_06237_),
    .ZN(_06238_)
  );
  OR2_X1 _13772_ (
    .A1(_06236_),
    .A2(_06238_),
    .ZN(_06239_)
  );
  AND2_X1 _13773_ (
    .A1(_03044_),
    .A2(_06239_),
    .ZN(_06240_)
  );
  AND2_X1 _13774_ (
    .A1(_06235_),
    .A2(_06240_),
    .ZN(_06241_)
  );
  OR2_X1 _13775_ (
    .A1(_03063_),
    .A2(_06241_),
    .ZN(_06242_)
  );
  OR2_X1 _13776_ (
    .A1(_06231_),
    .A2(_06242_),
    .ZN(_06243_)
  );
  OR2_X1 _13777_ (
    .A1(\rf[28] [31]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06244_)
  );
  OR2_X1 _13778_ (
    .A1(\rf[24] [31]),
    .A2(_03046_),
    .ZN(_06245_)
  );
  AND2_X1 _13779_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_06244_),
    .ZN(_06246_)
  );
  AND2_X1 _13780_ (
    .A1(_06245_),
    .A2(_06246_),
    .ZN(_06247_)
  );
  MUX2_X1 _13781_ (
    .A(\rf[30] [31]),
    .B(\rf[26] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06248_)
  );
  AND2_X1 _13782_ (
    .A1(_03045_),
    .A2(_06248_),
    .ZN(_06249_)
  );
  OR2_X1 _13783_ (
    .A1(_03044_),
    .A2(_06249_),
    .ZN(_06250_)
  );
  OR2_X1 _13784_ (
    .A1(_06247_),
    .A2(_06250_),
    .ZN(_06251_)
  );
  MUX2_X1 _13785_ (
    .A(\rf[29] [31]),
    .B(\rf[25] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06252_)
  );
  AND2_X1 _13786_ (
    .A1(\rf[27] [31]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06253_)
  );
  MUX2_X1 _13787_ (
    .A(_06252_),
    .B(_06253_),
    .S(_03045_),
    .Z(_06254_)
  );
  OR2_X1 _13788_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_06254_),
    .ZN(_06255_)
  );
  AND2_X1 _13789_ (
    .A1(_06251_),
    .A2(_06255_),
    .ZN(_06256_)
  );
  OR2_X1 _13790_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[4]),
    .A2(_06256_),
    .ZN(_06257_)
  );
  AND2_X1 _13791_ (
    .A1(_06243_),
    .A2(_06257_),
    .ZN(_06258_)
  );
  MUX2_X1 _13792_ (
    .A(_06221_),
    .B(_06258_),
    .S(_03047_),
    .Z(_06259_)
  );
  MUX2_X1 _13793_ (
    .A(_06259_),
    .B(_06192_),
    .S(_04074_),
    .Z(_06260_)
  );
  AND2_X1 _13794_ (
    .A1(_04044_),
    .A2(_06260_),
    .ZN(_06261_)
  );
  OR2_X1 _13795_ (
    .A1(_06189_),
    .A2(_06261_),
    .ZN(_06262_)
  );
  MUX2_X1 _13796_ (
    .A(ex_reg_rs_msb_0[29]),
    .B(_06262_),
    .S(_04042_),
    .Z(_00096_)
  );
  OR2_X1 _13797_ (
    .A1(ibuf_io_inst_0_bits_raw[0]),
    .A2(_03583_),
    .ZN(_06263_)
  );
  MUX2_X1 _13798_ (
    .A(wb_reg_wdata[0]),
    .B(csr_io_rw_rdata[0]),
    .S(_04077_),
    .Z(_06264_)
  );
  MUX2_X1 _13799_ (
    .A(div_io_resp_bits_data[0]),
    .B(_06264_),
    .S(_03114_),
    .Z(_06265_)
  );
  MUX2_X1 _13800_ (
    .A(_06265_),
    .B(io_dmem_resp_bits_data[0]),
    .S(_03097_),
    .Z(_06266_)
  );
  OR2_X1 _13801_ (
    .A1(_04075_),
    .A2(_06266_),
    .ZN(_06267_)
  );
  OR2_X1 _13802_ (
    .A1(\rf[17] [0]),
    .A2(_03046_),
    .ZN(_06268_)
  );
  OR2_X1 _13803_ (
    .A1(\rf[21] [0]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06269_)
  );
  AND2_X1 _13804_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_06269_),
    .ZN(_06270_)
  );
  AND2_X1 _13805_ (
    .A1(_06268_),
    .A2(_06270_),
    .ZN(_06271_)
  );
  MUX2_X1 _13806_ (
    .A(\rf[23] [0]),
    .B(\rf[19] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06272_)
  );
  AND2_X1 _13807_ (
    .A1(_03045_),
    .A2(_06272_),
    .ZN(_06273_)
  );
  OR2_X1 _13808_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_06273_),
    .ZN(_06274_)
  );
  OR2_X1 _13809_ (
    .A1(_06271_),
    .A2(_06274_),
    .ZN(_06275_)
  );
  OR2_X1 _13810_ (
    .A1(\rf[20] [0]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06276_)
  );
  OR2_X1 _13811_ (
    .A1(\rf[16] [0]),
    .A2(_03046_),
    .ZN(_06277_)
  );
  AND2_X1 _13812_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_06277_),
    .ZN(_06278_)
  );
  AND2_X1 _13813_ (
    .A1(_06276_),
    .A2(_06278_),
    .ZN(_06279_)
  );
  MUX2_X1 _13814_ (
    .A(\rf[22] [0]),
    .B(\rf[18] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06280_)
  );
  AND2_X1 _13815_ (
    .A1(_03045_),
    .A2(_06280_),
    .ZN(_06281_)
  );
  OR2_X1 _13816_ (
    .A1(_03044_),
    .A2(_06281_),
    .ZN(_06282_)
  );
  OR2_X1 _13817_ (
    .A1(_06279_),
    .A2(_06282_),
    .ZN(_06283_)
  );
  AND2_X1 _13818_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_06275_),
    .ZN(_06284_)
  );
  AND2_X1 _13819_ (
    .A1(_06283_),
    .A2(_06284_),
    .ZN(_06285_)
  );
  OR2_X1 _13820_ (
    .A1(\rf[28] [0]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06286_)
  );
  OR2_X1 _13821_ (
    .A1(\rf[24] [0]),
    .A2(_03046_),
    .ZN(_06287_)
  );
  AND2_X1 _13822_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_06286_),
    .ZN(_06288_)
  );
  AND2_X1 _13823_ (
    .A1(_06287_),
    .A2(_06288_),
    .ZN(_06289_)
  );
  MUX2_X1 _13824_ (
    .A(\rf[30] [0]),
    .B(\rf[26] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06290_)
  );
  AND2_X1 _13825_ (
    .A1(_03045_),
    .A2(_06290_),
    .ZN(_06291_)
  );
  OR2_X1 _13826_ (
    .A1(_03044_),
    .A2(_06291_),
    .ZN(_06292_)
  );
  OR2_X1 _13827_ (
    .A1(_06289_),
    .A2(_06292_),
    .ZN(_06293_)
  );
  MUX2_X1 _13828_ (
    .A(\rf[29] [0]),
    .B(\rf[25] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06294_)
  );
  AND2_X1 _13829_ (
    .A1(\rf[27] [0]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06295_)
  );
  MUX2_X1 _13830_ (
    .A(_06294_),
    .B(_06295_),
    .S(_03045_),
    .Z(_06296_)
  );
  OR2_X1 _13831_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_06296_),
    .ZN(_06297_)
  );
  AND2_X1 _13832_ (
    .A1(_03047_),
    .A2(_06297_),
    .ZN(_06298_)
  );
  AND2_X1 _13833_ (
    .A1(_06293_),
    .A2(_06298_),
    .ZN(_06299_)
  );
  OR2_X1 _13834_ (
    .A1(_06285_),
    .A2(_06299_),
    .ZN(_06300_)
  );
  OR2_X1 _13835_ (
    .A1(\rf[10] [0]),
    .A2(_03046_),
    .ZN(_06301_)
  );
  OR2_X1 _13836_ (
    .A1(\rf[14] [0]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06302_)
  );
  AND2_X1 _13837_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_06302_),
    .ZN(_06303_)
  );
  AND2_X1 _13838_ (
    .A1(_06301_),
    .A2(_06303_),
    .ZN(_06304_)
  );
  MUX2_X1 _13839_ (
    .A(\rf[15] [0]),
    .B(\rf[11] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06305_)
  );
  AND2_X1 _13840_ (
    .A1(_03044_),
    .A2(_06305_),
    .ZN(_06306_)
  );
  OR2_X1 _13841_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_06306_),
    .ZN(_06307_)
  );
  OR2_X1 _13842_ (
    .A1(_06304_),
    .A2(_06307_),
    .ZN(_06308_)
  );
  OR2_X1 _13843_ (
    .A1(\rf[12] [0]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06309_)
  );
  OR2_X1 _13844_ (
    .A1(\rf[8] [0]),
    .A2(_03046_),
    .ZN(_06310_)
  );
  AND2_X1 _13845_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_06309_),
    .ZN(_06311_)
  );
  AND2_X1 _13846_ (
    .A1(_06310_),
    .A2(_06311_),
    .ZN(_06312_)
  );
  MUX2_X1 _13847_ (
    .A(\rf[13] [0]),
    .B(\rf[9] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06313_)
  );
  AND2_X1 _13848_ (
    .A1(_03044_),
    .A2(_06313_),
    .ZN(_06314_)
  );
  OR2_X1 _13849_ (
    .A1(_03045_),
    .A2(_06314_),
    .ZN(_06315_)
  );
  OR2_X1 _13850_ (
    .A1(_06312_),
    .A2(_06315_),
    .ZN(_06316_)
  );
  AND2_X1 _13851_ (
    .A1(_03047_),
    .A2(_06316_),
    .ZN(_06317_)
  );
  AND2_X1 _13852_ (
    .A1(_06308_),
    .A2(_06317_),
    .ZN(_06318_)
  );
  MUX2_X1 _13853_ (
    .A(\rf[6] [0]),
    .B(\rf[2] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06319_)
  );
  AND2_X1 _13854_ (
    .A1(_03045_),
    .A2(_06319_),
    .ZN(_06320_)
  );
  MUX2_X1 _13855_ (
    .A(\rf[4] [0]),
    .B(\rf[0] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06321_)
  );
  AND2_X1 _13856_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_06321_),
    .ZN(_06322_)
  );
  OR2_X1 _13857_ (
    .A1(_03044_),
    .A2(_06322_),
    .ZN(_06323_)
  );
  OR2_X1 _13858_ (
    .A1(_06320_),
    .A2(_06323_),
    .ZN(_06324_)
  );
  MUX2_X1 _13859_ (
    .A(\rf[7] [0]),
    .B(\rf[3] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06325_)
  );
  AND2_X1 _13860_ (
    .A1(_03045_),
    .A2(_06325_),
    .ZN(_06326_)
  );
  MUX2_X1 _13861_ (
    .A(\rf[5] [0]),
    .B(\rf[1] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06327_)
  );
  AND2_X1 _13862_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_06327_),
    .ZN(_06328_)
  );
  OR2_X1 _13863_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_06328_),
    .ZN(_06329_)
  );
  OR2_X1 _13864_ (
    .A1(_06326_),
    .A2(_06329_),
    .ZN(_06330_)
  );
  AND2_X1 _13865_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_06330_),
    .ZN(_06331_)
  );
  AND2_X1 _13866_ (
    .A1(_06324_),
    .A2(_06331_),
    .ZN(_06332_)
  );
  OR2_X1 _13867_ (
    .A1(_06318_),
    .A2(_06332_),
    .ZN(_06333_)
  );
  MUX2_X1 _13868_ (
    .A(_06300_),
    .B(_06333_),
    .S(ibuf_io_inst_0_bits_inst_rs1[4]),
    .Z(_06334_)
  );
  OR2_X1 _13869_ (
    .A1(_04074_),
    .A2(_06334_),
    .ZN(_06335_)
  );
  AND2_X1 _13870_ (
    .A1(_03490_),
    .A2(_06335_),
    .ZN(_06336_)
  );
  AND2_X1 _13871_ (
    .A1(_06267_),
    .A2(_06336_),
    .ZN(_06337_)
  );
  OR2_X1 _13872_ (
    .A1(_03092_),
    .A2(_03472_),
    .ZN(_06338_)
  );
  OR2_X1 _13873_ (
    .A1(_03485_),
    .A2(_06338_),
    .ZN(_06339_)
  );
  OR2_X1 _13874_ (
    .A1(_03467_),
    .A2(_06339_),
    .ZN(_06340_)
  );
  AND2_X1 _13875_ (
    .A1(_03451_),
    .A2(_06340_),
    .ZN(_06341_)
  );
  OR2_X1 _13876_ (
    .A1(_03582_),
    .A2(_06341_),
    .ZN(_06342_)
  );
  AND2_X1 _13877_ (
    .A1(_04045_),
    .A2(_06342_),
    .ZN(_06343_)
  );
  OR2_X1 _13878_ (
    .A1(_06337_),
    .A2(_06343_),
    .ZN(_06344_)
  );
  AND2_X1 _13879_ (
    .A1(_06263_),
    .A2(_06344_),
    .ZN(_06345_)
  );
  MUX2_X1 _13880_ (
    .A(_06345_),
    .B(ex_reg_rs_lsb_0[0]),
    .S(_04146_),
    .Z(_00097_)
  );
  AND2_X1 _13881_ (
    .A1(_03469_),
    .A2(_03585_),
    .ZN(_06346_)
  );
  AND2_X1 _13882_ (
    .A1(ibuf_io_inst_0_bits_raw[1]),
    .A2(_03582_),
    .ZN(_06347_)
  );
  OR2_X1 _13883_ (
    .A1(_06346_),
    .A2(_06347_),
    .ZN(_06348_)
  );
  OR2_X1 _13884_ (
    .A1(\rf[10] [1]),
    .A2(_03046_),
    .ZN(_06349_)
  );
  OR2_X1 _13885_ (
    .A1(\rf[14] [1]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06350_)
  );
  AND2_X1 _13886_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_06350_),
    .ZN(_06351_)
  );
  AND2_X1 _13887_ (
    .A1(_06349_),
    .A2(_06351_),
    .ZN(_06352_)
  );
  MUX2_X1 _13888_ (
    .A(\rf[15] [1]),
    .B(\rf[11] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06353_)
  );
  AND2_X1 _13889_ (
    .A1(_03044_),
    .A2(_06353_),
    .ZN(_06354_)
  );
  OR2_X1 _13890_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_06354_),
    .ZN(_06355_)
  );
  OR2_X1 _13891_ (
    .A1(_06352_),
    .A2(_06355_),
    .ZN(_06356_)
  );
  OR2_X1 _13892_ (
    .A1(\rf[12] [1]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06357_)
  );
  OR2_X1 _13893_ (
    .A1(\rf[8] [1]),
    .A2(_03046_),
    .ZN(_06358_)
  );
  AND2_X1 _13894_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_06357_),
    .ZN(_06359_)
  );
  AND2_X1 _13895_ (
    .A1(_06358_),
    .A2(_06359_),
    .ZN(_06360_)
  );
  MUX2_X1 _13896_ (
    .A(\rf[13] [1]),
    .B(\rf[9] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06361_)
  );
  AND2_X1 _13897_ (
    .A1(_03044_),
    .A2(_06361_),
    .ZN(_06362_)
  );
  OR2_X1 _13898_ (
    .A1(_03045_),
    .A2(_06362_),
    .ZN(_06363_)
  );
  OR2_X1 _13899_ (
    .A1(_06360_),
    .A2(_06363_),
    .ZN(_06364_)
  );
  AND2_X1 _13900_ (
    .A1(_03047_),
    .A2(_06364_),
    .ZN(_06365_)
  );
  AND2_X1 _13901_ (
    .A1(_06356_),
    .A2(_06365_),
    .ZN(_06366_)
  );
  MUX2_X1 _13902_ (
    .A(\rf[7] [1]),
    .B(\rf[3] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06367_)
  );
  AND2_X1 _13903_ (
    .A1(_03044_),
    .A2(_06367_),
    .ZN(_06368_)
  );
  OR2_X1 _13904_ (
    .A1(\rf[2] [1]),
    .A2(_03046_),
    .ZN(_06369_)
  );
  OR2_X1 _13905_ (
    .A1(\rf[6] [1]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06370_)
  );
  AND2_X1 _13906_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_06370_),
    .ZN(_06371_)
  );
  AND2_X1 _13907_ (
    .A1(_06369_),
    .A2(_06371_),
    .ZN(_06372_)
  );
  OR2_X1 _13908_ (
    .A1(_06368_),
    .A2(_06372_),
    .ZN(_06373_)
  );
  OR2_X1 _13909_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_06373_),
    .ZN(_06374_)
  );
  OR2_X1 _13910_ (
    .A1(\rf[0] [1]),
    .A2(_03046_),
    .ZN(_06375_)
  );
  OR2_X1 _13911_ (
    .A1(\rf[4] [1]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06376_)
  );
  AND2_X1 _13912_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_06376_),
    .ZN(_06377_)
  );
  AND2_X1 _13913_ (
    .A1(_06375_),
    .A2(_06377_),
    .ZN(_06378_)
  );
  MUX2_X1 _13914_ (
    .A(\rf[5] [1]),
    .B(\rf[1] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06379_)
  );
  AND2_X1 _13915_ (
    .A1(_03044_),
    .A2(_06379_),
    .ZN(_06380_)
  );
  OR2_X1 _13916_ (
    .A1(_03045_),
    .A2(_06380_),
    .ZN(_06381_)
  );
  OR2_X1 _13917_ (
    .A1(_06378_),
    .A2(_06381_),
    .ZN(_06382_)
  );
  AND2_X1 _13918_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_06382_),
    .ZN(_06383_)
  );
  AND2_X1 _13919_ (
    .A1(_06374_),
    .A2(_06383_),
    .ZN(_06384_)
  );
  OR2_X1 _13920_ (
    .A1(_06366_),
    .A2(_06384_),
    .ZN(_06385_)
  );
  MUX2_X1 _13921_ (
    .A(\rf[29] [1]),
    .B(\rf[25] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06386_)
  );
  AND2_X1 _13922_ (
    .A1(_03044_),
    .A2(_06386_),
    .ZN(_06387_)
  );
  MUX2_X1 _13923_ (
    .A(\rf[28] [1]),
    .B(\rf[24] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06388_)
  );
  AND2_X1 _13924_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_06388_),
    .ZN(_06389_)
  );
  OR2_X1 _13925_ (
    .A1(_03045_),
    .A2(_06389_),
    .ZN(_06390_)
  );
  OR2_X1 _13926_ (
    .A1(_06387_),
    .A2(_06390_),
    .ZN(_06391_)
  );
  MUX2_X1 _13927_ (
    .A(\rf[30] [1]),
    .B(\rf[26] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06392_)
  );
  AND2_X1 _13928_ (
    .A1(\rf[27] [1]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06393_)
  );
  MUX2_X1 _13929_ (
    .A(_06392_),
    .B(_06393_),
    .S(_03044_),
    .Z(_06394_)
  );
  OR2_X1 _13930_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_06394_),
    .ZN(_06395_)
  );
  AND2_X1 _13931_ (
    .A1(_03047_),
    .A2(_06395_),
    .ZN(_06396_)
  );
  AND2_X1 _13932_ (
    .A1(_06391_),
    .A2(_06396_),
    .ZN(_06397_)
  );
  OR2_X1 _13933_ (
    .A1(\rf[18] [1]),
    .A2(_03046_),
    .ZN(_06398_)
  );
  OR2_X1 _13934_ (
    .A1(\rf[22] [1]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06399_)
  );
  AND2_X1 _13935_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_06399_),
    .ZN(_06400_)
  );
  AND2_X1 _13936_ (
    .A1(_06398_),
    .A2(_06400_),
    .ZN(_06401_)
  );
  MUX2_X1 _13937_ (
    .A(\rf[23] [1]),
    .B(\rf[19] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06402_)
  );
  AND2_X1 _13938_ (
    .A1(_03044_),
    .A2(_06402_),
    .ZN(_06403_)
  );
  OR2_X1 _13939_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[1]),
    .A2(_06403_),
    .ZN(_06404_)
  );
  OR2_X1 _13940_ (
    .A1(_06401_),
    .A2(_06404_),
    .ZN(_06405_)
  );
  MUX2_X1 _13941_ (
    .A(\rf[21] [1]),
    .B(\rf[17] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs1[2]),
    .Z(_06406_)
  );
  AND2_X1 _13942_ (
    .A1(_03044_),
    .A2(_06406_),
    .ZN(_06407_)
  );
  OR2_X1 _13943_ (
    .A1(\rf[20] [1]),
    .A2(ibuf_io_inst_0_bits_inst_rs1[2]),
    .ZN(_06408_)
  );
  OR2_X1 _13944_ (
    .A1(\rf[16] [1]),
    .A2(_03046_),
    .ZN(_06409_)
  );
  AND2_X1 _13945_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[0]),
    .A2(_06408_),
    .ZN(_06410_)
  );
  AND2_X1 _13946_ (
    .A1(_06409_),
    .A2(_06410_),
    .ZN(_06411_)
  );
  OR2_X1 _13947_ (
    .A1(_03045_),
    .A2(_06407_),
    .ZN(_06412_)
  );
  OR2_X1 _13948_ (
    .A1(_06411_),
    .A2(_06412_),
    .ZN(_06413_)
  );
  AND2_X1 _13949_ (
    .A1(ibuf_io_inst_0_bits_inst_rs1[3]),
    .A2(_06405_),
    .ZN(_06414_)
  );
  AND2_X1 _13950_ (
    .A1(_06413_),
    .A2(_06414_),
    .ZN(_06415_)
  );
  OR2_X1 _13951_ (
    .A1(_06397_),
    .A2(_06415_),
    .ZN(_06416_)
  );
  MUX2_X1 _13952_ (
    .A(_06385_),
    .B(_06416_),
    .S(_03063_),
    .Z(_06417_)
  );
  MUX2_X1 _13953_ (
    .A(wb_reg_wdata[1]),
    .B(csr_io_rw_rdata[1]),
    .S(_04077_),
    .Z(_06418_)
  );
  MUX2_X1 _13954_ (
    .A(div_io_resp_bits_data[1]),
    .B(_06418_),
    .S(_03114_),
    .Z(_06419_)
  );
  MUX2_X1 _13955_ (
    .A(_06419_),
    .B(io_dmem_resp_bits_data[1]),
    .S(_03097_),
    .Z(_06420_)
  );
  MUX2_X1 _13956_ (
    .A(_06417_),
    .B(_06420_),
    .S(_04074_),
    .Z(_06421_)
  );
  AND2_X1 _13957_ (
    .A1(_04044_),
    .A2(_06421_),
    .ZN(_06422_)
  );
  OR2_X1 _13958_ (
    .A1(_06348_),
    .A2(_06422_),
    .ZN(_06423_)
  );
  MUX2_X1 _13959_ (
    .A(_06423_),
    .B(ex_reg_rs_lsb_0[1]),
    .S(_04146_),
    .Z(_00098_)
  );
  AND2_X1 _13960_ (
    .A1(_03452_),
    .A2(_04002_),
    .ZN(_06424_)
  );
  INV_X1 _13961_ (
    .A(_06424_),
    .ZN(_06425_)
  );
  AND2_X1 _13962_ (
    .A1(_03811_),
    .A2(_06425_),
    .ZN(_06426_)
  );
  INV_X1 _13963_ (
    .A(_06426_),
    .ZN(_06427_)
  );
  OR2_X1 _13964_ (
    .A1(_03912_),
    .A2(_06427_),
    .ZN(_06428_)
  );
  MUX2_X1 _13965_ (
    .A(_06428_),
    .B(ex_reg_rs_bypass_1),
    .S(_04146_),
    .Z(_00099_)
  );
  AND2_X1 _13966_ (
    .A1(_03488_),
    .A2(_03583_),
    .ZN(_06429_)
  );
  MUX2_X1 _13967_ (
    .A(_06429_),
    .B(ex_reg_rs_bypass_0),
    .S(_04146_),
    .Z(_00100_)
  );
  OR2_X1 _13968_ (
    .A1(mem_reg_valid),
    .A2(mem_reg_replay),
    .ZN(_06430_)
  );
  INV_X1 _13969_ (
    .A(_06430_),
    .ZN(_06431_)
  );
  AND2_X1 _13970_ (
    .A1(_03094_),
    .A2(_06431_),
    .ZN(_06432_)
  );
  OR2_X1 _13971_ (
    .A1(mem_reg_xcpt_interrupt),
    .A2(_06430_),
    .ZN(_06433_)
  );
  MUX2_X1 _13972_ (
    .A(wb_reg_raw_inst[0]),
    .B(mem_reg_raw_inst[0]),
    .S(_06433_),
    .Z(_00101_)
  );
  MUX2_X1 _13973_ (
    .A(wb_reg_raw_inst[1]),
    .B(mem_reg_raw_inst[1]),
    .S(_06433_),
    .Z(_00102_)
  );
  MUX2_X1 _13974_ (
    .A(wb_reg_raw_inst[2]),
    .B(mem_reg_raw_inst[2]),
    .S(_06433_),
    .Z(_00103_)
  );
  MUX2_X1 _13975_ (
    .A(wb_reg_raw_inst[3]),
    .B(mem_reg_raw_inst[3]),
    .S(_06433_),
    .Z(_00104_)
  );
  MUX2_X1 _13976_ (
    .A(wb_reg_raw_inst[4]),
    .B(mem_reg_raw_inst[4]),
    .S(_06433_),
    .Z(_00105_)
  );
  MUX2_X1 _13977_ (
    .A(wb_reg_raw_inst[5]),
    .B(mem_reg_raw_inst[5]),
    .S(_06433_),
    .Z(_00106_)
  );
  MUX2_X1 _13978_ (
    .A(wb_reg_raw_inst[6]),
    .B(mem_reg_raw_inst[6]),
    .S(_06433_),
    .Z(_00107_)
  );
  MUX2_X1 _13979_ (
    .A(wb_reg_raw_inst[7]),
    .B(mem_reg_raw_inst[7]),
    .S(_06433_),
    .Z(_00108_)
  );
  MUX2_X1 _13980_ (
    .A(wb_reg_raw_inst[8]),
    .B(mem_reg_raw_inst[8]),
    .S(_06433_),
    .Z(_00109_)
  );
  MUX2_X1 _13981_ (
    .A(wb_reg_raw_inst[9]),
    .B(mem_reg_raw_inst[9]),
    .S(_06433_),
    .Z(_00110_)
  );
  MUX2_X1 _13982_ (
    .A(wb_reg_raw_inst[10]),
    .B(mem_reg_raw_inst[10]),
    .S(_06433_),
    .Z(_00111_)
  );
  MUX2_X1 _13983_ (
    .A(wb_reg_raw_inst[11]),
    .B(mem_reg_raw_inst[11]),
    .S(_06433_),
    .Z(_00112_)
  );
  MUX2_X1 _13984_ (
    .A(wb_reg_raw_inst[12]),
    .B(mem_reg_raw_inst[12]),
    .S(_06433_),
    .Z(_00113_)
  );
  MUX2_X1 _13985_ (
    .A(wb_reg_raw_inst[13]),
    .B(mem_reg_raw_inst[13]),
    .S(_06433_),
    .Z(_00114_)
  );
  MUX2_X1 _13986_ (
    .A(wb_reg_raw_inst[14]),
    .B(mem_reg_raw_inst[14]),
    .S(_06433_),
    .Z(_00115_)
  );
  MUX2_X1 _13987_ (
    .A(wb_reg_raw_inst[15]),
    .B(mem_reg_raw_inst[15]),
    .S(_06433_),
    .Z(_00116_)
  );
  MUX2_X1 _13988_ (
    .A(mem_reg_rvc),
    .B(mem_reg_inst[21]),
    .S(mem_ctrl_jal),
    .Z(_06434_)
  );
  MUX2_X1 _13989_ (
    .A(_06434_),
    .B(mem_reg_inst[8]),
    .S(_04030_),
    .Z(_06435_)
  );
  AND2_X1 _13990_ (
    .A1(mem_reg_pc[1]),
    .A2(_06435_),
    .ZN(_06436_)
  );
  XOR2_X1 _13991_ (
    .A(mem_reg_pc[1]),
    .B(_06435_),
    .Z(_06437_)
  );
  MUX2_X1 _13992_ (
    .A(mem_reg_wdata[1]),
    .B(_06437_),
    .S(_03030_),
    .Z(_06438_)
  );
  AND2_X1 _13993_ (
    .A1(_03079_),
    .A2(_06438_),
    .ZN(_06439_)
  );
  XOR2_X1 _13994_ (
    .A(mem_ctrl_jalr),
    .B(_06439_),
    .Z(_06440_)
  );
  XOR2_X1 _13995_ (
    .A(_03030_),
    .B(_06439_),
    .Z(_06441_)
  );
  AND2_X1 _13996_ (
    .A1(_take_pc_mem_T),
    .A2(_06440_),
    .ZN(_06442_)
  );
  OR2_X1 _13997_ (
    .A1(_03091_),
    .A2(_06441_),
    .ZN(_06443_)
  );
  MUX2_X1 _13998_ (
    .A(mem_reg_pc[0]),
    .B(mem_reg_wdata[0]),
    .S(_06443_),
    .Z(_06444_)
  );
  MUX2_X1 _13999_ (
    .A(wb_reg_wdata[0]),
    .B(_06444_),
    .S(_06433_),
    .Z(_00117_)
  );
  MUX2_X1 _14000_ (
    .A(mem_reg_wdata[1]),
    .B(_06437_),
    .S(_06442_),
    .Z(_06445_)
  );
  MUX2_X1 _14001_ (
    .A(wb_reg_wdata[1]),
    .B(_06445_),
    .S(_06433_),
    .Z(_00118_)
  );
  MUX2_X1 _14002_ (
    .A(_mem_br_target_T_6[2]),
    .B(mem_reg_inst[22]),
    .S(mem_ctrl_jal),
    .Z(_06446_)
  );
  MUX2_X1 _14003_ (
    .A(_06446_),
    .B(mem_reg_inst[9]),
    .S(_04030_),
    .Z(_06447_)
  );
  AND2_X1 _14004_ (
    .A1(mem_reg_pc[2]),
    .A2(_06447_),
    .ZN(_06448_)
  );
  XOR2_X1 _14005_ (
    .A(mem_reg_pc[2]),
    .B(_06447_),
    .Z(_06449_)
  );
  AND2_X1 _14006_ (
    .A1(_06436_),
    .A2(_06449_),
    .ZN(_06450_)
  );
  XOR2_X1 _14007_ (
    .A(_06436_),
    .B(_06449_),
    .Z(_06451_)
  );
  MUX2_X1 _14008_ (
    .A(mem_reg_wdata[2]),
    .B(_06451_),
    .S(_06442_),
    .Z(_06452_)
  );
  MUX2_X1 _14009_ (
    .A(wb_reg_wdata[2]),
    .B(_06452_),
    .S(_06433_),
    .Z(_00119_)
  );
  OR2_X1 _14010_ (
    .A1(_06448_),
    .A2(_06450_),
    .ZN(_06453_)
  );
  AND2_X1 _14011_ (
    .A1(mem_reg_inst[23]),
    .A2(mem_ctrl_jal),
    .ZN(_06454_)
  );
  MUX2_X1 _14012_ (
    .A(_06454_),
    .B(mem_reg_inst[10]),
    .S(_04030_),
    .Z(_06455_)
  );
  AND2_X1 _14013_ (
    .A1(mem_reg_pc[3]),
    .A2(_06455_),
    .ZN(_06456_)
  );
  OR2_X1 _14014_ (
    .A1(mem_reg_pc[3]),
    .A2(_06455_),
    .ZN(_06457_)
  );
  XOR2_X1 _14015_ (
    .A(mem_reg_pc[3]),
    .B(_06455_),
    .Z(_06458_)
  );
  XOR2_X1 _14016_ (
    .A(_06453_),
    .B(_06458_),
    .Z(_06459_)
  );
  MUX2_X1 _14017_ (
    .A(mem_reg_wdata[3]),
    .B(_06459_),
    .S(_06442_),
    .Z(_06460_)
  );
  MUX2_X1 _14018_ (
    .A(wb_reg_wdata[3]),
    .B(_06460_),
    .S(_06433_),
    .Z(_00120_)
  );
  AND2_X1 _14019_ (
    .A1(mem_reg_inst[24]),
    .A2(mem_ctrl_jal),
    .ZN(_06461_)
  );
  MUX2_X1 _14020_ (
    .A(_06461_),
    .B(mem_reg_inst[11]),
    .S(_04030_),
    .Z(_06462_)
  );
  AND2_X1 _14021_ (
    .A1(mem_reg_pc[4]),
    .A2(_06462_),
    .ZN(_06463_)
  );
  XOR2_X1 _14022_ (
    .A(mem_reg_pc[4]),
    .B(_06462_),
    .Z(_06464_)
  );
  AND2_X1 _14023_ (
    .A1(_06453_),
    .A2(_06457_),
    .ZN(_06465_)
  );
  OR2_X1 _14024_ (
    .A1(_06456_),
    .A2(_06465_),
    .ZN(_06466_)
  );
  AND2_X1 _14025_ (
    .A1(_06464_),
    .A2(_06466_),
    .ZN(_06467_)
  );
  XOR2_X1 _14026_ (
    .A(_06464_),
    .B(_06466_),
    .Z(_06468_)
  );
  MUX2_X1 _14027_ (
    .A(mem_reg_wdata[4]),
    .B(_06468_),
    .S(_06442_),
    .Z(_06469_)
  );
  MUX2_X1 _14028_ (
    .A(wb_reg_wdata[4]),
    .B(_06469_),
    .S(_06433_),
    .Z(_00121_)
  );
  AND2_X1 _14029_ (
    .A1(wb_reg_wdata[5]),
    .A2(_06432_),
    .ZN(_06470_)
  );
  OR2_X1 _14030_ (
    .A1(_06463_),
    .A2(_06467_),
    .ZN(_06471_)
  );
  AND2_X1 _14031_ (
    .A1(mem_reg_inst[25]),
    .A2(_04031_),
    .ZN(_06472_)
  );
  AND2_X1 _14032_ (
    .A1(mem_reg_pc[5]),
    .A2(_06472_),
    .ZN(_06473_)
  );
  XOR2_X1 _14033_ (
    .A(mem_reg_pc[5]),
    .B(_06472_),
    .Z(_06474_)
  );
  AND2_X1 _14034_ (
    .A1(_06471_),
    .A2(_06474_),
    .ZN(_06475_)
  );
  XOR2_X1 _14035_ (
    .A(_06471_),
    .B(_06474_),
    .Z(_06476_)
  );
  OR2_X1 _14036_ (
    .A1(_06443_),
    .A2(_06476_),
    .ZN(_06477_)
  );
  OR2_X1 _14037_ (
    .A1(mem_reg_wdata[5]),
    .A2(_06442_),
    .ZN(_06478_)
  );
  AND2_X1 _14038_ (
    .A1(_06433_),
    .A2(_06478_),
    .ZN(_06479_)
  );
  AND2_X1 _14039_ (
    .A1(_06477_),
    .A2(_06479_),
    .ZN(_06480_)
  );
  OR2_X1 _14040_ (
    .A1(_06470_),
    .A2(_06480_),
    .ZN(_00122_)
  );
  AND2_X1 _14041_ (
    .A1(wb_reg_wdata[6]),
    .A2(_06432_),
    .ZN(_06481_)
  );
  OR2_X1 _14042_ (
    .A1(_06473_),
    .A2(_06475_),
    .ZN(_06482_)
  );
  AND2_X1 _14043_ (
    .A1(mem_reg_inst[26]),
    .A2(_04031_),
    .ZN(_06483_)
  );
  AND2_X1 _14044_ (
    .A1(mem_reg_pc[6]),
    .A2(_06483_),
    .ZN(_06484_)
  );
  XOR2_X1 _14045_ (
    .A(mem_reg_pc[6]),
    .B(_06483_),
    .Z(_06485_)
  );
  AND2_X1 _14046_ (
    .A1(_06482_),
    .A2(_06485_),
    .ZN(_06486_)
  );
  XOR2_X1 _14047_ (
    .A(_06482_),
    .B(_06485_),
    .Z(_06487_)
  );
  OR2_X1 _14048_ (
    .A1(_06443_),
    .A2(_06487_),
    .ZN(_06488_)
  );
  OR2_X1 _14049_ (
    .A1(mem_reg_wdata[6]),
    .A2(_06442_),
    .ZN(_06489_)
  );
  AND2_X1 _14050_ (
    .A1(_06433_),
    .A2(_06489_),
    .ZN(_06490_)
  );
  AND2_X1 _14051_ (
    .A1(_06488_),
    .A2(_06490_),
    .ZN(_06491_)
  );
  OR2_X1 _14052_ (
    .A1(_06481_),
    .A2(_06491_),
    .ZN(_00123_)
  );
  AND2_X1 _14053_ (
    .A1(wb_reg_wdata[7]),
    .A2(_06432_),
    .ZN(_06492_)
  );
  OR2_X1 _14054_ (
    .A1(_06484_),
    .A2(_06486_),
    .ZN(_06493_)
  );
  AND2_X1 _14055_ (
    .A1(mem_reg_inst[27]),
    .A2(_04031_),
    .ZN(_06494_)
  );
  AND2_X1 _14056_ (
    .A1(mem_reg_pc[7]),
    .A2(_06494_),
    .ZN(_06495_)
  );
  OR2_X1 _14057_ (
    .A1(mem_reg_pc[7]),
    .A2(_06494_),
    .ZN(_06496_)
  );
  XOR2_X1 _14058_ (
    .A(mem_reg_pc[7]),
    .B(_06494_),
    .Z(_06497_)
  );
  XOR2_X1 _14059_ (
    .A(_06493_),
    .B(_06497_),
    .Z(_06498_)
  );
  OR2_X1 _14060_ (
    .A1(_06443_),
    .A2(_06498_),
    .ZN(_06499_)
  );
  OR2_X1 _14061_ (
    .A1(mem_reg_wdata[7]),
    .A2(_06442_),
    .ZN(_06500_)
  );
  AND2_X1 _14062_ (
    .A1(_06433_),
    .A2(_06500_),
    .ZN(_06501_)
  );
  AND2_X1 _14063_ (
    .A1(_06499_),
    .A2(_06501_),
    .ZN(_06502_)
  );
  OR2_X1 _14064_ (
    .A1(_06492_),
    .A2(_06502_),
    .ZN(_00124_)
  );
  AND2_X1 _14065_ (
    .A1(mem_reg_inst[28]),
    .A2(_04031_),
    .ZN(_06503_)
  );
  AND2_X1 _14066_ (
    .A1(mem_reg_pc[8]),
    .A2(_06503_),
    .ZN(_06504_)
  );
  XOR2_X1 _14067_ (
    .A(mem_reg_pc[8]),
    .B(_06503_),
    .Z(_06505_)
  );
  OR2_X1 _14068_ (
    .A1(_06493_),
    .A2(_06495_),
    .ZN(_06506_)
  );
  AND2_X1 _14069_ (
    .A1(_06496_),
    .A2(_06506_),
    .ZN(_06507_)
  );
  AND2_X1 _14070_ (
    .A1(_06505_),
    .A2(_06507_),
    .ZN(_06508_)
  );
  XOR2_X1 _14071_ (
    .A(_06505_),
    .B(_06507_),
    .Z(_06509_)
  );
  MUX2_X1 _14072_ (
    .A(mem_reg_wdata[8]),
    .B(_06509_),
    .S(_06442_),
    .Z(_06510_)
  );
  MUX2_X1 _14073_ (
    .A(wb_reg_wdata[8]),
    .B(_06510_),
    .S(_06433_),
    .Z(_00125_)
  );
  AND2_X1 _14074_ (
    .A1(wb_reg_wdata[9]),
    .A2(_06432_),
    .ZN(_06511_)
  );
  OR2_X1 _14075_ (
    .A1(_06504_),
    .A2(_06508_),
    .ZN(_06512_)
  );
  AND2_X1 _14076_ (
    .A1(mem_reg_inst[29]),
    .A2(_04031_),
    .ZN(_06513_)
  );
  AND2_X1 _14077_ (
    .A1(mem_reg_pc[9]),
    .A2(_06513_),
    .ZN(_06514_)
  );
  OR2_X1 _14078_ (
    .A1(mem_reg_pc[9]),
    .A2(_06513_),
    .ZN(_06515_)
  );
  XOR2_X1 _14079_ (
    .A(mem_reg_pc[9]),
    .B(_06513_),
    .Z(_06516_)
  );
  XOR2_X1 _14080_ (
    .A(_06512_),
    .B(_06516_),
    .Z(_06517_)
  );
  OR2_X1 _14081_ (
    .A1(_06443_),
    .A2(_06517_),
    .ZN(_06518_)
  );
  OR2_X1 _14082_ (
    .A1(mem_reg_wdata[9]),
    .A2(_06442_),
    .ZN(_06519_)
  );
  AND2_X1 _14083_ (
    .A1(_06433_),
    .A2(_06519_),
    .ZN(_06520_)
  );
  AND2_X1 _14084_ (
    .A1(_06518_),
    .A2(_06520_),
    .ZN(_06521_)
  );
  OR2_X1 _14085_ (
    .A1(_06511_),
    .A2(_06521_),
    .ZN(_00126_)
  );
  AND2_X1 _14086_ (
    .A1(wb_reg_wdata[10]),
    .A2(_06432_),
    .ZN(_06522_)
  );
  AND2_X1 _14087_ (
    .A1(mem_reg_inst[30]),
    .A2(_04031_),
    .ZN(_06523_)
  );
  AND2_X1 _14088_ (
    .A1(mem_reg_pc[10]),
    .A2(_06523_),
    .ZN(_06524_)
  );
  XOR2_X1 _14089_ (
    .A(mem_reg_pc[10]),
    .B(_06523_),
    .Z(_06525_)
  );
  OR2_X1 _14090_ (
    .A1(_06512_),
    .A2(_06514_),
    .ZN(_06526_)
  );
  AND2_X1 _14091_ (
    .A1(_06515_),
    .A2(_06526_),
    .ZN(_06527_)
  );
  AND2_X1 _14092_ (
    .A1(_06525_),
    .A2(_06527_),
    .ZN(_06528_)
  );
  XOR2_X1 _14093_ (
    .A(_06525_),
    .B(_06527_),
    .Z(_06529_)
  );
  OR2_X1 _14094_ (
    .A1(_06443_),
    .A2(_06529_),
    .ZN(_06530_)
  );
  OR2_X1 _14095_ (
    .A1(mem_reg_wdata[10]),
    .A2(_06442_),
    .ZN(_06531_)
  );
  AND2_X1 _14096_ (
    .A1(_06433_),
    .A2(_06531_),
    .ZN(_06532_)
  );
  AND2_X1 _14097_ (
    .A1(_06530_),
    .A2(_06532_),
    .ZN(_06533_)
  );
  OR2_X1 _14098_ (
    .A1(_06522_),
    .A2(_06533_),
    .ZN(_00127_)
  );
  AND2_X1 _14099_ (
    .A1(wb_reg_wdata[11]),
    .A2(_06432_),
    .ZN(_06534_)
  );
  OR2_X1 _14100_ (
    .A1(_06524_),
    .A2(_06528_),
    .ZN(_06535_)
  );
  AND2_X1 _14101_ (
    .A1(mem_reg_inst[20]),
    .A2(mem_ctrl_jal),
    .ZN(_06536_)
  );
  MUX2_X1 _14102_ (
    .A(_06536_),
    .B(mem_reg_inst[7]),
    .S(_04030_),
    .Z(_06537_)
  );
  AND2_X1 _14103_ (
    .A1(mem_reg_pc[11]),
    .A2(_06537_),
    .ZN(_06538_)
  );
  OR2_X1 _14104_ (
    .A1(mem_reg_pc[11]),
    .A2(_06537_),
    .ZN(_06539_)
  );
  XOR2_X1 _14105_ (
    .A(mem_reg_pc[11]),
    .B(_06537_),
    .Z(_06540_)
  );
  XOR2_X1 _14106_ (
    .A(_06535_),
    .B(_06540_),
    .Z(_06541_)
  );
  OR2_X1 _14107_ (
    .A1(_06443_),
    .A2(_06541_),
    .ZN(_06542_)
  );
  OR2_X1 _14108_ (
    .A1(mem_reg_wdata[11]),
    .A2(_06442_),
    .ZN(_06543_)
  );
  AND2_X1 _14109_ (
    .A1(_06433_),
    .A2(_06543_),
    .ZN(_06544_)
  );
  AND2_X1 _14110_ (
    .A1(_06542_),
    .A2(_06544_),
    .ZN(_06545_)
  );
  OR2_X1 _14111_ (
    .A1(_06534_),
    .A2(_06545_),
    .ZN(_00128_)
  );
  AND2_X1 _14112_ (
    .A1(wb_reg_wdata[12]),
    .A2(_06432_),
    .ZN(_06546_)
  );
  AND2_X1 _14113_ (
    .A1(mem_reg_inst[12]),
    .A2(mem_ctrl_jal),
    .ZN(_06547_)
  );
  MUX2_X1 _14114_ (
    .A(_06547_),
    .B(mem_reg_inst[31]),
    .S(_04030_),
    .Z(_06548_)
  );
  AND2_X1 _14115_ (
    .A1(mem_reg_pc[12]),
    .A2(_06548_),
    .ZN(_06549_)
  );
  XOR2_X1 _14116_ (
    .A(mem_reg_pc[12]),
    .B(_06548_),
    .Z(_06550_)
  );
  OR2_X1 _14117_ (
    .A1(_06535_),
    .A2(_06538_),
    .ZN(_06551_)
  );
  AND2_X1 _14118_ (
    .A1(_06539_),
    .A2(_06551_),
    .ZN(_06552_)
  );
  AND2_X1 _14119_ (
    .A1(_06550_),
    .A2(_06552_),
    .ZN(_06553_)
  );
  XOR2_X1 _14120_ (
    .A(_06550_),
    .B(_06552_),
    .Z(_06554_)
  );
  OR2_X1 _14121_ (
    .A1(_06443_),
    .A2(_06554_),
    .ZN(_06555_)
  );
  OR2_X1 _14122_ (
    .A1(mem_reg_wdata[12]),
    .A2(_06442_),
    .ZN(_06556_)
  );
  AND2_X1 _14123_ (
    .A1(_06433_),
    .A2(_06556_),
    .ZN(_06557_)
  );
  AND2_X1 _14124_ (
    .A1(_06555_),
    .A2(_06557_),
    .ZN(_06558_)
  );
  OR2_X1 _14125_ (
    .A1(_06546_),
    .A2(_06558_),
    .ZN(_00129_)
  );
  AND2_X1 _14126_ (
    .A1(wb_reg_wdata[13]),
    .A2(_06432_),
    .ZN(_06559_)
  );
  OR2_X1 _14127_ (
    .A1(_06549_),
    .A2(_06553_),
    .ZN(_06560_)
  );
  AND2_X1 _14128_ (
    .A1(mem_reg_inst[13]),
    .A2(mem_ctrl_jal),
    .ZN(_06561_)
  );
  MUX2_X1 _14129_ (
    .A(_06561_),
    .B(mem_reg_inst[31]),
    .S(_04030_),
    .Z(_06562_)
  );
  AND2_X1 _14130_ (
    .A1(mem_reg_pc[13]),
    .A2(_06562_),
    .ZN(_06563_)
  );
  OR2_X1 _14131_ (
    .A1(mem_reg_pc[13]),
    .A2(_06562_),
    .ZN(_06564_)
  );
  XOR2_X1 _14132_ (
    .A(mem_reg_pc[13]),
    .B(_06562_),
    .Z(_06565_)
  );
  XOR2_X1 _14133_ (
    .A(_06560_),
    .B(_06565_),
    .Z(_06566_)
  );
  OR2_X1 _14134_ (
    .A1(_06443_),
    .A2(_06566_),
    .ZN(_06567_)
  );
  OR2_X1 _14135_ (
    .A1(mem_reg_wdata[13]),
    .A2(_06442_),
    .ZN(_06568_)
  );
  AND2_X1 _14136_ (
    .A1(_06433_),
    .A2(_06568_),
    .ZN(_06569_)
  );
  AND2_X1 _14137_ (
    .A1(_06567_),
    .A2(_06569_),
    .ZN(_06570_)
  );
  OR2_X1 _14138_ (
    .A1(_06559_),
    .A2(_06570_),
    .ZN(_00130_)
  );
  AND2_X1 _14139_ (
    .A1(wb_reg_wdata[14]),
    .A2(_06432_),
    .ZN(_06571_)
  );
  AND2_X1 _14140_ (
    .A1(mem_reg_inst[14]),
    .A2(mem_ctrl_jal),
    .ZN(_06572_)
  );
  MUX2_X1 _14141_ (
    .A(_06572_),
    .B(mem_reg_inst[31]),
    .S(_04030_),
    .Z(_06573_)
  );
  AND2_X1 _14142_ (
    .A1(mem_reg_pc[14]),
    .A2(_06573_),
    .ZN(_06574_)
  );
  XOR2_X1 _14143_ (
    .A(mem_reg_pc[14]),
    .B(_06573_),
    .Z(_06575_)
  );
  OR2_X1 _14144_ (
    .A1(_06560_),
    .A2(_06563_),
    .ZN(_06576_)
  );
  AND2_X1 _14145_ (
    .A1(_06564_),
    .A2(_06576_),
    .ZN(_06577_)
  );
  AND2_X1 _14146_ (
    .A1(_06575_),
    .A2(_06577_),
    .ZN(_06578_)
  );
  XOR2_X1 _14147_ (
    .A(_06575_),
    .B(_06577_),
    .Z(_06579_)
  );
  OR2_X1 _14148_ (
    .A1(_06443_),
    .A2(_06579_),
    .ZN(_06580_)
  );
  OR2_X1 _14149_ (
    .A1(mem_reg_wdata[14]),
    .A2(_06442_),
    .ZN(_06581_)
  );
  AND2_X1 _14150_ (
    .A1(_06433_),
    .A2(_06581_),
    .ZN(_06582_)
  );
  AND2_X1 _14151_ (
    .A1(_06580_),
    .A2(_06582_),
    .ZN(_06583_)
  );
  OR2_X1 _14152_ (
    .A1(_06571_),
    .A2(_06583_),
    .ZN(_00131_)
  );
  AND2_X1 _14153_ (
    .A1(wb_reg_wdata[15]),
    .A2(_06432_),
    .ZN(_06584_)
  );
  OR2_X1 _14154_ (
    .A1(_06574_),
    .A2(_06578_),
    .ZN(_06585_)
  );
  AND2_X1 _14155_ (
    .A1(mem_reg_inst[15]),
    .A2(mem_ctrl_jal),
    .ZN(_06586_)
  );
  MUX2_X1 _14156_ (
    .A(_06586_),
    .B(mem_reg_inst[31]),
    .S(_04030_),
    .Z(_06587_)
  );
  AND2_X1 _14157_ (
    .A1(mem_reg_pc[15]),
    .A2(_06587_),
    .ZN(_06588_)
  );
  OR2_X1 _14158_ (
    .A1(mem_reg_pc[15]),
    .A2(_06587_),
    .ZN(_06589_)
  );
  XOR2_X1 _14159_ (
    .A(mem_reg_pc[15]),
    .B(_06587_),
    .Z(_06590_)
  );
  XOR2_X1 _14160_ (
    .A(_06585_),
    .B(_06590_),
    .Z(_06591_)
  );
  OR2_X1 _14161_ (
    .A1(_06443_),
    .A2(_06591_),
    .ZN(_06592_)
  );
  OR2_X1 _14162_ (
    .A1(mem_reg_wdata[15]),
    .A2(_06442_),
    .ZN(_06593_)
  );
  AND2_X1 _14163_ (
    .A1(_06433_),
    .A2(_06593_),
    .ZN(_06594_)
  );
  AND2_X1 _14164_ (
    .A1(_06592_),
    .A2(_06594_),
    .ZN(_06595_)
  );
  OR2_X1 _14165_ (
    .A1(_06584_),
    .A2(_06595_),
    .ZN(_00132_)
  );
  AND2_X1 _14166_ (
    .A1(wb_reg_wdata[16]),
    .A2(_06432_),
    .ZN(_06596_)
  );
  AND2_X1 _14167_ (
    .A1(mem_reg_inst[16]),
    .A2(mem_ctrl_jal),
    .ZN(_06597_)
  );
  MUX2_X1 _14168_ (
    .A(_06597_),
    .B(mem_reg_inst[31]),
    .S(_04030_),
    .Z(_06598_)
  );
  AND2_X1 _14169_ (
    .A1(mem_reg_pc[16]),
    .A2(_06598_),
    .ZN(_06599_)
  );
  XOR2_X1 _14170_ (
    .A(mem_reg_pc[16]),
    .B(_06598_),
    .Z(_06600_)
  );
  OR2_X1 _14171_ (
    .A1(_06585_),
    .A2(_06588_),
    .ZN(_06601_)
  );
  AND2_X1 _14172_ (
    .A1(_06589_),
    .A2(_06601_),
    .ZN(_06602_)
  );
  AND2_X1 _14173_ (
    .A1(_06600_),
    .A2(_06602_),
    .ZN(_06603_)
  );
  XOR2_X1 _14174_ (
    .A(_06600_),
    .B(_06602_),
    .Z(_06604_)
  );
  OR2_X1 _14175_ (
    .A1(_06443_),
    .A2(_06604_),
    .ZN(_06605_)
  );
  OR2_X1 _14176_ (
    .A1(mem_reg_wdata[16]),
    .A2(_06442_),
    .ZN(_06606_)
  );
  AND2_X1 _14177_ (
    .A1(_06433_),
    .A2(_06606_),
    .ZN(_06607_)
  );
  AND2_X1 _14178_ (
    .A1(_06605_),
    .A2(_06607_),
    .ZN(_06608_)
  );
  OR2_X1 _14179_ (
    .A1(_06596_),
    .A2(_06608_),
    .ZN(_00133_)
  );
  AND2_X1 _14180_ (
    .A1(wb_reg_wdata[17]),
    .A2(_06432_),
    .ZN(_06609_)
  );
  OR2_X1 _14181_ (
    .A1(_06599_),
    .A2(_06603_),
    .ZN(_06610_)
  );
  AND2_X1 _14182_ (
    .A1(mem_reg_inst[17]),
    .A2(mem_ctrl_jal),
    .ZN(_06611_)
  );
  MUX2_X1 _14183_ (
    .A(_06611_),
    .B(mem_reg_inst[31]),
    .S(_04030_),
    .Z(_06612_)
  );
  AND2_X1 _14184_ (
    .A1(mem_reg_pc[17]),
    .A2(_06612_),
    .ZN(_06613_)
  );
  OR2_X1 _14185_ (
    .A1(mem_reg_pc[17]),
    .A2(_06612_),
    .ZN(_06614_)
  );
  XOR2_X1 _14186_ (
    .A(mem_reg_pc[17]),
    .B(_06612_),
    .Z(_06615_)
  );
  XOR2_X1 _14187_ (
    .A(_06610_),
    .B(_06615_),
    .Z(_06616_)
  );
  OR2_X1 _14188_ (
    .A1(_06443_),
    .A2(_06616_),
    .ZN(_06617_)
  );
  OR2_X1 _14189_ (
    .A1(mem_reg_wdata[17]),
    .A2(_06442_),
    .ZN(_06618_)
  );
  AND2_X1 _14190_ (
    .A1(_06433_),
    .A2(_06618_),
    .ZN(_06619_)
  );
  AND2_X1 _14191_ (
    .A1(_06617_),
    .A2(_06619_),
    .ZN(_06620_)
  );
  OR2_X1 _14192_ (
    .A1(_06609_),
    .A2(_06620_),
    .ZN(_00134_)
  );
  AND2_X1 _14193_ (
    .A1(wb_reg_wdata[18]),
    .A2(_06432_),
    .ZN(_06621_)
  );
  AND2_X1 _14194_ (
    .A1(mem_reg_inst[18]),
    .A2(mem_ctrl_jal),
    .ZN(_06622_)
  );
  MUX2_X1 _14195_ (
    .A(_06622_),
    .B(mem_reg_inst[31]),
    .S(_04030_),
    .Z(_06623_)
  );
  AND2_X1 _14196_ (
    .A1(mem_reg_pc[18]),
    .A2(_06623_),
    .ZN(_06624_)
  );
  XOR2_X1 _14197_ (
    .A(mem_reg_pc[18]),
    .B(_06623_),
    .Z(_06625_)
  );
  OR2_X1 _14198_ (
    .A1(_06610_),
    .A2(_06613_),
    .ZN(_06626_)
  );
  AND2_X1 _14199_ (
    .A1(_06614_),
    .A2(_06626_),
    .ZN(_06627_)
  );
  AND2_X1 _14200_ (
    .A1(_06625_),
    .A2(_06627_),
    .ZN(_06628_)
  );
  XOR2_X1 _14201_ (
    .A(_06625_),
    .B(_06627_),
    .Z(_06629_)
  );
  OR2_X1 _14202_ (
    .A1(_06443_),
    .A2(_06629_),
    .ZN(_06630_)
  );
  OR2_X1 _14203_ (
    .A1(mem_reg_wdata[18]),
    .A2(_06442_),
    .ZN(_06631_)
  );
  AND2_X1 _14204_ (
    .A1(_06433_),
    .A2(_06631_),
    .ZN(_06632_)
  );
  AND2_X1 _14205_ (
    .A1(_06630_),
    .A2(_06632_),
    .ZN(_06633_)
  );
  OR2_X1 _14206_ (
    .A1(_06621_),
    .A2(_06633_),
    .ZN(_00135_)
  );
  AND2_X1 _14207_ (
    .A1(wb_reg_wdata[19]),
    .A2(_06432_),
    .ZN(_06634_)
  );
  OR2_X1 _14208_ (
    .A1(_06624_),
    .A2(_06628_),
    .ZN(_06635_)
  );
  AND2_X1 _14209_ (
    .A1(mem_reg_inst[19]),
    .A2(mem_ctrl_jal),
    .ZN(_06636_)
  );
  MUX2_X1 _14210_ (
    .A(_06636_),
    .B(mem_reg_inst[31]),
    .S(_04030_),
    .Z(_06637_)
  );
  AND2_X1 _14211_ (
    .A1(mem_reg_pc[19]),
    .A2(_06637_),
    .ZN(_06638_)
  );
  OR2_X1 _14212_ (
    .A1(mem_reg_pc[19]),
    .A2(_06637_),
    .ZN(_06639_)
  );
  XOR2_X1 _14213_ (
    .A(mem_reg_pc[19]),
    .B(_06637_),
    .Z(_06640_)
  );
  XOR2_X1 _14214_ (
    .A(_06635_),
    .B(_06640_),
    .Z(_06641_)
  );
  OR2_X1 _14215_ (
    .A1(_06443_),
    .A2(_06641_),
    .ZN(_06642_)
  );
  OR2_X1 _14216_ (
    .A1(mem_reg_wdata[19]),
    .A2(_06442_),
    .ZN(_06643_)
  );
  AND2_X1 _14217_ (
    .A1(_06433_),
    .A2(_06643_),
    .ZN(_06644_)
  );
  AND2_X1 _14218_ (
    .A1(_06642_),
    .A2(_06644_),
    .ZN(_06645_)
  );
  OR2_X1 _14219_ (
    .A1(_06634_),
    .A2(_06645_),
    .ZN(_00136_)
  );
  AND2_X1 _14220_ (
    .A1(wb_reg_wdata[20]),
    .A2(_06432_),
    .ZN(_06646_)
  );
  AND2_X1 _14221_ (
    .A1(mem_reg_inst[31]),
    .A2(_04031_),
    .ZN(_06647_)
  );
  AND2_X1 _14222_ (
    .A1(mem_reg_pc[20]),
    .A2(_06647_),
    .ZN(_06648_)
  );
  XOR2_X1 _14223_ (
    .A(mem_reg_pc[20]),
    .B(_06647_),
    .Z(_06649_)
  );
  OR2_X1 _14224_ (
    .A1(_06635_),
    .A2(_06638_),
    .ZN(_06650_)
  );
  AND2_X1 _14225_ (
    .A1(_06639_),
    .A2(_06650_),
    .ZN(_06651_)
  );
  AND2_X1 _14226_ (
    .A1(_06649_),
    .A2(_06651_),
    .ZN(_06652_)
  );
  XOR2_X1 _14227_ (
    .A(_06649_),
    .B(_06651_),
    .Z(_06653_)
  );
  OR2_X1 _14228_ (
    .A1(_06443_),
    .A2(_06653_),
    .ZN(_06654_)
  );
  OR2_X1 _14229_ (
    .A1(mem_reg_wdata[20]),
    .A2(_06442_),
    .ZN(_06655_)
  );
  AND2_X1 _14230_ (
    .A1(_06433_),
    .A2(_06655_),
    .ZN(_06656_)
  );
  AND2_X1 _14231_ (
    .A1(_06654_),
    .A2(_06656_),
    .ZN(_06657_)
  );
  OR2_X1 _14232_ (
    .A1(_06646_),
    .A2(_06657_),
    .ZN(_00137_)
  );
  AND2_X1 _14233_ (
    .A1(wb_reg_wdata[21]),
    .A2(_06432_),
    .ZN(_06658_)
  );
  OR2_X1 _14234_ (
    .A1(_06648_),
    .A2(_06652_),
    .ZN(_06659_)
  );
  AND2_X1 _14235_ (
    .A1(mem_reg_pc[21]),
    .A2(_06647_),
    .ZN(_06660_)
  );
  XOR2_X1 _14236_ (
    .A(mem_reg_pc[21]),
    .B(_06647_),
    .Z(_06661_)
  );
  XOR2_X1 _14237_ (
    .A(_06659_),
    .B(_06661_),
    .Z(_06662_)
  );
  OR2_X1 _14238_ (
    .A1(_06443_),
    .A2(_06662_),
    .ZN(_06663_)
  );
  OR2_X1 _14239_ (
    .A1(mem_reg_wdata[21]),
    .A2(_06442_),
    .ZN(_06664_)
  );
  AND2_X1 _14240_ (
    .A1(_06433_),
    .A2(_06664_),
    .ZN(_06665_)
  );
  AND2_X1 _14241_ (
    .A1(_06663_),
    .A2(_06665_),
    .ZN(_06666_)
  );
  OR2_X1 _14242_ (
    .A1(_06658_),
    .A2(_06666_),
    .ZN(_00138_)
  );
  AND2_X1 _14243_ (
    .A1(wb_reg_wdata[22]),
    .A2(_06432_),
    .ZN(_06667_)
  );
  OR2_X1 _14244_ (
    .A1(_06648_),
    .A2(_06660_),
    .ZN(_06668_)
  );
  AND2_X1 _14245_ (
    .A1(_06652_),
    .A2(_06661_),
    .ZN(_06669_)
  );
  OR2_X1 _14246_ (
    .A1(_06668_),
    .A2(_06669_),
    .ZN(_06670_)
  );
  AND2_X1 _14247_ (
    .A1(mem_reg_pc[22]),
    .A2(_06647_),
    .ZN(_06671_)
  );
  XOR2_X1 _14248_ (
    .A(mem_reg_pc[22]),
    .B(_06647_),
    .Z(_06672_)
  );
  AND2_X1 _14249_ (
    .A1(_06670_),
    .A2(_06672_),
    .ZN(_06673_)
  );
  XOR2_X1 _14250_ (
    .A(_06670_),
    .B(_06672_),
    .Z(_06674_)
  );
  OR2_X1 _14251_ (
    .A1(_06443_),
    .A2(_06674_),
    .ZN(_06675_)
  );
  OR2_X1 _14252_ (
    .A1(mem_reg_wdata[22]),
    .A2(_06442_),
    .ZN(_06676_)
  );
  AND2_X1 _14253_ (
    .A1(_06433_),
    .A2(_06676_),
    .ZN(_06677_)
  );
  AND2_X1 _14254_ (
    .A1(_06675_),
    .A2(_06677_),
    .ZN(_06678_)
  );
  OR2_X1 _14255_ (
    .A1(_06667_),
    .A2(_06678_),
    .ZN(_00139_)
  );
  AND2_X1 _14256_ (
    .A1(wb_reg_wdata[23]),
    .A2(_06432_),
    .ZN(_06679_)
  );
  OR2_X1 _14257_ (
    .A1(_06671_),
    .A2(_06673_),
    .ZN(_06680_)
  );
  AND2_X1 _14258_ (
    .A1(mem_reg_pc[23]),
    .A2(_06647_),
    .ZN(_06681_)
  );
  XOR2_X1 _14259_ (
    .A(mem_reg_pc[23]),
    .B(_06647_),
    .Z(_06682_)
  );
  XOR2_X1 _14260_ (
    .A(_06680_),
    .B(_06682_),
    .Z(_06683_)
  );
  OR2_X1 _14261_ (
    .A1(_06443_),
    .A2(_06683_),
    .ZN(_06684_)
  );
  OR2_X1 _14262_ (
    .A1(mem_reg_wdata[23]),
    .A2(_06442_),
    .ZN(_06685_)
  );
  AND2_X1 _14263_ (
    .A1(_06433_),
    .A2(_06685_),
    .ZN(_06686_)
  );
  AND2_X1 _14264_ (
    .A1(_06684_),
    .A2(_06686_),
    .ZN(_06687_)
  );
  OR2_X1 _14265_ (
    .A1(_06679_),
    .A2(_06687_),
    .ZN(_00140_)
  );
  AND2_X1 _14266_ (
    .A1(wb_reg_wdata[24]),
    .A2(_06432_),
    .ZN(_06688_)
  );
  AND2_X1 _14267_ (
    .A1(_06672_),
    .A2(_06682_),
    .ZN(_06689_)
  );
  AND2_X1 _14268_ (
    .A1(_06669_),
    .A2(_06689_),
    .ZN(_06690_)
  );
  AND2_X1 _14269_ (
    .A1(_06668_),
    .A2(_06689_),
    .ZN(_06691_)
  );
  OR2_X1 _14270_ (
    .A1(_06671_),
    .A2(_06681_),
    .ZN(_06692_)
  );
  OR2_X1 _14271_ (
    .A1(_06691_),
    .A2(_06692_),
    .ZN(_06693_)
  );
  OR2_X1 _14272_ (
    .A1(_06690_),
    .A2(_06693_),
    .ZN(_06694_)
  );
  AND2_X1 _14273_ (
    .A1(mem_reg_pc[24]),
    .A2(_06647_),
    .ZN(_06695_)
  );
  XOR2_X1 _14274_ (
    .A(mem_reg_pc[24]),
    .B(_06647_),
    .Z(_06696_)
  );
  AND2_X1 _14275_ (
    .A1(_06694_),
    .A2(_06696_),
    .ZN(_06697_)
  );
  XOR2_X1 _14276_ (
    .A(_06694_),
    .B(_06696_),
    .Z(_06698_)
  );
  OR2_X1 _14277_ (
    .A1(_06443_),
    .A2(_06698_),
    .ZN(_06699_)
  );
  OR2_X1 _14278_ (
    .A1(mem_reg_wdata[24]),
    .A2(_06442_),
    .ZN(_06700_)
  );
  AND2_X1 _14279_ (
    .A1(_06433_),
    .A2(_06700_),
    .ZN(_06701_)
  );
  AND2_X1 _14280_ (
    .A1(_06699_),
    .A2(_06701_),
    .ZN(_06702_)
  );
  OR2_X1 _14281_ (
    .A1(_06688_),
    .A2(_06702_),
    .ZN(_00141_)
  );
  AND2_X1 _14282_ (
    .A1(wb_reg_wdata[25]),
    .A2(_06432_),
    .ZN(_06703_)
  );
  OR2_X1 _14283_ (
    .A1(_06695_),
    .A2(_06697_),
    .ZN(_06704_)
  );
  AND2_X1 _14284_ (
    .A1(mem_reg_pc[25]),
    .A2(_06647_),
    .ZN(_06705_)
  );
  XOR2_X1 _14285_ (
    .A(mem_reg_pc[25]),
    .B(_06647_),
    .Z(_06706_)
  );
  XOR2_X1 _14286_ (
    .A(_06704_),
    .B(_06706_),
    .Z(_06707_)
  );
  OR2_X1 _14287_ (
    .A1(_06443_),
    .A2(_06707_),
    .ZN(_06708_)
  );
  OR2_X1 _14288_ (
    .A1(mem_reg_wdata[25]),
    .A2(_06442_),
    .ZN(_06709_)
  );
  AND2_X1 _14289_ (
    .A1(_06433_),
    .A2(_06709_),
    .ZN(_06710_)
  );
  AND2_X1 _14290_ (
    .A1(_06708_),
    .A2(_06710_),
    .ZN(_06711_)
  );
  OR2_X1 _14291_ (
    .A1(_06703_),
    .A2(_06711_),
    .ZN(_00142_)
  );
  AND2_X1 _14292_ (
    .A1(wb_reg_wdata[26]),
    .A2(_06432_),
    .ZN(_06712_)
  );
  OR2_X1 _14293_ (
    .A1(_06695_),
    .A2(_06705_),
    .ZN(_06713_)
  );
  AND2_X1 _14294_ (
    .A1(_06697_),
    .A2(_06706_),
    .ZN(_06714_)
  );
  OR2_X1 _14295_ (
    .A1(_06713_),
    .A2(_06714_),
    .ZN(_06715_)
  );
  AND2_X1 _14296_ (
    .A1(mem_reg_pc[26]),
    .A2(_06647_),
    .ZN(_06716_)
  );
  XOR2_X1 _14297_ (
    .A(mem_reg_pc[26]),
    .B(_06647_),
    .Z(_06717_)
  );
  AND2_X1 _14298_ (
    .A1(_06715_),
    .A2(_06717_),
    .ZN(_06718_)
  );
  XOR2_X1 _14299_ (
    .A(_06715_),
    .B(_06717_),
    .Z(_06719_)
  );
  OR2_X1 _14300_ (
    .A1(_06443_),
    .A2(_06719_),
    .ZN(_06720_)
  );
  OR2_X1 _14301_ (
    .A1(mem_reg_wdata[26]),
    .A2(_06442_),
    .ZN(_06721_)
  );
  AND2_X1 _14302_ (
    .A1(_06433_),
    .A2(_06721_),
    .ZN(_06722_)
  );
  AND2_X1 _14303_ (
    .A1(_06720_),
    .A2(_06722_),
    .ZN(_06723_)
  );
  OR2_X1 _14304_ (
    .A1(_06712_),
    .A2(_06723_),
    .ZN(_00143_)
  );
  AND2_X1 _14305_ (
    .A1(wb_reg_wdata[27]),
    .A2(_06432_),
    .ZN(_06724_)
  );
  OR2_X1 _14306_ (
    .A1(_06716_),
    .A2(_06718_),
    .ZN(_06725_)
  );
  AND2_X1 _14307_ (
    .A1(mem_reg_pc[27]),
    .A2(_06647_),
    .ZN(_06726_)
  );
  XOR2_X1 _14308_ (
    .A(mem_reg_pc[27]),
    .B(_06647_),
    .Z(_06727_)
  );
  XOR2_X1 _14309_ (
    .A(_06725_),
    .B(_06727_),
    .Z(_06728_)
  );
  OR2_X1 _14310_ (
    .A1(_06443_),
    .A2(_06728_),
    .ZN(_06729_)
  );
  OR2_X1 _14311_ (
    .A1(mem_reg_wdata[27]),
    .A2(_06442_),
    .ZN(_06730_)
  );
  AND2_X1 _14312_ (
    .A1(_06433_),
    .A2(_06730_),
    .ZN(_06731_)
  );
  AND2_X1 _14313_ (
    .A1(_06729_),
    .A2(_06731_),
    .ZN(_06732_)
  );
  OR2_X1 _14314_ (
    .A1(_06724_),
    .A2(_06732_),
    .ZN(_00144_)
  );
  AND2_X1 _14315_ (
    .A1(wb_reg_wdata[28]),
    .A2(_06432_),
    .ZN(_06733_)
  );
  AND2_X1 _14316_ (
    .A1(_06717_),
    .A2(_06727_),
    .ZN(_06734_)
  );
  AND2_X1 _14317_ (
    .A1(_06714_),
    .A2(_06734_),
    .ZN(_06735_)
  );
  AND2_X1 _14318_ (
    .A1(_06713_),
    .A2(_06734_),
    .ZN(_06736_)
  );
  OR2_X1 _14319_ (
    .A1(_06716_),
    .A2(_06726_),
    .ZN(_06737_)
  );
  OR2_X1 _14320_ (
    .A1(_06736_),
    .A2(_06737_),
    .ZN(_06738_)
  );
  OR2_X1 _14321_ (
    .A1(_06735_),
    .A2(_06738_),
    .ZN(_06739_)
  );
  AND2_X1 _14322_ (
    .A1(mem_reg_pc[28]),
    .A2(_06647_),
    .ZN(_06740_)
  );
  XOR2_X1 _14323_ (
    .A(mem_reg_pc[28]),
    .B(_06647_),
    .Z(_06741_)
  );
  INV_X1 _14324_ (
    .A(_06741_),
    .ZN(_06742_)
  );
  AND2_X1 _14325_ (
    .A1(_06739_),
    .A2(_06741_),
    .ZN(_06743_)
  );
  XOR2_X1 _14326_ (
    .A(_06739_),
    .B(_06741_),
    .Z(_06744_)
  );
  XOR2_X1 _14327_ (
    .A(_06739_),
    .B(_06742_),
    .Z(_06745_)
  );
  OR2_X1 _14328_ (
    .A1(_06443_),
    .A2(_06744_),
    .ZN(_06746_)
  );
  OR2_X1 _14329_ (
    .A1(mem_reg_wdata[28]),
    .A2(_06442_),
    .ZN(_06747_)
  );
  AND2_X1 _14330_ (
    .A1(_06433_),
    .A2(_06747_),
    .ZN(_06748_)
  );
  AND2_X1 _14331_ (
    .A1(_06746_),
    .A2(_06748_),
    .ZN(_06749_)
  );
  OR2_X1 _14332_ (
    .A1(_06733_),
    .A2(_06749_),
    .ZN(_00145_)
  );
  AND2_X1 _14333_ (
    .A1(wb_reg_wdata[29]),
    .A2(_06432_),
    .ZN(_06750_)
  );
  OR2_X1 _14334_ (
    .A1(_06740_),
    .A2(_06743_),
    .ZN(_06751_)
  );
  AND2_X1 _14335_ (
    .A1(mem_reg_pc[29]),
    .A2(_06647_),
    .ZN(_06752_)
  );
  OR2_X1 _14336_ (
    .A1(mem_reg_pc[29]),
    .A2(_06647_),
    .ZN(_06753_)
  );
  XOR2_X1 _14337_ (
    .A(mem_reg_pc[29]),
    .B(_06647_),
    .Z(_06754_)
  );
  XOR2_X1 _14338_ (
    .A(_06751_),
    .B(_06754_),
    .Z(_06755_)
  );
  OR2_X1 _14339_ (
    .A1(_06443_),
    .A2(_06755_),
    .ZN(_06756_)
  );
  OR2_X1 _14340_ (
    .A1(mem_reg_wdata[29]),
    .A2(_06442_),
    .ZN(_06757_)
  );
  AND2_X1 _14341_ (
    .A1(_06433_),
    .A2(_06757_),
    .ZN(_06758_)
  );
  AND2_X1 _14342_ (
    .A1(_06756_),
    .A2(_06758_),
    .ZN(_06759_)
  );
  OR2_X1 _14343_ (
    .A1(_06750_),
    .A2(_06759_),
    .ZN(_00146_)
  );
  AND2_X1 _14344_ (
    .A1(wb_reg_wdata[30]),
    .A2(_06432_),
    .ZN(_06760_)
  );
  AND2_X1 _14345_ (
    .A1(mem_reg_pc[30]),
    .A2(_06647_),
    .ZN(_06761_)
  );
  XOR2_X1 _14346_ (
    .A(mem_reg_pc[30]),
    .B(_06647_),
    .Z(_06762_)
  );
  AND2_X1 _14347_ (
    .A1(_06751_),
    .A2(_06753_),
    .ZN(_06763_)
  );
  OR2_X1 _14348_ (
    .A1(_06752_),
    .A2(_06763_),
    .ZN(_06764_)
  );
  AND2_X1 _14349_ (
    .A1(_06762_),
    .A2(_06764_),
    .ZN(_06765_)
  );
  XOR2_X1 _14350_ (
    .A(_06762_),
    .B(_06764_),
    .Z(_06766_)
  );
  OR2_X1 _14351_ (
    .A1(_06443_),
    .A2(_06766_),
    .ZN(_06767_)
  );
  OR2_X1 _14352_ (
    .A1(mem_reg_wdata[30]),
    .A2(_06442_),
    .ZN(_06768_)
  );
  AND2_X1 _14353_ (
    .A1(_06433_),
    .A2(_06768_),
    .ZN(_06769_)
  );
  AND2_X1 _14354_ (
    .A1(_06767_),
    .A2(_06769_),
    .ZN(_06770_)
  );
  OR2_X1 _14355_ (
    .A1(_06760_),
    .A2(_06770_),
    .ZN(_00147_)
  );
  AND2_X1 _14356_ (
    .A1(wb_reg_wdata[31]),
    .A2(_06432_),
    .ZN(_06771_)
  );
  OR2_X1 _14357_ (
    .A1(_06761_),
    .A2(_06765_),
    .ZN(_06772_)
  );
  XOR2_X1 _14358_ (
    .A(mem_reg_pc[31]),
    .B(_06647_),
    .Z(_06773_)
  );
  XOR2_X1 _14359_ (
    .A(_06772_),
    .B(_06773_),
    .Z(_06774_)
  );
  OR2_X1 _14360_ (
    .A1(_06443_),
    .A2(_06774_),
    .ZN(_06775_)
  );
  OR2_X1 _14361_ (
    .A1(mem_reg_wdata[31]),
    .A2(_06442_),
    .ZN(_06776_)
  );
  AND2_X1 _14362_ (
    .A1(_06433_),
    .A2(_06776_),
    .ZN(_06777_)
  );
  AND2_X1 _14363_ (
    .A1(_06775_),
    .A2(_06777_),
    .ZN(_06778_)
  );
  OR2_X1 _14364_ (
    .A1(_06771_),
    .A2(_06778_),
    .ZN(_00148_)
  );
  OR2_X1 _14365_ (
    .A1(_03807_),
    .A2(_06428_),
    .ZN(_06779_)
  );
  INV_X1 _14366_ (
    .A(_06779_),
    .ZN(_06780_)
  );
  AND2_X1 _14367_ (
    .A1(_ex_reg_valid_T),
    .A2(_06780_),
    .ZN(_06781_)
  );
  XOR2_X1 _14368_ (
    .A(_03064_),
    .B(_04054_),
    .Z(_06782_)
  );
  XOR2_X1 _14369_ (
    .A(ibuf_io_inst_0_bits_inst_rs2[2]),
    .B(_04052_),
    .Z(_06783_)
  );
  AND2_X1 _14370_ (
    .A1(_06782_),
    .A2(_06783_),
    .ZN(_06784_)
  );
  XOR2_X1 _14371_ (
    .A(_03049_),
    .B(_04047_),
    .Z(_06785_)
  );
  XOR2_X1 _14372_ (
    .A(_03048_),
    .B(_04049_),
    .Z(_06786_)
  );
  AND2_X1 _14373_ (
    .A1(_06785_),
    .A2(_06786_),
    .ZN(_06787_)
  );
  XOR2_X1 _14374_ (
    .A(_03051_),
    .B(_04056_),
    .Z(_06788_)
  );
  AND2_X1 _14375_ (
    .A1(_06787_),
    .A2(_06788_),
    .ZN(_06789_)
  );
  AND2_X1 _14376_ (
    .A1(_06784_),
    .A2(_06789_),
    .ZN(_06790_)
  );
  AND2_X1 _14377_ (
    .A1(_04062_),
    .A2(_06790_),
    .ZN(_06791_)
  );
  INV_X1 _14378_ (
    .A(_06791_),
    .ZN(_06792_)
  );
  MUX2_X1 _14379_ (
    .A(\rf[7] [2]),
    .B(\rf[3] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06793_)
  );
  AND2_X1 _14380_ (
    .A1(_03049_),
    .A2(_06793_),
    .ZN(_06794_)
  );
  MUX2_X1 _14381_ (
    .A(\rf[5] [2]),
    .B(\rf[1] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06795_)
  );
  AND2_X1 _14382_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_06795_),
    .ZN(_06796_)
  );
  OR2_X1 _14383_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_06796_),
    .ZN(_06797_)
  );
  OR2_X1 _14384_ (
    .A1(_06794_),
    .A2(_06797_),
    .ZN(_06798_)
  );
  MUX2_X1 _14385_ (
    .A(\rf[6] [2]),
    .B(\rf[2] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06799_)
  );
  AND2_X1 _14386_ (
    .A1(_03049_),
    .A2(_06799_),
    .ZN(_06800_)
  );
  MUX2_X1 _14387_ (
    .A(\rf[4] [2]),
    .B(\rf[0] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06801_)
  );
  AND2_X1 _14388_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_06801_),
    .ZN(_06802_)
  );
  OR2_X1 _14389_ (
    .A1(_03048_),
    .A2(_06802_),
    .ZN(_06803_)
  );
  OR2_X1 _14390_ (
    .A1(_06800_),
    .A2(_06803_),
    .ZN(_06804_)
  );
  AND2_X1 _14391_ (
    .A1(_06798_),
    .A2(_06804_),
    .ZN(_06805_)
  );
  AND2_X1 _14392_ (
    .A1(\rf[14] [2]),
    .A2(_03049_),
    .ZN(_06806_)
  );
  AND2_X1 _14393_ (
    .A1(\rf[12] [2]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_06807_)
  );
  OR2_X1 _14394_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[2]),
    .A2(_06807_),
    .ZN(_06808_)
  );
  OR2_X1 _14395_ (
    .A1(_06806_),
    .A2(_06808_),
    .ZN(_06809_)
  );
  AND2_X1 _14396_ (
    .A1(\rf[10] [2]),
    .A2(_03049_),
    .ZN(_06810_)
  );
  AND2_X1 _14397_ (
    .A1(\rf[8] [2]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_06811_)
  );
  OR2_X1 _14398_ (
    .A1(_03050_),
    .A2(_06811_),
    .ZN(_06812_)
  );
  OR2_X1 _14399_ (
    .A1(_06810_),
    .A2(_06812_),
    .ZN(_06813_)
  );
  AND2_X1 _14400_ (
    .A1(_06809_),
    .A2(_06813_),
    .ZN(_06814_)
  );
  AND2_X1 _14401_ (
    .A1(\rf[15] [2]),
    .A2(_03049_),
    .ZN(_06815_)
  );
  AND2_X1 _14402_ (
    .A1(\rf[13] [2]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_06816_)
  );
  OR2_X1 _14403_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[2]),
    .A2(_06816_),
    .ZN(_06817_)
  );
  OR2_X1 _14404_ (
    .A1(_06815_),
    .A2(_06817_),
    .ZN(_06818_)
  );
  AND2_X1 _14405_ (
    .A1(\rf[11] [2]),
    .A2(_03049_),
    .ZN(_06819_)
  );
  AND2_X1 _14406_ (
    .A1(\rf[9] [2]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_06820_)
  );
  OR2_X1 _14407_ (
    .A1(_03050_),
    .A2(_06820_),
    .ZN(_06821_)
  );
  OR2_X1 _14408_ (
    .A1(_06819_),
    .A2(_06821_),
    .ZN(_06822_)
  );
  AND2_X1 _14409_ (
    .A1(_06818_),
    .A2(_06822_),
    .ZN(_06823_)
  );
  MUX2_X1 _14410_ (
    .A(_06814_),
    .B(_06823_),
    .S(_03048_),
    .Z(_06824_)
  );
  MUX2_X1 _14411_ (
    .A(_06805_),
    .B(_06824_),
    .S(_03051_),
    .Z(_06825_)
  );
  AND2_X1 _14412_ (
    .A1(\rf[26] [2]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_06826_)
  );
  AND2_X1 _14413_ (
    .A1(\rf[30] [2]),
    .A2(_03050_),
    .ZN(_06827_)
  );
  OR2_X1 _14414_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_06827_),
    .ZN(_06828_)
  );
  OR2_X1 _14415_ (
    .A1(_06826_),
    .A2(_06828_),
    .ZN(_06829_)
  );
  AND2_X1 _14416_ (
    .A1(\rf[24] [2]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_06830_)
  );
  AND2_X1 _14417_ (
    .A1(\rf[28] [2]),
    .A2(_03050_),
    .ZN(_06831_)
  );
  OR2_X1 _14418_ (
    .A1(_03049_),
    .A2(_06831_),
    .ZN(_06832_)
  );
  OR2_X1 _14419_ (
    .A1(_06830_),
    .A2(_06832_),
    .ZN(_06833_)
  );
  AND2_X1 _14420_ (
    .A1(_06829_),
    .A2(_06833_),
    .ZN(_06834_)
  );
  MUX2_X1 _14421_ (
    .A(\rf[29] [2]),
    .B(\rf[25] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06835_)
  );
  AND2_X1 _14422_ (
    .A1(\rf[27] [2]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_06836_)
  );
  MUX2_X1 _14423_ (
    .A(_06835_),
    .B(_06836_),
    .S(_03049_),
    .Z(_06837_)
  );
  MUX2_X1 _14424_ (
    .A(_06834_),
    .B(_06837_),
    .S(_03048_),
    .Z(_06838_)
  );
  OR2_X1 _14425_ (
    .A1(\rf[20] [2]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_06839_)
  );
  OR2_X1 _14426_ (
    .A1(\rf[16] [2]),
    .A2(_03050_),
    .ZN(_06840_)
  );
  AND2_X1 _14427_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_06840_),
    .ZN(_06841_)
  );
  AND2_X1 _14428_ (
    .A1(_06839_),
    .A2(_06841_),
    .ZN(_06842_)
  );
  MUX2_X1 _14429_ (
    .A(\rf[22] [2]),
    .B(\rf[18] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06843_)
  );
  AND2_X1 _14430_ (
    .A1(_03049_),
    .A2(_06843_),
    .ZN(_06844_)
  );
  OR2_X1 _14431_ (
    .A1(_03048_),
    .A2(_06844_),
    .ZN(_06845_)
  );
  OR2_X1 _14432_ (
    .A1(_06842_),
    .A2(_06845_),
    .ZN(_06846_)
  );
  OR2_X1 _14433_ (
    .A1(\rf[17] [2]),
    .A2(_03050_),
    .ZN(_06847_)
  );
  OR2_X1 _14434_ (
    .A1(\rf[21] [2]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_06848_)
  );
  AND2_X1 _14435_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_06848_),
    .ZN(_06849_)
  );
  AND2_X1 _14436_ (
    .A1(_06847_),
    .A2(_06849_),
    .ZN(_06850_)
  );
  MUX2_X1 _14437_ (
    .A(\rf[23] [2]),
    .B(\rf[19] [2]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06851_)
  );
  AND2_X1 _14438_ (
    .A1(_03049_),
    .A2(_06851_),
    .ZN(_06852_)
  );
  OR2_X1 _14439_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_06852_),
    .ZN(_06853_)
  );
  OR2_X1 _14440_ (
    .A1(_06850_),
    .A2(_06853_),
    .ZN(_06854_)
  );
  AND2_X1 _14441_ (
    .A1(_06846_),
    .A2(_06854_),
    .ZN(_06855_)
  );
  MUX2_X1 _14442_ (
    .A(_06838_),
    .B(_06855_),
    .S(ibuf_io_inst_0_bits_inst_rs2[3]),
    .Z(_06856_)
  );
  MUX2_X1 _14443_ (
    .A(_06825_),
    .B(_06856_),
    .S(_03064_),
    .Z(_06857_)
  );
  MUX2_X1 _14444_ (
    .A(_06857_),
    .B(_04080_),
    .S(_06791_),
    .Z(_06858_)
  );
  MUX2_X1 _14445_ (
    .A(ex_reg_rs_msb_1[0]),
    .B(_06858_),
    .S(_06781_),
    .Z(_00149_)
  );
  MUX2_X1 _14446_ (
    .A(\rf[3] [3]),
    .B(\rf[2] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_06859_)
  );
  MUX2_X1 _14447_ (
    .A(\rf[7] [3]),
    .B(\rf[6] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_06860_)
  );
  MUX2_X1 _14448_ (
    .A(_06859_),
    .B(_06860_),
    .S(_03050_),
    .Z(_06861_)
  );
  OR2_X1 _14449_ (
    .A1(_03051_),
    .A2(_06861_),
    .ZN(_06862_)
  );
  OR2_X1 _14450_ (
    .A1(_03048_),
    .A2(ibuf_io_inst_0_bits_inst_rs2[3]),
    .ZN(_06863_)
  );
  MUX2_X1 _14451_ (
    .A(\rf[14] [3]),
    .B(\rf[10] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06864_)
  );
  OR2_X1 _14452_ (
    .A1(_06863_),
    .A2(_06864_),
    .ZN(_06865_)
  );
  MUX2_X1 _14453_ (
    .A(\rf[15] [3]),
    .B(\rf[11] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06866_)
  );
  OR2_X1 _14454_ (
    .A1(_03808_),
    .A2(_06866_),
    .ZN(_06867_)
  );
  AND2_X1 _14455_ (
    .A1(_03049_),
    .A2(_06867_),
    .ZN(_06868_)
  );
  AND2_X1 _14456_ (
    .A1(_06865_),
    .A2(_06868_),
    .ZN(_06869_)
  );
  AND2_X1 _14457_ (
    .A1(_06862_),
    .A2(_06869_),
    .ZN(_06870_)
  );
  MUX2_X1 _14458_ (
    .A(\rf[1] [3]),
    .B(\rf[0] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_06871_)
  );
  MUX2_X1 _14459_ (
    .A(\rf[5] [3]),
    .B(\rf[4] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_06872_)
  );
  MUX2_X1 _14460_ (
    .A(_06871_),
    .B(_06872_),
    .S(_03050_),
    .Z(_06873_)
  );
  OR2_X1 _14461_ (
    .A1(_03051_),
    .A2(_06873_),
    .ZN(_06874_)
  );
  MUX2_X1 _14462_ (
    .A(\rf[12] [3]),
    .B(\rf[8] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06875_)
  );
  OR2_X1 _14463_ (
    .A1(_06863_),
    .A2(_06875_),
    .ZN(_06876_)
  );
  MUX2_X1 _14464_ (
    .A(\rf[13] [3]),
    .B(\rf[9] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06877_)
  );
  OR2_X1 _14465_ (
    .A1(_03808_),
    .A2(_06877_),
    .ZN(_06878_)
  );
  AND2_X1 _14466_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_06878_),
    .ZN(_06879_)
  );
  AND2_X1 _14467_ (
    .A1(_06876_),
    .A2(_06879_),
    .ZN(_06880_)
  );
  AND2_X1 _14468_ (
    .A1(_06874_),
    .A2(_06880_),
    .ZN(_06881_)
  );
  OR2_X1 _14469_ (
    .A1(_06870_),
    .A2(_06881_),
    .ZN(_06882_)
  );
  OR2_X1 _14470_ (
    .A1(\rf[17] [3]),
    .A2(_03050_),
    .ZN(_06883_)
  );
  OR2_X1 _14471_ (
    .A1(\rf[21] [3]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_06884_)
  );
  AND2_X1 _14472_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_06884_),
    .ZN(_06885_)
  );
  AND2_X1 _14473_ (
    .A1(_06883_),
    .A2(_06885_),
    .ZN(_06886_)
  );
  MUX2_X1 _14474_ (
    .A(\rf[23] [3]),
    .B(\rf[19] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06887_)
  );
  AND2_X1 _14475_ (
    .A1(_03049_),
    .A2(_06887_),
    .ZN(_06888_)
  );
  OR2_X1 _14476_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_06888_),
    .ZN(_06889_)
  );
  OR2_X1 _14477_ (
    .A1(_06886_),
    .A2(_06889_),
    .ZN(_06890_)
  );
  OR2_X1 _14478_ (
    .A1(\rf[20] [3]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_06891_)
  );
  OR2_X1 _14479_ (
    .A1(\rf[16] [3]),
    .A2(_03050_),
    .ZN(_06892_)
  );
  AND2_X1 _14480_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_06892_),
    .ZN(_06893_)
  );
  AND2_X1 _14481_ (
    .A1(_06891_),
    .A2(_06893_),
    .ZN(_06894_)
  );
  MUX2_X1 _14482_ (
    .A(\rf[22] [3]),
    .B(\rf[18] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06895_)
  );
  AND2_X1 _14483_ (
    .A1(_03049_),
    .A2(_06895_),
    .ZN(_06896_)
  );
  OR2_X1 _14484_ (
    .A1(_03048_),
    .A2(_06896_),
    .ZN(_06897_)
  );
  OR2_X1 _14485_ (
    .A1(_06894_),
    .A2(_06897_),
    .ZN(_06898_)
  );
  AND2_X1 _14486_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_06890_),
    .ZN(_06899_)
  );
  AND2_X1 _14487_ (
    .A1(_06898_),
    .A2(_06899_),
    .ZN(_06900_)
  );
  OR2_X1 _14488_ (
    .A1(\rf[28] [3]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_06901_)
  );
  OR2_X1 _14489_ (
    .A1(\rf[24] [3]),
    .A2(_03050_),
    .ZN(_06902_)
  );
  AND2_X1 _14490_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_06901_),
    .ZN(_06903_)
  );
  AND2_X1 _14491_ (
    .A1(_06902_),
    .A2(_06903_),
    .ZN(_06904_)
  );
  MUX2_X1 _14492_ (
    .A(\rf[30] [3]),
    .B(\rf[26] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06905_)
  );
  AND2_X1 _14493_ (
    .A1(_03049_),
    .A2(_06905_),
    .ZN(_06906_)
  );
  OR2_X1 _14494_ (
    .A1(_03048_),
    .A2(_06906_),
    .ZN(_06907_)
  );
  OR2_X1 _14495_ (
    .A1(_06904_),
    .A2(_06907_),
    .ZN(_06908_)
  );
  MUX2_X1 _14496_ (
    .A(\rf[29] [3]),
    .B(\rf[25] [3]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06909_)
  );
  AND2_X1 _14497_ (
    .A1(\rf[27] [3]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_06910_)
  );
  MUX2_X1 _14498_ (
    .A(_06909_),
    .B(_06910_),
    .S(_03049_),
    .Z(_06911_)
  );
  OR2_X1 _14499_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_06911_),
    .ZN(_06912_)
  );
  AND2_X1 _14500_ (
    .A1(_03051_),
    .A2(_06912_),
    .ZN(_06913_)
  );
  AND2_X1 _14501_ (
    .A1(_06908_),
    .A2(_06913_),
    .ZN(_06914_)
  );
  OR2_X1 _14502_ (
    .A1(_06900_),
    .A2(_06914_),
    .ZN(_06915_)
  );
  MUX2_X1 _14503_ (
    .A(_06882_),
    .B(_06915_),
    .S(_03064_),
    .Z(_06916_)
  );
  MUX2_X1 _14504_ (
    .A(_06916_),
    .B(_04150_),
    .S(_06791_),
    .Z(_06917_)
  );
  MUX2_X1 _14505_ (
    .A(ex_reg_rs_msb_1[1]),
    .B(_06917_),
    .S(_06781_),
    .Z(_00150_)
  );
  MUX2_X1 _14506_ (
    .A(\rf[3] [4]),
    .B(\rf[2] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_06918_)
  );
  MUX2_X1 _14507_ (
    .A(\rf[7] [4]),
    .B(\rf[6] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_06919_)
  );
  MUX2_X1 _14508_ (
    .A(_06918_),
    .B(_06919_),
    .S(_03050_),
    .Z(_06920_)
  );
  OR2_X1 _14509_ (
    .A1(_03051_),
    .A2(_06920_),
    .ZN(_06921_)
  );
  MUX2_X1 _14510_ (
    .A(\rf[14] [4]),
    .B(\rf[10] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06922_)
  );
  OR2_X1 _14511_ (
    .A1(_06863_),
    .A2(_06922_),
    .ZN(_06923_)
  );
  MUX2_X1 _14512_ (
    .A(\rf[15] [4]),
    .B(\rf[11] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06924_)
  );
  OR2_X1 _14513_ (
    .A1(_03808_),
    .A2(_06924_),
    .ZN(_06925_)
  );
  AND2_X1 _14514_ (
    .A1(_03049_),
    .A2(_06925_),
    .ZN(_06926_)
  );
  AND2_X1 _14515_ (
    .A1(_06923_),
    .A2(_06926_),
    .ZN(_06927_)
  );
  AND2_X1 _14516_ (
    .A1(_06921_),
    .A2(_06927_),
    .ZN(_06928_)
  );
  MUX2_X1 _14517_ (
    .A(\rf[1] [4]),
    .B(\rf[0] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_06929_)
  );
  MUX2_X1 _14518_ (
    .A(\rf[5] [4]),
    .B(\rf[4] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_06930_)
  );
  MUX2_X1 _14519_ (
    .A(_06929_),
    .B(_06930_),
    .S(_03050_),
    .Z(_06931_)
  );
  OR2_X1 _14520_ (
    .A1(_03051_),
    .A2(_06931_),
    .ZN(_06932_)
  );
  MUX2_X1 _14521_ (
    .A(\rf[12] [4]),
    .B(\rf[8] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06933_)
  );
  OR2_X1 _14522_ (
    .A1(_06863_),
    .A2(_06933_),
    .ZN(_06934_)
  );
  MUX2_X1 _14523_ (
    .A(\rf[13] [4]),
    .B(\rf[9] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06935_)
  );
  OR2_X1 _14524_ (
    .A1(_03808_),
    .A2(_06935_),
    .ZN(_06936_)
  );
  AND2_X1 _14525_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_06936_),
    .ZN(_06937_)
  );
  AND2_X1 _14526_ (
    .A1(_06934_),
    .A2(_06937_),
    .ZN(_06938_)
  );
  AND2_X1 _14527_ (
    .A1(_06932_),
    .A2(_06938_),
    .ZN(_06939_)
  );
  OR2_X1 _14528_ (
    .A1(_06928_),
    .A2(_06939_),
    .ZN(_06940_)
  );
  OR2_X1 _14529_ (
    .A1(\rf[17] [4]),
    .A2(_03050_),
    .ZN(_06941_)
  );
  OR2_X1 _14530_ (
    .A1(\rf[21] [4]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_06942_)
  );
  AND2_X1 _14531_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_06942_),
    .ZN(_06943_)
  );
  AND2_X1 _14532_ (
    .A1(_06941_),
    .A2(_06943_),
    .ZN(_06944_)
  );
  MUX2_X1 _14533_ (
    .A(\rf[23] [4]),
    .B(\rf[19] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06945_)
  );
  AND2_X1 _14534_ (
    .A1(_03049_),
    .A2(_06945_),
    .ZN(_06946_)
  );
  OR2_X1 _14535_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_06946_),
    .ZN(_06947_)
  );
  OR2_X1 _14536_ (
    .A1(_06944_),
    .A2(_06947_),
    .ZN(_06948_)
  );
  OR2_X1 _14537_ (
    .A1(\rf[20] [4]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_06949_)
  );
  OR2_X1 _14538_ (
    .A1(\rf[16] [4]),
    .A2(_03050_),
    .ZN(_06950_)
  );
  AND2_X1 _14539_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_06950_),
    .ZN(_06951_)
  );
  AND2_X1 _14540_ (
    .A1(_06949_),
    .A2(_06951_),
    .ZN(_06952_)
  );
  MUX2_X1 _14541_ (
    .A(\rf[22] [4]),
    .B(\rf[18] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06953_)
  );
  AND2_X1 _14542_ (
    .A1(_03049_),
    .A2(_06953_),
    .ZN(_06954_)
  );
  OR2_X1 _14543_ (
    .A1(_03048_),
    .A2(_06954_),
    .ZN(_06955_)
  );
  OR2_X1 _14544_ (
    .A1(_06952_),
    .A2(_06955_),
    .ZN(_06956_)
  );
  AND2_X1 _14545_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_06948_),
    .ZN(_06957_)
  );
  AND2_X1 _14546_ (
    .A1(_06956_),
    .A2(_06957_),
    .ZN(_06958_)
  );
  OR2_X1 _14547_ (
    .A1(\rf[28] [4]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_06959_)
  );
  OR2_X1 _14548_ (
    .A1(\rf[24] [4]),
    .A2(_03050_),
    .ZN(_06960_)
  );
  AND2_X1 _14549_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_06959_),
    .ZN(_06961_)
  );
  AND2_X1 _14550_ (
    .A1(_06960_),
    .A2(_06961_),
    .ZN(_06962_)
  );
  MUX2_X1 _14551_ (
    .A(\rf[30] [4]),
    .B(\rf[26] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06963_)
  );
  AND2_X1 _14552_ (
    .A1(_03049_),
    .A2(_06963_),
    .ZN(_06964_)
  );
  OR2_X1 _14553_ (
    .A1(_03048_),
    .A2(_06964_),
    .ZN(_06965_)
  );
  OR2_X1 _14554_ (
    .A1(_06962_),
    .A2(_06965_),
    .ZN(_06966_)
  );
  MUX2_X1 _14555_ (
    .A(\rf[29] [4]),
    .B(\rf[25] [4]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06967_)
  );
  AND2_X1 _14556_ (
    .A1(\rf[27] [4]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_06968_)
  );
  MUX2_X1 _14557_ (
    .A(_06967_),
    .B(_06968_),
    .S(_03049_),
    .Z(_06969_)
  );
  OR2_X1 _14558_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_06969_),
    .ZN(_06970_)
  );
  AND2_X1 _14559_ (
    .A1(_03051_),
    .A2(_06970_),
    .ZN(_06971_)
  );
  AND2_X1 _14560_ (
    .A1(_06966_),
    .A2(_06971_),
    .ZN(_06972_)
  );
  OR2_X1 _14561_ (
    .A1(_06958_),
    .A2(_06972_),
    .ZN(_06973_)
  );
  MUX2_X1 _14562_ (
    .A(_06940_),
    .B(_06973_),
    .S(_03064_),
    .Z(_06974_)
  );
  MUX2_X1 _14563_ (
    .A(_06974_),
    .B(_04233_),
    .S(_06791_),
    .Z(_06975_)
  );
  MUX2_X1 _14564_ (
    .A(ex_reg_rs_msb_1[2]),
    .B(_06975_),
    .S(_06781_),
    .Z(_00151_)
  );
  MUX2_X1 _14565_ (
    .A(\rf[7] [5]),
    .B(\rf[3] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06976_)
  );
  AND2_X1 _14566_ (
    .A1(_03049_),
    .A2(_06976_),
    .ZN(_06977_)
  );
  MUX2_X1 _14567_ (
    .A(\rf[5] [5]),
    .B(\rf[1] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06978_)
  );
  AND2_X1 _14568_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_06978_),
    .ZN(_06979_)
  );
  OR2_X1 _14569_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_06979_),
    .ZN(_06980_)
  );
  OR2_X1 _14570_ (
    .A1(_06977_),
    .A2(_06980_),
    .ZN(_06981_)
  );
  MUX2_X1 _14571_ (
    .A(\rf[6] [5]),
    .B(\rf[2] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06982_)
  );
  AND2_X1 _14572_ (
    .A1(_03049_),
    .A2(_06982_),
    .ZN(_06983_)
  );
  MUX2_X1 _14573_ (
    .A(\rf[4] [5]),
    .B(\rf[0] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_06984_)
  );
  AND2_X1 _14574_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_06984_),
    .ZN(_06985_)
  );
  OR2_X1 _14575_ (
    .A1(_03048_),
    .A2(_06985_),
    .ZN(_06986_)
  );
  OR2_X1 _14576_ (
    .A1(_06983_),
    .A2(_06986_),
    .ZN(_06987_)
  );
  AND2_X1 _14577_ (
    .A1(_06981_),
    .A2(_06987_),
    .ZN(_06988_)
  );
  AND2_X1 _14578_ (
    .A1(\rf[14] [5]),
    .A2(_03049_),
    .ZN(_06989_)
  );
  AND2_X1 _14579_ (
    .A1(\rf[12] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_06990_)
  );
  OR2_X1 _14580_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[2]),
    .A2(_06990_),
    .ZN(_06991_)
  );
  OR2_X1 _14581_ (
    .A1(_06989_),
    .A2(_06991_),
    .ZN(_06992_)
  );
  AND2_X1 _14582_ (
    .A1(\rf[10] [5]),
    .A2(_03049_),
    .ZN(_06993_)
  );
  AND2_X1 _14583_ (
    .A1(\rf[8] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_06994_)
  );
  OR2_X1 _14584_ (
    .A1(_03050_),
    .A2(_06994_),
    .ZN(_06995_)
  );
  OR2_X1 _14585_ (
    .A1(_06993_),
    .A2(_06995_),
    .ZN(_06996_)
  );
  AND2_X1 _14586_ (
    .A1(_06992_),
    .A2(_06996_),
    .ZN(_06997_)
  );
  AND2_X1 _14587_ (
    .A1(\rf[15] [5]),
    .A2(_03049_),
    .ZN(_06998_)
  );
  AND2_X1 _14588_ (
    .A1(\rf[13] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_06999_)
  );
  OR2_X1 _14589_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[2]),
    .A2(_06999_),
    .ZN(_07000_)
  );
  OR2_X1 _14590_ (
    .A1(_06998_),
    .A2(_07000_),
    .ZN(_07001_)
  );
  AND2_X1 _14591_ (
    .A1(\rf[11] [5]),
    .A2(_03049_),
    .ZN(_07002_)
  );
  AND2_X1 _14592_ (
    .A1(\rf[9] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_07003_)
  );
  OR2_X1 _14593_ (
    .A1(_03050_),
    .A2(_07003_),
    .ZN(_07004_)
  );
  OR2_X1 _14594_ (
    .A1(_07002_),
    .A2(_07004_),
    .ZN(_07005_)
  );
  AND2_X1 _14595_ (
    .A1(_07001_),
    .A2(_07005_),
    .ZN(_07006_)
  );
  MUX2_X1 _14596_ (
    .A(_06997_),
    .B(_07006_),
    .S(_03048_),
    .Z(_07007_)
  );
  MUX2_X1 _14597_ (
    .A(_06988_),
    .B(_07007_),
    .S(_03051_),
    .Z(_07008_)
  );
  OR2_X1 _14598_ (
    .A1(\rf[28] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07009_)
  );
  OR2_X1 _14599_ (
    .A1(\rf[24] [5]),
    .A2(_03050_),
    .ZN(_07010_)
  );
  AND2_X1 _14600_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07009_),
    .ZN(_07011_)
  );
  AND2_X1 _14601_ (
    .A1(_07010_),
    .A2(_07011_),
    .ZN(_07012_)
  );
  MUX2_X1 _14602_ (
    .A(\rf[30] [5]),
    .B(\rf[26] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07013_)
  );
  AND2_X1 _14603_ (
    .A1(_03049_),
    .A2(_07013_),
    .ZN(_07014_)
  );
  OR2_X1 _14604_ (
    .A1(_03048_),
    .A2(_07014_),
    .ZN(_07015_)
  );
  OR2_X1 _14605_ (
    .A1(_07012_),
    .A2(_07015_),
    .ZN(_07016_)
  );
  MUX2_X1 _14606_ (
    .A(\rf[29] [5]),
    .B(\rf[25] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07017_)
  );
  AND2_X1 _14607_ (
    .A1(\rf[27] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07018_)
  );
  MUX2_X1 _14608_ (
    .A(_07017_),
    .B(_07018_),
    .S(_03049_),
    .Z(_07019_)
  );
  OR2_X1 _14609_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07019_),
    .ZN(_07020_)
  );
  AND2_X1 _14610_ (
    .A1(_07016_),
    .A2(_07020_),
    .ZN(_07021_)
  );
  OR2_X1 _14611_ (
    .A1(\rf[20] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07022_)
  );
  OR2_X1 _14612_ (
    .A1(\rf[16] [5]),
    .A2(_03050_),
    .ZN(_07023_)
  );
  AND2_X1 _14613_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07023_),
    .ZN(_07024_)
  );
  AND2_X1 _14614_ (
    .A1(_07022_),
    .A2(_07024_),
    .ZN(_07025_)
  );
  MUX2_X1 _14615_ (
    .A(\rf[22] [5]),
    .B(\rf[18] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07026_)
  );
  AND2_X1 _14616_ (
    .A1(_03049_),
    .A2(_07026_),
    .ZN(_07027_)
  );
  OR2_X1 _14617_ (
    .A1(_03048_),
    .A2(_07027_),
    .ZN(_07028_)
  );
  OR2_X1 _14618_ (
    .A1(_07025_),
    .A2(_07028_),
    .ZN(_07029_)
  );
  OR2_X1 _14619_ (
    .A1(\rf[17] [5]),
    .A2(_03050_),
    .ZN(_07030_)
  );
  OR2_X1 _14620_ (
    .A1(\rf[21] [5]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07031_)
  );
  AND2_X1 _14621_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07031_),
    .ZN(_07032_)
  );
  AND2_X1 _14622_ (
    .A1(_07030_),
    .A2(_07032_),
    .ZN(_07033_)
  );
  MUX2_X1 _14623_ (
    .A(\rf[23] [5]),
    .B(\rf[19] [5]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07034_)
  );
  AND2_X1 _14624_ (
    .A1(_03049_),
    .A2(_07034_),
    .ZN(_07035_)
  );
  OR2_X1 _14625_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07035_),
    .ZN(_07036_)
  );
  OR2_X1 _14626_ (
    .A1(_07033_),
    .A2(_07036_),
    .ZN(_07037_)
  );
  AND2_X1 _14627_ (
    .A1(_07029_),
    .A2(_07037_),
    .ZN(_07038_)
  );
  MUX2_X1 _14628_ (
    .A(_07021_),
    .B(_07038_),
    .S(ibuf_io_inst_0_bits_inst_rs2[3]),
    .Z(_07039_)
  );
  MUX2_X1 _14629_ (
    .A(_07008_),
    .B(_07039_),
    .S(_03064_),
    .Z(_07040_)
  );
  MUX2_X1 _14630_ (
    .A(_07040_),
    .B(_04305_),
    .S(_06791_),
    .Z(_07041_)
  );
  MUX2_X1 _14631_ (
    .A(ex_reg_rs_msb_1[3]),
    .B(_07041_),
    .S(_06781_),
    .Z(_00152_)
  );
  OR2_X1 _14632_ (
    .A1(\rf[10] [6]),
    .A2(_03050_),
    .ZN(_07042_)
  );
  OR2_X1 _14633_ (
    .A1(\rf[14] [6]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07043_)
  );
  AND2_X1 _14634_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07043_),
    .ZN(_07044_)
  );
  AND2_X1 _14635_ (
    .A1(_07042_),
    .A2(_07044_),
    .ZN(_07045_)
  );
  MUX2_X1 _14636_ (
    .A(\rf[15] [6]),
    .B(\rf[11] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07046_)
  );
  AND2_X1 _14637_ (
    .A1(_03048_),
    .A2(_07046_),
    .ZN(_07047_)
  );
  OR2_X1 _14638_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07047_),
    .ZN(_07048_)
  );
  OR2_X1 _14639_ (
    .A1(_07045_),
    .A2(_07048_),
    .ZN(_07049_)
  );
  OR2_X1 _14640_ (
    .A1(\rf[12] [6]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07050_)
  );
  OR2_X1 _14641_ (
    .A1(\rf[8] [6]),
    .A2(_03050_),
    .ZN(_07051_)
  );
  AND2_X1 _14642_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07050_),
    .ZN(_07052_)
  );
  AND2_X1 _14643_ (
    .A1(_07051_),
    .A2(_07052_),
    .ZN(_07053_)
  );
  MUX2_X1 _14644_ (
    .A(\rf[13] [6]),
    .B(\rf[9] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07054_)
  );
  AND2_X1 _14645_ (
    .A1(_03048_),
    .A2(_07054_),
    .ZN(_07055_)
  );
  OR2_X1 _14646_ (
    .A1(_03049_),
    .A2(_07055_),
    .ZN(_07056_)
  );
  OR2_X1 _14647_ (
    .A1(_07053_),
    .A2(_07056_),
    .ZN(_07057_)
  );
  AND2_X1 _14648_ (
    .A1(_03051_),
    .A2(_07057_),
    .ZN(_07058_)
  );
  AND2_X1 _14649_ (
    .A1(_07049_),
    .A2(_07058_),
    .ZN(_07059_)
  );
  MUX2_X1 _14650_ (
    .A(\rf[6] [6]),
    .B(\rf[2] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07060_)
  );
  AND2_X1 _14651_ (
    .A1(_03049_),
    .A2(_07060_),
    .ZN(_07061_)
  );
  MUX2_X1 _14652_ (
    .A(\rf[4] [6]),
    .B(\rf[0] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07062_)
  );
  AND2_X1 _14653_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07062_),
    .ZN(_07063_)
  );
  OR2_X1 _14654_ (
    .A1(_03048_),
    .A2(_07063_),
    .ZN(_07064_)
  );
  OR2_X1 _14655_ (
    .A1(_07061_),
    .A2(_07064_),
    .ZN(_07065_)
  );
  MUX2_X1 _14656_ (
    .A(\rf[7] [6]),
    .B(\rf[3] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07066_)
  );
  AND2_X1 _14657_ (
    .A1(_03049_),
    .A2(_07066_),
    .ZN(_07067_)
  );
  MUX2_X1 _14658_ (
    .A(\rf[5] [6]),
    .B(\rf[1] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07068_)
  );
  AND2_X1 _14659_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07068_),
    .ZN(_07069_)
  );
  OR2_X1 _14660_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07069_),
    .ZN(_07070_)
  );
  OR2_X1 _14661_ (
    .A1(_07067_),
    .A2(_07070_),
    .ZN(_07071_)
  );
  AND2_X1 _14662_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_07071_),
    .ZN(_07072_)
  );
  AND2_X1 _14663_ (
    .A1(_07065_),
    .A2(_07072_),
    .ZN(_07073_)
  );
  OR2_X1 _14664_ (
    .A1(_07059_),
    .A2(_07073_),
    .ZN(_07074_)
  );
  OR2_X1 _14665_ (
    .A1(\rf[17] [6]),
    .A2(_03050_),
    .ZN(_07075_)
  );
  OR2_X1 _14666_ (
    .A1(\rf[21] [6]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07076_)
  );
  AND2_X1 _14667_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07076_),
    .ZN(_07077_)
  );
  AND2_X1 _14668_ (
    .A1(_07075_),
    .A2(_07077_),
    .ZN(_07078_)
  );
  MUX2_X1 _14669_ (
    .A(\rf[23] [6]),
    .B(\rf[19] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07079_)
  );
  AND2_X1 _14670_ (
    .A1(_03049_),
    .A2(_07079_),
    .ZN(_07080_)
  );
  OR2_X1 _14671_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07080_),
    .ZN(_07081_)
  );
  OR2_X1 _14672_ (
    .A1(_07078_),
    .A2(_07081_),
    .ZN(_07082_)
  );
  OR2_X1 _14673_ (
    .A1(\rf[20] [6]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07083_)
  );
  OR2_X1 _14674_ (
    .A1(\rf[16] [6]),
    .A2(_03050_),
    .ZN(_07084_)
  );
  AND2_X1 _14675_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07084_),
    .ZN(_07085_)
  );
  AND2_X1 _14676_ (
    .A1(_07083_),
    .A2(_07085_),
    .ZN(_07086_)
  );
  MUX2_X1 _14677_ (
    .A(\rf[22] [6]),
    .B(\rf[18] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07087_)
  );
  AND2_X1 _14678_ (
    .A1(_03049_),
    .A2(_07087_),
    .ZN(_07088_)
  );
  OR2_X1 _14679_ (
    .A1(_03048_),
    .A2(_07088_),
    .ZN(_07089_)
  );
  OR2_X1 _14680_ (
    .A1(_07086_),
    .A2(_07089_),
    .ZN(_07090_)
  );
  AND2_X1 _14681_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_07082_),
    .ZN(_07091_)
  );
  AND2_X1 _14682_ (
    .A1(_07090_),
    .A2(_07091_),
    .ZN(_07092_)
  );
  OR2_X1 _14683_ (
    .A1(\rf[28] [6]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07093_)
  );
  OR2_X1 _14684_ (
    .A1(\rf[24] [6]),
    .A2(_03050_),
    .ZN(_07094_)
  );
  AND2_X1 _14685_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07093_),
    .ZN(_07095_)
  );
  AND2_X1 _14686_ (
    .A1(_07094_),
    .A2(_07095_),
    .ZN(_07096_)
  );
  MUX2_X1 _14687_ (
    .A(\rf[30] [6]),
    .B(\rf[26] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07097_)
  );
  AND2_X1 _14688_ (
    .A1(_03049_),
    .A2(_07097_),
    .ZN(_07098_)
  );
  OR2_X1 _14689_ (
    .A1(_03048_),
    .A2(_07098_),
    .ZN(_07099_)
  );
  OR2_X1 _14690_ (
    .A1(_07096_),
    .A2(_07099_),
    .ZN(_07100_)
  );
  MUX2_X1 _14691_ (
    .A(\rf[29] [6]),
    .B(\rf[25] [6]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07101_)
  );
  AND2_X1 _14692_ (
    .A1(\rf[27] [6]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07102_)
  );
  MUX2_X1 _14693_ (
    .A(_07101_),
    .B(_07102_),
    .S(_03049_),
    .Z(_07103_)
  );
  OR2_X1 _14694_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07103_),
    .ZN(_07104_)
  );
  AND2_X1 _14695_ (
    .A1(_03051_),
    .A2(_07104_),
    .ZN(_07105_)
  );
  AND2_X1 _14696_ (
    .A1(_07100_),
    .A2(_07105_),
    .ZN(_07106_)
  );
  OR2_X1 _14697_ (
    .A1(_07092_),
    .A2(_07106_),
    .ZN(_07107_)
  );
  MUX2_X1 _14698_ (
    .A(_07074_),
    .B(_07107_),
    .S(_03064_),
    .Z(_07108_)
  );
  MUX2_X1 _14699_ (
    .A(_07108_),
    .B(_04379_),
    .S(_06791_),
    .Z(_07109_)
  );
  MUX2_X1 _14700_ (
    .A(ex_reg_rs_msb_1[4]),
    .B(_07109_),
    .S(_06781_),
    .Z(_00153_)
  );
  MUX2_X1 _14701_ (
    .A(\rf[1] [7]),
    .B(\rf[0] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_07110_)
  );
  MUX2_X1 _14702_ (
    .A(\rf[5] [7]),
    .B(\rf[4] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_07111_)
  );
  MUX2_X1 _14703_ (
    .A(_07110_),
    .B(_07111_),
    .S(_03050_),
    .Z(_07112_)
  );
  OR2_X1 _14704_ (
    .A1(_03051_),
    .A2(_07112_),
    .ZN(_07113_)
  );
  MUX2_X1 _14705_ (
    .A(\rf[12] [7]),
    .B(\rf[8] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07114_)
  );
  OR2_X1 _14706_ (
    .A1(_06863_),
    .A2(_07114_),
    .ZN(_07115_)
  );
  MUX2_X1 _14707_ (
    .A(\rf[13] [7]),
    .B(\rf[9] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07116_)
  );
  OR2_X1 _14708_ (
    .A1(_03808_),
    .A2(_07116_),
    .ZN(_07117_)
  );
  AND2_X1 _14709_ (
    .A1(_07115_),
    .A2(_07117_),
    .ZN(_07118_)
  );
  AND2_X1 _14710_ (
    .A1(_07113_),
    .A2(_07118_),
    .ZN(_07119_)
  );
  MUX2_X1 _14711_ (
    .A(\rf[3] [7]),
    .B(\rf[2] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_07120_)
  );
  MUX2_X1 _14712_ (
    .A(\rf[7] [7]),
    .B(\rf[6] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_07121_)
  );
  MUX2_X1 _14713_ (
    .A(_07120_),
    .B(_07121_),
    .S(_03050_),
    .Z(_07122_)
  );
  OR2_X1 _14714_ (
    .A1(_03051_),
    .A2(_07122_),
    .ZN(_07123_)
  );
  MUX2_X1 _14715_ (
    .A(\rf[15] [7]),
    .B(\rf[11] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07124_)
  );
  OR2_X1 _14716_ (
    .A1(_03808_),
    .A2(_07124_),
    .ZN(_07125_)
  );
  MUX2_X1 _14717_ (
    .A(\rf[14] [7]),
    .B(\rf[10] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07126_)
  );
  OR2_X1 _14718_ (
    .A1(_06863_),
    .A2(_07126_),
    .ZN(_07127_)
  );
  AND2_X1 _14719_ (
    .A1(_07125_),
    .A2(_07127_),
    .ZN(_07128_)
  );
  AND2_X1 _14720_ (
    .A1(_07123_),
    .A2(_07128_),
    .ZN(_07129_)
  );
  MUX2_X1 _14721_ (
    .A(_07119_),
    .B(_07129_),
    .S(_03049_),
    .Z(_07130_)
  );
  OR2_X1 _14722_ (
    .A1(\rf[17] [7]),
    .A2(_03050_),
    .ZN(_07131_)
  );
  OR2_X1 _14723_ (
    .A1(\rf[21] [7]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07132_)
  );
  AND2_X1 _14724_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07132_),
    .ZN(_07133_)
  );
  AND2_X1 _14725_ (
    .A1(_07131_),
    .A2(_07133_),
    .ZN(_07134_)
  );
  MUX2_X1 _14726_ (
    .A(\rf[23] [7]),
    .B(\rf[19] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07135_)
  );
  AND2_X1 _14727_ (
    .A1(_03049_),
    .A2(_07135_),
    .ZN(_07136_)
  );
  OR2_X1 _14728_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07136_),
    .ZN(_07137_)
  );
  OR2_X1 _14729_ (
    .A1(_07134_),
    .A2(_07137_),
    .ZN(_07138_)
  );
  OR2_X1 _14730_ (
    .A1(\rf[20] [7]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07139_)
  );
  OR2_X1 _14731_ (
    .A1(\rf[16] [7]),
    .A2(_03050_),
    .ZN(_07140_)
  );
  AND2_X1 _14732_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07140_),
    .ZN(_07141_)
  );
  AND2_X1 _14733_ (
    .A1(_07139_),
    .A2(_07141_),
    .ZN(_07142_)
  );
  MUX2_X1 _14734_ (
    .A(\rf[22] [7]),
    .B(\rf[18] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07143_)
  );
  AND2_X1 _14735_ (
    .A1(_03049_),
    .A2(_07143_),
    .ZN(_07144_)
  );
  OR2_X1 _14736_ (
    .A1(_03048_),
    .A2(_07144_),
    .ZN(_07145_)
  );
  OR2_X1 _14737_ (
    .A1(_07142_),
    .A2(_07145_),
    .ZN(_07146_)
  );
  AND2_X1 _14738_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_07138_),
    .ZN(_07147_)
  );
  AND2_X1 _14739_ (
    .A1(_07146_),
    .A2(_07147_),
    .ZN(_07148_)
  );
  OR2_X1 _14740_ (
    .A1(\rf[28] [7]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07149_)
  );
  OR2_X1 _14741_ (
    .A1(\rf[24] [7]),
    .A2(_03050_),
    .ZN(_07150_)
  );
  AND2_X1 _14742_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07149_),
    .ZN(_07151_)
  );
  AND2_X1 _14743_ (
    .A1(_07150_),
    .A2(_07151_),
    .ZN(_07152_)
  );
  MUX2_X1 _14744_ (
    .A(\rf[30] [7]),
    .B(\rf[26] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07153_)
  );
  AND2_X1 _14745_ (
    .A1(_03049_),
    .A2(_07153_),
    .ZN(_07154_)
  );
  OR2_X1 _14746_ (
    .A1(_03048_),
    .A2(_07154_),
    .ZN(_07155_)
  );
  OR2_X1 _14747_ (
    .A1(_07152_),
    .A2(_07155_),
    .ZN(_07156_)
  );
  MUX2_X1 _14748_ (
    .A(\rf[29] [7]),
    .B(\rf[25] [7]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07157_)
  );
  AND2_X1 _14749_ (
    .A1(\rf[27] [7]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07158_)
  );
  MUX2_X1 _14750_ (
    .A(_07157_),
    .B(_07158_),
    .S(_03049_),
    .Z(_07159_)
  );
  OR2_X1 _14751_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07159_),
    .ZN(_07160_)
  );
  AND2_X1 _14752_ (
    .A1(_03051_),
    .A2(_07160_),
    .ZN(_07161_)
  );
  AND2_X1 _14753_ (
    .A1(_07156_),
    .A2(_07161_),
    .ZN(_07162_)
  );
  OR2_X1 _14754_ (
    .A1(_07148_),
    .A2(_07162_),
    .ZN(_07163_)
  );
  MUX2_X1 _14755_ (
    .A(_07130_),
    .B(_07163_),
    .S(_03064_),
    .Z(_07164_)
  );
  MUX2_X1 _14756_ (
    .A(_07164_),
    .B(_04450_),
    .S(_06791_),
    .Z(_07165_)
  );
  MUX2_X1 _14757_ (
    .A(ex_reg_rs_msb_1[5]),
    .B(_07165_),
    .S(_06781_),
    .Z(_00154_)
  );
  OR2_X1 _14758_ (
    .A1(\rf[10] [8]),
    .A2(_03050_),
    .ZN(_07166_)
  );
  OR2_X1 _14759_ (
    .A1(\rf[14] [8]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07167_)
  );
  AND2_X1 _14760_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07167_),
    .ZN(_07168_)
  );
  AND2_X1 _14761_ (
    .A1(_07166_),
    .A2(_07168_),
    .ZN(_07169_)
  );
  MUX2_X1 _14762_ (
    .A(\rf[15] [8]),
    .B(\rf[11] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07170_)
  );
  AND2_X1 _14763_ (
    .A1(_03048_),
    .A2(_07170_),
    .ZN(_07171_)
  );
  OR2_X1 _14764_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07171_),
    .ZN(_07172_)
  );
  OR2_X1 _14765_ (
    .A1(_07169_),
    .A2(_07172_),
    .ZN(_07173_)
  );
  OR2_X1 _14766_ (
    .A1(\rf[12] [8]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07174_)
  );
  OR2_X1 _14767_ (
    .A1(\rf[8] [8]),
    .A2(_03050_),
    .ZN(_07175_)
  );
  AND2_X1 _14768_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07174_),
    .ZN(_07176_)
  );
  AND2_X1 _14769_ (
    .A1(_07175_),
    .A2(_07176_),
    .ZN(_07177_)
  );
  MUX2_X1 _14770_ (
    .A(\rf[13] [8]),
    .B(\rf[9] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07178_)
  );
  AND2_X1 _14771_ (
    .A1(_03048_),
    .A2(_07178_),
    .ZN(_07179_)
  );
  OR2_X1 _14772_ (
    .A1(_03049_),
    .A2(_07179_),
    .ZN(_07180_)
  );
  OR2_X1 _14773_ (
    .A1(_07177_),
    .A2(_07180_),
    .ZN(_07181_)
  );
  AND2_X1 _14774_ (
    .A1(_03051_),
    .A2(_07181_),
    .ZN(_07182_)
  );
  AND2_X1 _14775_ (
    .A1(_07173_),
    .A2(_07182_),
    .ZN(_07183_)
  );
  MUX2_X1 _14776_ (
    .A(\rf[6] [8]),
    .B(\rf[2] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07184_)
  );
  AND2_X1 _14777_ (
    .A1(_03049_),
    .A2(_07184_),
    .ZN(_07185_)
  );
  MUX2_X1 _14778_ (
    .A(\rf[4] [8]),
    .B(\rf[0] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07186_)
  );
  AND2_X1 _14779_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07186_),
    .ZN(_07187_)
  );
  OR2_X1 _14780_ (
    .A1(_03048_),
    .A2(_07187_),
    .ZN(_07188_)
  );
  OR2_X1 _14781_ (
    .A1(_07185_),
    .A2(_07188_),
    .ZN(_07189_)
  );
  MUX2_X1 _14782_ (
    .A(\rf[7] [8]),
    .B(\rf[3] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07190_)
  );
  AND2_X1 _14783_ (
    .A1(_03049_),
    .A2(_07190_),
    .ZN(_07191_)
  );
  MUX2_X1 _14784_ (
    .A(\rf[5] [8]),
    .B(\rf[1] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07192_)
  );
  AND2_X1 _14785_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07192_),
    .ZN(_07193_)
  );
  OR2_X1 _14786_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07193_),
    .ZN(_07194_)
  );
  OR2_X1 _14787_ (
    .A1(_07191_),
    .A2(_07194_),
    .ZN(_07195_)
  );
  AND2_X1 _14788_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_07195_),
    .ZN(_07196_)
  );
  AND2_X1 _14789_ (
    .A1(_07189_),
    .A2(_07196_),
    .ZN(_07197_)
  );
  OR2_X1 _14790_ (
    .A1(_07183_),
    .A2(_07197_),
    .ZN(_07198_)
  );
  OR2_X1 _14791_ (
    .A1(\rf[17] [8]),
    .A2(_03050_),
    .ZN(_07199_)
  );
  OR2_X1 _14792_ (
    .A1(\rf[21] [8]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07200_)
  );
  AND2_X1 _14793_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07200_),
    .ZN(_07201_)
  );
  AND2_X1 _14794_ (
    .A1(_07199_),
    .A2(_07201_),
    .ZN(_07202_)
  );
  MUX2_X1 _14795_ (
    .A(\rf[23] [8]),
    .B(\rf[19] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07203_)
  );
  AND2_X1 _14796_ (
    .A1(_03049_),
    .A2(_07203_),
    .ZN(_07204_)
  );
  OR2_X1 _14797_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07204_),
    .ZN(_07205_)
  );
  OR2_X1 _14798_ (
    .A1(_07202_),
    .A2(_07205_),
    .ZN(_07206_)
  );
  OR2_X1 _14799_ (
    .A1(\rf[20] [8]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07207_)
  );
  OR2_X1 _14800_ (
    .A1(\rf[16] [8]),
    .A2(_03050_),
    .ZN(_07208_)
  );
  AND2_X1 _14801_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07208_),
    .ZN(_07209_)
  );
  AND2_X1 _14802_ (
    .A1(_07207_),
    .A2(_07209_),
    .ZN(_07210_)
  );
  MUX2_X1 _14803_ (
    .A(\rf[22] [8]),
    .B(\rf[18] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07211_)
  );
  AND2_X1 _14804_ (
    .A1(_03049_),
    .A2(_07211_),
    .ZN(_07212_)
  );
  OR2_X1 _14805_ (
    .A1(_03048_),
    .A2(_07212_),
    .ZN(_07213_)
  );
  OR2_X1 _14806_ (
    .A1(_07210_),
    .A2(_07213_),
    .ZN(_07214_)
  );
  AND2_X1 _14807_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_07206_),
    .ZN(_07215_)
  );
  AND2_X1 _14808_ (
    .A1(_07214_),
    .A2(_07215_),
    .ZN(_07216_)
  );
  OR2_X1 _14809_ (
    .A1(\rf[28] [8]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07217_)
  );
  OR2_X1 _14810_ (
    .A1(\rf[24] [8]),
    .A2(_03050_),
    .ZN(_07218_)
  );
  AND2_X1 _14811_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07217_),
    .ZN(_07219_)
  );
  AND2_X1 _14812_ (
    .A1(_07218_),
    .A2(_07219_),
    .ZN(_07220_)
  );
  MUX2_X1 _14813_ (
    .A(\rf[30] [8]),
    .B(\rf[26] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07221_)
  );
  AND2_X1 _14814_ (
    .A1(_03049_),
    .A2(_07221_),
    .ZN(_07222_)
  );
  OR2_X1 _14815_ (
    .A1(_03048_),
    .A2(_07222_),
    .ZN(_07223_)
  );
  OR2_X1 _14816_ (
    .A1(_07220_),
    .A2(_07223_),
    .ZN(_07224_)
  );
  MUX2_X1 _14817_ (
    .A(\rf[29] [8]),
    .B(\rf[25] [8]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07225_)
  );
  AND2_X1 _14818_ (
    .A1(\rf[27] [8]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07226_)
  );
  MUX2_X1 _14819_ (
    .A(_07225_),
    .B(_07226_),
    .S(_03049_),
    .Z(_07227_)
  );
  OR2_X1 _14820_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07227_),
    .ZN(_07228_)
  );
  AND2_X1 _14821_ (
    .A1(_03051_),
    .A2(_07228_),
    .ZN(_07229_)
  );
  AND2_X1 _14822_ (
    .A1(_07224_),
    .A2(_07229_),
    .ZN(_07230_)
  );
  OR2_X1 _14823_ (
    .A1(_07216_),
    .A2(_07230_),
    .ZN(_07231_)
  );
  MUX2_X1 _14824_ (
    .A(_07198_),
    .B(_07231_),
    .S(_03064_),
    .Z(_07232_)
  );
  MUX2_X1 _14825_ (
    .A(_07232_),
    .B(_04521_),
    .S(_06791_),
    .Z(_07233_)
  );
  MUX2_X1 _14826_ (
    .A(ex_reg_rs_msb_1[6]),
    .B(_07233_),
    .S(_06781_),
    .Z(_00155_)
  );
  OR2_X1 _14827_ (
    .A1(\rf[10] [9]),
    .A2(_03050_),
    .ZN(_07234_)
  );
  OR2_X1 _14828_ (
    .A1(\rf[14] [9]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07235_)
  );
  AND2_X1 _14829_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07235_),
    .ZN(_07236_)
  );
  AND2_X1 _14830_ (
    .A1(_07234_),
    .A2(_07236_),
    .ZN(_07237_)
  );
  MUX2_X1 _14831_ (
    .A(\rf[15] [9]),
    .B(\rf[11] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07238_)
  );
  AND2_X1 _14832_ (
    .A1(_03048_),
    .A2(_07238_),
    .ZN(_07239_)
  );
  OR2_X1 _14833_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07239_),
    .ZN(_07240_)
  );
  OR2_X1 _14834_ (
    .A1(_07237_),
    .A2(_07240_),
    .ZN(_07241_)
  );
  OR2_X1 _14835_ (
    .A1(\rf[12] [9]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07242_)
  );
  OR2_X1 _14836_ (
    .A1(\rf[8] [9]),
    .A2(_03050_),
    .ZN(_07243_)
  );
  AND2_X1 _14837_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07242_),
    .ZN(_07244_)
  );
  AND2_X1 _14838_ (
    .A1(_07243_),
    .A2(_07244_),
    .ZN(_07245_)
  );
  MUX2_X1 _14839_ (
    .A(\rf[13] [9]),
    .B(\rf[9] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07246_)
  );
  AND2_X1 _14840_ (
    .A1(_03048_),
    .A2(_07246_),
    .ZN(_07247_)
  );
  OR2_X1 _14841_ (
    .A1(_03049_),
    .A2(_07247_),
    .ZN(_07248_)
  );
  OR2_X1 _14842_ (
    .A1(_07245_),
    .A2(_07248_),
    .ZN(_07249_)
  );
  AND2_X1 _14843_ (
    .A1(_03051_),
    .A2(_07249_),
    .ZN(_07250_)
  );
  AND2_X1 _14844_ (
    .A1(_07241_),
    .A2(_07250_),
    .ZN(_07251_)
  );
  MUX2_X1 _14845_ (
    .A(\rf[6] [9]),
    .B(\rf[2] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07252_)
  );
  AND2_X1 _14846_ (
    .A1(_03049_),
    .A2(_07252_),
    .ZN(_07253_)
  );
  MUX2_X1 _14847_ (
    .A(\rf[4] [9]),
    .B(\rf[0] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07254_)
  );
  AND2_X1 _14848_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07254_),
    .ZN(_07255_)
  );
  OR2_X1 _14849_ (
    .A1(_03048_),
    .A2(_07255_),
    .ZN(_07256_)
  );
  OR2_X1 _14850_ (
    .A1(_07253_),
    .A2(_07256_),
    .ZN(_07257_)
  );
  MUX2_X1 _14851_ (
    .A(\rf[7] [9]),
    .B(\rf[3] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07258_)
  );
  AND2_X1 _14852_ (
    .A1(_03049_),
    .A2(_07258_),
    .ZN(_07259_)
  );
  MUX2_X1 _14853_ (
    .A(\rf[5] [9]),
    .B(\rf[1] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07260_)
  );
  AND2_X1 _14854_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07260_),
    .ZN(_07261_)
  );
  OR2_X1 _14855_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07261_),
    .ZN(_07262_)
  );
  OR2_X1 _14856_ (
    .A1(_07259_),
    .A2(_07262_),
    .ZN(_07263_)
  );
  AND2_X1 _14857_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_07263_),
    .ZN(_07264_)
  );
  AND2_X1 _14858_ (
    .A1(_07257_),
    .A2(_07264_),
    .ZN(_07265_)
  );
  OR2_X1 _14859_ (
    .A1(_07251_),
    .A2(_07265_),
    .ZN(_07266_)
  );
  OR2_X1 _14860_ (
    .A1(\rf[17] [9]),
    .A2(_03050_),
    .ZN(_07267_)
  );
  OR2_X1 _14861_ (
    .A1(\rf[21] [9]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07268_)
  );
  AND2_X1 _14862_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07268_),
    .ZN(_07269_)
  );
  AND2_X1 _14863_ (
    .A1(_07267_),
    .A2(_07269_),
    .ZN(_07270_)
  );
  MUX2_X1 _14864_ (
    .A(\rf[23] [9]),
    .B(\rf[19] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07271_)
  );
  AND2_X1 _14865_ (
    .A1(_03049_),
    .A2(_07271_),
    .ZN(_07272_)
  );
  OR2_X1 _14866_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07272_),
    .ZN(_07273_)
  );
  OR2_X1 _14867_ (
    .A1(_07270_),
    .A2(_07273_),
    .ZN(_07274_)
  );
  OR2_X1 _14868_ (
    .A1(\rf[20] [9]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07275_)
  );
  OR2_X1 _14869_ (
    .A1(\rf[16] [9]),
    .A2(_03050_),
    .ZN(_07276_)
  );
  AND2_X1 _14870_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07276_),
    .ZN(_07277_)
  );
  AND2_X1 _14871_ (
    .A1(_07275_),
    .A2(_07277_),
    .ZN(_07278_)
  );
  MUX2_X1 _14872_ (
    .A(\rf[22] [9]),
    .B(\rf[18] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07279_)
  );
  AND2_X1 _14873_ (
    .A1(_03049_),
    .A2(_07279_),
    .ZN(_07280_)
  );
  OR2_X1 _14874_ (
    .A1(_03048_),
    .A2(_07280_),
    .ZN(_07281_)
  );
  OR2_X1 _14875_ (
    .A1(_07278_),
    .A2(_07281_),
    .ZN(_07282_)
  );
  AND2_X1 _14876_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_07274_),
    .ZN(_07283_)
  );
  AND2_X1 _14877_ (
    .A1(_07282_),
    .A2(_07283_),
    .ZN(_07284_)
  );
  OR2_X1 _14878_ (
    .A1(\rf[28] [9]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07285_)
  );
  OR2_X1 _14879_ (
    .A1(\rf[24] [9]),
    .A2(_03050_),
    .ZN(_07286_)
  );
  AND2_X1 _14880_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07285_),
    .ZN(_07287_)
  );
  AND2_X1 _14881_ (
    .A1(_07286_),
    .A2(_07287_),
    .ZN(_07288_)
  );
  MUX2_X1 _14882_ (
    .A(\rf[30] [9]),
    .B(\rf[26] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07289_)
  );
  AND2_X1 _14883_ (
    .A1(_03049_),
    .A2(_07289_),
    .ZN(_07290_)
  );
  OR2_X1 _14884_ (
    .A1(_03048_),
    .A2(_07290_),
    .ZN(_07291_)
  );
  OR2_X1 _14885_ (
    .A1(_07288_),
    .A2(_07291_),
    .ZN(_07292_)
  );
  MUX2_X1 _14886_ (
    .A(\rf[29] [9]),
    .B(\rf[25] [9]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07293_)
  );
  AND2_X1 _14887_ (
    .A1(\rf[27] [9]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07294_)
  );
  MUX2_X1 _14888_ (
    .A(_07293_),
    .B(_07294_),
    .S(_03049_),
    .Z(_07295_)
  );
  OR2_X1 _14889_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07295_),
    .ZN(_07296_)
  );
  AND2_X1 _14890_ (
    .A1(_03051_),
    .A2(_07296_),
    .ZN(_07297_)
  );
  AND2_X1 _14891_ (
    .A1(_07292_),
    .A2(_07297_),
    .ZN(_07298_)
  );
  OR2_X1 _14892_ (
    .A1(_07284_),
    .A2(_07298_),
    .ZN(_07299_)
  );
  MUX2_X1 _14893_ (
    .A(_07266_),
    .B(_07299_),
    .S(_03064_),
    .Z(_07300_)
  );
  MUX2_X1 _14894_ (
    .A(_07300_),
    .B(_04590_),
    .S(_06791_),
    .Z(_07301_)
  );
  MUX2_X1 _14895_ (
    .A(ex_reg_rs_msb_1[7]),
    .B(_07301_),
    .S(_06781_),
    .Z(_00156_)
  );
  MUX2_X1 _14896_ (
    .A(\rf[3] [10]),
    .B(\rf[2] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_07302_)
  );
  MUX2_X1 _14897_ (
    .A(\rf[7] [10]),
    .B(\rf[6] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_07303_)
  );
  MUX2_X1 _14898_ (
    .A(_07302_),
    .B(_07303_),
    .S(_03050_),
    .Z(_07304_)
  );
  OR2_X1 _14899_ (
    .A1(_03051_),
    .A2(_07304_),
    .ZN(_07305_)
  );
  MUX2_X1 _14900_ (
    .A(\rf[15] [10]),
    .B(\rf[11] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07306_)
  );
  OR2_X1 _14901_ (
    .A1(_03808_),
    .A2(_07306_),
    .ZN(_07307_)
  );
  MUX2_X1 _14902_ (
    .A(\rf[14] [10]),
    .B(\rf[10] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07308_)
  );
  OR2_X1 _14903_ (
    .A1(_06863_),
    .A2(_07308_),
    .ZN(_07309_)
  );
  AND2_X1 _14904_ (
    .A1(_07307_),
    .A2(_07309_),
    .ZN(_07310_)
  );
  AND2_X1 _14905_ (
    .A1(_07305_),
    .A2(_07310_),
    .ZN(_07311_)
  );
  MUX2_X1 _14906_ (
    .A(\rf[1] [10]),
    .B(\rf[0] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_07312_)
  );
  MUX2_X1 _14907_ (
    .A(\rf[5] [10]),
    .B(\rf[4] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_07313_)
  );
  MUX2_X1 _14908_ (
    .A(_07312_),
    .B(_07313_),
    .S(_03050_),
    .Z(_07314_)
  );
  OR2_X1 _14909_ (
    .A1(_03051_),
    .A2(_07314_),
    .ZN(_07315_)
  );
  MUX2_X1 _14910_ (
    .A(\rf[12] [10]),
    .B(\rf[8] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07316_)
  );
  OR2_X1 _14911_ (
    .A1(_06863_),
    .A2(_07316_),
    .ZN(_07317_)
  );
  MUX2_X1 _14912_ (
    .A(\rf[13] [10]),
    .B(\rf[9] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07318_)
  );
  OR2_X1 _14913_ (
    .A1(_03808_),
    .A2(_07318_),
    .ZN(_07319_)
  );
  AND2_X1 _14914_ (
    .A1(_07317_),
    .A2(_07319_),
    .ZN(_07320_)
  );
  AND2_X1 _14915_ (
    .A1(_07315_),
    .A2(_07320_),
    .ZN(_07321_)
  );
  OR2_X1 _14916_ (
    .A1(\rf[28] [10]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07322_)
  );
  OR2_X1 _14917_ (
    .A1(\rf[24] [10]),
    .A2(_03050_),
    .ZN(_07323_)
  );
  AND2_X1 _14918_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07322_),
    .ZN(_07324_)
  );
  AND2_X1 _14919_ (
    .A1(_07323_),
    .A2(_07324_),
    .ZN(_07325_)
  );
  MUX2_X1 _14920_ (
    .A(\rf[30] [10]),
    .B(\rf[26] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07326_)
  );
  AND2_X1 _14921_ (
    .A1(_03049_),
    .A2(_07326_),
    .ZN(_07327_)
  );
  OR2_X1 _14922_ (
    .A1(_03048_),
    .A2(_07327_),
    .ZN(_07328_)
  );
  OR2_X1 _14923_ (
    .A1(_07325_),
    .A2(_07328_),
    .ZN(_07329_)
  );
  MUX2_X1 _14924_ (
    .A(\rf[29] [10]),
    .B(\rf[25] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07330_)
  );
  AND2_X1 _14925_ (
    .A1(\rf[27] [10]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07331_)
  );
  MUX2_X1 _14926_ (
    .A(_07330_),
    .B(_07331_),
    .S(_03049_),
    .Z(_07332_)
  );
  OR2_X1 _14927_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07332_),
    .ZN(_07333_)
  );
  AND2_X1 _14928_ (
    .A1(_07329_),
    .A2(_07333_),
    .ZN(_07334_)
  );
  OR2_X1 _14929_ (
    .A1(\rf[20] [10]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07335_)
  );
  OR2_X1 _14930_ (
    .A1(\rf[16] [10]),
    .A2(_03050_),
    .ZN(_07336_)
  );
  AND2_X1 _14931_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07336_),
    .ZN(_07337_)
  );
  AND2_X1 _14932_ (
    .A1(_07335_),
    .A2(_07337_),
    .ZN(_07338_)
  );
  MUX2_X1 _14933_ (
    .A(\rf[22] [10]),
    .B(\rf[18] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07339_)
  );
  AND2_X1 _14934_ (
    .A1(_03049_),
    .A2(_07339_),
    .ZN(_07340_)
  );
  OR2_X1 _14935_ (
    .A1(_03048_),
    .A2(_07340_),
    .ZN(_07341_)
  );
  OR2_X1 _14936_ (
    .A1(_07338_),
    .A2(_07341_),
    .ZN(_07342_)
  );
  OR2_X1 _14937_ (
    .A1(\rf[17] [10]),
    .A2(_03050_),
    .ZN(_07343_)
  );
  OR2_X1 _14938_ (
    .A1(\rf[21] [10]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07344_)
  );
  AND2_X1 _14939_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07344_),
    .ZN(_07345_)
  );
  AND2_X1 _14940_ (
    .A1(_07343_),
    .A2(_07345_),
    .ZN(_07346_)
  );
  MUX2_X1 _14941_ (
    .A(\rf[23] [10]),
    .B(\rf[19] [10]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07347_)
  );
  AND2_X1 _14942_ (
    .A1(_03049_),
    .A2(_07347_),
    .ZN(_07348_)
  );
  OR2_X1 _14943_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07348_),
    .ZN(_07349_)
  );
  OR2_X1 _14944_ (
    .A1(_07346_),
    .A2(_07349_),
    .ZN(_07350_)
  );
  AND2_X1 _14945_ (
    .A1(_07342_),
    .A2(_07350_),
    .ZN(_07351_)
  );
  MUX2_X1 _14946_ (
    .A(_07334_),
    .B(_07351_),
    .S(ibuf_io_inst_0_bits_inst_rs2[3]),
    .Z(_07352_)
  );
  MUX2_X1 _14947_ (
    .A(_07311_),
    .B(_07321_),
    .S(ibuf_io_inst_0_bits_inst_rs2[1]),
    .Z(_07353_)
  );
  MUX2_X1 _14948_ (
    .A(_07352_),
    .B(_07353_),
    .S(ibuf_io_inst_0_bits_inst_rs2[4]),
    .Z(_07354_)
  );
  MUX2_X1 _14949_ (
    .A(_07354_),
    .B(_04659_),
    .S(_06791_),
    .Z(_07355_)
  );
  MUX2_X1 _14950_ (
    .A(ex_reg_rs_msb_1[8]),
    .B(_07355_),
    .S(_06781_),
    .Z(_00157_)
  );
  OR2_X1 _14951_ (
    .A1(\rf[10] [11]),
    .A2(_03050_),
    .ZN(_07356_)
  );
  OR2_X1 _14952_ (
    .A1(\rf[14] [11]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07357_)
  );
  AND2_X1 _14953_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07357_),
    .ZN(_07358_)
  );
  AND2_X1 _14954_ (
    .A1(_07356_),
    .A2(_07358_),
    .ZN(_07359_)
  );
  MUX2_X1 _14955_ (
    .A(\rf[15] [11]),
    .B(\rf[11] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07360_)
  );
  AND2_X1 _14956_ (
    .A1(_03048_),
    .A2(_07360_),
    .ZN(_07361_)
  );
  OR2_X1 _14957_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07361_),
    .ZN(_07362_)
  );
  OR2_X1 _14958_ (
    .A1(_07359_),
    .A2(_07362_),
    .ZN(_07363_)
  );
  OR2_X1 _14959_ (
    .A1(\rf[12] [11]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07364_)
  );
  OR2_X1 _14960_ (
    .A1(\rf[8] [11]),
    .A2(_03050_),
    .ZN(_07365_)
  );
  AND2_X1 _14961_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07364_),
    .ZN(_07366_)
  );
  AND2_X1 _14962_ (
    .A1(_07365_),
    .A2(_07366_),
    .ZN(_07367_)
  );
  MUX2_X1 _14963_ (
    .A(\rf[13] [11]),
    .B(\rf[9] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07368_)
  );
  AND2_X1 _14964_ (
    .A1(_03048_),
    .A2(_07368_),
    .ZN(_07369_)
  );
  OR2_X1 _14965_ (
    .A1(_03049_),
    .A2(_07369_),
    .ZN(_07370_)
  );
  OR2_X1 _14966_ (
    .A1(_07367_),
    .A2(_07370_),
    .ZN(_07371_)
  );
  AND2_X1 _14967_ (
    .A1(_03051_),
    .A2(_07371_),
    .ZN(_07372_)
  );
  AND2_X1 _14968_ (
    .A1(_07363_),
    .A2(_07372_),
    .ZN(_07373_)
  );
  MUX2_X1 _14969_ (
    .A(\rf[6] [11]),
    .B(\rf[2] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07374_)
  );
  AND2_X1 _14970_ (
    .A1(_03049_),
    .A2(_07374_),
    .ZN(_07375_)
  );
  MUX2_X1 _14971_ (
    .A(\rf[4] [11]),
    .B(\rf[0] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07376_)
  );
  AND2_X1 _14972_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07376_),
    .ZN(_07377_)
  );
  OR2_X1 _14973_ (
    .A1(_03048_),
    .A2(_07377_),
    .ZN(_07378_)
  );
  OR2_X1 _14974_ (
    .A1(_07375_),
    .A2(_07378_),
    .ZN(_07379_)
  );
  MUX2_X1 _14975_ (
    .A(\rf[7] [11]),
    .B(\rf[3] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07380_)
  );
  AND2_X1 _14976_ (
    .A1(_03049_),
    .A2(_07380_),
    .ZN(_07381_)
  );
  MUX2_X1 _14977_ (
    .A(\rf[5] [11]),
    .B(\rf[1] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07382_)
  );
  AND2_X1 _14978_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07382_),
    .ZN(_07383_)
  );
  OR2_X1 _14979_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07383_),
    .ZN(_07384_)
  );
  OR2_X1 _14980_ (
    .A1(_07381_),
    .A2(_07384_),
    .ZN(_07385_)
  );
  AND2_X1 _14981_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_07385_),
    .ZN(_07386_)
  );
  AND2_X1 _14982_ (
    .A1(_07379_),
    .A2(_07386_),
    .ZN(_07387_)
  );
  OR2_X1 _14983_ (
    .A1(_07373_),
    .A2(_07387_),
    .ZN(_07388_)
  );
  OR2_X1 _14984_ (
    .A1(\rf[17] [11]),
    .A2(_03050_),
    .ZN(_07389_)
  );
  OR2_X1 _14985_ (
    .A1(\rf[21] [11]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07390_)
  );
  AND2_X1 _14986_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07390_),
    .ZN(_07391_)
  );
  AND2_X1 _14987_ (
    .A1(_07389_),
    .A2(_07391_),
    .ZN(_07392_)
  );
  MUX2_X1 _14988_ (
    .A(\rf[23] [11]),
    .B(\rf[19] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07393_)
  );
  AND2_X1 _14989_ (
    .A1(_03049_),
    .A2(_07393_),
    .ZN(_07394_)
  );
  OR2_X1 _14990_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07394_),
    .ZN(_07395_)
  );
  OR2_X1 _14991_ (
    .A1(_07392_),
    .A2(_07395_),
    .ZN(_07396_)
  );
  OR2_X1 _14992_ (
    .A1(\rf[20] [11]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07397_)
  );
  OR2_X1 _14993_ (
    .A1(\rf[16] [11]),
    .A2(_03050_),
    .ZN(_07398_)
  );
  AND2_X1 _14994_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07398_),
    .ZN(_07399_)
  );
  AND2_X1 _14995_ (
    .A1(_07397_),
    .A2(_07399_),
    .ZN(_07400_)
  );
  MUX2_X1 _14996_ (
    .A(\rf[22] [11]),
    .B(\rf[18] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07401_)
  );
  AND2_X1 _14997_ (
    .A1(_03049_),
    .A2(_07401_),
    .ZN(_07402_)
  );
  OR2_X1 _14998_ (
    .A1(_03048_),
    .A2(_07402_),
    .ZN(_07403_)
  );
  OR2_X1 _14999_ (
    .A1(_07400_),
    .A2(_07403_),
    .ZN(_07404_)
  );
  AND2_X1 _15000_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_07396_),
    .ZN(_07405_)
  );
  AND2_X1 _15001_ (
    .A1(_07404_),
    .A2(_07405_),
    .ZN(_07406_)
  );
  OR2_X1 _15002_ (
    .A1(\rf[28] [11]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07407_)
  );
  OR2_X1 _15003_ (
    .A1(\rf[24] [11]),
    .A2(_03050_),
    .ZN(_07408_)
  );
  AND2_X1 _15004_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07407_),
    .ZN(_07409_)
  );
  AND2_X1 _15005_ (
    .A1(_07408_),
    .A2(_07409_),
    .ZN(_07410_)
  );
  MUX2_X1 _15006_ (
    .A(\rf[30] [11]),
    .B(\rf[26] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07411_)
  );
  AND2_X1 _15007_ (
    .A1(_03049_),
    .A2(_07411_),
    .ZN(_07412_)
  );
  OR2_X1 _15008_ (
    .A1(_03048_),
    .A2(_07412_),
    .ZN(_07413_)
  );
  OR2_X1 _15009_ (
    .A1(_07410_),
    .A2(_07413_),
    .ZN(_07414_)
  );
  MUX2_X1 _15010_ (
    .A(\rf[29] [11]),
    .B(\rf[25] [11]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07415_)
  );
  AND2_X1 _15011_ (
    .A1(\rf[27] [11]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07416_)
  );
  MUX2_X1 _15012_ (
    .A(_07415_),
    .B(_07416_),
    .S(_03049_),
    .Z(_07417_)
  );
  OR2_X1 _15013_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07417_),
    .ZN(_07418_)
  );
  AND2_X1 _15014_ (
    .A1(_03051_),
    .A2(_07418_),
    .ZN(_07419_)
  );
  AND2_X1 _15015_ (
    .A1(_07414_),
    .A2(_07419_),
    .ZN(_07420_)
  );
  OR2_X1 _15016_ (
    .A1(_07406_),
    .A2(_07420_),
    .ZN(_07421_)
  );
  MUX2_X1 _15017_ (
    .A(_07388_),
    .B(_07421_),
    .S(_03064_),
    .Z(_07422_)
  );
  MUX2_X1 _15018_ (
    .A(_07422_),
    .B(_04742_),
    .S(_06791_),
    .Z(_07423_)
  );
  MUX2_X1 _15019_ (
    .A(ex_reg_rs_msb_1[9]),
    .B(_07423_),
    .S(_06781_),
    .Z(_00158_)
  );
  MUX2_X1 _15020_ (
    .A(\rf[7] [12]),
    .B(\rf[3] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07424_)
  );
  AND2_X1 _15021_ (
    .A1(_03049_),
    .A2(_07424_),
    .ZN(_07425_)
  );
  MUX2_X1 _15022_ (
    .A(\rf[5] [12]),
    .B(\rf[1] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07426_)
  );
  AND2_X1 _15023_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07426_),
    .ZN(_07427_)
  );
  OR2_X1 _15024_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07427_),
    .ZN(_07428_)
  );
  OR2_X1 _15025_ (
    .A1(_07425_),
    .A2(_07428_),
    .ZN(_07429_)
  );
  MUX2_X1 _15026_ (
    .A(\rf[6] [12]),
    .B(\rf[2] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07430_)
  );
  AND2_X1 _15027_ (
    .A1(_03049_),
    .A2(_07430_),
    .ZN(_07431_)
  );
  MUX2_X1 _15028_ (
    .A(\rf[4] [12]),
    .B(\rf[0] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07432_)
  );
  AND2_X1 _15029_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07432_),
    .ZN(_07433_)
  );
  OR2_X1 _15030_ (
    .A1(_03048_),
    .A2(_07433_),
    .ZN(_07434_)
  );
  OR2_X1 _15031_ (
    .A1(_07431_),
    .A2(_07434_),
    .ZN(_07435_)
  );
  AND2_X1 _15032_ (
    .A1(_07429_),
    .A2(_07435_),
    .ZN(_07436_)
  );
  AND2_X1 _15033_ (
    .A1(\rf[14] [12]),
    .A2(_03049_),
    .ZN(_07437_)
  );
  AND2_X1 _15034_ (
    .A1(\rf[12] [12]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_07438_)
  );
  OR2_X1 _15035_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[2]),
    .A2(_07438_),
    .ZN(_07439_)
  );
  OR2_X1 _15036_ (
    .A1(_07437_),
    .A2(_07439_),
    .ZN(_07440_)
  );
  AND2_X1 _15037_ (
    .A1(\rf[10] [12]),
    .A2(_03049_),
    .ZN(_07441_)
  );
  AND2_X1 _15038_ (
    .A1(\rf[8] [12]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_07442_)
  );
  OR2_X1 _15039_ (
    .A1(_03050_),
    .A2(_07442_),
    .ZN(_07443_)
  );
  OR2_X1 _15040_ (
    .A1(_07441_),
    .A2(_07443_),
    .ZN(_07444_)
  );
  AND2_X1 _15041_ (
    .A1(_07440_),
    .A2(_07444_),
    .ZN(_07445_)
  );
  AND2_X1 _15042_ (
    .A1(\rf[15] [12]),
    .A2(_03049_),
    .ZN(_07446_)
  );
  AND2_X1 _15043_ (
    .A1(\rf[13] [12]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_07447_)
  );
  OR2_X1 _15044_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[2]),
    .A2(_07447_),
    .ZN(_07448_)
  );
  OR2_X1 _15045_ (
    .A1(_07446_),
    .A2(_07448_),
    .ZN(_07449_)
  );
  AND2_X1 _15046_ (
    .A1(\rf[11] [12]),
    .A2(_03049_),
    .ZN(_07450_)
  );
  AND2_X1 _15047_ (
    .A1(\rf[9] [12]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_07451_)
  );
  OR2_X1 _15048_ (
    .A1(_03050_),
    .A2(_07451_),
    .ZN(_07452_)
  );
  OR2_X1 _15049_ (
    .A1(_07450_),
    .A2(_07452_),
    .ZN(_07453_)
  );
  AND2_X1 _15050_ (
    .A1(_07449_),
    .A2(_07453_),
    .ZN(_07454_)
  );
  MUX2_X1 _15051_ (
    .A(_07445_),
    .B(_07454_),
    .S(_03048_),
    .Z(_07455_)
  );
  MUX2_X1 _15052_ (
    .A(_07436_),
    .B(_07455_),
    .S(_03051_),
    .Z(_07456_)
  );
  OR2_X1 _15053_ (
    .A1(\rf[28] [12]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07457_)
  );
  OR2_X1 _15054_ (
    .A1(\rf[24] [12]),
    .A2(_03050_),
    .ZN(_07458_)
  );
  AND2_X1 _15055_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07457_),
    .ZN(_07459_)
  );
  AND2_X1 _15056_ (
    .A1(_07458_),
    .A2(_07459_),
    .ZN(_07460_)
  );
  MUX2_X1 _15057_ (
    .A(\rf[30] [12]),
    .B(\rf[26] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07461_)
  );
  AND2_X1 _15058_ (
    .A1(_03049_),
    .A2(_07461_),
    .ZN(_07462_)
  );
  OR2_X1 _15059_ (
    .A1(_03048_),
    .A2(_07462_),
    .ZN(_07463_)
  );
  OR2_X1 _15060_ (
    .A1(_07460_),
    .A2(_07463_),
    .ZN(_07464_)
  );
  MUX2_X1 _15061_ (
    .A(\rf[29] [12]),
    .B(\rf[25] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07465_)
  );
  AND2_X1 _15062_ (
    .A1(\rf[27] [12]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07466_)
  );
  MUX2_X1 _15063_ (
    .A(_07465_),
    .B(_07466_),
    .S(_03049_),
    .Z(_07467_)
  );
  OR2_X1 _15064_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07467_),
    .ZN(_07468_)
  );
  AND2_X1 _15065_ (
    .A1(_07464_),
    .A2(_07468_),
    .ZN(_07469_)
  );
  OR2_X1 _15066_ (
    .A1(\rf[20] [12]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07470_)
  );
  OR2_X1 _15067_ (
    .A1(\rf[16] [12]),
    .A2(_03050_),
    .ZN(_07471_)
  );
  AND2_X1 _15068_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07471_),
    .ZN(_07472_)
  );
  AND2_X1 _15069_ (
    .A1(_07470_),
    .A2(_07472_),
    .ZN(_07473_)
  );
  MUX2_X1 _15070_ (
    .A(\rf[22] [12]),
    .B(\rf[18] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07474_)
  );
  AND2_X1 _15071_ (
    .A1(_03049_),
    .A2(_07474_),
    .ZN(_07475_)
  );
  OR2_X1 _15072_ (
    .A1(_03048_),
    .A2(_07475_),
    .ZN(_07476_)
  );
  OR2_X1 _15073_ (
    .A1(_07473_),
    .A2(_07476_),
    .ZN(_07477_)
  );
  OR2_X1 _15074_ (
    .A1(\rf[17] [12]),
    .A2(_03050_),
    .ZN(_07478_)
  );
  OR2_X1 _15075_ (
    .A1(\rf[21] [12]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07479_)
  );
  AND2_X1 _15076_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07479_),
    .ZN(_07480_)
  );
  AND2_X1 _15077_ (
    .A1(_07478_),
    .A2(_07480_),
    .ZN(_07481_)
  );
  MUX2_X1 _15078_ (
    .A(\rf[23] [12]),
    .B(\rf[19] [12]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07482_)
  );
  AND2_X1 _15079_ (
    .A1(_03049_),
    .A2(_07482_),
    .ZN(_07483_)
  );
  OR2_X1 _15080_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07483_),
    .ZN(_07484_)
  );
  OR2_X1 _15081_ (
    .A1(_07481_),
    .A2(_07484_),
    .ZN(_07485_)
  );
  AND2_X1 _15082_ (
    .A1(_07477_),
    .A2(_07485_),
    .ZN(_07486_)
  );
  MUX2_X1 _15083_ (
    .A(_07469_),
    .B(_07486_),
    .S(ibuf_io_inst_0_bits_inst_rs2[3]),
    .Z(_07487_)
  );
  MUX2_X1 _15084_ (
    .A(_07456_),
    .B(_07487_),
    .S(_03064_),
    .Z(_07488_)
  );
  MUX2_X1 _15085_ (
    .A(_07488_),
    .B(_04811_),
    .S(_06791_),
    .Z(_07489_)
  );
  MUX2_X1 _15086_ (
    .A(ex_reg_rs_msb_1[10]),
    .B(_07489_),
    .S(_06781_),
    .Z(_00159_)
  );
  MUX2_X1 _15087_ (
    .A(\rf[7] [13]),
    .B(\rf[3] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07490_)
  );
  AND2_X1 _15088_ (
    .A1(_03049_),
    .A2(_07490_),
    .ZN(_07491_)
  );
  MUX2_X1 _15089_ (
    .A(\rf[5] [13]),
    .B(\rf[1] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07492_)
  );
  AND2_X1 _15090_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07492_),
    .ZN(_07493_)
  );
  OR2_X1 _15091_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07493_),
    .ZN(_07494_)
  );
  OR2_X1 _15092_ (
    .A1(_07491_),
    .A2(_07494_),
    .ZN(_07495_)
  );
  MUX2_X1 _15093_ (
    .A(\rf[6] [13]),
    .B(\rf[2] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07496_)
  );
  AND2_X1 _15094_ (
    .A1(_03049_),
    .A2(_07496_),
    .ZN(_07497_)
  );
  MUX2_X1 _15095_ (
    .A(\rf[4] [13]),
    .B(\rf[0] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07498_)
  );
  AND2_X1 _15096_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07498_),
    .ZN(_07499_)
  );
  OR2_X1 _15097_ (
    .A1(_03048_),
    .A2(_07499_),
    .ZN(_07500_)
  );
  OR2_X1 _15098_ (
    .A1(_07497_),
    .A2(_07500_),
    .ZN(_07501_)
  );
  AND2_X1 _15099_ (
    .A1(_07495_),
    .A2(_07501_),
    .ZN(_07502_)
  );
  AND2_X1 _15100_ (
    .A1(\rf[14] [13]),
    .A2(_03049_),
    .ZN(_07503_)
  );
  AND2_X1 _15101_ (
    .A1(\rf[12] [13]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_07504_)
  );
  OR2_X1 _15102_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[2]),
    .A2(_07504_),
    .ZN(_07505_)
  );
  OR2_X1 _15103_ (
    .A1(_07503_),
    .A2(_07505_),
    .ZN(_07506_)
  );
  AND2_X1 _15104_ (
    .A1(\rf[10] [13]),
    .A2(_03049_),
    .ZN(_07507_)
  );
  AND2_X1 _15105_ (
    .A1(\rf[8] [13]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_07508_)
  );
  OR2_X1 _15106_ (
    .A1(_03050_),
    .A2(_07508_),
    .ZN(_07509_)
  );
  OR2_X1 _15107_ (
    .A1(_07507_),
    .A2(_07509_),
    .ZN(_07510_)
  );
  AND2_X1 _15108_ (
    .A1(_07506_),
    .A2(_07510_),
    .ZN(_07511_)
  );
  AND2_X1 _15109_ (
    .A1(\rf[15] [13]),
    .A2(_03049_),
    .ZN(_07512_)
  );
  AND2_X1 _15110_ (
    .A1(\rf[13] [13]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_07513_)
  );
  OR2_X1 _15111_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[2]),
    .A2(_07513_),
    .ZN(_07514_)
  );
  OR2_X1 _15112_ (
    .A1(_07512_),
    .A2(_07514_),
    .ZN(_07515_)
  );
  AND2_X1 _15113_ (
    .A1(\rf[11] [13]),
    .A2(_03049_),
    .ZN(_07516_)
  );
  AND2_X1 _15114_ (
    .A1(\rf[9] [13]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_07517_)
  );
  OR2_X1 _15115_ (
    .A1(_03050_),
    .A2(_07517_),
    .ZN(_07518_)
  );
  OR2_X1 _15116_ (
    .A1(_07516_),
    .A2(_07518_),
    .ZN(_07519_)
  );
  AND2_X1 _15117_ (
    .A1(_07515_),
    .A2(_07519_),
    .ZN(_07520_)
  );
  MUX2_X1 _15118_ (
    .A(_07511_),
    .B(_07520_),
    .S(_03048_),
    .Z(_07521_)
  );
  MUX2_X1 _15119_ (
    .A(_07502_),
    .B(_07521_),
    .S(_03051_),
    .Z(_07522_)
  );
  OR2_X1 _15120_ (
    .A1(\rf[28] [13]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07523_)
  );
  OR2_X1 _15121_ (
    .A1(\rf[24] [13]),
    .A2(_03050_),
    .ZN(_07524_)
  );
  AND2_X1 _15122_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07523_),
    .ZN(_07525_)
  );
  AND2_X1 _15123_ (
    .A1(_07524_),
    .A2(_07525_),
    .ZN(_07526_)
  );
  MUX2_X1 _15124_ (
    .A(\rf[30] [13]),
    .B(\rf[26] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07527_)
  );
  AND2_X1 _15125_ (
    .A1(_03049_),
    .A2(_07527_),
    .ZN(_07528_)
  );
  OR2_X1 _15126_ (
    .A1(_03048_),
    .A2(_07528_),
    .ZN(_07529_)
  );
  OR2_X1 _15127_ (
    .A1(_07526_),
    .A2(_07529_),
    .ZN(_07530_)
  );
  MUX2_X1 _15128_ (
    .A(\rf[29] [13]),
    .B(\rf[25] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07531_)
  );
  AND2_X1 _15129_ (
    .A1(\rf[27] [13]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07532_)
  );
  MUX2_X1 _15130_ (
    .A(_07531_),
    .B(_07532_),
    .S(_03049_),
    .Z(_07533_)
  );
  OR2_X1 _15131_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07533_),
    .ZN(_07534_)
  );
  AND2_X1 _15132_ (
    .A1(_07530_),
    .A2(_07534_),
    .ZN(_07535_)
  );
  OR2_X1 _15133_ (
    .A1(\rf[20] [13]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07536_)
  );
  OR2_X1 _15134_ (
    .A1(\rf[16] [13]),
    .A2(_03050_),
    .ZN(_07537_)
  );
  AND2_X1 _15135_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07537_),
    .ZN(_07538_)
  );
  AND2_X1 _15136_ (
    .A1(_07536_),
    .A2(_07538_),
    .ZN(_07539_)
  );
  MUX2_X1 _15137_ (
    .A(\rf[22] [13]),
    .B(\rf[18] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07540_)
  );
  AND2_X1 _15138_ (
    .A1(_03049_),
    .A2(_07540_),
    .ZN(_07541_)
  );
  OR2_X1 _15139_ (
    .A1(_03048_),
    .A2(_07541_),
    .ZN(_07542_)
  );
  OR2_X1 _15140_ (
    .A1(_07539_),
    .A2(_07542_),
    .ZN(_07543_)
  );
  OR2_X1 _15141_ (
    .A1(\rf[17] [13]),
    .A2(_03050_),
    .ZN(_07544_)
  );
  OR2_X1 _15142_ (
    .A1(\rf[21] [13]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07545_)
  );
  AND2_X1 _15143_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07545_),
    .ZN(_07546_)
  );
  AND2_X1 _15144_ (
    .A1(_07544_),
    .A2(_07546_),
    .ZN(_07547_)
  );
  MUX2_X1 _15145_ (
    .A(\rf[23] [13]),
    .B(\rf[19] [13]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07548_)
  );
  AND2_X1 _15146_ (
    .A1(_03049_),
    .A2(_07548_),
    .ZN(_07549_)
  );
  OR2_X1 _15147_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07549_),
    .ZN(_07550_)
  );
  OR2_X1 _15148_ (
    .A1(_07547_),
    .A2(_07550_),
    .ZN(_07551_)
  );
  AND2_X1 _15149_ (
    .A1(_07543_),
    .A2(_07551_),
    .ZN(_07552_)
  );
  MUX2_X1 _15150_ (
    .A(_07535_),
    .B(_07552_),
    .S(ibuf_io_inst_0_bits_inst_rs2[3]),
    .Z(_07553_)
  );
  MUX2_X1 _15151_ (
    .A(_07522_),
    .B(_07553_),
    .S(_03064_),
    .Z(_07554_)
  );
  MUX2_X1 _15152_ (
    .A(_07554_),
    .B(_04882_),
    .S(_06791_),
    .Z(_07555_)
  );
  MUX2_X1 _15153_ (
    .A(ex_reg_rs_msb_1[11]),
    .B(_07555_),
    .S(_06781_),
    .Z(_00160_)
  );
  OR2_X1 _15154_ (
    .A1(\rf[10] [14]),
    .A2(_03050_),
    .ZN(_07556_)
  );
  OR2_X1 _15155_ (
    .A1(\rf[14] [14]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07557_)
  );
  AND2_X1 _15156_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07557_),
    .ZN(_07558_)
  );
  AND2_X1 _15157_ (
    .A1(_07556_),
    .A2(_07558_),
    .ZN(_07559_)
  );
  MUX2_X1 _15158_ (
    .A(\rf[15] [14]),
    .B(\rf[11] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07560_)
  );
  AND2_X1 _15159_ (
    .A1(_03048_),
    .A2(_07560_),
    .ZN(_07561_)
  );
  OR2_X1 _15160_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07561_),
    .ZN(_07562_)
  );
  OR2_X1 _15161_ (
    .A1(_07559_),
    .A2(_07562_),
    .ZN(_07563_)
  );
  OR2_X1 _15162_ (
    .A1(\rf[12] [14]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07564_)
  );
  OR2_X1 _15163_ (
    .A1(\rf[8] [14]),
    .A2(_03050_),
    .ZN(_07565_)
  );
  AND2_X1 _15164_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07564_),
    .ZN(_07566_)
  );
  AND2_X1 _15165_ (
    .A1(_07565_),
    .A2(_07566_),
    .ZN(_07567_)
  );
  MUX2_X1 _15166_ (
    .A(\rf[13] [14]),
    .B(\rf[9] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07568_)
  );
  AND2_X1 _15167_ (
    .A1(_03048_),
    .A2(_07568_),
    .ZN(_07569_)
  );
  OR2_X1 _15168_ (
    .A1(_03049_),
    .A2(_07569_),
    .ZN(_07570_)
  );
  OR2_X1 _15169_ (
    .A1(_07567_),
    .A2(_07570_),
    .ZN(_07571_)
  );
  AND2_X1 _15170_ (
    .A1(_03051_),
    .A2(_07571_),
    .ZN(_07572_)
  );
  AND2_X1 _15171_ (
    .A1(_07563_),
    .A2(_07572_),
    .ZN(_07573_)
  );
  MUX2_X1 _15172_ (
    .A(\rf[6] [14]),
    .B(\rf[2] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07574_)
  );
  AND2_X1 _15173_ (
    .A1(_03049_),
    .A2(_07574_),
    .ZN(_07575_)
  );
  MUX2_X1 _15174_ (
    .A(\rf[4] [14]),
    .B(\rf[0] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07576_)
  );
  AND2_X1 _15175_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07576_),
    .ZN(_07577_)
  );
  OR2_X1 _15176_ (
    .A1(_03048_),
    .A2(_07577_),
    .ZN(_07578_)
  );
  OR2_X1 _15177_ (
    .A1(_07575_),
    .A2(_07578_),
    .ZN(_07579_)
  );
  MUX2_X1 _15178_ (
    .A(\rf[7] [14]),
    .B(\rf[3] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07580_)
  );
  AND2_X1 _15179_ (
    .A1(_03049_),
    .A2(_07580_),
    .ZN(_07581_)
  );
  MUX2_X1 _15180_ (
    .A(\rf[5] [14]),
    .B(\rf[1] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07582_)
  );
  AND2_X1 _15181_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07582_),
    .ZN(_07583_)
  );
  OR2_X1 _15182_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07583_),
    .ZN(_07584_)
  );
  OR2_X1 _15183_ (
    .A1(_07581_),
    .A2(_07584_),
    .ZN(_07585_)
  );
  AND2_X1 _15184_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_07585_),
    .ZN(_07586_)
  );
  AND2_X1 _15185_ (
    .A1(_07579_),
    .A2(_07586_),
    .ZN(_07587_)
  );
  OR2_X1 _15186_ (
    .A1(_07573_),
    .A2(_07587_),
    .ZN(_07588_)
  );
  OR2_X1 _15187_ (
    .A1(\rf[17] [14]),
    .A2(_03050_),
    .ZN(_07589_)
  );
  OR2_X1 _15188_ (
    .A1(\rf[21] [14]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07590_)
  );
  AND2_X1 _15189_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07590_),
    .ZN(_07591_)
  );
  AND2_X1 _15190_ (
    .A1(_07589_),
    .A2(_07591_),
    .ZN(_07592_)
  );
  MUX2_X1 _15191_ (
    .A(\rf[23] [14]),
    .B(\rf[19] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07593_)
  );
  AND2_X1 _15192_ (
    .A1(_03049_),
    .A2(_07593_),
    .ZN(_07594_)
  );
  OR2_X1 _15193_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07594_),
    .ZN(_07595_)
  );
  OR2_X1 _15194_ (
    .A1(_07592_),
    .A2(_07595_),
    .ZN(_07596_)
  );
  OR2_X1 _15195_ (
    .A1(\rf[20] [14]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07597_)
  );
  OR2_X1 _15196_ (
    .A1(\rf[16] [14]),
    .A2(_03050_),
    .ZN(_07598_)
  );
  AND2_X1 _15197_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07598_),
    .ZN(_07599_)
  );
  AND2_X1 _15198_ (
    .A1(_07597_),
    .A2(_07599_),
    .ZN(_07600_)
  );
  MUX2_X1 _15199_ (
    .A(\rf[22] [14]),
    .B(\rf[18] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07601_)
  );
  AND2_X1 _15200_ (
    .A1(_03049_),
    .A2(_07601_),
    .ZN(_07602_)
  );
  OR2_X1 _15201_ (
    .A1(_03048_),
    .A2(_07602_),
    .ZN(_07603_)
  );
  OR2_X1 _15202_ (
    .A1(_07600_),
    .A2(_07603_),
    .ZN(_07604_)
  );
  AND2_X1 _15203_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_07596_),
    .ZN(_07605_)
  );
  AND2_X1 _15204_ (
    .A1(_07604_),
    .A2(_07605_),
    .ZN(_07606_)
  );
  OR2_X1 _15205_ (
    .A1(\rf[28] [14]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07607_)
  );
  OR2_X1 _15206_ (
    .A1(\rf[24] [14]),
    .A2(_03050_),
    .ZN(_07608_)
  );
  AND2_X1 _15207_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07607_),
    .ZN(_07609_)
  );
  AND2_X1 _15208_ (
    .A1(_07608_),
    .A2(_07609_),
    .ZN(_07610_)
  );
  MUX2_X1 _15209_ (
    .A(\rf[30] [14]),
    .B(\rf[26] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07611_)
  );
  AND2_X1 _15210_ (
    .A1(_03049_),
    .A2(_07611_),
    .ZN(_07612_)
  );
  OR2_X1 _15211_ (
    .A1(_03048_),
    .A2(_07612_),
    .ZN(_07613_)
  );
  OR2_X1 _15212_ (
    .A1(_07610_),
    .A2(_07613_),
    .ZN(_07614_)
  );
  MUX2_X1 _15213_ (
    .A(\rf[29] [14]),
    .B(\rf[25] [14]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07615_)
  );
  AND2_X1 _15214_ (
    .A1(\rf[27] [14]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07616_)
  );
  MUX2_X1 _15215_ (
    .A(_07615_),
    .B(_07616_),
    .S(_03049_),
    .Z(_07617_)
  );
  OR2_X1 _15216_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07617_),
    .ZN(_07618_)
  );
  AND2_X1 _15217_ (
    .A1(_03051_),
    .A2(_07618_),
    .ZN(_07619_)
  );
  AND2_X1 _15218_ (
    .A1(_07614_),
    .A2(_07619_),
    .ZN(_07620_)
  );
  OR2_X1 _15219_ (
    .A1(_07606_),
    .A2(_07620_),
    .ZN(_07621_)
  );
  MUX2_X1 _15220_ (
    .A(_07588_),
    .B(_07621_),
    .S(_03064_),
    .Z(_07622_)
  );
  MUX2_X1 _15221_ (
    .A(_07622_),
    .B(_04953_),
    .S(_06791_),
    .Z(_07623_)
  );
  MUX2_X1 _15222_ (
    .A(ex_reg_rs_msb_1[12]),
    .B(_07623_),
    .S(_06781_),
    .Z(_00161_)
  );
  MUX2_X1 _15223_ (
    .A(\rf[7] [15]),
    .B(\rf[3] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07624_)
  );
  AND2_X1 _15224_ (
    .A1(_03049_),
    .A2(_07624_),
    .ZN(_07625_)
  );
  MUX2_X1 _15225_ (
    .A(\rf[5] [15]),
    .B(\rf[1] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07626_)
  );
  AND2_X1 _15226_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07626_),
    .ZN(_07627_)
  );
  OR2_X1 _15227_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07627_),
    .ZN(_07628_)
  );
  OR2_X1 _15228_ (
    .A1(_07625_),
    .A2(_07628_),
    .ZN(_07629_)
  );
  MUX2_X1 _15229_ (
    .A(\rf[6] [15]),
    .B(\rf[2] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07630_)
  );
  AND2_X1 _15230_ (
    .A1(_03049_),
    .A2(_07630_),
    .ZN(_07631_)
  );
  MUX2_X1 _15231_ (
    .A(\rf[4] [15]),
    .B(\rf[0] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07632_)
  );
  AND2_X1 _15232_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07632_),
    .ZN(_07633_)
  );
  OR2_X1 _15233_ (
    .A1(_03048_),
    .A2(_07633_),
    .ZN(_07634_)
  );
  OR2_X1 _15234_ (
    .A1(_07631_),
    .A2(_07634_),
    .ZN(_07635_)
  );
  AND2_X1 _15235_ (
    .A1(_07629_),
    .A2(_07635_),
    .ZN(_07636_)
  );
  AND2_X1 _15236_ (
    .A1(\rf[14] [15]),
    .A2(_03049_),
    .ZN(_07637_)
  );
  AND2_X1 _15237_ (
    .A1(\rf[12] [15]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_07638_)
  );
  OR2_X1 _15238_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[2]),
    .A2(_07638_),
    .ZN(_07639_)
  );
  OR2_X1 _15239_ (
    .A1(_07637_),
    .A2(_07639_),
    .ZN(_07640_)
  );
  AND2_X1 _15240_ (
    .A1(\rf[10] [15]),
    .A2(_03049_),
    .ZN(_07641_)
  );
  AND2_X1 _15241_ (
    .A1(\rf[8] [15]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_07642_)
  );
  OR2_X1 _15242_ (
    .A1(_03050_),
    .A2(_07642_),
    .ZN(_07643_)
  );
  OR2_X1 _15243_ (
    .A1(_07641_),
    .A2(_07643_),
    .ZN(_07644_)
  );
  AND2_X1 _15244_ (
    .A1(_07640_),
    .A2(_07644_),
    .ZN(_07645_)
  );
  AND2_X1 _15245_ (
    .A1(\rf[15] [15]),
    .A2(_03049_),
    .ZN(_07646_)
  );
  AND2_X1 _15246_ (
    .A1(\rf[13] [15]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_07647_)
  );
  OR2_X1 _15247_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[2]),
    .A2(_07647_),
    .ZN(_07648_)
  );
  OR2_X1 _15248_ (
    .A1(_07646_),
    .A2(_07648_),
    .ZN(_07649_)
  );
  AND2_X1 _15249_ (
    .A1(\rf[11] [15]),
    .A2(_03049_),
    .ZN(_07650_)
  );
  AND2_X1 _15250_ (
    .A1(\rf[9] [15]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_07651_)
  );
  OR2_X1 _15251_ (
    .A1(_03050_),
    .A2(_07651_),
    .ZN(_07652_)
  );
  OR2_X1 _15252_ (
    .A1(_07650_),
    .A2(_07652_),
    .ZN(_07653_)
  );
  AND2_X1 _15253_ (
    .A1(_07649_),
    .A2(_07653_),
    .ZN(_07654_)
  );
  MUX2_X1 _15254_ (
    .A(_07645_),
    .B(_07654_),
    .S(_03048_),
    .Z(_07655_)
  );
  MUX2_X1 _15255_ (
    .A(_07636_),
    .B(_07655_),
    .S(_03051_),
    .Z(_07656_)
  );
  OR2_X1 _15256_ (
    .A1(\rf[28] [15]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07657_)
  );
  OR2_X1 _15257_ (
    .A1(\rf[24] [15]),
    .A2(_03050_),
    .ZN(_07658_)
  );
  AND2_X1 _15258_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07657_),
    .ZN(_07659_)
  );
  AND2_X1 _15259_ (
    .A1(_07658_),
    .A2(_07659_),
    .ZN(_07660_)
  );
  MUX2_X1 _15260_ (
    .A(\rf[30] [15]),
    .B(\rf[26] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07661_)
  );
  AND2_X1 _15261_ (
    .A1(_03049_),
    .A2(_07661_),
    .ZN(_07662_)
  );
  OR2_X1 _15262_ (
    .A1(_03048_),
    .A2(_07662_),
    .ZN(_07663_)
  );
  OR2_X1 _15263_ (
    .A1(_07660_),
    .A2(_07663_),
    .ZN(_07664_)
  );
  MUX2_X1 _15264_ (
    .A(\rf[29] [15]),
    .B(\rf[25] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07665_)
  );
  AND2_X1 _15265_ (
    .A1(\rf[27] [15]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07666_)
  );
  MUX2_X1 _15266_ (
    .A(_07665_),
    .B(_07666_),
    .S(_03049_),
    .Z(_07667_)
  );
  OR2_X1 _15267_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07667_),
    .ZN(_07668_)
  );
  AND2_X1 _15268_ (
    .A1(_07664_),
    .A2(_07668_),
    .ZN(_07669_)
  );
  OR2_X1 _15269_ (
    .A1(\rf[20] [15]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07670_)
  );
  OR2_X1 _15270_ (
    .A1(\rf[16] [15]),
    .A2(_03050_),
    .ZN(_07671_)
  );
  AND2_X1 _15271_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07671_),
    .ZN(_07672_)
  );
  AND2_X1 _15272_ (
    .A1(_07670_),
    .A2(_07672_),
    .ZN(_07673_)
  );
  MUX2_X1 _15273_ (
    .A(\rf[22] [15]),
    .B(\rf[18] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07674_)
  );
  AND2_X1 _15274_ (
    .A1(_03049_),
    .A2(_07674_),
    .ZN(_07675_)
  );
  OR2_X1 _15275_ (
    .A1(_03048_),
    .A2(_07675_),
    .ZN(_07676_)
  );
  OR2_X1 _15276_ (
    .A1(_07673_),
    .A2(_07676_),
    .ZN(_07677_)
  );
  OR2_X1 _15277_ (
    .A1(\rf[17] [15]),
    .A2(_03050_),
    .ZN(_07678_)
  );
  OR2_X1 _15278_ (
    .A1(\rf[21] [15]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07679_)
  );
  AND2_X1 _15279_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07679_),
    .ZN(_07680_)
  );
  AND2_X1 _15280_ (
    .A1(_07678_),
    .A2(_07680_),
    .ZN(_07681_)
  );
  MUX2_X1 _15281_ (
    .A(\rf[23] [15]),
    .B(\rf[19] [15]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07682_)
  );
  AND2_X1 _15282_ (
    .A1(_03049_),
    .A2(_07682_),
    .ZN(_07683_)
  );
  OR2_X1 _15283_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07683_),
    .ZN(_07684_)
  );
  OR2_X1 _15284_ (
    .A1(_07681_),
    .A2(_07684_),
    .ZN(_07685_)
  );
  AND2_X1 _15285_ (
    .A1(_07677_),
    .A2(_07685_),
    .ZN(_07686_)
  );
  MUX2_X1 _15286_ (
    .A(_07669_),
    .B(_07686_),
    .S(ibuf_io_inst_0_bits_inst_rs2[3]),
    .Z(_07687_)
  );
  MUX2_X1 _15287_ (
    .A(_07656_),
    .B(_07687_),
    .S(_03064_),
    .Z(_07688_)
  );
  MUX2_X1 _15288_ (
    .A(_07688_),
    .B(_05027_),
    .S(_06791_),
    .Z(_07689_)
  );
  MUX2_X1 _15289_ (
    .A(ex_reg_rs_msb_1[13]),
    .B(_07689_),
    .S(_06781_),
    .Z(_00162_)
  );
  MUX2_X1 _15290_ (
    .A(\rf[1] [16]),
    .B(\rf[0] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_07690_)
  );
  MUX2_X1 _15291_ (
    .A(\rf[5] [16]),
    .B(\rf[4] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_07691_)
  );
  MUX2_X1 _15292_ (
    .A(_07690_),
    .B(_07691_),
    .S(_03050_),
    .Z(_07692_)
  );
  OR2_X1 _15293_ (
    .A1(_03051_),
    .A2(_07692_),
    .ZN(_07693_)
  );
  MUX2_X1 _15294_ (
    .A(\rf[12] [16]),
    .B(\rf[8] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07694_)
  );
  OR2_X1 _15295_ (
    .A1(_06863_),
    .A2(_07694_),
    .ZN(_07695_)
  );
  MUX2_X1 _15296_ (
    .A(\rf[13] [16]),
    .B(\rf[9] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07696_)
  );
  OR2_X1 _15297_ (
    .A1(_03808_),
    .A2(_07696_),
    .ZN(_07697_)
  );
  AND2_X1 _15298_ (
    .A1(_07695_),
    .A2(_07697_),
    .ZN(_07698_)
  );
  AND2_X1 _15299_ (
    .A1(_07693_),
    .A2(_07698_),
    .ZN(_07699_)
  );
  MUX2_X1 _15300_ (
    .A(\rf[3] [16]),
    .B(\rf[2] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_07700_)
  );
  MUX2_X1 _15301_ (
    .A(\rf[7] [16]),
    .B(\rf[6] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_07701_)
  );
  MUX2_X1 _15302_ (
    .A(_07700_),
    .B(_07701_),
    .S(_03050_),
    .Z(_07702_)
  );
  OR2_X1 _15303_ (
    .A1(_03051_),
    .A2(_07702_),
    .ZN(_07703_)
  );
  MUX2_X1 _15304_ (
    .A(\rf[14] [16]),
    .B(\rf[10] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07704_)
  );
  OR2_X1 _15305_ (
    .A1(_06863_),
    .A2(_07704_),
    .ZN(_07705_)
  );
  MUX2_X1 _15306_ (
    .A(\rf[15] [16]),
    .B(\rf[11] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07706_)
  );
  OR2_X1 _15307_ (
    .A1(_03808_),
    .A2(_07706_),
    .ZN(_07707_)
  );
  AND2_X1 _15308_ (
    .A1(_07705_),
    .A2(_07707_),
    .ZN(_07708_)
  );
  AND2_X1 _15309_ (
    .A1(_07703_),
    .A2(_07708_),
    .ZN(_07709_)
  );
  MUX2_X1 _15310_ (
    .A(_07699_),
    .B(_07709_),
    .S(_03049_),
    .Z(_07710_)
  );
  OR2_X1 _15311_ (
    .A1(\rf[17] [16]),
    .A2(_03050_),
    .ZN(_07711_)
  );
  OR2_X1 _15312_ (
    .A1(\rf[21] [16]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07712_)
  );
  AND2_X1 _15313_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07712_),
    .ZN(_07713_)
  );
  AND2_X1 _15314_ (
    .A1(_07711_),
    .A2(_07713_),
    .ZN(_07714_)
  );
  MUX2_X1 _15315_ (
    .A(\rf[23] [16]),
    .B(\rf[19] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07715_)
  );
  AND2_X1 _15316_ (
    .A1(_03049_),
    .A2(_07715_),
    .ZN(_07716_)
  );
  OR2_X1 _15317_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07716_),
    .ZN(_07717_)
  );
  OR2_X1 _15318_ (
    .A1(_07714_),
    .A2(_07717_),
    .ZN(_07718_)
  );
  OR2_X1 _15319_ (
    .A1(\rf[20] [16]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07719_)
  );
  OR2_X1 _15320_ (
    .A1(\rf[16] [16]),
    .A2(_03050_),
    .ZN(_07720_)
  );
  AND2_X1 _15321_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07720_),
    .ZN(_07721_)
  );
  AND2_X1 _15322_ (
    .A1(_07719_),
    .A2(_07721_),
    .ZN(_07722_)
  );
  MUX2_X1 _15323_ (
    .A(\rf[22] [16]),
    .B(\rf[18] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07723_)
  );
  AND2_X1 _15324_ (
    .A1(_03049_),
    .A2(_07723_),
    .ZN(_07724_)
  );
  OR2_X1 _15325_ (
    .A1(_03048_),
    .A2(_07724_),
    .ZN(_07725_)
  );
  OR2_X1 _15326_ (
    .A1(_07722_),
    .A2(_07725_),
    .ZN(_07726_)
  );
  AND2_X1 _15327_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_07718_),
    .ZN(_07727_)
  );
  AND2_X1 _15328_ (
    .A1(_07726_),
    .A2(_07727_),
    .ZN(_07728_)
  );
  OR2_X1 _15329_ (
    .A1(\rf[28] [16]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07729_)
  );
  OR2_X1 _15330_ (
    .A1(\rf[24] [16]),
    .A2(_03050_),
    .ZN(_07730_)
  );
  AND2_X1 _15331_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07729_),
    .ZN(_07731_)
  );
  AND2_X1 _15332_ (
    .A1(_07730_),
    .A2(_07731_),
    .ZN(_07732_)
  );
  MUX2_X1 _15333_ (
    .A(\rf[30] [16]),
    .B(\rf[26] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07733_)
  );
  AND2_X1 _15334_ (
    .A1(_03049_),
    .A2(_07733_),
    .ZN(_07734_)
  );
  OR2_X1 _15335_ (
    .A1(_03048_),
    .A2(_07734_),
    .ZN(_07735_)
  );
  OR2_X1 _15336_ (
    .A1(_07732_),
    .A2(_07735_),
    .ZN(_07736_)
  );
  MUX2_X1 _15337_ (
    .A(\rf[29] [16]),
    .B(\rf[25] [16]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07737_)
  );
  AND2_X1 _15338_ (
    .A1(\rf[27] [16]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07738_)
  );
  MUX2_X1 _15339_ (
    .A(_07737_),
    .B(_07738_),
    .S(_03049_),
    .Z(_07739_)
  );
  OR2_X1 _15340_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07739_),
    .ZN(_07740_)
  );
  AND2_X1 _15341_ (
    .A1(_03051_),
    .A2(_07740_),
    .ZN(_07741_)
  );
  AND2_X1 _15342_ (
    .A1(_07736_),
    .A2(_07741_),
    .ZN(_07742_)
  );
  OR2_X1 _15343_ (
    .A1(_07728_),
    .A2(_07742_),
    .ZN(_07743_)
  );
  MUX2_X1 _15344_ (
    .A(_07710_),
    .B(_07743_),
    .S(_03064_),
    .Z(_07744_)
  );
  MUX2_X1 _15345_ (
    .A(_07744_),
    .B(_05095_),
    .S(_06791_),
    .Z(_07745_)
  );
  MUX2_X1 _15346_ (
    .A(ex_reg_rs_msb_1[14]),
    .B(_07745_),
    .S(_06781_),
    .Z(_00163_)
  );
  MUX2_X1 _15347_ (
    .A(\rf[1] [17]),
    .B(\rf[0] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_07746_)
  );
  MUX2_X1 _15348_ (
    .A(\rf[5] [17]),
    .B(\rf[4] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_07747_)
  );
  MUX2_X1 _15349_ (
    .A(_07746_),
    .B(_07747_),
    .S(_03050_),
    .Z(_07748_)
  );
  OR2_X1 _15350_ (
    .A1(_03051_),
    .A2(_07748_),
    .ZN(_07749_)
  );
  MUX2_X1 _15351_ (
    .A(\rf[12] [17]),
    .B(\rf[8] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07750_)
  );
  OR2_X1 _15352_ (
    .A1(_06863_),
    .A2(_07750_),
    .ZN(_07751_)
  );
  MUX2_X1 _15353_ (
    .A(\rf[13] [17]),
    .B(\rf[9] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07752_)
  );
  OR2_X1 _15354_ (
    .A1(_03808_),
    .A2(_07752_),
    .ZN(_07753_)
  );
  AND2_X1 _15355_ (
    .A1(_07751_),
    .A2(_07753_),
    .ZN(_07754_)
  );
  AND2_X1 _15356_ (
    .A1(_07749_),
    .A2(_07754_),
    .ZN(_07755_)
  );
  MUX2_X1 _15357_ (
    .A(\rf[3] [17]),
    .B(\rf[2] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_07756_)
  );
  MUX2_X1 _15358_ (
    .A(\rf[7] [17]),
    .B(\rf[6] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_07757_)
  );
  MUX2_X1 _15359_ (
    .A(_07756_),
    .B(_07757_),
    .S(_03050_),
    .Z(_07758_)
  );
  OR2_X1 _15360_ (
    .A1(_03051_),
    .A2(_07758_),
    .ZN(_07759_)
  );
  MUX2_X1 _15361_ (
    .A(\rf[14] [17]),
    .B(\rf[10] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07760_)
  );
  OR2_X1 _15362_ (
    .A1(_06863_),
    .A2(_07760_),
    .ZN(_07761_)
  );
  MUX2_X1 _15363_ (
    .A(\rf[15] [17]),
    .B(\rf[11] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07762_)
  );
  OR2_X1 _15364_ (
    .A1(_03808_),
    .A2(_07762_),
    .ZN(_07763_)
  );
  AND2_X1 _15365_ (
    .A1(_07761_),
    .A2(_07763_),
    .ZN(_07764_)
  );
  AND2_X1 _15366_ (
    .A1(_07759_),
    .A2(_07764_),
    .ZN(_07765_)
  );
  MUX2_X1 _15367_ (
    .A(_07755_),
    .B(_07765_),
    .S(_03049_),
    .Z(_07766_)
  );
  OR2_X1 _15368_ (
    .A1(\rf[17] [17]),
    .A2(_03050_),
    .ZN(_07767_)
  );
  OR2_X1 _15369_ (
    .A1(\rf[21] [17]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07768_)
  );
  AND2_X1 _15370_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07768_),
    .ZN(_07769_)
  );
  AND2_X1 _15371_ (
    .A1(_07767_),
    .A2(_07769_),
    .ZN(_07770_)
  );
  MUX2_X1 _15372_ (
    .A(\rf[23] [17]),
    .B(\rf[19] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07771_)
  );
  AND2_X1 _15373_ (
    .A1(_03049_),
    .A2(_07771_),
    .ZN(_07772_)
  );
  OR2_X1 _15374_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07772_),
    .ZN(_07773_)
  );
  OR2_X1 _15375_ (
    .A1(_07770_),
    .A2(_07773_),
    .ZN(_07774_)
  );
  OR2_X1 _15376_ (
    .A1(\rf[20] [17]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07775_)
  );
  OR2_X1 _15377_ (
    .A1(\rf[16] [17]),
    .A2(_03050_),
    .ZN(_07776_)
  );
  AND2_X1 _15378_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07776_),
    .ZN(_07777_)
  );
  AND2_X1 _15379_ (
    .A1(_07775_),
    .A2(_07777_),
    .ZN(_07778_)
  );
  MUX2_X1 _15380_ (
    .A(\rf[22] [17]),
    .B(\rf[18] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07779_)
  );
  AND2_X1 _15381_ (
    .A1(_03049_),
    .A2(_07779_),
    .ZN(_07780_)
  );
  OR2_X1 _15382_ (
    .A1(_03048_),
    .A2(_07780_),
    .ZN(_07781_)
  );
  OR2_X1 _15383_ (
    .A1(_07778_),
    .A2(_07781_),
    .ZN(_07782_)
  );
  AND2_X1 _15384_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_07774_),
    .ZN(_07783_)
  );
  AND2_X1 _15385_ (
    .A1(_07782_),
    .A2(_07783_),
    .ZN(_07784_)
  );
  OR2_X1 _15386_ (
    .A1(\rf[28] [17]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07785_)
  );
  OR2_X1 _15387_ (
    .A1(\rf[24] [17]),
    .A2(_03050_),
    .ZN(_07786_)
  );
  AND2_X1 _15388_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07785_),
    .ZN(_07787_)
  );
  AND2_X1 _15389_ (
    .A1(_07786_),
    .A2(_07787_),
    .ZN(_07788_)
  );
  MUX2_X1 _15390_ (
    .A(\rf[30] [17]),
    .B(\rf[26] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07789_)
  );
  AND2_X1 _15391_ (
    .A1(_03049_),
    .A2(_07789_),
    .ZN(_07790_)
  );
  OR2_X1 _15392_ (
    .A1(_03048_),
    .A2(_07790_),
    .ZN(_07791_)
  );
  OR2_X1 _15393_ (
    .A1(_07788_),
    .A2(_07791_),
    .ZN(_07792_)
  );
  MUX2_X1 _15394_ (
    .A(\rf[29] [17]),
    .B(\rf[25] [17]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07793_)
  );
  AND2_X1 _15395_ (
    .A1(\rf[27] [17]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07794_)
  );
  MUX2_X1 _15396_ (
    .A(_07793_),
    .B(_07794_),
    .S(_03049_),
    .Z(_07795_)
  );
  OR2_X1 _15397_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07795_),
    .ZN(_07796_)
  );
  AND2_X1 _15398_ (
    .A1(_03051_),
    .A2(_07796_),
    .ZN(_07797_)
  );
  AND2_X1 _15399_ (
    .A1(_07792_),
    .A2(_07797_),
    .ZN(_07798_)
  );
  OR2_X1 _15400_ (
    .A1(_07784_),
    .A2(_07798_),
    .ZN(_07799_)
  );
  MUX2_X1 _15401_ (
    .A(_07766_),
    .B(_07799_),
    .S(_03064_),
    .Z(_07800_)
  );
  MUX2_X1 _15402_ (
    .A(_07800_),
    .B(_05170_),
    .S(_06791_),
    .Z(_07801_)
  );
  MUX2_X1 _15403_ (
    .A(ex_reg_rs_msb_1[15]),
    .B(_07801_),
    .S(_06781_),
    .Z(_00164_)
  );
  OR2_X1 _15404_ (
    .A1(\rf[10] [18]),
    .A2(_03050_),
    .ZN(_07802_)
  );
  OR2_X1 _15405_ (
    .A1(\rf[14] [18]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07803_)
  );
  AND2_X1 _15406_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07803_),
    .ZN(_07804_)
  );
  AND2_X1 _15407_ (
    .A1(_07802_),
    .A2(_07804_),
    .ZN(_07805_)
  );
  MUX2_X1 _15408_ (
    .A(\rf[15] [18]),
    .B(\rf[11] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07806_)
  );
  AND2_X1 _15409_ (
    .A1(_03048_),
    .A2(_07806_),
    .ZN(_07807_)
  );
  OR2_X1 _15410_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07807_),
    .ZN(_07808_)
  );
  OR2_X1 _15411_ (
    .A1(_07805_),
    .A2(_07808_),
    .ZN(_07809_)
  );
  OR2_X1 _15412_ (
    .A1(\rf[12] [18]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07810_)
  );
  OR2_X1 _15413_ (
    .A1(\rf[8] [18]),
    .A2(_03050_),
    .ZN(_07811_)
  );
  AND2_X1 _15414_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07810_),
    .ZN(_07812_)
  );
  AND2_X1 _15415_ (
    .A1(_07811_),
    .A2(_07812_),
    .ZN(_07813_)
  );
  MUX2_X1 _15416_ (
    .A(\rf[13] [18]),
    .B(\rf[9] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07814_)
  );
  AND2_X1 _15417_ (
    .A1(_03048_),
    .A2(_07814_),
    .ZN(_07815_)
  );
  OR2_X1 _15418_ (
    .A1(_03049_),
    .A2(_07815_),
    .ZN(_07816_)
  );
  OR2_X1 _15419_ (
    .A1(_07813_),
    .A2(_07816_),
    .ZN(_07817_)
  );
  AND2_X1 _15420_ (
    .A1(_03051_),
    .A2(_07817_),
    .ZN(_07818_)
  );
  AND2_X1 _15421_ (
    .A1(_07809_),
    .A2(_07818_),
    .ZN(_07819_)
  );
  MUX2_X1 _15422_ (
    .A(\rf[6] [18]),
    .B(\rf[2] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07820_)
  );
  AND2_X1 _15423_ (
    .A1(_03049_),
    .A2(_07820_),
    .ZN(_07821_)
  );
  MUX2_X1 _15424_ (
    .A(\rf[4] [18]),
    .B(\rf[0] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07822_)
  );
  AND2_X1 _15425_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07822_),
    .ZN(_07823_)
  );
  OR2_X1 _15426_ (
    .A1(_03048_),
    .A2(_07823_),
    .ZN(_07824_)
  );
  OR2_X1 _15427_ (
    .A1(_07821_),
    .A2(_07824_),
    .ZN(_07825_)
  );
  MUX2_X1 _15428_ (
    .A(\rf[7] [18]),
    .B(\rf[3] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07826_)
  );
  AND2_X1 _15429_ (
    .A1(_03049_),
    .A2(_07826_),
    .ZN(_07827_)
  );
  MUX2_X1 _15430_ (
    .A(\rf[5] [18]),
    .B(\rf[1] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07828_)
  );
  AND2_X1 _15431_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07828_),
    .ZN(_07829_)
  );
  OR2_X1 _15432_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07829_),
    .ZN(_07830_)
  );
  OR2_X1 _15433_ (
    .A1(_07827_),
    .A2(_07830_),
    .ZN(_07831_)
  );
  AND2_X1 _15434_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_07831_),
    .ZN(_07832_)
  );
  AND2_X1 _15435_ (
    .A1(_07825_),
    .A2(_07832_),
    .ZN(_07833_)
  );
  OR2_X1 _15436_ (
    .A1(_07819_),
    .A2(_07833_),
    .ZN(_07834_)
  );
  OR2_X1 _15437_ (
    .A1(\rf[17] [18]),
    .A2(_03050_),
    .ZN(_07835_)
  );
  OR2_X1 _15438_ (
    .A1(\rf[21] [18]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07836_)
  );
  AND2_X1 _15439_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07836_),
    .ZN(_07837_)
  );
  AND2_X1 _15440_ (
    .A1(_07835_),
    .A2(_07837_),
    .ZN(_07838_)
  );
  MUX2_X1 _15441_ (
    .A(\rf[23] [18]),
    .B(\rf[19] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07839_)
  );
  AND2_X1 _15442_ (
    .A1(_03049_),
    .A2(_07839_),
    .ZN(_07840_)
  );
  OR2_X1 _15443_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07840_),
    .ZN(_07841_)
  );
  OR2_X1 _15444_ (
    .A1(_07838_),
    .A2(_07841_),
    .ZN(_07842_)
  );
  OR2_X1 _15445_ (
    .A1(\rf[20] [18]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07843_)
  );
  OR2_X1 _15446_ (
    .A1(\rf[16] [18]),
    .A2(_03050_),
    .ZN(_07844_)
  );
  AND2_X1 _15447_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07844_),
    .ZN(_07845_)
  );
  AND2_X1 _15448_ (
    .A1(_07843_),
    .A2(_07845_),
    .ZN(_07846_)
  );
  MUX2_X1 _15449_ (
    .A(\rf[22] [18]),
    .B(\rf[18] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07847_)
  );
  AND2_X1 _15450_ (
    .A1(_03049_),
    .A2(_07847_),
    .ZN(_07848_)
  );
  OR2_X1 _15451_ (
    .A1(_03048_),
    .A2(_07848_),
    .ZN(_07849_)
  );
  OR2_X1 _15452_ (
    .A1(_07846_),
    .A2(_07849_),
    .ZN(_07850_)
  );
  AND2_X1 _15453_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_07842_),
    .ZN(_07851_)
  );
  AND2_X1 _15454_ (
    .A1(_07850_),
    .A2(_07851_),
    .ZN(_07852_)
  );
  OR2_X1 _15455_ (
    .A1(\rf[28] [18]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07853_)
  );
  OR2_X1 _15456_ (
    .A1(\rf[24] [18]),
    .A2(_03050_),
    .ZN(_07854_)
  );
  AND2_X1 _15457_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07853_),
    .ZN(_07855_)
  );
  AND2_X1 _15458_ (
    .A1(_07854_),
    .A2(_07855_),
    .ZN(_07856_)
  );
  MUX2_X1 _15459_ (
    .A(\rf[30] [18]),
    .B(\rf[26] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07857_)
  );
  AND2_X1 _15460_ (
    .A1(_03049_),
    .A2(_07857_),
    .ZN(_07858_)
  );
  OR2_X1 _15461_ (
    .A1(_03048_),
    .A2(_07858_),
    .ZN(_07859_)
  );
  OR2_X1 _15462_ (
    .A1(_07856_),
    .A2(_07859_),
    .ZN(_07860_)
  );
  MUX2_X1 _15463_ (
    .A(\rf[29] [18]),
    .B(\rf[25] [18]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07861_)
  );
  AND2_X1 _15464_ (
    .A1(\rf[27] [18]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07862_)
  );
  MUX2_X1 _15465_ (
    .A(_07861_),
    .B(_07862_),
    .S(_03049_),
    .Z(_07863_)
  );
  OR2_X1 _15466_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07863_),
    .ZN(_07864_)
  );
  AND2_X1 _15467_ (
    .A1(_03051_),
    .A2(_07864_),
    .ZN(_07865_)
  );
  AND2_X1 _15468_ (
    .A1(_07860_),
    .A2(_07865_),
    .ZN(_07866_)
  );
  OR2_X1 _15469_ (
    .A1(_07852_),
    .A2(_07866_),
    .ZN(_07867_)
  );
  MUX2_X1 _15470_ (
    .A(_07834_),
    .B(_07867_),
    .S(_03064_),
    .Z(_07868_)
  );
  MUX2_X1 _15471_ (
    .A(_07868_),
    .B(_05302_),
    .S(_06791_),
    .Z(_07869_)
  );
  MUX2_X1 _15472_ (
    .A(ex_reg_rs_msb_1[16]),
    .B(_07869_),
    .S(_06781_),
    .Z(_00165_)
  );
  MUX2_X1 _15473_ (
    .A(\rf[7] [19]),
    .B(\rf[3] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07870_)
  );
  AND2_X1 _15474_ (
    .A1(_03049_),
    .A2(_07870_),
    .ZN(_07871_)
  );
  MUX2_X1 _15475_ (
    .A(\rf[5] [19]),
    .B(\rf[1] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07872_)
  );
  AND2_X1 _15476_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07872_),
    .ZN(_07873_)
  );
  OR2_X1 _15477_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07873_),
    .ZN(_07874_)
  );
  OR2_X1 _15478_ (
    .A1(_07871_),
    .A2(_07874_),
    .ZN(_07875_)
  );
  MUX2_X1 _15479_ (
    .A(\rf[6] [19]),
    .B(\rf[2] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07876_)
  );
  AND2_X1 _15480_ (
    .A1(_03049_),
    .A2(_07876_),
    .ZN(_07877_)
  );
  MUX2_X1 _15481_ (
    .A(\rf[4] [19]),
    .B(\rf[0] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07878_)
  );
  AND2_X1 _15482_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07878_),
    .ZN(_07879_)
  );
  OR2_X1 _15483_ (
    .A1(_03048_),
    .A2(_07879_),
    .ZN(_07880_)
  );
  OR2_X1 _15484_ (
    .A1(_07877_),
    .A2(_07880_),
    .ZN(_07881_)
  );
  AND2_X1 _15485_ (
    .A1(_07875_),
    .A2(_07881_),
    .ZN(_07882_)
  );
  AND2_X1 _15486_ (
    .A1(\rf[14] [19]),
    .A2(_03049_),
    .ZN(_07883_)
  );
  AND2_X1 _15487_ (
    .A1(\rf[12] [19]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_07884_)
  );
  OR2_X1 _15488_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[2]),
    .A2(_07884_),
    .ZN(_07885_)
  );
  OR2_X1 _15489_ (
    .A1(_07883_),
    .A2(_07885_),
    .ZN(_07886_)
  );
  AND2_X1 _15490_ (
    .A1(\rf[10] [19]),
    .A2(_03049_),
    .ZN(_07887_)
  );
  AND2_X1 _15491_ (
    .A1(\rf[8] [19]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_07888_)
  );
  OR2_X1 _15492_ (
    .A1(_03050_),
    .A2(_07888_),
    .ZN(_07889_)
  );
  OR2_X1 _15493_ (
    .A1(_07887_),
    .A2(_07889_),
    .ZN(_07890_)
  );
  AND2_X1 _15494_ (
    .A1(_07886_),
    .A2(_07890_),
    .ZN(_07891_)
  );
  AND2_X1 _15495_ (
    .A1(\rf[15] [19]),
    .A2(_03049_),
    .ZN(_07892_)
  );
  AND2_X1 _15496_ (
    .A1(\rf[13] [19]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_07893_)
  );
  OR2_X1 _15497_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[2]),
    .A2(_07893_),
    .ZN(_07894_)
  );
  OR2_X1 _15498_ (
    .A1(_07892_),
    .A2(_07894_),
    .ZN(_07895_)
  );
  AND2_X1 _15499_ (
    .A1(\rf[11] [19]),
    .A2(_03049_),
    .ZN(_07896_)
  );
  AND2_X1 _15500_ (
    .A1(\rf[9] [19]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[1]),
    .ZN(_07897_)
  );
  OR2_X1 _15501_ (
    .A1(_03050_),
    .A2(_07897_),
    .ZN(_07898_)
  );
  OR2_X1 _15502_ (
    .A1(_07896_),
    .A2(_07898_),
    .ZN(_07899_)
  );
  AND2_X1 _15503_ (
    .A1(_07895_),
    .A2(_07899_),
    .ZN(_07900_)
  );
  MUX2_X1 _15504_ (
    .A(_07891_),
    .B(_07900_),
    .S(_03048_),
    .Z(_07901_)
  );
  MUX2_X1 _15505_ (
    .A(_07882_),
    .B(_07901_),
    .S(_03051_),
    .Z(_07902_)
  );
  OR2_X1 _15506_ (
    .A1(\rf[28] [19]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07903_)
  );
  OR2_X1 _15507_ (
    .A1(\rf[24] [19]),
    .A2(_03050_),
    .ZN(_07904_)
  );
  AND2_X1 _15508_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07903_),
    .ZN(_07905_)
  );
  AND2_X1 _15509_ (
    .A1(_07904_),
    .A2(_07905_),
    .ZN(_07906_)
  );
  MUX2_X1 _15510_ (
    .A(\rf[30] [19]),
    .B(\rf[26] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07907_)
  );
  AND2_X1 _15511_ (
    .A1(_03049_),
    .A2(_07907_),
    .ZN(_07908_)
  );
  OR2_X1 _15512_ (
    .A1(_03048_),
    .A2(_07908_),
    .ZN(_07909_)
  );
  OR2_X1 _15513_ (
    .A1(_07906_),
    .A2(_07909_),
    .ZN(_07910_)
  );
  MUX2_X1 _15514_ (
    .A(\rf[29] [19]),
    .B(\rf[25] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07911_)
  );
  AND2_X1 _15515_ (
    .A1(\rf[27] [19]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07912_)
  );
  MUX2_X1 _15516_ (
    .A(_07911_),
    .B(_07912_),
    .S(_03049_),
    .Z(_07913_)
  );
  OR2_X1 _15517_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07913_),
    .ZN(_07914_)
  );
  AND2_X1 _15518_ (
    .A1(_07910_),
    .A2(_07914_),
    .ZN(_07915_)
  );
  OR2_X1 _15519_ (
    .A1(\rf[20] [19]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07916_)
  );
  OR2_X1 _15520_ (
    .A1(\rf[16] [19]),
    .A2(_03050_),
    .ZN(_07917_)
  );
  AND2_X1 _15521_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07917_),
    .ZN(_07918_)
  );
  AND2_X1 _15522_ (
    .A1(_07916_),
    .A2(_07918_),
    .ZN(_07919_)
  );
  MUX2_X1 _15523_ (
    .A(\rf[22] [19]),
    .B(\rf[18] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07920_)
  );
  AND2_X1 _15524_ (
    .A1(_03049_),
    .A2(_07920_),
    .ZN(_07921_)
  );
  OR2_X1 _15525_ (
    .A1(_03048_),
    .A2(_07921_),
    .ZN(_07922_)
  );
  OR2_X1 _15526_ (
    .A1(_07919_),
    .A2(_07922_),
    .ZN(_07923_)
  );
  OR2_X1 _15527_ (
    .A1(\rf[17] [19]),
    .A2(_03050_),
    .ZN(_07924_)
  );
  OR2_X1 _15528_ (
    .A1(\rf[21] [19]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07925_)
  );
  AND2_X1 _15529_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07925_),
    .ZN(_07926_)
  );
  AND2_X1 _15530_ (
    .A1(_07924_),
    .A2(_07926_),
    .ZN(_07927_)
  );
  MUX2_X1 _15531_ (
    .A(\rf[23] [19]),
    .B(\rf[19] [19]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07928_)
  );
  AND2_X1 _15532_ (
    .A1(_03049_),
    .A2(_07928_),
    .ZN(_07929_)
  );
  OR2_X1 _15533_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07929_),
    .ZN(_07930_)
  );
  OR2_X1 _15534_ (
    .A1(_07927_),
    .A2(_07930_),
    .ZN(_07931_)
  );
  AND2_X1 _15535_ (
    .A1(_07923_),
    .A2(_07931_),
    .ZN(_07932_)
  );
  MUX2_X1 _15536_ (
    .A(_07915_),
    .B(_07932_),
    .S(ibuf_io_inst_0_bits_inst_rs2[3]),
    .Z(_07933_)
  );
  MUX2_X1 _15537_ (
    .A(_07902_),
    .B(_07933_),
    .S(_03064_),
    .Z(_07934_)
  );
  MUX2_X1 _15538_ (
    .A(_07934_),
    .B(_05310_),
    .S(_06791_),
    .Z(_07935_)
  );
  MUX2_X1 _15539_ (
    .A(ex_reg_rs_msb_1[17]),
    .B(_07935_),
    .S(_06781_),
    .Z(_00166_)
  );
  OR2_X1 _15540_ (
    .A1(\rf[10] [20]),
    .A2(_03050_),
    .ZN(_07936_)
  );
  OR2_X1 _15541_ (
    .A1(\rf[14] [20]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07937_)
  );
  AND2_X1 _15542_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07937_),
    .ZN(_07938_)
  );
  AND2_X1 _15543_ (
    .A1(_07936_),
    .A2(_07938_),
    .ZN(_07939_)
  );
  MUX2_X1 _15544_ (
    .A(\rf[15] [20]),
    .B(\rf[11] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07940_)
  );
  AND2_X1 _15545_ (
    .A1(_03048_),
    .A2(_07940_),
    .ZN(_07941_)
  );
  OR2_X1 _15546_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07941_),
    .ZN(_07942_)
  );
  OR2_X1 _15547_ (
    .A1(_07939_),
    .A2(_07942_),
    .ZN(_07943_)
  );
  OR2_X1 _15548_ (
    .A1(\rf[12] [20]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07944_)
  );
  OR2_X1 _15549_ (
    .A1(\rf[8] [20]),
    .A2(_03050_),
    .ZN(_07945_)
  );
  AND2_X1 _15550_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07944_),
    .ZN(_07946_)
  );
  AND2_X1 _15551_ (
    .A1(_07945_),
    .A2(_07946_),
    .ZN(_07947_)
  );
  MUX2_X1 _15552_ (
    .A(\rf[13] [20]),
    .B(\rf[9] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07948_)
  );
  AND2_X1 _15553_ (
    .A1(_03048_),
    .A2(_07948_),
    .ZN(_07949_)
  );
  OR2_X1 _15554_ (
    .A1(_03049_),
    .A2(_07949_),
    .ZN(_07950_)
  );
  OR2_X1 _15555_ (
    .A1(_07947_),
    .A2(_07950_),
    .ZN(_07951_)
  );
  AND2_X1 _15556_ (
    .A1(_03051_),
    .A2(_07951_),
    .ZN(_07952_)
  );
  AND2_X1 _15557_ (
    .A1(_07943_),
    .A2(_07952_),
    .ZN(_07953_)
  );
  MUX2_X1 _15558_ (
    .A(\rf[6] [20]),
    .B(\rf[2] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07954_)
  );
  AND2_X1 _15559_ (
    .A1(_03049_),
    .A2(_07954_),
    .ZN(_07955_)
  );
  MUX2_X1 _15560_ (
    .A(\rf[4] [20]),
    .B(\rf[0] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07956_)
  );
  AND2_X1 _15561_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07956_),
    .ZN(_07957_)
  );
  OR2_X1 _15562_ (
    .A1(_03048_),
    .A2(_07957_),
    .ZN(_07958_)
  );
  OR2_X1 _15563_ (
    .A1(_07955_),
    .A2(_07958_),
    .ZN(_07959_)
  );
  MUX2_X1 _15564_ (
    .A(\rf[7] [20]),
    .B(\rf[3] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07960_)
  );
  AND2_X1 _15565_ (
    .A1(_03049_),
    .A2(_07960_),
    .ZN(_07961_)
  );
  MUX2_X1 _15566_ (
    .A(\rf[5] [20]),
    .B(\rf[1] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07962_)
  );
  AND2_X1 _15567_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07962_),
    .ZN(_07963_)
  );
  OR2_X1 _15568_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07963_),
    .ZN(_07964_)
  );
  OR2_X1 _15569_ (
    .A1(_07961_),
    .A2(_07964_),
    .ZN(_07965_)
  );
  AND2_X1 _15570_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_07965_),
    .ZN(_07966_)
  );
  AND2_X1 _15571_ (
    .A1(_07959_),
    .A2(_07966_),
    .ZN(_07967_)
  );
  OR2_X1 _15572_ (
    .A1(_07953_),
    .A2(_07967_),
    .ZN(_07968_)
  );
  OR2_X1 _15573_ (
    .A1(\rf[17] [20]),
    .A2(_03050_),
    .ZN(_07969_)
  );
  OR2_X1 _15574_ (
    .A1(\rf[21] [20]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07970_)
  );
  AND2_X1 _15575_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07970_),
    .ZN(_07971_)
  );
  AND2_X1 _15576_ (
    .A1(_07969_),
    .A2(_07971_),
    .ZN(_07972_)
  );
  MUX2_X1 _15577_ (
    .A(\rf[23] [20]),
    .B(\rf[19] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07973_)
  );
  AND2_X1 _15578_ (
    .A1(_03049_),
    .A2(_07973_),
    .ZN(_07974_)
  );
  OR2_X1 _15579_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07974_),
    .ZN(_07975_)
  );
  OR2_X1 _15580_ (
    .A1(_07972_),
    .A2(_07975_),
    .ZN(_07976_)
  );
  OR2_X1 _15581_ (
    .A1(\rf[20] [20]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07977_)
  );
  OR2_X1 _15582_ (
    .A1(\rf[16] [20]),
    .A2(_03050_),
    .ZN(_07978_)
  );
  AND2_X1 _15583_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07978_),
    .ZN(_07979_)
  );
  AND2_X1 _15584_ (
    .A1(_07977_),
    .A2(_07979_),
    .ZN(_07980_)
  );
  MUX2_X1 _15585_ (
    .A(\rf[22] [20]),
    .B(\rf[18] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07981_)
  );
  AND2_X1 _15586_ (
    .A1(_03049_),
    .A2(_07981_),
    .ZN(_07982_)
  );
  OR2_X1 _15587_ (
    .A1(_03048_),
    .A2(_07982_),
    .ZN(_07983_)
  );
  OR2_X1 _15588_ (
    .A1(_07980_),
    .A2(_07983_),
    .ZN(_07984_)
  );
  AND2_X1 _15589_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_07976_),
    .ZN(_07985_)
  );
  AND2_X1 _15590_ (
    .A1(_07984_),
    .A2(_07985_),
    .ZN(_07986_)
  );
  OR2_X1 _15591_ (
    .A1(\rf[28] [20]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07987_)
  );
  OR2_X1 _15592_ (
    .A1(\rf[24] [20]),
    .A2(_03050_),
    .ZN(_07988_)
  );
  AND2_X1 _15593_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_07987_),
    .ZN(_07989_)
  );
  AND2_X1 _15594_ (
    .A1(_07988_),
    .A2(_07989_),
    .ZN(_07990_)
  );
  MUX2_X1 _15595_ (
    .A(\rf[30] [20]),
    .B(\rf[26] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07991_)
  );
  AND2_X1 _15596_ (
    .A1(_03049_),
    .A2(_07991_),
    .ZN(_07992_)
  );
  OR2_X1 _15597_ (
    .A1(_03048_),
    .A2(_07992_),
    .ZN(_07993_)
  );
  OR2_X1 _15598_ (
    .A1(_07990_),
    .A2(_07993_),
    .ZN(_07994_)
  );
  MUX2_X1 _15599_ (
    .A(\rf[29] [20]),
    .B(\rf[25] [20]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_07995_)
  );
  AND2_X1 _15600_ (
    .A1(\rf[27] [20]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_07996_)
  );
  MUX2_X1 _15601_ (
    .A(_07995_),
    .B(_07996_),
    .S(_03049_),
    .Z(_07997_)
  );
  OR2_X1 _15602_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_07997_),
    .ZN(_07998_)
  );
  AND2_X1 _15603_ (
    .A1(_03051_),
    .A2(_07998_),
    .ZN(_07999_)
  );
  AND2_X1 _15604_ (
    .A1(_07994_),
    .A2(_07999_),
    .ZN(_08000_)
  );
  OR2_X1 _15605_ (
    .A1(_07986_),
    .A2(_08000_),
    .ZN(_08001_)
  );
  MUX2_X1 _15606_ (
    .A(_07968_),
    .B(_08001_),
    .S(_03064_),
    .Z(_08002_)
  );
  MUX2_X1 _15607_ (
    .A(_08002_),
    .B(_05442_),
    .S(_06791_),
    .Z(_08003_)
  );
  MUX2_X1 _15608_ (
    .A(ex_reg_rs_msb_1[18]),
    .B(_08003_),
    .S(_06781_),
    .Z(_00167_)
  );
  OR2_X1 _15609_ (
    .A1(\rf[10] [21]),
    .A2(_03050_),
    .ZN(_08004_)
  );
  OR2_X1 _15610_ (
    .A1(\rf[14] [21]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08005_)
  );
  AND2_X1 _15611_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08005_),
    .ZN(_08006_)
  );
  AND2_X1 _15612_ (
    .A1(_08004_),
    .A2(_08006_),
    .ZN(_08007_)
  );
  MUX2_X1 _15613_ (
    .A(\rf[15] [21]),
    .B(\rf[11] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08008_)
  );
  AND2_X1 _15614_ (
    .A1(_03048_),
    .A2(_08008_),
    .ZN(_08009_)
  );
  OR2_X1 _15615_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08009_),
    .ZN(_08010_)
  );
  OR2_X1 _15616_ (
    .A1(_08007_),
    .A2(_08010_),
    .ZN(_08011_)
  );
  OR2_X1 _15617_ (
    .A1(\rf[12] [21]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08012_)
  );
  OR2_X1 _15618_ (
    .A1(\rf[8] [21]),
    .A2(_03050_),
    .ZN(_08013_)
  );
  AND2_X1 _15619_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08012_),
    .ZN(_08014_)
  );
  AND2_X1 _15620_ (
    .A1(_08013_),
    .A2(_08014_),
    .ZN(_08015_)
  );
  MUX2_X1 _15621_ (
    .A(\rf[13] [21]),
    .B(\rf[9] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08016_)
  );
  AND2_X1 _15622_ (
    .A1(_03048_),
    .A2(_08016_),
    .ZN(_08017_)
  );
  OR2_X1 _15623_ (
    .A1(_03049_),
    .A2(_08017_),
    .ZN(_08018_)
  );
  OR2_X1 _15624_ (
    .A1(_08015_),
    .A2(_08018_),
    .ZN(_08019_)
  );
  AND2_X1 _15625_ (
    .A1(_03051_),
    .A2(_08019_),
    .ZN(_08020_)
  );
  AND2_X1 _15626_ (
    .A1(_08011_),
    .A2(_08020_),
    .ZN(_08021_)
  );
  MUX2_X1 _15627_ (
    .A(\rf[6] [21]),
    .B(\rf[2] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08022_)
  );
  AND2_X1 _15628_ (
    .A1(_03049_),
    .A2(_08022_),
    .ZN(_08023_)
  );
  MUX2_X1 _15629_ (
    .A(\rf[4] [21]),
    .B(\rf[0] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08024_)
  );
  AND2_X1 _15630_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08024_),
    .ZN(_08025_)
  );
  OR2_X1 _15631_ (
    .A1(_03048_),
    .A2(_08025_),
    .ZN(_08026_)
  );
  OR2_X1 _15632_ (
    .A1(_08023_),
    .A2(_08026_),
    .ZN(_08027_)
  );
  MUX2_X1 _15633_ (
    .A(\rf[7] [21]),
    .B(\rf[3] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08028_)
  );
  AND2_X1 _15634_ (
    .A1(_03049_),
    .A2(_08028_),
    .ZN(_08029_)
  );
  MUX2_X1 _15635_ (
    .A(\rf[5] [21]),
    .B(\rf[1] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08030_)
  );
  AND2_X1 _15636_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08030_),
    .ZN(_08031_)
  );
  OR2_X1 _15637_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08031_),
    .ZN(_08032_)
  );
  OR2_X1 _15638_ (
    .A1(_08029_),
    .A2(_08032_),
    .ZN(_08033_)
  );
  AND2_X1 _15639_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_08033_),
    .ZN(_08034_)
  );
  AND2_X1 _15640_ (
    .A1(_08027_),
    .A2(_08034_),
    .ZN(_08035_)
  );
  OR2_X1 _15641_ (
    .A1(_08021_),
    .A2(_08035_),
    .ZN(_08036_)
  );
  OR2_X1 _15642_ (
    .A1(\rf[17] [21]),
    .A2(_03050_),
    .ZN(_08037_)
  );
  OR2_X1 _15643_ (
    .A1(\rf[21] [21]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08038_)
  );
  AND2_X1 _15644_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08038_),
    .ZN(_08039_)
  );
  AND2_X1 _15645_ (
    .A1(_08037_),
    .A2(_08039_),
    .ZN(_08040_)
  );
  MUX2_X1 _15646_ (
    .A(\rf[23] [21]),
    .B(\rf[19] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08041_)
  );
  AND2_X1 _15647_ (
    .A1(_03049_),
    .A2(_08041_),
    .ZN(_08042_)
  );
  OR2_X1 _15648_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08042_),
    .ZN(_08043_)
  );
  OR2_X1 _15649_ (
    .A1(_08040_),
    .A2(_08043_),
    .ZN(_08044_)
  );
  OR2_X1 _15650_ (
    .A1(\rf[20] [21]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08045_)
  );
  OR2_X1 _15651_ (
    .A1(\rf[16] [21]),
    .A2(_03050_),
    .ZN(_08046_)
  );
  AND2_X1 _15652_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08046_),
    .ZN(_08047_)
  );
  AND2_X1 _15653_ (
    .A1(_08045_),
    .A2(_08047_),
    .ZN(_08048_)
  );
  MUX2_X1 _15654_ (
    .A(\rf[22] [21]),
    .B(\rf[18] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08049_)
  );
  AND2_X1 _15655_ (
    .A1(_03049_),
    .A2(_08049_),
    .ZN(_08050_)
  );
  OR2_X1 _15656_ (
    .A1(_03048_),
    .A2(_08050_),
    .ZN(_08051_)
  );
  OR2_X1 _15657_ (
    .A1(_08048_),
    .A2(_08051_),
    .ZN(_08052_)
  );
  AND2_X1 _15658_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_08044_),
    .ZN(_08053_)
  );
  AND2_X1 _15659_ (
    .A1(_08052_),
    .A2(_08053_),
    .ZN(_08054_)
  );
  OR2_X1 _15660_ (
    .A1(\rf[28] [21]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08055_)
  );
  OR2_X1 _15661_ (
    .A1(\rf[24] [21]),
    .A2(_03050_),
    .ZN(_08056_)
  );
  AND2_X1 _15662_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08055_),
    .ZN(_08057_)
  );
  AND2_X1 _15663_ (
    .A1(_08056_),
    .A2(_08057_),
    .ZN(_08058_)
  );
  MUX2_X1 _15664_ (
    .A(\rf[30] [21]),
    .B(\rf[26] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08059_)
  );
  AND2_X1 _15665_ (
    .A1(_03049_),
    .A2(_08059_),
    .ZN(_08060_)
  );
  OR2_X1 _15666_ (
    .A1(_03048_),
    .A2(_08060_),
    .ZN(_08061_)
  );
  OR2_X1 _15667_ (
    .A1(_08058_),
    .A2(_08061_),
    .ZN(_08062_)
  );
  MUX2_X1 _15668_ (
    .A(\rf[29] [21]),
    .B(\rf[25] [21]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08063_)
  );
  AND2_X1 _15669_ (
    .A1(\rf[27] [21]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08064_)
  );
  MUX2_X1 _15670_ (
    .A(_08063_),
    .B(_08064_),
    .S(_03049_),
    .Z(_08065_)
  );
  OR2_X1 _15671_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08065_),
    .ZN(_08066_)
  );
  AND2_X1 _15672_ (
    .A1(_03051_),
    .A2(_08066_),
    .ZN(_08067_)
  );
  AND2_X1 _15673_ (
    .A1(_08062_),
    .A2(_08067_),
    .ZN(_08068_)
  );
  OR2_X1 _15674_ (
    .A1(_08054_),
    .A2(_08068_),
    .ZN(_08069_)
  );
  MUX2_X1 _15675_ (
    .A(_08036_),
    .B(_08069_),
    .S(_03064_),
    .Z(_08070_)
  );
  MUX2_X1 _15676_ (
    .A(_08070_),
    .B(_05450_),
    .S(_06791_),
    .Z(_08071_)
  );
  MUX2_X1 _15677_ (
    .A(ex_reg_rs_msb_1[19]),
    .B(_08071_),
    .S(_06781_),
    .Z(_00168_)
  );
  OR2_X1 _15678_ (
    .A1(\rf[10] [22]),
    .A2(_03050_),
    .ZN(_08072_)
  );
  OR2_X1 _15679_ (
    .A1(\rf[14] [22]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08073_)
  );
  AND2_X1 _15680_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08073_),
    .ZN(_08074_)
  );
  AND2_X1 _15681_ (
    .A1(_08072_),
    .A2(_08074_),
    .ZN(_08075_)
  );
  MUX2_X1 _15682_ (
    .A(\rf[15] [22]),
    .B(\rf[11] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08076_)
  );
  AND2_X1 _15683_ (
    .A1(_03048_),
    .A2(_08076_),
    .ZN(_08077_)
  );
  OR2_X1 _15684_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08077_),
    .ZN(_08078_)
  );
  OR2_X1 _15685_ (
    .A1(_08075_),
    .A2(_08078_),
    .ZN(_08079_)
  );
  OR2_X1 _15686_ (
    .A1(\rf[12] [22]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08080_)
  );
  OR2_X1 _15687_ (
    .A1(\rf[8] [22]),
    .A2(_03050_),
    .ZN(_08081_)
  );
  AND2_X1 _15688_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08080_),
    .ZN(_08082_)
  );
  AND2_X1 _15689_ (
    .A1(_08081_),
    .A2(_08082_),
    .ZN(_08083_)
  );
  MUX2_X1 _15690_ (
    .A(\rf[13] [22]),
    .B(\rf[9] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08084_)
  );
  AND2_X1 _15691_ (
    .A1(_03048_),
    .A2(_08084_),
    .ZN(_08085_)
  );
  OR2_X1 _15692_ (
    .A1(_03049_),
    .A2(_08085_),
    .ZN(_08086_)
  );
  OR2_X1 _15693_ (
    .A1(_08083_),
    .A2(_08086_),
    .ZN(_08087_)
  );
  AND2_X1 _15694_ (
    .A1(_03051_),
    .A2(_08087_),
    .ZN(_08088_)
  );
  AND2_X1 _15695_ (
    .A1(_08079_),
    .A2(_08088_),
    .ZN(_08089_)
  );
  MUX2_X1 _15696_ (
    .A(\rf[6] [22]),
    .B(\rf[2] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08090_)
  );
  AND2_X1 _15697_ (
    .A1(_03049_),
    .A2(_08090_),
    .ZN(_08091_)
  );
  MUX2_X1 _15698_ (
    .A(\rf[4] [22]),
    .B(\rf[0] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08092_)
  );
  AND2_X1 _15699_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08092_),
    .ZN(_08093_)
  );
  OR2_X1 _15700_ (
    .A1(_03048_),
    .A2(_08093_),
    .ZN(_08094_)
  );
  OR2_X1 _15701_ (
    .A1(_08091_),
    .A2(_08094_),
    .ZN(_08095_)
  );
  MUX2_X1 _15702_ (
    .A(\rf[7] [22]),
    .B(\rf[3] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08096_)
  );
  AND2_X1 _15703_ (
    .A1(_03049_),
    .A2(_08096_),
    .ZN(_08097_)
  );
  MUX2_X1 _15704_ (
    .A(\rf[5] [22]),
    .B(\rf[1] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08098_)
  );
  AND2_X1 _15705_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08098_),
    .ZN(_08099_)
  );
  OR2_X1 _15706_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08099_),
    .ZN(_08100_)
  );
  OR2_X1 _15707_ (
    .A1(_08097_),
    .A2(_08100_),
    .ZN(_08101_)
  );
  AND2_X1 _15708_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_08101_),
    .ZN(_08102_)
  );
  AND2_X1 _15709_ (
    .A1(_08095_),
    .A2(_08102_),
    .ZN(_08103_)
  );
  OR2_X1 _15710_ (
    .A1(_08089_),
    .A2(_08103_),
    .ZN(_08104_)
  );
  OR2_X1 _15711_ (
    .A1(\rf[17] [22]),
    .A2(_03050_),
    .ZN(_08105_)
  );
  OR2_X1 _15712_ (
    .A1(\rf[21] [22]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08106_)
  );
  AND2_X1 _15713_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08106_),
    .ZN(_08107_)
  );
  AND2_X1 _15714_ (
    .A1(_08105_),
    .A2(_08107_),
    .ZN(_08108_)
  );
  MUX2_X1 _15715_ (
    .A(\rf[23] [22]),
    .B(\rf[19] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08109_)
  );
  AND2_X1 _15716_ (
    .A1(_03049_),
    .A2(_08109_),
    .ZN(_08110_)
  );
  OR2_X1 _15717_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08110_),
    .ZN(_08111_)
  );
  OR2_X1 _15718_ (
    .A1(_08108_),
    .A2(_08111_),
    .ZN(_08112_)
  );
  OR2_X1 _15719_ (
    .A1(\rf[20] [22]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08113_)
  );
  OR2_X1 _15720_ (
    .A1(\rf[16] [22]),
    .A2(_03050_),
    .ZN(_08114_)
  );
  AND2_X1 _15721_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08114_),
    .ZN(_08115_)
  );
  AND2_X1 _15722_ (
    .A1(_08113_),
    .A2(_08115_),
    .ZN(_08116_)
  );
  MUX2_X1 _15723_ (
    .A(\rf[22] [22]),
    .B(\rf[18] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08117_)
  );
  AND2_X1 _15724_ (
    .A1(_03049_),
    .A2(_08117_),
    .ZN(_08118_)
  );
  OR2_X1 _15725_ (
    .A1(_03048_),
    .A2(_08118_),
    .ZN(_08119_)
  );
  OR2_X1 _15726_ (
    .A1(_08116_),
    .A2(_08119_),
    .ZN(_08120_)
  );
  AND2_X1 _15727_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_08112_),
    .ZN(_08121_)
  );
  AND2_X1 _15728_ (
    .A1(_08120_),
    .A2(_08121_),
    .ZN(_08122_)
  );
  OR2_X1 _15729_ (
    .A1(\rf[28] [22]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08123_)
  );
  OR2_X1 _15730_ (
    .A1(\rf[24] [22]),
    .A2(_03050_),
    .ZN(_08124_)
  );
  AND2_X1 _15731_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08123_),
    .ZN(_08125_)
  );
  AND2_X1 _15732_ (
    .A1(_08124_),
    .A2(_08125_),
    .ZN(_08126_)
  );
  MUX2_X1 _15733_ (
    .A(\rf[30] [22]),
    .B(\rf[26] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08127_)
  );
  AND2_X1 _15734_ (
    .A1(_03049_),
    .A2(_08127_),
    .ZN(_08128_)
  );
  OR2_X1 _15735_ (
    .A1(_03048_),
    .A2(_08128_),
    .ZN(_08129_)
  );
  OR2_X1 _15736_ (
    .A1(_08126_),
    .A2(_08129_),
    .ZN(_08130_)
  );
  MUX2_X1 _15737_ (
    .A(\rf[29] [22]),
    .B(\rf[25] [22]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08131_)
  );
  AND2_X1 _15738_ (
    .A1(\rf[27] [22]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08132_)
  );
  MUX2_X1 _15739_ (
    .A(_08131_),
    .B(_08132_),
    .S(_03049_),
    .Z(_08133_)
  );
  OR2_X1 _15740_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08133_),
    .ZN(_08134_)
  );
  AND2_X1 _15741_ (
    .A1(_03051_),
    .A2(_08134_),
    .ZN(_08135_)
  );
  AND2_X1 _15742_ (
    .A1(_08130_),
    .A2(_08135_),
    .ZN(_08136_)
  );
  OR2_X1 _15743_ (
    .A1(_08122_),
    .A2(_08136_),
    .ZN(_08137_)
  );
  MUX2_X1 _15744_ (
    .A(_08104_),
    .B(_08137_),
    .S(_03064_),
    .Z(_08138_)
  );
  MUX2_X1 _15745_ (
    .A(_08138_),
    .B(_05592_),
    .S(_06791_),
    .Z(_08139_)
  );
  MUX2_X1 _15746_ (
    .A(ex_reg_rs_msb_1[20]),
    .B(_08139_),
    .S(_06781_),
    .Z(_00169_)
  );
  MUX2_X1 _15747_ (
    .A(\rf[3] [23]),
    .B(\rf[2] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_08140_)
  );
  MUX2_X1 _15748_ (
    .A(\rf[7] [23]),
    .B(\rf[6] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_08141_)
  );
  MUX2_X1 _15749_ (
    .A(_08140_),
    .B(_08141_),
    .S(_03050_),
    .Z(_08142_)
  );
  OR2_X1 _15750_ (
    .A1(_03051_),
    .A2(_08142_),
    .ZN(_08143_)
  );
  MUX2_X1 _15751_ (
    .A(\rf[14] [23]),
    .B(\rf[10] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08144_)
  );
  OR2_X1 _15752_ (
    .A1(_06863_),
    .A2(_08144_),
    .ZN(_08145_)
  );
  MUX2_X1 _15753_ (
    .A(\rf[15] [23]),
    .B(\rf[11] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08146_)
  );
  OR2_X1 _15754_ (
    .A1(_03808_),
    .A2(_08146_),
    .ZN(_08147_)
  );
  AND2_X1 _15755_ (
    .A1(_08145_),
    .A2(_08147_),
    .ZN(_08148_)
  );
  AND2_X1 _15756_ (
    .A1(_08143_),
    .A2(_08148_),
    .ZN(_08149_)
  );
  MUX2_X1 _15757_ (
    .A(\rf[1] [23]),
    .B(\rf[0] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_08150_)
  );
  MUX2_X1 _15758_ (
    .A(\rf[5] [23]),
    .B(\rf[4] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_08151_)
  );
  MUX2_X1 _15759_ (
    .A(_08150_),
    .B(_08151_),
    .S(_03050_),
    .Z(_08152_)
  );
  OR2_X1 _15760_ (
    .A1(_03051_),
    .A2(_08152_),
    .ZN(_08153_)
  );
  MUX2_X1 _15761_ (
    .A(\rf[12] [23]),
    .B(\rf[8] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08154_)
  );
  OR2_X1 _15762_ (
    .A1(_06863_),
    .A2(_08154_),
    .ZN(_08155_)
  );
  MUX2_X1 _15763_ (
    .A(\rf[13] [23]),
    .B(\rf[9] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08156_)
  );
  OR2_X1 _15764_ (
    .A1(_03808_),
    .A2(_08156_),
    .ZN(_08157_)
  );
  AND2_X1 _15765_ (
    .A1(_08155_),
    .A2(_08157_),
    .ZN(_08158_)
  );
  AND2_X1 _15766_ (
    .A1(_08153_),
    .A2(_08158_),
    .ZN(_08159_)
  );
  OR2_X1 _15767_ (
    .A1(\rf[28] [23]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08160_)
  );
  OR2_X1 _15768_ (
    .A1(\rf[24] [23]),
    .A2(_03050_),
    .ZN(_08161_)
  );
  AND2_X1 _15769_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08160_),
    .ZN(_08162_)
  );
  AND2_X1 _15770_ (
    .A1(_08161_),
    .A2(_08162_),
    .ZN(_08163_)
  );
  MUX2_X1 _15771_ (
    .A(\rf[30] [23]),
    .B(\rf[26] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08164_)
  );
  AND2_X1 _15772_ (
    .A1(_03049_),
    .A2(_08164_),
    .ZN(_08165_)
  );
  OR2_X1 _15773_ (
    .A1(_03048_),
    .A2(_08165_),
    .ZN(_08166_)
  );
  OR2_X1 _15774_ (
    .A1(_08163_),
    .A2(_08166_),
    .ZN(_08167_)
  );
  MUX2_X1 _15775_ (
    .A(\rf[29] [23]),
    .B(\rf[25] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08168_)
  );
  AND2_X1 _15776_ (
    .A1(\rf[27] [23]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08169_)
  );
  MUX2_X1 _15777_ (
    .A(_08168_),
    .B(_08169_),
    .S(_03049_),
    .Z(_08170_)
  );
  OR2_X1 _15778_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08170_),
    .ZN(_08171_)
  );
  AND2_X1 _15779_ (
    .A1(_08167_),
    .A2(_08171_),
    .ZN(_08172_)
  );
  OR2_X1 _15780_ (
    .A1(\rf[20] [23]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08173_)
  );
  OR2_X1 _15781_ (
    .A1(\rf[16] [23]),
    .A2(_03050_),
    .ZN(_08174_)
  );
  AND2_X1 _15782_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08174_),
    .ZN(_08175_)
  );
  AND2_X1 _15783_ (
    .A1(_08173_),
    .A2(_08175_),
    .ZN(_08176_)
  );
  MUX2_X1 _15784_ (
    .A(\rf[22] [23]),
    .B(\rf[18] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08177_)
  );
  AND2_X1 _15785_ (
    .A1(_03049_),
    .A2(_08177_),
    .ZN(_08178_)
  );
  OR2_X1 _15786_ (
    .A1(_03048_),
    .A2(_08178_),
    .ZN(_08179_)
  );
  OR2_X1 _15787_ (
    .A1(_08176_),
    .A2(_08179_),
    .ZN(_08180_)
  );
  OR2_X1 _15788_ (
    .A1(\rf[17] [23]),
    .A2(_03050_),
    .ZN(_08181_)
  );
  OR2_X1 _15789_ (
    .A1(\rf[21] [23]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08182_)
  );
  AND2_X1 _15790_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08182_),
    .ZN(_08183_)
  );
  AND2_X1 _15791_ (
    .A1(_08181_),
    .A2(_08183_),
    .ZN(_08184_)
  );
  MUX2_X1 _15792_ (
    .A(\rf[23] [23]),
    .B(\rf[19] [23]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08185_)
  );
  AND2_X1 _15793_ (
    .A1(_03049_),
    .A2(_08185_),
    .ZN(_08186_)
  );
  OR2_X1 _15794_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08186_),
    .ZN(_08187_)
  );
  OR2_X1 _15795_ (
    .A1(_08184_),
    .A2(_08187_),
    .ZN(_08188_)
  );
  AND2_X1 _15796_ (
    .A1(_08180_),
    .A2(_08188_),
    .ZN(_08189_)
  );
  MUX2_X1 _15797_ (
    .A(_08172_),
    .B(_08189_),
    .S(ibuf_io_inst_0_bits_inst_rs2[3]),
    .Z(_08190_)
  );
  MUX2_X1 _15798_ (
    .A(_08149_),
    .B(_08159_),
    .S(ibuf_io_inst_0_bits_inst_rs2[1]),
    .Z(_08191_)
  );
  MUX2_X1 _15799_ (
    .A(_08190_),
    .B(_08191_),
    .S(ibuf_io_inst_0_bits_inst_rs2[4]),
    .Z(_08192_)
  );
  MUX2_X1 _15800_ (
    .A(_08192_),
    .B(_05657_),
    .S(_06791_),
    .Z(_08193_)
  );
  MUX2_X1 _15801_ (
    .A(ex_reg_rs_msb_1[21]),
    .B(_08193_),
    .S(_06781_),
    .Z(_00170_)
  );
  OR2_X1 _15802_ (
    .A1(\rf[10] [24]),
    .A2(_03050_),
    .ZN(_08194_)
  );
  OR2_X1 _15803_ (
    .A1(\rf[14] [24]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08195_)
  );
  AND2_X1 _15804_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08195_),
    .ZN(_08196_)
  );
  AND2_X1 _15805_ (
    .A1(_08194_),
    .A2(_08196_),
    .ZN(_08197_)
  );
  MUX2_X1 _15806_ (
    .A(\rf[15] [24]),
    .B(\rf[11] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08198_)
  );
  AND2_X1 _15807_ (
    .A1(_03048_),
    .A2(_08198_),
    .ZN(_08199_)
  );
  OR2_X1 _15808_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08199_),
    .ZN(_08200_)
  );
  OR2_X1 _15809_ (
    .A1(_08197_),
    .A2(_08200_),
    .ZN(_08201_)
  );
  OR2_X1 _15810_ (
    .A1(\rf[12] [24]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08202_)
  );
  OR2_X1 _15811_ (
    .A1(\rf[8] [24]),
    .A2(_03050_),
    .ZN(_08203_)
  );
  AND2_X1 _15812_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08202_),
    .ZN(_08204_)
  );
  AND2_X1 _15813_ (
    .A1(_08203_),
    .A2(_08204_),
    .ZN(_08205_)
  );
  MUX2_X1 _15814_ (
    .A(\rf[13] [24]),
    .B(\rf[9] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08206_)
  );
  AND2_X1 _15815_ (
    .A1(_03048_),
    .A2(_08206_),
    .ZN(_08207_)
  );
  OR2_X1 _15816_ (
    .A1(_03049_),
    .A2(_08207_),
    .ZN(_08208_)
  );
  OR2_X1 _15817_ (
    .A1(_08205_),
    .A2(_08208_),
    .ZN(_08209_)
  );
  AND2_X1 _15818_ (
    .A1(_03051_),
    .A2(_08209_),
    .ZN(_08210_)
  );
  AND2_X1 _15819_ (
    .A1(_08201_),
    .A2(_08210_),
    .ZN(_08211_)
  );
  MUX2_X1 _15820_ (
    .A(\rf[6] [24]),
    .B(\rf[2] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08212_)
  );
  AND2_X1 _15821_ (
    .A1(_03049_),
    .A2(_08212_),
    .ZN(_08213_)
  );
  MUX2_X1 _15822_ (
    .A(\rf[4] [24]),
    .B(\rf[0] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08214_)
  );
  AND2_X1 _15823_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08214_),
    .ZN(_08215_)
  );
  OR2_X1 _15824_ (
    .A1(_03048_),
    .A2(_08215_),
    .ZN(_08216_)
  );
  OR2_X1 _15825_ (
    .A1(_08213_),
    .A2(_08216_),
    .ZN(_08217_)
  );
  MUX2_X1 _15826_ (
    .A(\rf[7] [24]),
    .B(\rf[3] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08218_)
  );
  AND2_X1 _15827_ (
    .A1(_03049_),
    .A2(_08218_),
    .ZN(_08219_)
  );
  MUX2_X1 _15828_ (
    .A(\rf[5] [24]),
    .B(\rf[1] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08220_)
  );
  AND2_X1 _15829_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08220_),
    .ZN(_08221_)
  );
  OR2_X1 _15830_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08221_),
    .ZN(_08222_)
  );
  OR2_X1 _15831_ (
    .A1(_08219_),
    .A2(_08222_),
    .ZN(_08223_)
  );
  AND2_X1 _15832_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_08223_),
    .ZN(_08224_)
  );
  AND2_X1 _15833_ (
    .A1(_08217_),
    .A2(_08224_),
    .ZN(_08225_)
  );
  OR2_X1 _15834_ (
    .A1(_08211_),
    .A2(_08225_),
    .ZN(_08226_)
  );
  OR2_X1 _15835_ (
    .A1(\rf[17] [24]),
    .A2(_03050_),
    .ZN(_08227_)
  );
  OR2_X1 _15836_ (
    .A1(\rf[21] [24]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08228_)
  );
  AND2_X1 _15837_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08228_),
    .ZN(_08229_)
  );
  AND2_X1 _15838_ (
    .A1(_08227_),
    .A2(_08229_),
    .ZN(_08230_)
  );
  MUX2_X1 _15839_ (
    .A(\rf[23] [24]),
    .B(\rf[19] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08231_)
  );
  AND2_X1 _15840_ (
    .A1(_03049_),
    .A2(_08231_),
    .ZN(_08232_)
  );
  OR2_X1 _15841_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08232_),
    .ZN(_08233_)
  );
  OR2_X1 _15842_ (
    .A1(_08230_),
    .A2(_08233_),
    .ZN(_08234_)
  );
  OR2_X1 _15843_ (
    .A1(\rf[20] [24]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08235_)
  );
  OR2_X1 _15844_ (
    .A1(\rf[16] [24]),
    .A2(_03050_),
    .ZN(_08236_)
  );
  AND2_X1 _15845_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08236_),
    .ZN(_08237_)
  );
  AND2_X1 _15846_ (
    .A1(_08235_),
    .A2(_08237_),
    .ZN(_08238_)
  );
  MUX2_X1 _15847_ (
    .A(\rf[22] [24]),
    .B(\rf[18] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08239_)
  );
  AND2_X1 _15848_ (
    .A1(_03049_),
    .A2(_08239_),
    .ZN(_08240_)
  );
  OR2_X1 _15849_ (
    .A1(_03048_),
    .A2(_08240_),
    .ZN(_08241_)
  );
  OR2_X1 _15850_ (
    .A1(_08238_),
    .A2(_08241_),
    .ZN(_08242_)
  );
  AND2_X1 _15851_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_08234_),
    .ZN(_08243_)
  );
  AND2_X1 _15852_ (
    .A1(_08242_),
    .A2(_08243_),
    .ZN(_08244_)
  );
  OR2_X1 _15853_ (
    .A1(\rf[28] [24]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08245_)
  );
  OR2_X1 _15854_ (
    .A1(\rf[24] [24]),
    .A2(_03050_),
    .ZN(_08246_)
  );
  AND2_X1 _15855_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08245_),
    .ZN(_08247_)
  );
  AND2_X1 _15856_ (
    .A1(_08246_),
    .A2(_08247_),
    .ZN(_08248_)
  );
  MUX2_X1 _15857_ (
    .A(\rf[30] [24]),
    .B(\rf[26] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08249_)
  );
  AND2_X1 _15858_ (
    .A1(_03049_),
    .A2(_08249_),
    .ZN(_08250_)
  );
  OR2_X1 _15859_ (
    .A1(_03048_),
    .A2(_08250_),
    .ZN(_08251_)
  );
  OR2_X1 _15860_ (
    .A1(_08248_),
    .A2(_08251_),
    .ZN(_08252_)
  );
  MUX2_X1 _15861_ (
    .A(\rf[29] [24]),
    .B(\rf[25] [24]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08253_)
  );
  AND2_X1 _15862_ (
    .A1(\rf[27] [24]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08254_)
  );
  MUX2_X1 _15863_ (
    .A(_08253_),
    .B(_08254_),
    .S(_03049_),
    .Z(_08255_)
  );
  OR2_X1 _15864_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08255_),
    .ZN(_08256_)
  );
  AND2_X1 _15865_ (
    .A1(_03051_),
    .A2(_08256_),
    .ZN(_08257_)
  );
  AND2_X1 _15866_ (
    .A1(_08252_),
    .A2(_08257_),
    .ZN(_08258_)
  );
  OR2_X1 _15867_ (
    .A1(_08244_),
    .A2(_08258_),
    .ZN(_08259_)
  );
  MUX2_X1 _15868_ (
    .A(_08226_),
    .B(_08259_),
    .S(_03064_),
    .Z(_08260_)
  );
  MUX2_X1 _15869_ (
    .A(_08260_),
    .B(_05665_),
    .S(_06791_),
    .Z(_08261_)
  );
  MUX2_X1 _15870_ (
    .A(ex_reg_rs_msb_1[22]),
    .B(_08261_),
    .S(_06781_),
    .Z(_00171_)
  );
  OR2_X1 _15871_ (
    .A1(\rf[10] [25]),
    .A2(_03050_),
    .ZN(_08262_)
  );
  OR2_X1 _15872_ (
    .A1(\rf[14] [25]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08263_)
  );
  AND2_X1 _15873_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08263_),
    .ZN(_08264_)
  );
  AND2_X1 _15874_ (
    .A1(_08262_),
    .A2(_08264_),
    .ZN(_08265_)
  );
  MUX2_X1 _15875_ (
    .A(\rf[15] [25]),
    .B(\rf[11] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08266_)
  );
  AND2_X1 _15876_ (
    .A1(_03048_),
    .A2(_08266_),
    .ZN(_08267_)
  );
  OR2_X1 _15877_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08267_),
    .ZN(_08268_)
  );
  OR2_X1 _15878_ (
    .A1(_08265_),
    .A2(_08268_),
    .ZN(_08269_)
  );
  OR2_X1 _15879_ (
    .A1(\rf[12] [25]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08270_)
  );
  OR2_X1 _15880_ (
    .A1(\rf[8] [25]),
    .A2(_03050_),
    .ZN(_08271_)
  );
  AND2_X1 _15881_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08270_),
    .ZN(_08272_)
  );
  AND2_X1 _15882_ (
    .A1(_08271_),
    .A2(_08272_),
    .ZN(_08273_)
  );
  MUX2_X1 _15883_ (
    .A(\rf[13] [25]),
    .B(\rf[9] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08274_)
  );
  AND2_X1 _15884_ (
    .A1(_03048_),
    .A2(_08274_),
    .ZN(_08275_)
  );
  OR2_X1 _15885_ (
    .A1(_03049_),
    .A2(_08275_),
    .ZN(_08276_)
  );
  OR2_X1 _15886_ (
    .A1(_08273_),
    .A2(_08276_),
    .ZN(_08277_)
  );
  AND2_X1 _15887_ (
    .A1(_03051_),
    .A2(_08277_),
    .ZN(_08278_)
  );
  AND2_X1 _15888_ (
    .A1(_08269_),
    .A2(_08278_),
    .ZN(_08279_)
  );
  MUX2_X1 _15889_ (
    .A(\rf[6] [25]),
    .B(\rf[2] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08280_)
  );
  AND2_X1 _15890_ (
    .A1(_03049_),
    .A2(_08280_),
    .ZN(_08281_)
  );
  MUX2_X1 _15891_ (
    .A(\rf[4] [25]),
    .B(\rf[0] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08282_)
  );
  AND2_X1 _15892_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08282_),
    .ZN(_08283_)
  );
  OR2_X1 _15893_ (
    .A1(_03048_),
    .A2(_08283_),
    .ZN(_08284_)
  );
  OR2_X1 _15894_ (
    .A1(_08281_),
    .A2(_08284_),
    .ZN(_08285_)
  );
  MUX2_X1 _15895_ (
    .A(\rf[7] [25]),
    .B(\rf[3] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08286_)
  );
  AND2_X1 _15896_ (
    .A1(_03049_),
    .A2(_08286_),
    .ZN(_08287_)
  );
  MUX2_X1 _15897_ (
    .A(\rf[5] [25]),
    .B(\rf[1] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08288_)
  );
  AND2_X1 _15898_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08288_),
    .ZN(_08289_)
  );
  OR2_X1 _15899_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08289_),
    .ZN(_08290_)
  );
  OR2_X1 _15900_ (
    .A1(_08287_),
    .A2(_08290_),
    .ZN(_08291_)
  );
  AND2_X1 _15901_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_08291_),
    .ZN(_08292_)
  );
  AND2_X1 _15902_ (
    .A1(_08285_),
    .A2(_08292_),
    .ZN(_08293_)
  );
  OR2_X1 _15903_ (
    .A1(_08279_),
    .A2(_08293_),
    .ZN(_08294_)
  );
  OR2_X1 _15904_ (
    .A1(\rf[17] [25]),
    .A2(_03050_),
    .ZN(_08295_)
  );
  OR2_X1 _15905_ (
    .A1(\rf[21] [25]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08296_)
  );
  AND2_X1 _15906_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08296_),
    .ZN(_08297_)
  );
  AND2_X1 _15907_ (
    .A1(_08295_),
    .A2(_08297_),
    .ZN(_08298_)
  );
  MUX2_X1 _15908_ (
    .A(\rf[23] [25]),
    .B(\rf[19] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08299_)
  );
  AND2_X1 _15909_ (
    .A1(_03049_),
    .A2(_08299_),
    .ZN(_08300_)
  );
  OR2_X1 _15910_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08300_),
    .ZN(_08301_)
  );
  OR2_X1 _15911_ (
    .A1(_08298_),
    .A2(_08301_),
    .ZN(_08302_)
  );
  OR2_X1 _15912_ (
    .A1(\rf[20] [25]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08303_)
  );
  OR2_X1 _15913_ (
    .A1(\rf[16] [25]),
    .A2(_03050_),
    .ZN(_08304_)
  );
  AND2_X1 _15914_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08304_),
    .ZN(_08305_)
  );
  AND2_X1 _15915_ (
    .A1(_08303_),
    .A2(_08305_),
    .ZN(_08306_)
  );
  MUX2_X1 _15916_ (
    .A(\rf[22] [25]),
    .B(\rf[18] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08307_)
  );
  AND2_X1 _15917_ (
    .A1(_03049_),
    .A2(_08307_),
    .ZN(_08308_)
  );
  OR2_X1 _15918_ (
    .A1(_03048_),
    .A2(_08308_),
    .ZN(_08309_)
  );
  OR2_X1 _15919_ (
    .A1(_08306_),
    .A2(_08309_),
    .ZN(_08310_)
  );
  AND2_X1 _15920_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_08302_),
    .ZN(_08311_)
  );
  AND2_X1 _15921_ (
    .A1(_08310_),
    .A2(_08311_),
    .ZN(_08312_)
  );
  OR2_X1 _15922_ (
    .A1(\rf[28] [25]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08313_)
  );
  OR2_X1 _15923_ (
    .A1(\rf[24] [25]),
    .A2(_03050_),
    .ZN(_08314_)
  );
  AND2_X1 _15924_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08313_),
    .ZN(_08315_)
  );
  AND2_X1 _15925_ (
    .A1(_08314_),
    .A2(_08315_),
    .ZN(_08316_)
  );
  MUX2_X1 _15926_ (
    .A(\rf[30] [25]),
    .B(\rf[26] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08317_)
  );
  AND2_X1 _15927_ (
    .A1(_03049_),
    .A2(_08317_),
    .ZN(_08318_)
  );
  OR2_X1 _15928_ (
    .A1(_03048_),
    .A2(_08318_),
    .ZN(_08319_)
  );
  OR2_X1 _15929_ (
    .A1(_08316_),
    .A2(_08319_),
    .ZN(_08320_)
  );
  MUX2_X1 _15930_ (
    .A(\rf[29] [25]),
    .B(\rf[25] [25]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08321_)
  );
  AND2_X1 _15931_ (
    .A1(\rf[27] [25]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08322_)
  );
  MUX2_X1 _15932_ (
    .A(_08321_),
    .B(_08322_),
    .S(_03049_),
    .Z(_08323_)
  );
  OR2_X1 _15933_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08323_),
    .ZN(_08324_)
  );
  AND2_X1 _15934_ (
    .A1(_03051_),
    .A2(_08324_),
    .ZN(_08325_)
  );
  AND2_X1 _15935_ (
    .A1(_08320_),
    .A2(_08325_),
    .ZN(_08326_)
  );
  OR2_X1 _15936_ (
    .A1(_08312_),
    .A2(_08326_),
    .ZN(_08327_)
  );
  MUX2_X1 _15937_ (
    .A(_08294_),
    .B(_08327_),
    .S(_03064_),
    .Z(_08328_)
  );
  MUX2_X1 _15938_ (
    .A(_08328_),
    .B(_05740_),
    .S(_06791_),
    .Z(_08329_)
  );
  MUX2_X1 _15939_ (
    .A(ex_reg_rs_msb_1[23]),
    .B(_08329_),
    .S(_06781_),
    .Z(_00172_)
  );
  MUX2_X1 _15940_ (
    .A(\rf[1] [26]),
    .B(\rf[0] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_08330_)
  );
  MUX2_X1 _15941_ (
    .A(\rf[5] [26]),
    .B(\rf[4] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_08331_)
  );
  MUX2_X1 _15942_ (
    .A(_08330_),
    .B(_08331_),
    .S(_03050_),
    .Z(_08332_)
  );
  OR2_X1 _15943_ (
    .A1(_03051_),
    .A2(_08332_),
    .ZN(_08333_)
  );
  MUX2_X1 _15944_ (
    .A(\rf[13] [26]),
    .B(\rf[9] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08334_)
  );
  OR2_X1 _15945_ (
    .A1(_03808_),
    .A2(_08334_),
    .ZN(_08335_)
  );
  MUX2_X1 _15946_ (
    .A(\rf[12] [26]),
    .B(\rf[8] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08336_)
  );
  OR2_X1 _15947_ (
    .A1(_06863_),
    .A2(_08336_),
    .ZN(_08337_)
  );
  AND2_X1 _15948_ (
    .A1(_08335_),
    .A2(_08337_),
    .ZN(_08338_)
  );
  AND2_X1 _15949_ (
    .A1(_08333_),
    .A2(_08338_),
    .ZN(_08339_)
  );
  MUX2_X1 _15950_ (
    .A(\rf[3] [26]),
    .B(\rf[2] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_08340_)
  );
  MUX2_X1 _15951_ (
    .A(\rf[7] [26]),
    .B(\rf[6] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_08341_)
  );
  MUX2_X1 _15952_ (
    .A(_08340_),
    .B(_08341_),
    .S(_03050_),
    .Z(_08342_)
  );
  OR2_X1 _15953_ (
    .A1(_03051_),
    .A2(_08342_),
    .ZN(_08343_)
  );
  MUX2_X1 _15954_ (
    .A(\rf[14] [26]),
    .B(\rf[10] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08344_)
  );
  OR2_X1 _15955_ (
    .A1(_06863_),
    .A2(_08344_),
    .ZN(_08345_)
  );
  MUX2_X1 _15956_ (
    .A(\rf[15] [26]),
    .B(\rf[11] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08346_)
  );
  OR2_X1 _15957_ (
    .A1(_03808_),
    .A2(_08346_),
    .ZN(_08347_)
  );
  AND2_X1 _15958_ (
    .A1(_08345_),
    .A2(_08347_),
    .ZN(_08348_)
  );
  AND2_X1 _15959_ (
    .A1(_08343_),
    .A2(_08348_),
    .ZN(_08349_)
  );
  MUX2_X1 _15960_ (
    .A(_08339_),
    .B(_08349_),
    .S(_03049_),
    .Z(_08350_)
  );
  OR2_X1 _15961_ (
    .A1(\rf[17] [26]),
    .A2(_03050_),
    .ZN(_08351_)
  );
  OR2_X1 _15962_ (
    .A1(\rf[21] [26]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08352_)
  );
  AND2_X1 _15963_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08352_),
    .ZN(_08353_)
  );
  AND2_X1 _15964_ (
    .A1(_08351_),
    .A2(_08353_),
    .ZN(_08354_)
  );
  MUX2_X1 _15965_ (
    .A(\rf[23] [26]),
    .B(\rf[19] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08355_)
  );
  AND2_X1 _15966_ (
    .A1(_03049_),
    .A2(_08355_),
    .ZN(_08356_)
  );
  OR2_X1 _15967_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08356_),
    .ZN(_08357_)
  );
  OR2_X1 _15968_ (
    .A1(_08354_),
    .A2(_08357_),
    .ZN(_08358_)
  );
  OR2_X1 _15969_ (
    .A1(\rf[20] [26]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08359_)
  );
  OR2_X1 _15970_ (
    .A1(\rf[16] [26]),
    .A2(_03050_),
    .ZN(_08360_)
  );
  AND2_X1 _15971_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08360_),
    .ZN(_08361_)
  );
  AND2_X1 _15972_ (
    .A1(_08359_),
    .A2(_08361_),
    .ZN(_08362_)
  );
  MUX2_X1 _15973_ (
    .A(\rf[22] [26]),
    .B(\rf[18] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08363_)
  );
  AND2_X1 _15974_ (
    .A1(_03049_),
    .A2(_08363_),
    .ZN(_08364_)
  );
  OR2_X1 _15975_ (
    .A1(_03048_),
    .A2(_08364_),
    .ZN(_08365_)
  );
  OR2_X1 _15976_ (
    .A1(_08362_),
    .A2(_08365_),
    .ZN(_08366_)
  );
  AND2_X1 _15977_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_08358_),
    .ZN(_08367_)
  );
  AND2_X1 _15978_ (
    .A1(_08366_),
    .A2(_08367_),
    .ZN(_08368_)
  );
  OR2_X1 _15979_ (
    .A1(\rf[28] [26]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08369_)
  );
  OR2_X1 _15980_ (
    .A1(\rf[24] [26]),
    .A2(_03050_),
    .ZN(_08370_)
  );
  AND2_X1 _15981_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08369_),
    .ZN(_08371_)
  );
  AND2_X1 _15982_ (
    .A1(_08370_),
    .A2(_08371_),
    .ZN(_08372_)
  );
  MUX2_X1 _15983_ (
    .A(\rf[30] [26]),
    .B(\rf[26] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08373_)
  );
  AND2_X1 _15984_ (
    .A1(_03049_),
    .A2(_08373_),
    .ZN(_08374_)
  );
  OR2_X1 _15985_ (
    .A1(_03048_),
    .A2(_08374_),
    .ZN(_08375_)
  );
  OR2_X1 _15986_ (
    .A1(_08372_),
    .A2(_08375_),
    .ZN(_08376_)
  );
  MUX2_X1 _15987_ (
    .A(\rf[29] [26]),
    .B(\rf[25] [26]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08377_)
  );
  AND2_X1 _15988_ (
    .A1(\rf[27] [26]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08378_)
  );
  MUX2_X1 _15989_ (
    .A(_08377_),
    .B(_08378_),
    .S(_03049_),
    .Z(_08379_)
  );
  OR2_X1 _15990_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08379_),
    .ZN(_08380_)
  );
  AND2_X1 _15991_ (
    .A1(_03051_),
    .A2(_08380_),
    .ZN(_08381_)
  );
  AND2_X1 _15992_ (
    .A1(_08376_),
    .A2(_08381_),
    .ZN(_08382_)
  );
  OR2_X1 _15993_ (
    .A1(_08368_),
    .A2(_08382_),
    .ZN(_08383_)
  );
  MUX2_X1 _15994_ (
    .A(_08350_),
    .B(_08383_),
    .S(_03064_),
    .Z(_08384_)
  );
  MUX2_X1 _15995_ (
    .A(_08384_),
    .B(_05882_),
    .S(_06791_),
    .Z(_08385_)
  );
  MUX2_X1 _15996_ (
    .A(ex_reg_rs_msb_1[24]),
    .B(_08385_),
    .S(_06781_),
    .Z(_00173_)
  );
  OR2_X1 _15997_ (
    .A1(\rf[10] [27]),
    .A2(_03050_),
    .ZN(_08386_)
  );
  OR2_X1 _15998_ (
    .A1(\rf[14] [27]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08387_)
  );
  AND2_X1 _15999_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08387_),
    .ZN(_08388_)
  );
  AND2_X1 _16000_ (
    .A1(_08386_),
    .A2(_08388_),
    .ZN(_08389_)
  );
  MUX2_X1 _16001_ (
    .A(\rf[15] [27]),
    .B(\rf[11] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08390_)
  );
  AND2_X1 _16002_ (
    .A1(_03048_),
    .A2(_08390_),
    .ZN(_08391_)
  );
  OR2_X1 _16003_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08391_),
    .ZN(_08392_)
  );
  OR2_X1 _16004_ (
    .A1(_08389_),
    .A2(_08392_),
    .ZN(_08393_)
  );
  OR2_X1 _16005_ (
    .A1(\rf[12] [27]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08394_)
  );
  OR2_X1 _16006_ (
    .A1(\rf[8] [27]),
    .A2(_03050_),
    .ZN(_08395_)
  );
  AND2_X1 _16007_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08394_),
    .ZN(_08396_)
  );
  AND2_X1 _16008_ (
    .A1(_08395_),
    .A2(_08396_),
    .ZN(_08397_)
  );
  MUX2_X1 _16009_ (
    .A(\rf[13] [27]),
    .B(\rf[9] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08398_)
  );
  AND2_X1 _16010_ (
    .A1(_03048_),
    .A2(_08398_),
    .ZN(_08399_)
  );
  OR2_X1 _16011_ (
    .A1(_03049_),
    .A2(_08399_),
    .ZN(_08400_)
  );
  OR2_X1 _16012_ (
    .A1(_08397_),
    .A2(_08400_),
    .ZN(_08401_)
  );
  AND2_X1 _16013_ (
    .A1(_03051_),
    .A2(_08401_),
    .ZN(_08402_)
  );
  AND2_X1 _16014_ (
    .A1(_08393_),
    .A2(_08402_),
    .ZN(_08403_)
  );
  MUX2_X1 _16015_ (
    .A(\rf[6] [27]),
    .B(\rf[2] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08404_)
  );
  AND2_X1 _16016_ (
    .A1(_03049_),
    .A2(_08404_),
    .ZN(_08405_)
  );
  MUX2_X1 _16017_ (
    .A(\rf[4] [27]),
    .B(\rf[0] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08406_)
  );
  AND2_X1 _16018_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08406_),
    .ZN(_08407_)
  );
  OR2_X1 _16019_ (
    .A1(_03048_),
    .A2(_08407_),
    .ZN(_08408_)
  );
  OR2_X1 _16020_ (
    .A1(_08405_),
    .A2(_08408_),
    .ZN(_08409_)
  );
  MUX2_X1 _16021_ (
    .A(\rf[7] [27]),
    .B(\rf[3] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08410_)
  );
  AND2_X1 _16022_ (
    .A1(_03049_),
    .A2(_08410_),
    .ZN(_08411_)
  );
  MUX2_X1 _16023_ (
    .A(\rf[5] [27]),
    .B(\rf[1] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08412_)
  );
  AND2_X1 _16024_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08412_),
    .ZN(_08413_)
  );
  OR2_X1 _16025_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08413_),
    .ZN(_08414_)
  );
  OR2_X1 _16026_ (
    .A1(_08411_),
    .A2(_08414_),
    .ZN(_08415_)
  );
  AND2_X1 _16027_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_08415_),
    .ZN(_08416_)
  );
  AND2_X1 _16028_ (
    .A1(_08409_),
    .A2(_08416_),
    .ZN(_08417_)
  );
  OR2_X1 _16029_ (
    .A1(_08403_),
    .A2(_08417_),
    .ZN(_08418_)
  );
  OR2_X1 _16030_ (
    .A1(\rf[17] [27]),
    .A2(_03050_),
    .ZN(_08419_)
  );
  OR2_X1 _16031_ (
    .A1(\rf[21] [27]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08420_)
  );
  AND2_X1 _16032_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08420_),
    .ZN(_08421_)
  );
  AND2_X1 _16033_ (
    .A1(_08419_),
    .A2(_08421_),
    .ZN(_08422_)
  );
  MUX2_X1 _16034_ (
    .A(\rf[23] [27]),
    .B(\rf[19] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08423_)
  );
  AND2_X1 _16035_ (
    .A1(_03049_),
    .A2(_08423_),
    .ZN(_08424_)
  );
  OR2_X1 _16036_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08424_),
    .ZN(_08425_)
  );
  OR2_X1 _16037_ (
    .A1(_08422_),
    .A2(_08425_),
    .ZN(_08426_)
  );
  OR2_X1 _16038_ (
    .A1(\rf[20] [27]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08427_)
  );
  OR2_X1 _16039_ (
    .A1(\rf[16] [27]),
    .A2(_03050_),
    .ZN(_08428_)
  );
  AND2_X1 _16040_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08428_),
    .ZN(_08429_)
  );
  AND2_X1 _16041_ (
    .A1(_08427_),
    .A2(_08429_),
    .ZN(_08430_)
  );
  MUX2_X1 _16042_ (
    .A(\rf[22] [27]),
    .B(\rf[18] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08431_)
  );
  AND2_X1 _16043_ (
    .A1(_03049_),
    .A2(_08431_),
    .ZN(_08432_)
  );
  OR2_X1 _16044_ (
    .A1(_03048_),
    .A2(_08432_),
    .ZN(_08433_)
  );
  OR2_X1 _16045_ (
    .A1(_08430_),
    .A2(_08433_),
    .ZN(_08434_)
  );
  AND2_X1 _16046_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_08426_),
    .ZN(_08435_)
  );
  AND2_X1 _16047_ (
    .A1(_08434_),
    .A2(_08435_),
    .ZN(_08436_)
  );
  OR2_X1 _16048_ (
    .A1(\rf[28] [27]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08437_)
  );
  OR2_X1 _16049_ (
    .A1(\rf[24] [27]),
    .A2(_03050_),
    .ZN(_08438_)
  );
  AND2_X1 _16050_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08437_),
    .ZN(_08439_)
  );
  AND2_X1 _16051_ (
    .A1(_08438_),
    .A2(_08439_),
    .ZN(_08440_)
  );
  MUX2_X1 _16052_ (
    .A(\rf[30] [27]),
    .B(\rf[26] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08441_)
  );
  AND2_X1 _16053_ (
    .A1(_03049_),
    .A2(_08441_),
    .ZN(_08442_)
  );
  OR2_X1 _16054_ (
    .A1(_03048_),
    .A2(_08442_),
    .ZN(_08443_)
  );
  OR2_X1 _16055_ (
    .A1(_08440_),
    .A2(_08443_),
    .ZN(_08444_)
  );
  MUX2_X1 _16056_ (
    .A(\rf[29] [27]),
    .B(\rf[25] [27]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08445_)
  );
  AND2_X1 _16057_ (
    .A1(\rf[27] [27]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08446_)
  );
  MUX2_X1 _16058_ (
    .A(_08445_),
    .B(_08446_),
    .S(_03049_),
    .Z(_08447_)
  );
  OR2_X1 _16059_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08447_),
    .ZN(_08448_)
  );
  AND2_X1 _16060_ (
    .A1(_03051_),
    .A2(_08448_),
    .ZN(_08449_)
  );
  AND2_X1 _16061_ (
    .A1(_08444_),
    .A2(_08449_),
    .ZN(_08450_)
  );
  OR2_X1 _16062_ (
    .A1(_08436_),
    .A2(_08450_),
    .ZN(_08451_)
  );
  MUX2_X1 _16063_ (
    .A(_08418_),
    .B(_08451_),
    .S(_03064_),
    .Z(_08452_)
  );
  MUX2_X1 _16064_ (
    .A(_08452_),
    .B(_05957_),
    .S(_06791_),
    .Z(_08453_)
  );
  MUX2_X1 _16065_ (
    .A(ex_reg_rs_msb_1[25]),
    .B(_08453_),
    .S(_06781_),
    .Z(_00174_)
  );
  OR2_X1 _16066_ (
    .A1(\rf[10] [28]),
    .A2(_03050_),
    .ZN(_08454_)
  );
  OR2_X1 _16067_ (
    .A1(\rf[14] [28]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08455_)
  );
  AND2_X1 _16068_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08455_),
    .ZN(_08456_)
  );
  AND2_X1 _16069_ (
    .A1(_08454_),
    .A2(_08456_),
    .ZN(_08457_)
  );
  MUX2_X1 _16070_ (
    .A(\rf[15] [28]),
    .B(\rf[11] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08458_)
  );
  AND2_X1 _16071_ (
    .A1(_03048_),
    .A2(_08458_),
    .ZN(_08459_)
  );
  OR2_X1 _16072_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08459_),
    .ZN(_08460_)
  );
  OR2_X1 _16073_ (
    .A1(_08457_),
    .A2(_08460_),
    .ZN(_08461_)
  );
  OR2_X1 _16074_ (
    .A1(\rf[12] [28]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08462_)
  );
  OR2_X1 _16075_ (
    .A1(\rf[8] [28]),
    .A2(_03050_),
    .ZN(_08463_)
  );
  AND2_X1 _16076_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08462_),
    .ZN(_08464_)
  );
  AND2_X1 _16077_ (
    .A1(_08463_),
    .A2(_08464_),
    .ZN(_08465_)
  );
  MUX2_X1 _16078_ (
    .A(\rf[13] [28]),
    .B(\rf[9] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08466_)
  );
  AND2_X1 _16079_ (
    .A1(_03048_),
    .A2(_08466_),
    .ZN(_08467_)
  );
  OR2_X1 _16080_ (
    .A1(_03049_),
    .A2(_08467_),
    .ZN(_08468_)
  );
  OR2_X1 _16081_ (
    .A1(_08465_),
    .A2(_08468_),
    .ZN(_08469_)
  );
  AND2_X1 _16082_ (
    .A1(_03051_),
    .A2(_08469_),
    .ZN(_08470_)
  );
  AND2_X1 _16083_ (
    .A1(_08461_),
    .A2(_08470_),
    .ZN(_08471_)
  );
  MUX2_X1 _16084_ (
    .A(\rf[6] [28]),
    .B(\rf[2] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08472_)
  );
  AND2_X1 _16085_ (
    .A1(_03049_),
    .A2(_08472_),
    .ZN(_08473_)
  );
  MUX2_X1 _16086_ (
    .A(\rf[4] [28]),
    .B(\rf[0] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08474_)
  );
  AND2_X1 _16087_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08474_),
    .ZN(_08475_)
  );
  OR2_X1 _16088_ (
    .A1(_03048_),
    .A2(_08475_),
    .ZN(_08476_)
  );
  OR2_X1 _16089_ (
    .A1(_08473_),
    .A2(_08476_),
    .ZN(_08477_)
  );
  MUX2_X1 _16090_ (
    .A(\rf[7] [28]),
    .B(\rf[3] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08478_)
  );
  AND2_X1 _16091_ (
    .A1(_03049_),
    .A2(_08478_),
    .ZN(_08479_)
  );
  MUX2_X1 _16092_ (
    .A(\rf[5] [28]),
    .B(\rf[1] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08480_)
  );
  AND2_X1 _16093_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08480_),
    .ZN(_08481_)
  );
  OR2_X1 _16094_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08481_),
    .ZN(_08482_)
  );
  OR2_X1 _16095_ (
    .A1(_08479_),
    .A2(_08482_),
    .ZN(_08483_)
  );
  AND2_X1 _16096_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_08483_),
    .ZN(_08484_)
  );
  AND2_X1 _16097_ (
    .A1(_08477_),
    .A2(_08484_),
    .ZN(_08485_)
  );
  OR2_X1 _16098_ (
    .A1(_08471_),
    .A2(_08485_),
    .ZN(_08486_)
  );
  OR2_X1 _16099_ (
    .A1(\rf[17] [28]),
    .A2(_03050_),
    .ZN(_08487_)
  );
  OR2_X1 _16100_ (
    .A1(\rf[21] [28]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08488_)
  );
  AND2_X1 _16101_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08488_),
    .ZN(_08489_)
  );
  AND2_X1 _16102_ (
    .A1(_08487_),
    .A2(_08489_),
    .ZN(_08490_)
  );
  MUX2_X1 _16103_ (
    .A(\rf[23] [28]),
    .B(\rf[19] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08491_)
  );
  AND2_X1 _16104_ (
    .A1(_03049_),
    .A2(_08491_),
    .ZN(_08492_)
  );
  OR2_X1 _16105_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08492_),
    .ZN(_08493_)
  );
  OR2_X1 _16106_ (
    .A1(_08490_),
    .A2(_08493_),
    .ZN(_08494_)
  );
  OR2_X1 _16107_ (
    .A1(\rf[20] [28]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08495_)
  );
  OR2_X1 _16108_ (
    .A1(\rf[16] [28]),
    .A2(_03050_),
    .ZN(_08496_)
  );
  AND2_X1 _16109_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08496_),
    .ZN(_08497_)
  );
  AND2_X1 _16110_ (
    .A1(_08495_),
    .A2(_08497_),
    .ZN(_08498_)
  );
  MUX2_X1 _16111_ (
    .A(\rf[22] [28]),
    .B(\rf[18] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08499_)
  );
  AND2_X1 _16112_ (
    .A1(_03049_),
    .A2(_08499_),
    .ZN(_08500_)
  );
  OR2_X1 _16113_ (
    .A1(_03048_),
    .A2(_08500_),
    .ZN(_08501_)
  );
  OR2_X1 _16114_ (
    .A1(_08498_),
    .A2(_08501_),
    .ZN(_08502_)
  );
  AND2_X1 _16115_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_08494_),
    .ZN(_08503_)
  );
  AND2_X1 _16116_ (
    .A1(_08502_),
    .A2(_08503_),
    .ZN(_08504_)
  );
  OR2_X1 _16117_ (
    .A1(\rf[28] [28]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08505_)
  );
  OR2_X1 _16118_ (
    .A1(\rf[24] [28]),
    .A2(_03050_),
    .ZN(_08506_)
  );
  AND2_X1 _16119_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08505_),
    .ZN(_08507_)
  );
  AND2_X1 _16120_ (
    .A1(_08506_),
    .A2(_08507_),
    .ZN(_08508_)
  );
  MUX2_X1 _16121_ (
    .A(\rf[30] [28]),
    .B(\rf[26] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08509_)
  );
  AND2_X1 _16122_ (
    .A1(_03049_),
    .A2(_08509_),
    .ZN(_08510_)
  );
  OR2_X1 _16123_ (
    .A1(_03048_),
    .A2(_08510_),
    .ZN(_08511_)
  );
  OR2_X1 _16124_ (
    .A1(_08508_),
    .A2(_08511_),
    .ZN(_08512_)
  );
  MUX2_X1 _16125_ (
    .A(\rf[29] [28]),
    .B(\rf[25] [28]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08513_)
  );
  AND2_X1 _16126_ (
    .A1(\rf[27] [28]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08514_)
  );
  MUX2_X1 _16127_ (
    .A(_08513_),
    .B(_08514_),
    .S(_03049_),
    .Z(_08515_)
  );
  OR2_X1 _16128_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08515_),
    .ZN(_08516_)
  );
  AND2_X1 _16129_ (
    .A1(_03051_),
    .A2(_08516_),
    .ZN(_08517_)
  );
  AND2_X1 _16130_ (
    .A1(_08512_),
    .A2(_08517_),
    .ZN(_08518_)
  );
  OR2_X1 _16131_ (
    .A1(_08504_),
    .A2(_08518_),
    .ZN(_08519_)
  );
  MUX2_X1 _16132_ (
    .A(_08486_),
    .B(_08519_),
    .S(_03064_),
    .Z(_08520_)
  );
  MUX2_X1 _16133_ (
    .A(_08520_),
    .B(_06032_),
    .S(_06791_),
    .Z(_08521_)
  );
  MUX2_X1 _16134_ (
    .A(ex_reg_rs_msb_1[26]),
    .B(_08521_),
    .S(_06781_),
    .Z(_00175_)
  );
  MUX2_X1 _16135_ (
    .A(\rf[1] [29]),
    .B(\rf[0] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_08522_)
  );
  MUX2_X1 _16136_ (
    .A(\rf[5] [29]),
    .B(\rf[4] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_08523_)
  );
  MUX2_X1 _16137_ (
    .A(_08522_),
    .B(_08523_),
    .S(_03050_),
    .Z(_08524_)
  );
  OR2_X1 _16138_ (
    .A1(_03051_),
    .A2(_08524_),
    .ZN(_08525_)
  );
  MUX2_X1 _16139_ (
    .A(\rf[12] [29]),
    .B(\rf[8] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08526_)
  );
  OR2_X1 _16140_ (
    .A1(_06863_),
    .A2(_08526_),
    .ZN(_08527_)
  );
  MUX2_X1 _16141_ (
    .A(\rf[13] [29]),
    .B(\rf[9] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08528_)
  );
  OR2_X1 _16142_ (
    .A1(_03808_),
    .A2(_08528_),
    .ZN(_08529_)
  );
  AND2_X1 _16143_ (
    .A1(_08527_),
    .A2(_08529_),
    .ZN(_08530_)
  );
  AND2_X1 _16144_ (
    .A1(_08525_),
    .A2(_08530_),
    .ZN(_08531_)
  );
  MUX2_X1 _16145_ (
    .A(\rf[3] [29]),
    .B(\rf[2] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_08532_)
  );
  MUX2_X1 _16146_ (
    .A(\rf[7] [29]),
    .B(\rf[6] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs2[0]),
    .Z(_08533_)
  );
  MUX2_X1 _16147_ (
    .A(_08532_),
    .B(_08533_),
    .S(_03050_),
    .Z(_08534_)
  );
  OR2_X1 _16148_ (
    .A1(_03051_),
    .A2(_08534_),
    .ZN(_08535_)
  );
  MUX2_X1 _16149_ (
    .A(\rf[14] [29]),
    .B(\rf[10] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08536_)
  );
  OR2_X1 _16150_ (
    .A1(_06863_),
    .A2(_08536_),
    .ZN(_08537_)
  );
  MUX2_X1 _16151_ (
    .A(\rf[15] [29]),
    .B(\rf[11] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08538_)
  );
  OR2_X1 _16152_ (
    .A1(_03808_),
    .A2(_08538_),
    .ZN(_08539_)
  );
  AND2_X1 _16153_ (
    .A1(_08537_),
    .A2(_08539_),
    .ZN(_08540_)
  );
  AND2_X1 _16154_ (
    .A1(_08535_),
    .A2(_08540_),
    .ZN(_08541_)
  );
  MUX2_X1 _16155_ (
    .A(_08531_),
    .B(_08541_),
    .S(_03049_),
    .Z(_08542_)
  );
  OR2_X1 _16156_ (
    .A1(\rf[17] [29]),
    .A2(_03050_),
    .ZN(_08543_)
  );
  OR2_X1 _16157_ (
    .A1(\rf[21] [29]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08544_)
  );
  AND2_X1 _16158_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08544_),
    .ZN(_08545_)
  );
  AND2_X1 _16159_ (
    .A1(_08543_),
    .A2(_08545_),
    .ZN(_08546_)
  );
  MUX2_X1 _16160_ (
    .A(\rf[23] [29]),
    .B(\rf[19] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08547_)
  );
  AND2_X1 _16161_ (
    .A1(_03049_),
    .A2(_08547_),
    .ZN(_08548_)
  );
  OR2_X1 _16162_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08548_),
    .ZN(_08549_)
  );
  OR2_X1 _16163_ (
    .A1(_08546_),
    .A2(_08549_),
    .ZN(_08550_)
  );
  OR2_X1 _16164_ (
    .A1(\rf[20] [29]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08551_)
  );
  OR2_X1 _16165_ (
    .A1(\rf[16] [29]),
    .A2(_03050_),
    .ZN(_08552_)
  );
  AND2_X1 _16166_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08552_),
    .ZN(_08553_)
  );
  AND2_X1 _16167_ (
    .A1(_08551_),
    .A2(_08553_),
    .ZN(_08554_)
  );
  MUX2_X1 _16168_ (
    .A(\rf[22] [29]),
    .B(\rf[18] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08555_)
  );
  AND2_X1 _16169_ (
    .A1(_03049_),
    .A2(_08555_),
    .ZN(_08556_)
  );
  OR2_X1 _16170_ (
    .A1(_03048_),
    .A2(_08556_),
    .ZN(_08557_)
  );
  OR2_X1 _16171_ (
    .A1(_08554_),
    .A2(_08557_),
    .ZN(_08558_)
  );
  AND2_X1 _16172_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_08550_),
    .ZN(_08559_)
  );
  AND2_X1 _16173_ (
    .A1(_08558_),
    .A2(_08559_),
    .ZN(_08560_)
  );
  OR2_X1 _16174_ (
    .A1(\rf[28] [29]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08561_)
  );
  OR2_X1 _16175_ (
    .A1(\rf[24] [29]),
    .A2(_03050_),
    .ZN(_08562_)
  );
  AND2_X1 _16176_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08561_),
    .ZN(_08563_)
  );
  AND2_X1 _16177_ (
    .A1(_08562_),
    .A2(_08563_),
    .ZN(_08564_)
  );
  MUX2_X1 _16178_ (
    .A(\rf[30] [29]),
    .B(\rf[26] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08565_)
  );
  AND2_X1 _16179_ (
    .A1(_03049_),
    .A2(_08565_),
    .ZN(_08566_)
  );
  OR2_X1 _16180_ (
    .A1(_03048_),
    .A2(_08566_),
    .ZN(_08567_)
  );
  OR2_X1 _16181_ (
    .A1(_08564_),
    .A2(_08567_),
    .ZN(_08568_)
  );
  MUX2_X1 _16182_ (
    .A(\rf[29] [29]),
    .B(\rf[25] [29]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08569_)
  );
  AND2_X1 _16183_ (
    .A1(\rf[27] [29]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08570_)
  );
  MUX2_X1 _16184_ (
    .A(_08569_),
    .B(_08570_),
    .S(_03049_),
    .Z(_08571_)
  );
  OR2_X1 _16185_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08571_),
    .ZN(_08572_)
  );
  AND2_X1 _16186_ (
    .A1(_03051_),
    .A2(_08572_),
    .ZN(_08573_)
  );
  AND2_X1 _16187_ (
    .A1(_08568_),
    .A2(_08573_),
    .ZN(_08574_)
  );
  OR2_X1 _16188_ (
    .A1(_08560_),
    .A2(_08574_),
    .ZN(_08575_)
  );
  MUX2_X1 _16189_ (
    .A(_08542_),
    .B(_08575_),
    .S(_03064_),
    .Z(_08576_)
  );
  MUX2_X1 _16190_ (
    .A(_08576_),
    .B(_06109_),
    .S(_06791_),
    .Z(_08577_)
  );
  MUX2_X1 _16191_ (
    .A(ex_reg_rs_msb_1[27]),
    .B(_08577_),
    .S(_06781_),
    .Z(_00176_)
  );
  OR2_X1 _16192_ (
    .A1(\rf[10] [30]),
    .A2(_03050_),
    .ZN(_08578_)
  );
  OR2_X1 _16193_ (
    .A1(\rf[14] [30]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08579_)
  );
  AND2_X1 _16194_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08579_),
    .ZN(_08580_)
  );
  AND2_X1 _16195_ (
    .A1(_08578_),
    .A2(_08580_),
    .ZN(_08581_)
  );
  MUX2_X1 _16196_ (
    .A(\rf[15] [30]),
    .B(\rf[11] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08582_)
  );
  AND2_X1 _16197_ (
    .A1(_03048_),
    .A2(_08582_),
    .ZN(_08583_)
  );
  OR2_X1 _16198_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08583_),
    .ZN(_08584_)
  );
  OR2_X1 _16199_ (
    .A1(_08581_),
    .A2(_08584_),
    .ZN(_08585_)
  );
  OR2_X1 _16200_ (
    .A1(\rf[12] [30]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08586_)
  );
  OR2_X1 _16201_ (
    .A1(\rf[8] [30]),
    .A2(_03050_),
    .ZN(_08587_)
  );
  AND2_X1 _16202_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08586_),
    .ZN(_08588_)
  );
  AND2_X1 _16203_ (
    .A1(_08587_),
    .A2(_08588_),
    .ZN(_08589_)
  );
  MUX2_X1 _16204_ (
    .A(\rf[13] [30]),
    .B(\rf[9] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08590_)
  );
  AND2_X1 _16205_ (
    .A1(_03048_),
    .A2(_08590_),
    .ZN(_08591_)
  );
  OR2_X1 _16206_ (
    .A1(_03049_),
    .A2(_08591_),
    .ZN(_08592_)
  );
  OR2_X1 _16207_ (
    .A1(_08589_),
    .A2(_08592_),
    .ZN(_08593_)
  );
  AND2_X1 _16208_ (
    .A1(_03051_),
    .A2(_08593_),
    .ZN(_08594_)
  );
  AND2_X1 _16209_ (
    .A1(_08585_),
    .A2(_08594_),
    .ZN(_08595_)
  );
  MUX2_X1 _16210_ (
    .A(\rf[6] [30]),
    .B(\rf[2] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08596_)
  );
  AND2_X1 _16211_ (
    .A1(_03049_),
    .A2(_08596_),
    .ZN(_08597_)
  );
  MUX2_X1 _16212_ (
    .A(\rf[4] [30]),
    .B(\rf[0] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08598_)
  );
  AND2_X1 _16213_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08598_),
    .ZN(_08599_)
  );
  OR2_X1 _16214_ (
    .A1(_03048_),
    .A2(_08599_),
    .ZN(_08600_)
  );
  OR2_X1 _16215_ (
    .A1(_08597_),
    .A2(_08600_),
    .ZN(_08601_)
  );
  MUX2_X1 _16216_ (
    .A(\rf[7] [30]),
    .B(\rf[3] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08602_)
  );
  AND2_X1 _16217_ (
    .A1(_03049_),
    .A2(_08602_),
    .ZN(_08603_)
  );
  MUX2_X1 _16218_ (
    .A(\rf[5] [30]),
    .B(\rf[1] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08604_)
  );
  AND2_X1 _16219_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08604_),
    .ZN(_08605_)
  );
  OR2_X1 _16220_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08605_),
    .ZN(_08606_)
  );
  OR2_X1 _16221_ (
    .A1(_08603_),
    .A2(_08606_),
    .ZN(_08607_)
  );
  AND2_X1 _16222_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_08607_),
    .ZN(_08608_)
  );
  AND2_X1 _16223_ (
    .A1(_08601_),
    .A2(_08608_),
    .ZN(_08609_)
  );
  OR2_X1 _16224_ (
    .A1(_08595_),
    .A2(_08609_),
    .ZN(_08610_)
  );
  OR2_X1 _16225_ (
    .A1(\rf[17] [30]),
    .A2(_03050_),
    .ZN(_08611_)
  );
  OR2_X1 _16226_ (
    .A1(\rf[21] [30]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08612_)
  );
  AND2_X1 _16227_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08612_),
    .ZN(_08613_)
  );
  AND2_X1 _16228_ (
    .A1(_08611_),
    .A2(_08613_),
    .ZN(_08614_)
  );
  MUX2_X1 _16229_ (
    .A(\rf[23] [30]),
    .B(\rf[19] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08615_)
  );
  AND2_X1 _16230_ (
    .A1(_03049_),
    .A2(_08615_),
    .ZN(_08616_)
  );
  OR2_X1 _16231_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08616_),
    .ZN(_08617_)
  );
  OR2_X1 _16232_ (
    .A1(_08614_),
    .A2(_08617_),
    .ZN(_08618_)
  );
  OR2_X1 _16233_ (
    .A1(\rf[20] [30]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08619_)
  );
  OR2_X1 _16234_ (
    .A1(\rf[16] [30]),
    .A2(_03050_),
    .ZN(_08620_)
  );
  AND2_X1 _16235_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08620_),
    .ZN(_08621_)
  );
  AND2_X1 _16236_ (
    .A1(_08619_),
    .A2(_08621_),
    .ZN(_08622_)
  );
  MUX2_X1 _16237_ (
    .A(\rf[22] [30]),
    .B(\rf[18] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08623_)
  );
  AND2_X1 _16238_ (
    .A1(_03049_),
    .A2(_08623_),
    .ZN(_08624_)
  );
  OR2_X1 _16239_ (
    .A1(_03048_),
    .A2(_08624_),
    .ZN(_08625_)
  );
  OR2_X1 _16240_ (
    .A1(_08622_),
    .A2(_08625_),
    .ZN(_08626_)
  );
  AND2_X1 _16241_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_08618_),
    .ZN(_08627_)
  );
  AND2_X1 _16242_ (
    .A1(_08626_),
    .A2(_08627_),
    .ZN(_08628_)
  );
  OR2_X1 _16243_ (
    .A1(\rf[28] [30]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08629_)
  );
  OR2_X1 _16244_ (
    .A1(\rf[24] [30]),
    .A2(_03050_),
    .ZN(_08630_)
  );
  AND2_X1 _16245_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08629_),
    .ZN(_08631_)
  );
  AND2_X1 _16246_ (
    .A1(_08630_),
    .A2(_08631_),
    .ZN(_08632_)
  );
  MUX2_X1 _16247_ (
    .A(\rf[30] [30]),
    .B(\rf[26] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08633_)
  );
  AND2_X1 _16248_ (
    .A1(_03049_),
    .A2(_08633_),
    .ZN(_08634_)
  );
  OR2_X1 _16249_ (
    .A1(_03048_),
    .A2(_08634_),
    .ZN(_08635_)
  );
  OR2_X1 _16250_ (
    .A1(_08632_),
    .A2(_08635_),
    .ZN(_08636_)
  );
  MUX2_X1 _16251_ (
    .A(\rf[29] [30]),
    .B(\rf[25] [30]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08637_)
  );
  AND2_X1 _16252_ (
    .A1(\rf[27] [30]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08638_)
  );
  MUX2_X1 _16253_ (
    .A(_08637_),
    .B(_08638_),
    .S(_03049_),
    .Z(_08639_)
  );
  OR2_X1 _16254_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08639_),
    .ZN(_08640_)
  );
  AND2_X1 _16255_ (
    .A1(_03051_),
    .A2(_08640_),
    .ZN(_08641_)
  );
  AND2_X1 _16256_ (
    .A1(_08636_),
    .A2(_08641_),
    .ZN(_08642_)
  );
  OR2_X1 _16257_ (
    .A1(_08628_),
    .A2(_08642_),
    .ZN(_08643_)
  );
  MUX2_X1 _16258_ (
    .A(_08610_),
    .B(_08643_),
    .S(_03064_),
    .Z(_08644_)
  );
  MUX2_X1 _16259_ (
    .A(_08644_),
    .B(_06117_),
    .S(_06791_),
    .Z(_08645_)
  );
  MUX2_X1 _16260_ (
    .A(ex_reg_rs_msb_1[28]),
    .B(_08645_),
    .S(_06781_),
    .Z(_00177_)
  );
  OR2_X1 _16261_ (
    .A1(\rf[10] [31]),
    .A2(_03050_),
    .ZN(_08646_)
  );
  OR2_X1 _16262_ (
    .A1(\rf[14] [31]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08647_)
  );
  AND2_X1 _16263_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08647_),
    .ZN(_08648_)
  );
  AND2_X1 _16264_ (
    .A1(_08646_),
    .A2(_08648_),
    .ZN(_08649_)
  );
  MUX2_X1 _16265_ (
    .A(\rf[15] [31]),
    .B(\rf[11] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08650_)
  );
  AND2_X1 _16266_ (
    .A1(_03048_),
    .A2(_08650_),
    .ZN(_08651_)
  );
  OR2_X1 _16267_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08651_),
    .ZN(_08652_)
  );
  OR2_X1 _16268_ (
    .A1(_08649_),
    .A2(_08652_),
    .ZN(_08653_)
  );
  OR2_X1 _16269_ (
    .A1(\rf[12] [31]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08654_)
  );
  OR2_X1 _16270_ (
    .A1(\rf[8] [31]),
    .A2(_03050_),
    .ZN(_08655_)
  );
  AND2_X1 _16271_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08654_),
    .ZN(_08656_)
  );
  AND2_X1 _16272_ (
    .A1(_08655_),
    .A2(_08656_),
    .ZN(_08657_)
  );
  MUX2_X1 _16273_ (
    .A(\rf[13] [31]),
    .B(\rf[9] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08658_)
  );
  AND2_X1 _16274_ (
    .A1(_03048_),
    .A2(_08658_),
    .ZN(_08659_)
  );
  OR2_X1 _16275_ (
    .A1(_03049_),
    .A2(_08659_),
    .ZN(_08660_)
  );
  OR2_X1 _16276_ (
    .A1(_08657_),
    .A2(_08660_),
    .ZN(_08661_)
  );
  AND2_X1 _16277_ (
    .A1(_03051_),
    .A2(_08661_),
    .ZN(_08662_)
  );
  AND2_X1 _16278_ (
    .A1(_08653_),
    .A2(_08662_),
    .ZN(_08663_)
  );
  MUX2_X1 _16279_ (
    .A(\rf[6] [31]),
    .B(\rf[2] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08664_)
  );
  AND2_X1 _16280_ (
    .A1(_03049_),
    .A2(_08664_),
    .ZN(_08665_)
  );
  MUX2_X1 _16281_ (
    .A(\rf[4] [31]),
    .B(\rf[0] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08666_)
  );
  AND2_X1 _16282_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08666_),
    .ZN(_08667_)
  );
  OR2_X1 _16283_ (
    .A1(_03048_),
    .A2(_08667_),
    .ZN(_08668_)
  );
  OR2_X1 _16284_ (
    .A1(_08665_),
    .A2(_08668_),
    .ZN(_08669_)
  );
  MUX2_X1 _16285_ (
    .A(\rf[7] [31]),
    .B(\rf[3] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08670_)
  );
  AND2_X1 _16286_ (
    .A1(_03049_),
    .A2(_08670_),
    .ZN(_08671_)
  );
  MUX2_X1 _16287_ (
    .A(\rf[5] [31]),
    .B(\rf[1] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08672_)
  );
  AND2_X1 _16288_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08672_),
    .ZN(_08673_)
  );
  OR2_X1 _16289_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08673_),
    .ZN(_08674_)
  );
  OR2_X1 _16290_ (
    .A1(_08671_),
    .A2(_08674_),
    .ZN(_08675_)
  );
  AND2_X1 _16291_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_08675_),
    .ZN(_08676_)
  );
  AND2_X1 _16292_ (
    .A1(_08669_),
    .A2(_08676_),
    .ZN(_08677_)
  );
  OR2_X1 _16293_ (
    .A1(_08663_),
    .A2(_08677_),
    .ZN(_08678_)
  );
  OR2_X1 _16294_ (
    .A1(\rf[17] [31]),
    .A2(_03050_),
    .ZN(_08679_)
  );
  OR2_X1 _16295_ (
    .A1(\rf[21] [31]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08680_)
  );
  AND2_X1 _16296_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08680_),
    .ZN(_08681_)
  );
  AND2_X1 _16297_ (
    .A1(_08679_),
    .A2(_08681_),
    .ZN(_08682_)
  );
  MUX2_X1 _16298_ (
    .A(\rf[23] [31]),
    .B(\rf[19] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08683_)
  );
  AND2_X1 _16299_ (
    .A1(_03049_),
    .A2(_08683_),
    .ZN(_08684_)
  );
  OR2_X1 _16300_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08684_),
    .ZN(_08685_)
  );
  OR2_X1 _16301_ (
    .A1(_08682_),
    .A2(_08685_),
    .ZN(_08686_)
  );
  OR2_X1 _16302_ (
    .A1(\rf[20] [31]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08687_)
  );
  OR2_X1 _16303_ (
    .A1(\rf[16] [31]),
    .A2(_03050_),
    .ZN(_08688_)
  );
  AND2_X1 _16304_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08688_),
    .ZN(_08689_)
  );
  AND2_X1 _16305_ (
    .A1(_08687_),
    .A2(_08689_),
    .ZN(_08690_)
  );
  MUX2_X1 _16306_ (
    .A(\rf[22] [31]),
    .B(\rf[18] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08691_)
  );
  AND2_X1 _16307_ (
    .A1(_03049_),
    .A2(_08691_),
    .ZN(_08692_)
  );
  OR2_X1 _16308_ (
    .A1(_03048_),
    .A2(_08692_),
    .ZN(_08693_)
  );
  OR2_X1 _16309_ (
    .A1(_08690_),
    .A2(_08693_),
    .ZN(_08694_)
  );
  AND2_X1 _16310_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_08686_),
    .ZN(_08695_)
  );
  AND2_X1 _16311_ (
    .A1(_08694_),
    .A2(_08695_),
    .ZN(_08696_)
  );
  OR2_X1 _16312_ (
    .A1(\rf[28] [31]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08697_)
  );
  OR2_X1 _16313_ (
    .A1(\rf[24] [31]),
    .A2(_03050_),
    .ZN(_08698_)
  );
  AND2_X1 _16314_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_08697_),
    .ZN(_08699_)
  );
  AND2_X1 _16315_ (
    .A1(_08698_),
    .A2(_08699_),
    .ZN(_08700_)
  );
  MUX2_X1 _16316_ (
    .A(\rf[30] [31]),
    .B(\rf[26] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08701_)
  );
  AND2_X1 _16317_ (
    .A1(_03049_),
    .A2(_08701_),
    .ZN(_08702_)
  );
  OR2_X1 _16318_ (
    .A1(_03048_),
    .A2(_08702_),
    .ZN(_08703_)
  );
  OR2_X1 _16319_ (
    .A1(_08700_),
    .A2(_08703_),
    .ZN(_08704_)
  );
  MUX2_X1 _16320_ (
    .A(\rf[29] [31]),
    .B(\rf[25] [31]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_08705_)
  );
  AND2_X1 _16321_ (
    .A1(\rf[27] [31]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_08706_)
  );
  MUX2_X1 _16322_ (
    .A(_08705_),
    .B(_08706_),
    .S(_03049_),
    .Z(_08707_)
  );
  OR2_X1 _16323_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_08707_),
    .ZN(_08708_)
  );
  AND2_X1 _16324_ (
    .A1(_03051_),
    .A2(_08708_),
    .ZN(_08709_)
  );
  AND2_X1 _16325_ (
    .A1(_08704_),
    .A2(_08709_),
    .ZN(_08710_)
  );
  OR2_X1 _16326_ (
    .A1(_08696_),
    .A2(_08710_),
    .ZN(_08711_)
  );
  MUX2_X1 _16327_ (
    .A(_08678_),
    .B(_08711_),
    .S(_03064_),
    .Z(_08712_)
  );
  MUX2_X1 _16328_ (
    .A(_08712_),
    .B(_06192_),
    .S(_06791_),
    .Z(_08713_)
  );
  MUX2_X1 _16329_ (
    .A(ex_reg_rs_msb_1[29]),
    .B(_08713_),
    .S(_06781_),
    .Z(_00178_)
  );
  OR2_X1 _16330_ (
    .A1(ibuf_io_inst_0_bits_xcpt1_ae_inst),
    .A2(ibuf_io_inst_0_bits_xcpt1_gf_inst),
    .ZN(_08714_)
  );
  OR2_X1 _16331_ (
    .A1(ibuf_io_inst_0_bits_xcpt1_pf_inst),
    .A2(_08714_),
    .ZN(_08715_)
  );
  INV_X1 _16332_ (
    .A(_08715_),
    .ZN(_08716_)
  );
  OR2_X1 _16333_ (
    .A1(ibuf_io_inst_0_bits_rvc),
    .A2(_08715_),
    .ZN(_08717_)
  );
  MUX2_X1 _16334_ (
    .A(_08717_),
    .B(ex_reg_rvc),
    .S(_04146_),
    .Z(_00179_)
  );
  OR2_X1 _16335_ (
    .A1(mem_reg_xcpt),
    .A2(mem_reg_xcpt_interrupt),
    .ZN(_08718_)
  );
  INV_X1 _16336_ (
    .A(_08718_),
    .ZN(_08719_)
  );
  AND2_X1 _16337_ (
    .A1(mem_reg_cause[4]),
    .A2(_08718_),
    .ZN(_08720_)
  );
  MUX2_X1 _16338_ (
    .A(wb_reg_cause[4]),
    .B(_08720_),
    .S(_06433_),
    .Z(_00180_)
  );
  AND2_X1 _16339_ (
    .A1(mem_reg_cause[5]),
    .A2(_08718_),
    .ZN(_08721_)
  );
  MUX2_X1 _16340_ (
    .A(wb_reg_cause[5]),
    .B(_08721_),
    .S(_06433_),
    .Z(_00181_)
  );
  AND2_X1 _16341_ (
    .A1(mem_reg_cause[6]),
    .A2(_08718_),
    .ZN(_08722_)
  );
  MUX2_X1 _16342_ (
    .A(wb_reg_cause[6]),
    .B(_08722_),
    .S(_06433_),
    .Z(_00182_)
  );
  AND2_X1 _16343_ (
    .A1(mem_reg_cause[7]),
    .A2(_08718_),
    .ZN(_08723_)
  );
  MUX2_X1 _16344_ (
    .A(wb_reg_cause[7]),
    .B(_08723_),
    .S(_06433_),
    .Z(_00183_)
  );
  AND2_X1 _16345_ (
    .A1(mem_reg_cause[8]),
    .A2(_08718_),
    .ZN(_08724_)
  );
  MUX2_X1 _16346_ (
    .A(wb_reg_cause[8]),
    .B(_08724_),
    .S(_06433_),
    .Z(_00184_)
  );
  AND2_X1 _16347_ (
    .A1(mem_reg_cause[9]),
    .A2(_08718_),
    .ZN(_08725_)
  );
  MUX2_X1 _16348_ (
    .A(wb_reg_cause[9]),
    .B(_08725_),
    .S(_06433_),
    .Z(_00185_)
  );
  AND2_X1 _16349_ (
    .A1(mem_reg_cause[10]),
    .A2(_08718_),
    .ZN(_08726_)
  );
  MUX2_X1 _16350_ (
    .A(wb_reg_cause[10]),
    .B(_08726_),
    .S(_06433_),
    .Z(_00186_)
  );
  AND2_X1 _16351_ (
    .A1(mem_reg_cause[11]),
    .A2(_08718_),
    .ZN(_08727_)
  );
  MUX2_X1 _16352_ (
    .A(wb_reg_cause[11]),
    .B(_08727_),
    .S(_06433_),
    .Z(_00187_)
  );
  AND2_X1 _16353_ (
    .A1(mem_reg_cause[12]),
    .A2(_08718_),
    .ZN(_08728_)
  );
  MUX2_X1 _16354_ (
    .A(wb_reg_cause[12]),
    .B(_08728_),
    .S(_06433_),
    .Z(_00188_)
  );
  AND2_X1 _16355_ (
    .A1(mem_reg_cause[13]),
    .A2(_08718_),
    .ZN(_08729_)
  );
  MUX2_X1 _16356_ (
    .A(wb_reg_cause[13]),
    .B(_08729_),
    .S(_06433_),
    .Z(_00189_)
  );
  AND2_X1 _16357_ (
    .A1(mem_reg_cause[14]),
    .A2(_08718_),
    .ZN(_08730_)
  );
  MUX2_X1 _16358_ (
    .A(wb_reg_cause[14]),
    .B(_08730_),
    .S(_06433_),
    .Z(_00190_)
  );
  AND2_X1 _16359_ (
    .A1(mem_reg_cause[15]),
    .A2(_08718_),
    .ZN(_08731_)
  );
  MUX2_X1 _16360_ (
    .A(wb_reg_cause[15]),
    .B(_08731_),
    .S(_06433_),
    .Z(_00191_)
  );
  AND2_X1 _16361_ (
    .A1(mem_reg_cause[16]),
    .A2(_08718_),
    .ZN(_08732_)
  );
  MUX2_X1 _16362_ (
    .A(wb_reg_cause[16]),
    .B(_08732_),
    .S(_06433_),
    .Z(_00192_)
  );
  AND2_X1 _16363_ (
    .A1(mem_reg_cause[17]),
    .A2(_08718_),
    .ZN(_08733_)
  );
  MUX2_X1 _16364_ (
    .A(wb_reg_cause[17]),
    .B(_08733_),
    .S(_06433_),
    .Z(_00193_)
  );
  AND2_X1 _16365_ (
    .A1(mem_reg_cause[18]),
    .A2(_08718_),
    .ZN(_08734_)
  );
  MUX2_X1 _16366_ (
    .A(wb_reg_cause[18]),
    .B(_08734_),
    .S(_06433_),
    .Z(_00194_)
  );
  AND2_X1 _16367_ (
    .A1(mem_reg_cause[19]),
    .A2(_08718_),
    .ZN(_08735_)
  );
  MUX2_X1 _16368_ (
    .A(wb_reg_cause[19]),
    .B(_08735_),
    .S(_06433_),
    .Z(_00195_)
  );
  AND2_X1 _16369_ (
    .A1(mem_reg_cause[20]),
    .A2(_08718_),
    .ZN(_08736_)
  );
  MUX2_X1 _16370_ (
    .A(wb_reg_cause[20]),
    .B(_08736_),
    .S(_06433_),
    .Z(_00196_)
  );
  AND2_X1 _16371_ (
    .A1(mem_reg_cause[21]),
    .A2(_08718_),
    .ZN(_08737_)
  );
  MUX2_X1 _16372_ (
    .A(wb_reg_cause[21]),
    .B(_08737_),
    .S(_06433_),
    .Z(_00197_)
  );
  AND2_X1 _16373_ (
    .A1(mem_reg_cause[22]),
    .A2(_08718_),
    .ZN(_08738_)
  );
  MUX2_X1 _16374_ (
    .A(wb_reg_cause[22]),
    .B(_08738_),
    .S(_06433_),
    .Z(_00198_)
  );
  AND2_X1 _16375_ (
    .A1(mem_reg_cause[23]),
    .A2(_08718_),
    .ZN(_08739_)
  );
  MUX2_X1 _16376_ (
    .A(wb_reg_cause[23]),
    .B(_08739_),
    .S(_06433_),
    .Z(_00199_)
  );
  AND2_X1 _16377_ (
    .A1(mem_reg_cause[24]),
    .A2(_08718_),
    .ZN(_08740_)
  );
  MUX2_X1 _16378_ (
    .A(wb_reg_cause[24]),
    .B(_08740_),
    .S(_06433_),
    .Z(_00200_)
  );
  AND2_X1 _16379_ (
    .A1(mem_reg_cause[25]),
    .A2(_08718_),
    .ZN(_08741_)
  );
  MUX2_X1 _16380_ (
    .A(wb_reg_cause[25]),
    .B(_08741_),
    .S(_06433_),
    .Z(_00201_)
  );
  AND2_X1 _16381_ (
    .A1(mem_reg_cause[26]),
    .A2(_08718_),
    .ZN(_08742_)
  );
  MUX2_X1 _16382_ (
    .A(wb_reg_cause[26]),
    .B(_08742_),
    .S(_06433_),
    .Z(_00202_)
  );
  AND2_X1 _16383_ (
    .A1(mem_reg_cause[27]),
    .A2(_08718_),
    .ZN(_08743_)
  );
  MUX2_X1 _16384_ (
    .A(wb_reg_cause[27]),
    .B(_08743_),
    .S(_06433_),
    .Z(_00203_)
  );
  AND2_X1 _16385_ (
    .A1(mem_reg_cause[28]),
    .A2(_08718_),
    .ZN(_08744_)
  );
  MUX2_X1 _16386_ (
    .A(wb_reg_cause[28]),
    .B(_08744_),
    .S(_06433_),
    .Z(_00204_)
  );
  AND2_X1 _16387_ (
    .A1(mem_reg_cause[29]),
    .A2(_08718_),
    .ZN(_08745_)
  );
  MUX2_X1 _16388_ (
    .A(wb_reg_cause[29]),
    .B(_08745_),
    .S(_06433_),
    .Z(_00205_)
  );
  AND2_X1 _16389_ (
    .A1(mem_reg_cause[30]),
    .A2(_08718_),
    .ZN(_08746_)
  );
  MUX2_X1 _16390_ (
    .A(wb_reg_cause[30]),
    .B(_08746_),
    .S(_06433_),
    .Z(_00206_)
  );
  AND2_X1 _16391_ (
    .A1(mem_reg_cause[31]),
    .A2(_08718_),
    .ZN(_08747_)
  );
  MUX2_X1 _16392_ (
    .A(wb_reg_cause[31]),
    .B(_08747_),
    .S(_06433_),
    .Z(_00207_)
  );
  MUX2_X1 _16393_ (
    .A(wb_reg_pc[0]),
    .B(mem_reg_pc[0]),
    .S(_06433_),
    .Z(_00208_)
  );
  MUX2_X1 _16394_ (
    .A(wb_reg_pc[1]),
    .B(mem_reg_pc[1]),
    .S(_06433_),
    .Z(_00209_)
  );
  MUX2_X1 _16395_ (
    .A(wb_reg_pc[2]),
    .B(mem_reg_pc[2]),
    .S(_06433_),
    .Z(_00210_)
  );
  MUX2_X1 _16396_ (
    .A(wb_reg_pc[3]),
    .B(mem_reg_pc[3]),
    .S(_06433_),
    .Z(_00211_)
  );
  MUX2_X1 _16397_ (
    .A(wb_reg_pc[4]),
    .B(mem_reg_pc[4]),
    .S(_06433_),
    .Z(_00212_)
  );
  MUX2_X1 _16398_ (
    .A(wb_reg_pc[5]),
    .B(mem_reg_pc[5]),
    .S(_06433_),
    .Z(_00213_)
  );
  MUX2_X1 _16399_ (
    .A(wb_reg_pc[6]),
    .B(mem_reg_pc[6]),
    .S(_06433_),
    .Z(_00214_)
  );
  MUX2_X1 _16400_ (
    .A(wb_reg_pc[7]),
    .B(mem_reg_pc[7]),
    .S(_06433_),
    .Z(_00215_)
  );
  MUX2_X1 _16401_ (
    .A(wb_reg_pc[8]),
    .B(mem_reg_pc[8]),
    .S(_06433_),
    .Z(_00216_)
  );
  MUX2_X1 _16402_ (
    .A(wb_reg_pc[9]),
    .B(mem_reg_pc[9]),
    .S(_06433_),
    .Z(_00217_)
  );
  MUX2_X1 _16403_ (
    .A(wb_reg_pc[10]),
    .B(mem_reg_pc[10]),
    .S(_06433_),
    .Z(_00218_)
  );
  MUX2_X1 _16404_ (
    .A(wb_reg_pc[11]),
    .B(mem_reg_pc[11]),
    .S(_06433_),
    .Z(_00219_)
  );
  MUX2_X1 _16405_ (
    .A(wb_reg_pc[12]),
    .B(mem_reg_pc[12]),
    .S(_06433_),
    .Z(_00220_)
  );
  MUX2_X1 _16406_ (
    .A(wb_reg_pc[13]),
    .B(mem_reg_pc[13]),
    .S(_06433_),
    .Z(_00221_)
  );
  MUX2_X1 _16407_ (
    .A(wb_reg_pc[14]),
    .B(mem_reg_pc[14]),
    .S(_06433_),
    .Z(_00222_)
  );
  MUX2_X1 _16408_ (
    .A(wb_reg_pc[15]),
    .B(mem_reg_pc[15]),
    .S(_06433_),
    .Z(_00223_)
  );
  MUX2_X1 _16409_ (
    .A(wb_reg_pc[16]),
    .B(mem_reg_pc[16]),
    .S(_06433_),
    .Z(_00224_)
  );
  MUX2_X1 _16410_ (
    .A(wb_reg_pc[17]),
    .B(mem_reg_pc[17]),
    .S(_06433_),
    .Z(_00225_)
  );
  MUX2_X1 _16411_ (
    .A(wb_reg_pc[18]),
    .B(mem_reg_pc[18]),
    .S(_06433_),
    .Z(_00226_)
  );
  MUX2_X1 _16412_ (
    .A(wb_reg_pc[19]),
    .B(mem_reg_pc[19]),
    .S(_06433_),
    .Z(_00227_)
  );
  MUX2_X1 _16413_ (
    .A(wb_reg_pc[20]),
    .B(mem_reg_pc[20]),
    .S(_06433_),
    .Z(_00228_)
  );
  MUX2_X1 _16414_ (
    .A(wb_reg_pc[21]),
    .B(mem_reg_pc[21]),
    .S(_06433_),
    .Z(_00229_)
  );
  MUX2_X1 _16415_ (
    .A(wb_reg_pc[22]),
    .B(mem_reg_pc[22]),
    .S(_06433_),
    .Z(_00230_)
  );
  MUX2_X1 _16416_ (
    .A(wb_reg_pc[23]),
    .B(mem_reg_pc[23]),
    .S(_06433_),
    .Z(_00231_)
  );
  MUX2_X1 _16417_ (
    .A(wb_reg_pc[24]),
    .B(mem_reg_pc[24]),
    .S(_06433_),
    .Z(_00232_)
  );
  MUX2_X1 _16418_ (
    .A(wb_reg_pc[25]),
    .B(mem_reg_pc[25]),
    .S(_06433_),
    .Z(_00233_)
  );
  MUX2_X1 _16419_ (
    .A(wb_reg_pc[26]),
    .B(mem_reg_pc[26]),
    .S(_06433_),
    .Z(_00234_)
  );
  MUX2_X1 _16420_ (
    .A(wb_reg_pc[27]),
    .B(mem_reg_pc[27]),
    .S(_06433_),
    .Z(_00235_)
  );
  MUX2_X1 _16421_ (
    .A(wb_reg_pc[28]),
    .B(mem_reg_pc[28]),
    .S(_06433_),
    .Z(_00236_)
  );
  MUX2_X1 _16422_ (
    .A(wb_reg_pc[29]),
    .B(mem_reg_pc[29]),
    .S(_06433_),
    .Z(_00237_)
  );
  MUX2_X1 _16423_ (
    .A(wb_reg_pc[30]),
    .B(mem_reg_pc[30]),
    .S(_06433_),
    .Z(_00238_)
  );
  MUX2_X1 _16424_ (
    .A(wb_reg_pc[31]),
    .B(mem_reg_pc[31]),
    .S(_06433_),
    .Z(_00239_)
  );
  OR2_X1 _16425_ (
    .A1(ex_reg_valid),
    .A2(ex_reg_replay),
    .ZN(_08748_)
  );
  OR2_X1 _16426_ (
    .A1(ex_reg_xcpt_interrupt),
    .A2(_08748_),
    .ZN(_08749_)
  );
  INV_X1 _16427_ (
    .A(_08749_),
    .ZN(_08750_)
  );
  AND2_X1 _16428_ (
    .A1(mem_reg_flush_pipe),
    .A2(mem_reg_valid),
    .ZN(_08751_)
  );
  OR2_X1 _16429_ (
    .A1(_08750_),
    .A2(_08751_),
    .ZN(_08752_)
  );
  INV_X1 _16430_ (
    .A(_08752_),
    .ZN(_08753_)
  );
  MUX2_X1 _16431_ (
    .A(alu_io_cmp_out),
    .B(mem_br_taken),
    .S(_08752_),
    .Z(_00240_)
  );
  OR2_X1 _16432_ (
    .A1(_00017_),
    .A2(_00035_),
    .ZN(_08754_)
  );
  AND2_X1 _16433_ (
    .A1(_03035_),
    .A2(_03062_),
    .ZN(_08755_)
  );
  INV_X1 _16434_ (
    .A(_08755_),
    .ZN(_08756_)
  );
  OR2_X1 _16435_ (
    .A1(ex_reg_rs_lsb_1[1]),
    .A2(_00017_),
    .ZN(_08757_)
  );
  INV_X1 _16436_ (
    .A(_08757_),
    .ZN(_08758_)
  );
  AND2_X1 _16437_ (
    .A1(_08756_),
    .A2(_08758_),
    .ZN(_08759_)
  );
  AND2_X1 _16438_ (
    .A1(mem_reg_wdata[0]),
    .A2(_08759_),
    .ZN(_08760_)
  );
  AND2_X1 _16439_ (
    .A1(wb_reg_wdata[0]),
    .A2(_08755_),
    .ZN(_08761_)
  );
  OR2_X1 _16440_ (
    .A1(_08760_),
    .A2(_08761_),
    .ZN(_08762_)
  );
  MUX2_X1 _16441_ (
    .A(io_dmem_resp_bits_data_word_bypass[0]),
    .B(_08762_),
    .S(_08754_),
    .Z(_08763_)
  );
  MUX2_X1 _16442_ (
    .A(ex_reg_rs_lsb_1[0]),
    .B(_08763_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[0])
  );
  AND2_X1 _16443_ (
    .A1(ex_ctrl_mem),
    .A2(_08753_),
    .ZN(_08764_)
  );
  INV_X1 _16444_ (
    .A(_08764_),
    .ZN(_08765_)
  );
  AND2_X1 _16445_ (
    .A1(ex_ctrl_rxs2),
    .A2(_08764_),
    .ZN(_08766_)
  );
  OR2_X1 _16446_ (
    .A1(_03034_),
    .A2(_08765_),
    .ZN(_08767_)
  );
  OR2_X1 _16447_ (
    .A1(_ex_op2_T[0]),
    .A2(_08767_),
    .ZN(_08768_)
  );
  MUX2_X1 _16448_ (
    .A(mem_reg_rs2[0]),
    .B(_ex_op2_T[0]),
    .S(_08766_),
    .Z(_00241_)
  );
  AND2_X1 _16449_ (
    .A1(mem_reg_wdata[1]),
    .A2(_08759_),
    .ZN(_08769_)
  );
  AND2_X1 _16450_ (
    .A1(wb_reg_wdata[1]),
    .A2(_08755_),
    .ZN(_08770_)
  );
  OR2_X1 _16451_ (
    .A1(_08769_),
    .A2(_08770_),
    .ZN(_08771_)
  );
  MUX2_X1 _16452_ (
    .A(io_dmem_resp_bits_data_word_bypass[1]),
    .B(_08771_),
    .S(_08754_),
    .Z(_08772_)
  );
  MUX2_X1 _16453_ (
    .A(ex_reg_rs_lsb_1[1]),
    .B(_08772_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[1])
  );
  OR2_X1 _16454_ (
    .A1(_08767_),
    .A2(_ex_op2_T[1]),
    .ZN(_08773_)
  );
  MUX2_X1 _16455_ (
    .A(mem_reg_rs2[1]),
    .B(_ex_op2_T[1]),
    .S(_08766_),
    .Z(_00242_)
  );
  AND2_X1 _16456_ (
    .A1(mem_reg_wdata[2]),
    .A2(_08759_),
    .ZN(_08774_)
  );
  AND2_X1 _16457_ (
    .A1(wb_reg_wdata[2]),
    .A2(_08755_),
    .ZN(_08775_)
  );
  OR2_X1 _16458_ (
    .A1(_08774_),
    .A2(_08775_),
    .ZN(_08776_)
  );
  MUX2_X1 _16459_ (
    .A(io_dmem_resp_bits_data_word_bypass[2]),
    .B(_08776_),
    .S(_08754_),
    .Z(_08777_)
  );
  MUX2_X1 _16460_ (
    .A(ex_reg_rs_msb_1[0]),
    .B(_08777_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[2])
  );
  OR2_X1 _16461_ (
    .A1(_08767_),
    .A2(_ex_op2_T[2]),
    .ZN(_08778_)
  );
  MUX2_X1 _16462_ (
    .A(mem_reg_rs2[2]),
    .B(_ex_op2_T[2]),
    .S(_08766_),
    .Z(_00243_)
  );
  AND2_X1 _16463_ (
    .A1(mem_reg_wdata[3]),
    .A2(_08759_),
    .ZN(_08779_)
  );
  AND2_X1 _16464_ (
    .A1(wb_reg_wdata[3]),
    .A2(_08755_),
    .ZN(_08780_)
  );
  OR2_X1 _16465_ (
    .A1(_08779_),
    .A2(_08780_),
    .ZN(_08781_)
  );
  MUX2_X1 _16466_ (
    .A(io_dmem_resp_bits_data_word_bypass[3]),
    .B(_08781_),
    .S(_08754_),
    .Z(_08782_)
  );
  MUX2_X1 _16467_ (
    .A(ex_reg_rs_msb_1[1]),
    .B(_08782_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[3])
  );
  OR2_X1 _16468_ (
    .A1(_08767_),
    .A2(_ex_op2_T[3]),
    .ZN(_08783_)
  );
  MUX2_X1 _16469_ (
    .A(mem_reg_rs2[3]),
    .B(_ex_op2_T[3]),
    .S(_08766_),
    .Z(_00244_)
  );
  AND2_X1 _16470_ (
    .A1(mem_reg_wdata[4]),
    .A2(_08759_),
    .ZN(_08784_)
  );
  AND2_X1 _16471_ (
    .A1(wb_reg_wdata[4]),
    .A2(_08755_),
    .ZN(_08785_)
  );
  OR2_X1 _16472_ (
    .A1(_08784_),
    .A2(_08785_),
    .ZN(_08786_)
  );
  MUX2_X1 _16473_ (
    .A(io_dmem_resp_bits_data_word_bypass[4]),
    .B(_08786_),
    .S(_08754_),
    .Z(_08787_)
  );
  MUX2_X1 _16474_ (
    .A(ex_reg_rs_msb_1[2]),
    .B(_08787_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[4])
  );
  OR2_X1 _16475_ (
    .A1(_08767_),
    .A2(_ex_op2_T[4]),
    .ZN(_08788_)
  );
  MUX2_X1 _16476_ (
    .A(mem_reg_rs2[4]),
    .B(_ex_op2_T[4]),
    .S(_08766_),
    .Z(_00245_)
  );
  AND2_X1 _16477_ (
    .A1(mem_reg_wdata[5]),
    .A2(_08759_),
    .ZN(_08789_)
  );
  AND2_X1 _16478_ (
    .A1(wb_reg_wdata[5]),
    .A2(_08755_),
    .ZN(_08790_)
  );
  OR2_X1 _16479_ (
    .A1(_08789_),
    .A2(_08790_),
    .ZN(_08791_)
  );
  MUX2_X1 _16480_ (
    .A(io_dmem_resp_bits_data_word_bypass[5]),
    .B(_08791_),
    .S(_08754_),
    .Z(_08792_)
  );
  MUX2_X1 _16481_ (
    .A(ex_reg_rs_msb_1[3]),
    .B(_08792_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[5])
  );
  OR2_X1 _16482_ (
    .A1(_08767_),
    .A2(_ex_op2_T[5]),
    .ZN(_08793_)
  );
  MUX2_X1 _16483_ (
    .A(mem_reg_rs2[5]),
    .B(_ex_op2_T[5]),
    .S(_08766_),
    .Z(_00246_)
  );
  AND2_X1 _16484_ (
    .A1(mem_reg_wdata[6]),
    .A2(_08759_),
    .ZN(_08794_)
  );
  AND2_X1 _16485_ (
    .A1(wb_reg_wdata[6]),
    .A2(_08755_),
    .ZN(_08795_)
  );
  OR2_X1 _16486_ (
    .A1(_08794_),
    .A2(_08795_),
    .ZN(_08796_)
  );
  MUX2_X1 _16487_ (
    .A(io_dmem_resp_bits_data_word_bypass[6]),
    .B(_08796_),
    .S(_08754_),
    .Z(_08797_)
  );
  MUX2_X1 _16488_ (
    .A(ex_reg_rs_msb_1[4]),
    .B(_08797_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[6])
  );
  MUX2_X1 _16489_ (
    .A(mem_reg_rs2[6]),
    .B(_ex_op2_T[6]),
    .S(_08766_),
    .Z(_00247_)
  );
  AND2_X1 _16490_ (
    .A1(mem_reg_wdata[7]),
    .A2(_08759_),
    .ZN(_08798_)
  );
  AND2_X1 _16491_ (
    .A1(wb_reg_wdata[7]),
    .A2(_08755_),
    .ZN(_08799_)
  );
  OR2_X1 _16492_ (
    .A1(_08798_),
    .A2(_08799_),
    .ZN(_08800_)
  );
  MUX2_X1 _16493_ (
    .A(io_dmem_resp_bits_data_word_bypass[7]),
    .B(_08800_),
    .S(_08754_),
    .Z(_08801_)
  );
  MUX2_X1 _16494_ (
    .A(ex_reg_rs_msb_1[5]),
    .B(_08801_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[7])
  );
  MUX2_X1 _16495_ (
    .A(mem_reg_rs2[7]),
    .B(_ex_op2_T[7]),
    .S(_08766_),
    .Z(_00248_)
  );
  OR2_X1 _16496_ (
    .A1(ex_reg_mem_size[0]),
    .A2(ex_reg_mem_size[1]),
    .ZN(_08802_)
  );
  INV_X1 _16497_ (
    .A(_08802_),
    .ZN(_08803_)
  );
  AND2_X1 _16498_ (
    .A1(mem_reg_wdata[8]),
    .A2(_08759_),
    .ZN(_08804_)
  );
  AND2_X1 _16499_ (
    .A1(wb_reg_wdata[8]),
    .A2(_08755_),
    .ZN(_08805_)
  );
  OR2_X1 _16500_ (
    .A1(_08804_),
    .A2(_08805_),
    .ZN(_08806_)
  );
  MUX2_X1 _16501_ (
    .A(io_dmem_resp_bits_data_word_bypass[8]),
    .B(_08806_),
    .S(_08754_),
    .Z(_08807_)
  );
  MUX2_X1 _16502_ (
    .A(ex_reg_rs_msb_1[6]),
    .B(_08807_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[8])
  );
  AND2_X1 _16503_ (
    .A1(_08802_),
    .A2(_ex_op2_T[8]),
    .ZN(_08808_)
  );
  OR2_X1 _16504_ (
    .A1(_08767_),
    .A2(_08803_),
    .ZN(_08809_)
  );
  AND2_X1 _16505_ (
    .A1(_08768_),
    .A2(_08809_),
    .ZN(_08810_)
  );
  OR2_X1 _16506_ (
    .A1(_08808_),
    .A2(_08810_),
    .ZN(_08811_)
  );
  OR2_X1 _16507_ (
    .A1(mem_reg_rs2[8]),
    .A2(_08766_),
    .ZN(_08812_)
  );
  AND2_X1 _16508_ (
    .A1(_08811_),
    .A2(_08812_),
    .ZN(_00249_)
  );
  AND2_X1 _16509_ (
    .A1(mem_reg_wdata[9]),
    .A2(_08759_),
    .ZN(_08813_)
  );
  AND2_X1 _16510_ (
    .A1(wb_reg_wdata[9]),
    .A2(_08755_),
    .ZN(_08814_)
  );
  OR2_X1 _16511_ (
    .A1(_08813_),
    .A2(_08814_),
    .ZN(_08815_)
  );
  MUX2_X1 _16512_ (
    .A(io_dmem_resp_bits_data_word_bypass[9]),
    .B(_08815_),
    .S(_08754_),
    .Z(_08816_)
  );
  MUX2_X1 _16513_ (
    .A(ex_reg_rs_msb_1[7]),
    .B(_08816_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[9])
  );
  AND2_X1 _16514_ (
    .A1(_08802_),
    .A2(_ex_op2_T[9]),
    .ZN(_08817_)
  );
  AND2_X1 _16515_ (
    .A1(_08773_),
    .A2(_08809_),
    .ZN(_08818_)
  );
  OR2_X1 _16516_ (
    .A1(_08817_),
    .A2(_08818_),
    .ZN(_08819_)
  );
  OR2_X1 _16517_ (
    .A1(mem_reg_rs2[9]),
    .A2(_08766_),
    .ZN(_08820_)
  );
  AND2_X1 _16518_ (
    .A1(_08819_),
    .A2(_08820_),
    .ZN(_00250_)
  );
  AND2_X1 _16519_ (
    .A1(mem_reg_wdata[10]),
    .A2(_08759_),
    .ZN(_08821_)
  );
  AND2_X1 _16520_ (
    .A1(wb_reg_wdata[10]),
    .A2(_08755_),
    .ZN(_08822_)
  );
  OR2_X1 _16521_ (
    .A1(_08821_),
    .A2(_08822_),
    .ZN(_08823_)
  );
  MUX2_X1 _16522_ (
    .A(io_dmem_resp_bits_data_word_bypass[10]),
    .B(_08823_),
    .S(_08754_),
    .Z(_08824_)
  );
  MUX2_X1 _16523_ (
    .A(ex_reg_rs_msb_1[8]),
    .B(_08824_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[10])
  );
  AND2_X1 _16524_ (
    .A1(_08802_),
    .A2(_ex_op2_T[10]),
    .ZN(_08825_)
  );
  AND2_X1 _16525_ (
    .A1(_08778_),
    .A2(_08809_),
    .ZN(_08826_)
  );
  OR2_X1 _16526_ (
    .A1(_08825_),
    .A2(_08826_),
    .ZN(_08827_)
  );
  OR2_X1 _16527_ (
    .A1(mem_reg_rs2[10]),
    .A2(_08766_),
    .ZN(_08828_)
  );
  AND2_X1 _16528_ (
    .A1(_08827_),
    .A2(_08828_),
    .ZN(_00251_)
  );
  AND2_X1 _16529_ (
    .A1(mem_reg_wdata[11]),
    .A2(_08759_),
    .ZN(_08829_)
  );
  AND2_X1 _16530_ (
    .A1(wb_reg_wdata[11]),
    .A2(_08755_),
    .ZN(_08830_)
  );
  OR2_X1 _16531_ (
    .A1(_08829_),
    .A2(_08830_),
    .ZN(_08831_)
  );
  MUX2_X1 _16532_ (
    .A(io_dmem_resp_bits_data_word_bypass[11]),
    .B(_08831_),
    .S(_08754_),
    .Z(_08832_)
  );
  MUX2_X1 _16533_ (
    .A(ex_reg_rs_msb_1[9]),
    .B(_08832_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[11])
  );
  AND2_X1 _16534_ (
    .A1(_08802_),
    .A2(_ex_op2_T[11]),
    .ZN(_08833_)
  );
  AND2_X1 _16535_ (
    .A1(_08783_),
    .A2(_08809_),
    .ZN(_08834_)
  );
  OR2_X1 _16536_ (
    .A1(_08833_),
    .A2(_08834_),
    .ZN(_08835_)
  );
  OR2_X1 _16537_ (
    .A1(mem_reg_rs2[11]),
    .A2(_08766_),
    .ZN(_08836_)
  );
  AND2_X1 _16538_ (
    .A1(_08835_),
    .A2(_08836_),
    .ZN(_00252_)
  );
  AND2_X1 _16539_ (
    .A1(mem_reg_wdata[12]),
    .A2(_08759_),
    .ZN(_08837_)
  );
  AND2_X1 _16540_ (
    .A1(wb_reg_wdata[12]),
    .A2(_08755_),
    .ZN(_08838_)
  );
  OR2_X1 _16541_ (
    .A1(_08837_),
    .A2(_08838_),
    .ZN(_08839_)
  );
  MUX2_X1 _16542_ (
    .A(io_dmem_resp_bits_data_word_bypass[12]),
    .B(_08839_),
    .S(_08754_),
    .Z(_08840_)
  );
  MUX2_X1 _16543_ (
    .A(ex_reg_rs_msb_1[10]),
    .B(_08840_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[12])
  );
  AND2_X1 _16544_ (
    .A1(_08802_),
    .A2(_ex_op2_T[12]),
    .ZN(_08841_)
  );
  AND2_X1 _16545_ (
    .A1(_08788_),
    .A2(_08809_),
    .ZN(_08842_)
  );
  OR2_X1 _16546_ (
    .A1(_08841_),
    .A2(_08842_),
    .ZN(_08843_)
  );
  OR2_X1 _16547_ (
    .A1(mem_reg_rs2[12]),
    .A2(_08766_),
    .ZN(_08844_)
  );
  AND2_X1 _16548_ (
    .A1(_08843_),
    .A2(_08844_),
    .ZN(_00253_)
  );
  AND2_X1 _16549_ (
    .A1(mem_reg_wdata[13]),
    .A2(_08759_),
    .ZN(_08845_)
  );
  AND2_X1 _16550_ (
    .A1(wb_reg_wdata[13]),
    .A2(_08755_),
    .ZN(_08846_)
  );
  OR2_X1 _16551_ (
    .A1(_08845_),
    .A2(_08846_),
    .ZN(_08847_)
  );
  MUX2_X1 _16552_ (
    .A(io_dmem_resp_bits_data_word_bypass[13]),
    .B(_08847_),
    .S(_08754_),
    .Z(_08848_)
  );
  MUX2_X1 _16553_ (
    .A(ex_reg_rs_msb_1[11]),
    .B(_08848_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[13])
  );
  AND2_X1 _16554_ (
    .A1(_08802_),
    .A2(_ex_op2_T[13]),
    .ZN(_08849_)
  );
  AND2_X1 _16555_ (
    .A1(_08793_),
    .A2(_08809_),
    .ZN(_08850_)
  );
  OR2_X1 _16556_ (
    .A1(_08849_),
    .A2(_08850_),
    .ZN(_08851_)
  );
  OR2_X1 _16557_ (
    .A1(mem_reg_rs2[13]),
    .A2(_08766_),
    .ZN(_08852_)
  );
  AND2_X1 _16558_ (
    .A1(_08851_),
    .A2(_08852_),
    .ZN(_00254_)
  );
  AND2_X1 _16559_ (
    .A1(mem_reg_wdata[14]),
    .A2(_08759_),
    .ZN(_08853_)
  );
  AND2_X1 _16560_ (
    .A1(wb_reg_wdata[14]),
    .A2(_08755_),
    .ZN(_08854_)
  );
  OR2_X1 _16561_ (
    .A1(_08853_),
    .A2(_08854_),
    .ZN(_08855_)
  );
  MUX2_X1 _16562_ (
    .A(io_dmem_resp_bits_data_word_bypass[14]),
    .B(_08855_),
    .S(_08754_),
    .Z(_08856_)
  );
  MUX2_X1 _16563_ (
    .A(ex_reg_rs_msb_1[12]),
    .B(_08856_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[14])
  );
  AND2_X1 _16564_ (
    .A1(_08802_),
    .A2(_ex_op2_T[14]),
    .ZN(_08857_)
  );
  AND2_X1 _16565_ (
    .A1(_ex_op2_T[6]),
    .A2(_08803_),
    .ZN(_08858_)
  );
  OR2_X1 _16566_ (
    .A1(_08857_),
    .A2(_08858_),
    .ZN(_08859_)
  );
  MUX2_X1 _16567_ (
    .A(mem_reg_rs2[14]),
    .B(_08859_),
    .S(_08766_),
    .Z(_00255_)
  );
  AND2_X1 _16568_ (
    .A1(mem_reg_wdata[15]),
    .A2(_08759_),
    .ZN(_08860_)
  );
  AND2_X1 _16569_ (
    .A1(wb_reg_wdata[15]),
    .A2(_08755_),
    .ZN(_08861_)
  );
  OR2_X1 _16570_ (
    .A1(_08860_),
    .A2(_08861_),
    .ZN(_08862_)
  );
  MUX2_X1 _16571_ (
    .A(io_dmem_resp_bits_data_word_bypass[15]),
    .B(_08862_),
    .S(_08754_),
    .Z(_08863_)
  );
  MUX2_X1 _16572_ (
    .A(ex_reg_rs_msb_1[13]),
    .B(_08863_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[15])
  );
  AND2_X1 _16573_ (
    .A1(_08802_),
    .A2(_ex_op2_T[15]),
    .ZN(_08864_)
  );
  AND2_X1 _16574_ (
    .A1(_ex_op2_T[7]),
    .A2(_08803_),
    .ZN(_08865_)
  );
  OR2_X1 _16575_ (
    .A1(_08864_),
    .A2(_08865_),
    .ZN(_08866_)
  );
  MUX2_X1 _16576_ (
    .A(mem_reg_rs2[15]),
    .B(_08866_),
    .S(_08766_),
    .Z(_00256_)
  );
  AND2_X1 _16577_ (
    .A1(_03010_),
    .A2(_03058_),
    .ZN(_08867_)
  );
  INV_X1 _16578_ (
    .A(_08867_),
    .ZN(_08868_)
  );
  AND2_X1 _16579_ (
    .A1(_08802_),
    .A2(_08868_),
    .ZN(_08869_)
  );
  AND2_X1 _16580_ (
    .A1(mem_reg_wdata[16]),
    .A2(_08759_),
    .ZN(_08870_)
  );
  AND2_X1 _16581_ (
    .A1(wb_reg_wdata[16]),
    .A2(_08755_),
    .ZN(_08871_)
  );
  OR2_X1 _16582_ (
    .A1(_08870_),
    .A2(_08871_),
    .ZN(_08872_)
  );
  MUX2_X1 _16583_ (
    .A(io_dmem_resp_bits_data_word_bypass[16]),
    .B(_08872_),
    .S(_08754_),
    .Z(_08873_)
  );
  MUX2_X1 _16584_ (
    .A(ex_reg_rs_msb_1[14]),
    .B(_08873_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[16])
  );
  MUX2_X1 _16585_ (
    .A(_ex_op2_T[0]),
    .B(_ex_op2_T[16]),
    .S(_08869_),
    .Z(_08874_)
  );
  MUX2_X1 _16586_ (
    .A(mem_reg_rs2[16]),
    .B(_08874_),
    .S(_08766_),
    .Z(_00257_)
  );
  AND2_X1 _16587_ (
    .A1(mem_reg_wdata[17]),
    .A2(_08759_),
    .ZN(_08875_)
  );
  AND2_X1 _16588_ (
    .A1(wb_reg_wdata[17]),
    .A2(_08755_),
    .ZN(_08876_)
  );
  OR2_X1 _16589_ (
    .A1(_08875_),
    .A2(_08876_),
    .ZN(_08877_)
  );
  MUX2_X1 _16590_ (
    .A(io_dmem_resp_bits_data_word_bypass[17]),
    .B(_08877_),
    .S(_08754_),
    .Z(_08878_)
  );
  MUX2_X1 _16591_ (
    .A(ex_reg_rs_msb_1[15]),
    .B(_08878_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[17])
  );
  MUX2_X1 _16592_ (
    .A(_ex_op2_T[1]),
    .B(_ex_op2_T[17]),
    .S(_08869_),
    .Z(_08879_)
  );
  MUX2_X1 _16593_ (
    .A(mem_reg_rs2[17]),
    .B(_08879_),
    .S(_08766_),
    .Z(_00258_)
  );
  AND2_X1 _16594_ (
    .A1(mem_reg_wdata[18]),
    .A2(_08759_),
    .ZN(_08880_)
  );
  AND2_X1 _16595_ (
    .A1(wb_reg_wdata[18]),
    .A2(_08755_),
    .ZN(_08881_)
  );
  OR2_X1 _16596_ (
    .A1(_08880_),
    .A2(_08881_),
    .ZN(_08882_)
  );
  MUX2_X1 _16597_ (
    .A(io_dmem_resp_bits_data_word_bypass[18]),
    .B(_08882_),
    .S(_08754_),
    .Z(_08883_)
  );
  MUX2_X1 _16598_ (
    .A(ex_reg_rs_msb_1[16]),
    .B(_08883_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[18])
  );
  MUX2_X1 _16599_ (
    .A(_ex_op2_T[2]),
    .B(_ex_op2_T[18]),
    .S(_08869_),
    .Z(_08884_)
  );
  MUX2_X1 _16600_ (
    .A(mem_reg_rs2[18]),
    .B(_08884_),
    .S(_08766_),
    .Z(_00259_)
  );
  AND2_X1 _16601_ (
    .A1(mem_reg_wdata[19]),
    .A2(_08759_),
    .ZN(_08885_)
  );
  AND2_X1 _16602_ (
    .A1(wb_reg_wdata[19]),
    .A2(_08755_),
    .ZN(_08886_)
  );
  OR2_X1 _16603_ (
    .A1(_08885_),
    .A2(_08886_),
    .ZN(_08887_)
  );
  MUX2_X1 _16604_ (
    .A(io_dmem_resp_bits_data_word_bypass[19]),
    .B(_08887_),
    .S(_08754_),
    .Z(_08888_)
  );
  MUX2_X1 _16605_ (
    .A(ex_reg_rs_msb_1[17]),
    .B(_08888_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[19])
  );
  MUX2_X1 _16606_ (
    .A(_ex_op2_T[3]),
    .B(_ex_op2_T[19]),
    .S(_08869_),
    .Z(_08889_)
  );
  MUX2_X1 _16607_ (
    .A(mem_reg_rs2[19]),
    .B(_08889_),
    .S(_08766_),
    .Z(_00260_)
  );
  AND2_X1 _16608_ (
    .A1(mem_reg_wdata[20]),
    .A2(_08759_),
    .ZN(_08890_)
  );
  AND2_X1 _16609_ (
    .A1(wb_reg_wdata[20]),
    .A2(_08755_),
    .ZN(_08891_)
  );
  OR2_X1 _16610_ (
    .A1(_08890_),
    .A2(_08891_),
    .ZN(_08892_)
  );
  MUX2_X1 _16611_ (
    .A(io_dmem_resp_bits_data_word_bypass[20]),
    .B(_08892_),
    .S(_08754_),
    .Z(_08893_)
  );
  MUX2_X1 _16612_ (
    .A(ex_reg_rs_msb_1[18]),
    .B(_08893_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[20])
  );
  MUX2_X1 _16613_ (
    .A(_ex_op2_T[4]),
    .B(_ex_op2_T[20]),
    .S(_08869_),
    .Z(_08894_)
  );
  MUX2_X1 _16614_ (
    .A(mem_reg_rs2[20]),
    .B(_08894_),
    .S(_08766_),
    .Z(_00261_)
  );
  AND2_X1 _16615_ (
    .A1(mem_reg_wdata[21]),
    .A2(_08759_),
    .ZN(_08895_)
  );
  AND2_X1 _16616_ (
    .A1(wb_reg_wdata[21]),
    .A2(_08755_),
    .ZN(_08896_)
  );
  OR2_X1 _16617_ (
    .A1(_08895_),
    .A2(_08896_),
    .ZN(_08897_)
  );
  MUX2_X1 _16618_ (
    .A(io_dmem_resp_bits_data_word_bypass[21]),
    .B(_08897_),
    .S(_08754_),
    .Z(_08898_)
  );
  MUX2_X1 _16619_ (
    .A(ex_reg_rs_msb_1[19]),
    .B(_08898_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[21])
  );
  MUX2_X1 _16620_ (
    .A(_ex_op2_T[5]),
    .B(_ex_op2_T[21]),
    .S(_08869_),
    .Z(_08899_)
  );
  MUX2_X1 _16621_ (
    .A(mem_reg_rs2[21]),
    .B(_08899_),
    .S(_08766_),
    .Z(_00262_)
  );
  AND2_X1 _16622_ (
    .A1(mem_reg_wdata[22]),
    .A2(_08759_),
    .ZN(_08900_)
  );
  AND2_X1 _16623_ (
    .A1(wb_reg_wdata[22]),
    .A2(_08755_),
    .ZN(_08901_)
  );
  OR2_X1 _16624_ (
    .A1(_08900_),
    .A2(_08901_),
    .ZN(_08902_)
  );
  MUX2_X1 _16625_ (
    .A(io_dmem_resp_bits_data_word_bypass[22]),
    .B(_08902_),
    .S(_08754_),
    .Z(_08903_)
  );
  MUX2_X1 _16626_ (
    .A(ex_reg_rs_msb_1[20]),
    .B(_08903_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[22])
  );
  MUX2_X1 _16627_ (
    .A(_ex_op2_T[6]),
    .B(_ex_op2_T[22]),
    .S(_08869_),
    .Z(_08904_)
  );
  MUX2_X1 _16628_ (
    .A(mem_reg_rs2[22]),
    .B(_08904_),
    .S(_08766_),
    .Z(_00263_)
  );
  AND2_X1 _16629_ (
    .A1(mem_reg_wdata[23]),
    .A2(_08759_),
    .ZN(_01588_)
  );
  AND2_X1 _16630_ (
    .A1(wb_reg_wdata[23]),
    .A2(_08755_),
    .ZN(_01589_)
  );
  OR2_X1 _16631_ (
    .A1(_01588_),
    .A2(_01589_),
    .ZN(_01590_)
  );
  MUX2_X1 _16632_ (
    .A(io_dmem_resp_bits_data_word_bypass[23]),
    .B(_01590_),
    .S(_08754_),
    .Z(_01591_)
  );
  MUX2_X1 _16633_ (
    .A(ex_reg_rs_msb_1[21]),
    .B(_01591_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[23])
  );
  MUX2_X1 _16634_ (
    .A(_ex_op2_T[7]),
    .B(_ex_op2_T[23]),
    .S(_08869_),
    .Z(_01592_)
  );
  MUX2_X1 _16635_ (
    .A(mem_reg_rs2[23]),
    .B(_01592_),
    .S(_08766_),
    .Z(_00264_)
  );
  OR2_X1 _16636_ (
    .A1(_08811_),
    .A2(_08869_),
    .ZN(_01593_)
  );
  AND2_X1 _16637_ (
    .A1(mem_reg_wdata[24]),
    .A2(_08759_),
    .ZN(_01594_)
  );
  AND2_X1 _16638_ (
    .A1(wb_reg_wdata[24]),
    .A2(_08755_),
    .ZN(_01595_)
  );
  OR2_X1 _16639_ (
    .A1(_01594_),
    .A2(_01595_),
    .ZN(_01596_)
  );
  MUX2_X1 _16640_ (
    .A(io_dmem_resp_bits_data_word_bypass[24]),
    .B(_01596_),
    .S(_08754_),
    .Z(_01597_)
  );
  MUX2_X1 _16641_ (
    .A(ex_reg_rs_msb_1[22]),
    .B(_01597_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[24])
  );
  OR2_X1 _16642_ (
    .A1(_08867_),
    .A2(_ex_op2_T[24]),
    .ZN(_01598_)
  );
  OR2_X1 _16643_ (
    .A1(_08810_),
    .A2(_01598_),
    .ZN(_01599_)
  );
  OR2_X1 _16644_ (
    .A1(mem_reg_rs2[24]),
    .A2(_08766_),
    .ZN(_01600_)
  );
  AND2_X1 _16645_ (
    .A1(_01599_),
    .A2(_01600_),
    .ZN(_01601_)
  );
  AND2_X1 _16646_ (
    .A1(_01593_),
    .A2(_01601_),
    .ZN(_00265_)
  );
  OR2_X1 _16647_ (
    .A1(_08819_),
    .A2(_08869_),
    .ZN(_01602_)
  );
  OR2_X1 _16648_ (
    .A1(mem_reg_rs2[25]),
    .A2(_08766_),
    .ZN(_01603_)
  );
  AND2_X1 _16649_ (
    .A1(mem_reg_wdata[25]),
    .A2(_08759_),
    .ZN(_01604_)
  );
  AND2_X1 _16650_ (
    .A1(wb_reg_wdata[25]),
    .A2(_08755_),
    .ZN(_01605_)
  );
  OR2_X1 _16651_ (
    .A1(_01604_),
    .A2(_01605_),
    .ZN(_01606_)
  );
  MUX2_X1 _16652_ (
    .A(io_dmem_resp_bits_data_word_bypass[25]),
    .B(_01606_),
    .S(_08754_),
    .Z(_01607_)
  );
  MUX2_X1 _16653_ (
    .A(ex_reg_rs_msb_1[23]),
    .B(_01607_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[25])
  );
  OR2_X1 _16654_ (
    .A1(_08867_),
    .A2(_ex_op2_T[25]),
    .ZN(_01608_)
  );
  OR2_X1 _16655_ (
    .A1(_08818_),
    .A2(_01608_),
    .ZN(_01609_)
  );
  AND2_X1 _16656_ (
    .A1(_01603_),
    .A2(_01609_),
    .ZN(_01610_)
  );
  AND2_X1 _16657_ (
    .A1(_01602_),
    .A2(_01610_),
    .ZN(_00266_)
  );
  OR2_X1 _16658_ (
    .A1(_08827_),
    .A2(_08869_),
    .ZN(_01611_)
  );
  AND2_X1 _16659_ (
    .A1(mem_reg_wdata[26]),
    .A2(_08759_),
    .ZN(_01612_)
  );
  AND2_X1 _16660_ (
    .A1(wb_reg_wdata[26]),
    .A2(_08755_),
    .ZN(_01613_)
  );
  OR2_X1 _16661_ (
    .A1(_01612_),
    .A2(_01613_),
    .ZN(_01614_)
  );
  MUX2_X1 _16662_ (
    .A(io_dmem_resp_bits_data_word_bypass[26]),
    .B(_01614_),
    .S(_08754_),
    .Z(_01615_)
  );
  MUX2_X1 _16663_ (
    .A(ex_reg_rs_msb_1[24]),
    .B(_01615_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[26])
  );
  OR2_X1 _16664_ (
    .A1(_08867_),
    .A2(_ex_op2_T[26]),
    .ZN(_01616_)
  );
  OR2_X1 _16665_ (
    .A1(_08826_),
    .A2(_01616_),
    .ZN(_01617_)
  );
  OR2_X1 _16666_ (
    .A1(mem_reg_rs2[26]),
    .A2(_08766_),
    .ZN(_01618_)
  );
  AND2_X1 _16667_ (
    .A1(_01617_),
    .A2(_01618_),
    .ZN(_01619_)
  );
  AND2_X1 _16668_ (
    .A1(_01611_),
    .A2(_01619_),
    .ZN(_00267_)
  );
  OR2_X1 _16669_ (
    .A1(_08835_),
    .A2(_08869_),
    .ZN(_01620_)
  );
  AND2_X1 _16670_ (
    .A1(mem_reg_wdata[27]),
    .A2(_08759_),
    .ZN(_01621_)
  );
  AND2_X1 _16671_ (
    .A1(wb_reg_wdata[27]),
    .A2(_08755_),
    .ZN(_01622_)
  );
  OR2_X1 _16672_ (
    .A1(_01621_),
    .A2(_01622_),
    .ZN(_01623_)
  );
  MUX2_X1 _16673_ (
    .A(io_dmem_resp_bits_data_word_bypass[27]),
    .B(_01623_),
    .S(_08754_),
    .Z(_01624_)
  );
  MUX2_X1 _16674_ (
    .A(ex_reg_rs_msb_1[25]),
    .B(_01624_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[27])
  );
  OR2_X1 _16675_ (
    .A1(_08867_),
    .A2(_ex_op2_T[27]),
    .ZN(_01625_)
  );
  OR2_X1 _16676_ (
    .A1(_08834_),
    .A2(_01625_),
    .ZN(_01626_)
  );
  OR2_X1 _16677_ (
    .A1(mem_reg_rs2[27]),
    .A2(_08766_),
    .ZN(_01627_)
  );
  AND2_X1 _16678_ (
    .A1(_01626_),
    .A2(_01627_),
    .ZN(_01628_)
  );
  AND2_X1 _16679_ (
    .A1(_01620_),
    .A2(_01628_),
    .ZN(_00268_)
  );
  OR2_X1 _16680_ (
    .A1(_08843_),
    .A2(_08869_),
    .ZN(_01629_)
  );
  AND2_X1 _16681_ (
    .A1(mem_reg_wdata[28]),
    .A2(_08759_),
    .ZN(_01630_)
  );
  AND2_X1 _16682_ (
    .A1(wb_reg_wdata[28]),
    .A2(_08755_),
    .ZN(_01631_)
  );
  OR2_X1 _16683_ (
    .A1(_01630_),
    .A2(_01631_),
    .ZN(_01632_)
  );
  MUX2_X1 _16684_ (
    .A(io_dmem_resp_bits_data_word_bypass[28]),
    .B(_01632_),
    .S(_08754_),
    .Z(_01633_)
  );
  MUX2_X1 _16685_ (
    .A(ex_reg_rs_msb_1[26]),
    .B(_01633_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[28])
  );
  OR2_X1 _16686_ (
    .A1(_08867_),
    .A2(_ex_op2_T[28]),
    .ZN(_01634_)
  );
  OR2_X1 _16687_ (
    .A1(_08842_),
    .A2(_01634_),
    .ZN(_01635_)
  );
  OR2_X1 _16688_ (
    .A1(mem_reg_rs2[28]),
    .A2(_08766_),
    .ZN(_01636_)
  );
  AND2_X1 _16689_ (
    .A1(_01635_),
    .A2(_01636_),
    .ZN(_01637_)
  );
  AND2_X1 _16690_ (
    .A1(_01629_),
    .A2(_01637_),
    .ZN(_00269_)
  );
  OR2_X1 _16691_ (
    .A1(_08851_),
    .A2(_08869_),
    .ZN(_01638_)
  );
  AND2_X1 _16692_ (
    .A1(mem_reg_wdata[29]),
    .A2(_08759_),
    .ZN(_01639_)
  );
  AND2_X1 _16693_ (
    .A1(wb_reg_wdata[29]),
    .A2(_08755_),
    .ZN(_01640_)
  );
  OR2_X1 _16694_ (
    .A1(_01639_),
    .A2(_01640_),
    .ZN(_01641_)
  );
  MUX2_X1 _16695_ (
    .A(io_dmem_resp_bits_data_word_bypass[29]),
    .B(_01641_),
    .S(_08754_),
    .Z(_01642_)
  );
  MUX2_X1 _16696_ (
    .A(ex_reg_rs_msb_1[27]),
    .B(_01642_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[29])
  );
  OR2_X1 _16697_ (
    .A1(_08867_),
    .A2(_ex_op2_T[29]),
    .ZN(_01643_)
  );
  OR2_X1 _16698_ (
    .A1(_08850_),
    .A2(_01643_),
    .ZN(_01644_)
  );
  OR2_X1 _16699_ (
    .A1(mem_reg_rs2[29]),
    .A2(_08766_),
    .ZN(_01645_)
  );
  AND2_X1 _16700_ (
    .A1(_01644_),
    .A2(_01645_),
    .ZN(_01646_)
  );
  AND2_X1 _16701_ (
    .A1(_01638_),
    .A2(_01646_),
    .ZN(_00270_)
  );
  OR2_X1 _16702_ (
    .A1(mem_reg_rs2[30]),
    .A2(_08766_),
    .ZN(_01647_)
  );
  AND2_X1 _16703_ (
    .A1(mem_reg_wdata[30]),
    .A2(_08759_),
    .ZN(_01648_)
  );
  AND2_X1 _16704_ (
    .A1(wb_reg_wdata[30]),
    .A2(_08755_),
    .ZN(_01649_)
  );
  OR2_X1 _16705_ (
    .A1(_01648_),
    .A2(_01649_),
    .ZN(_01650_)
  );
  MUX2_X1 _16706_ (
    .A(io_dmem_resp_bits_data_word_bypass[30]),
    .B(_01650_),
    .S(_08754_),
    .Z(_01651_)
  );
  MUX2_X1 _16707_ (
    .A(ex_reg_rs_msb_1[28]),
    .B(_01651_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[30])
  );
  OR2_X1 _16708_ (
    .A1(_08867_),
    .A2(_ex_op2_T[30]),
    .ZN(_01652_)
  );
  OR2_X1 _16709_ (
    .A1(_08857_),
    .A2(_08869_),
    .ZN(_01653_)
  );
  AND2_X1 _16710_ (
    .A1(_01652_),
    .A2(_01653_),
    .ZN(_01654_)
  );
  OR2_X1 _16711_ (
    .A1(_08767_),
    .A2(_01654_),
    .ZN(_01655_)
  );
  OR2_X1 _16712_ (
    .A1(_08858_),
    .A2(_01655_),
    .ZN(_01656_)
  );
  AND2_X1 _16713_ (
    .A1(_01647_),
    .A2(_01656_),
    .ZN(_00271_)
  );
  OR2_X1 _16714_ (
    .A1(mem_reg_rs2[31]),
    .A2(_08766_),
    .ZN(_01657_)
  );
  AND2_X1 _16715_ (
    .A1(mem_reg_wdata[31]),
    .A2(_08759_),
    .ZN(_01658_)
  );
  AND2_X1 _16716_ (
    .A1(wb_reg_wdata[31]),
    .A2(_08755_),
    .ZN(_01659_)
  );
  OR2_X1 _16717_ (
    .A1(_01658_),
    .A2(_01659_),
    .ZN(_01660_)
  );
  MUX2_X1 _16718_ (
    .A(io_dmem_resp_bits_data_word_bypass[31]),
    .B(_01660_),
    .S(_08754_),
    .Z(_01661_)
  );
  MUX2_X1 _16719_ (
    .A(ex_reg_rs_msb_1[29]),
    .B(_01661_),
    .S(ex_reg_rs_bypass_1),
    .Z(_ex_op2_T[31])
  );
  OR2_X1 _16720_ (
    .A1(_08867_),
    .A2(_ex_op2_T[31]),
    .ZN(_01662_)
  );
  OR2_X1 _16721_ (
    .A1(_08864_),
    .A2(_08869_),
    .ZN(_01663_)
  );
  AND2_X1 _16722_ (
    .A1(_01662_),
    .A2(_01663_),
    .ZN(_01664_)
  );
  OR2_X1 _16723_ (
    .A1(_08767_),
    .A2(_01664_),
    .ZN(_01665_)
  );
  OR2_X1 _16724_ (
    .A1(_08865_),
    .A2(_01665_),
    .ZN(_01666_)
  );
  AND2_X1 _16725_ (
    .A1(_01657_),
    .A2(_01666_),
    .ZN(_00272_)
  );
  MUX2_X1 _16726_ (
    .A(alu_io_out[0]),
    .B(mem_reg_wdata[0]),
    .S(_08752_),
    .Z(_00273_)
  );
  MUX2_X1 _16727_ (
    .A(alu_io_out[1]),
    .B(mem_reg_wdata[1]),
    .S(_08752_),
    .Z(_00274_)
  );
  MUX2_X1 _16728_ (
    .A(alu_io_out[2]),
    .B(mem_reg_wdata[2]),
    .S(_08752_),
    .Z(_00275_)
  );
  MUX2_X1 _16729_ (
    .A(alu_io_out[3]),
    .B(mem_reg_wdata[3]),
    .S(_08752_),
    .Z(_00276_)
  );
  MUX2_X1 _16730_ (
    .A(alu_io_out[4]),
    .B(mem_reg_wdata[4]),
    .S(_08752_),
    .Z(_00277_)
  );
  MUX2_X1 _16731_ (
    .A(alu_io_out[5]),
    .B(mem_reg_wdata[5]),
    .S(_08752_),
    .Z(_00278_)
  );
  MUX2_X1 _16732_ (
    .A(alu_io_out[6]),
    .B(mem_reg_wdata[6]),
    .S(_08752_),
    .Z(_00279_)
  );
  MUX2_X1 _16733_ (
    .A(alu_io_out[7]),
    .B(mem_reg_wdata[7]),
    .S(_08752_),
    .Z(_00280_)
  );
  MUX2_X1 _16734_ (
    .A(alu_io_out[8]),
    .B(mem_reg_wdata[8]),
    .S(_08752_),
    .Z(_00281_)
  );
  MUX2_X1 _16735_ (
    .A(alu_io_out[9]),
    .B(mem_reg_wdata[9]),
    .S(_08752_),
    .Z(_00282_)
  );
  MUX2_X1 _16736_ (
    .A(alu_io_out[10]),
    .B(mem_reg_wdata[10]),
    .S(_08752_),
    .Z(_00283_)
  );
  MUX2_X1 _16737_ (
    .A(alu_io_out[11]),
    .B(mem_reg_wdata[11]),
    .S(_08752_),
    .Z(_00284_)
  );
  MUX2_X1 _16738_ (
    .A(alu_io_out[12]),
    .B(mem_reg_wdata[12]),
    .S(_08752_),
    .Z(_00285_)
  );
  MUX2_X1 _16739_ (
    .A(alu_io_out[13]),
    .B(mem_reg_wdata[13]),
    .S(_08752_),
    .Z(_00286_)
  );
  MUX2_X1 _16740_ (
    .A(alu_io_out[14]),
    .B(mem_reg_wdata[14]),
    .S(_08752_),
    .Z(_00287_)
  );
  MUX2_X1 _16741_ (
    .A(alu_io_out[15]),
    .B(mem_reg_wdata[15]),
    .S(_08752_),
    .Z(_00288_)
  );
  MUX2_X1 _16742_ (
    .A(alu_io_out[16]),
    .B(mem_reg_wdata[16]),
    .S(_08752_),
    .Z(_00289_)
  );
  MUX2_X1 _16743_ (
    .A(alu_io_out[17]),
    .B(mem_reg_wdata[17]),
    .S(_08752_),
    .Z(_00290_)
  );
  MUX2_X1 _16744_ (
    .A(alu_io_out[18]),
    .B(mem_reg_wdata[18]),
    .S(_08752_),
    .Z(_00291_)
  );
  MUX2_X1 _16745_ (
    .A(alu_io_out[19]),
    .B(mem_reg_wdata[19]),
    .S(_08752_),
    .Z(_00292_)
  );
  MUX2_X1 _16746_ (
    .A(alu_io_out[20]),
    .B(mem_reg_wdata[20]),
    .S(_08752_),
    .Z(_00293_)
  );
  MUX2_X1 _16747_ (
    .A(alu_io_out[21]),
    .B(mem_reg_wdata[21]),
    .S(_08752_),
    .Z(_00294_)
  );
  MUX2_X1 _16748_ (
    .A(alu_io_out[22]),
    .B(mem_reg_wdata[22]),
    .S(_08752_),
    .Z(_00295_)
  );
  MUX2_X1 _16749_ (
    .A(alu_io_out[23]),
    .B(mem_reg_wdata[23]),
    .S(_08752_),
    .Z(_00296_)
  );
  MUX2_X1 _16750_ (
    .A(alu_io_out[24]),
    .B(mem_reg_wdata[24]),
    .S(_08752_),
    .Z(_00297_)
  );
  MUX2_X1 _16751_ (
    .A(alu_io_out[25]),
    .B(mem_reg_wdata[25]),
    .S(_08752_),
    .Z(_00298_)
  );
  MUX2_X1 _16752_ (
    .A(alu_io_out[26]),
    .B(mem_reg_wdata[26]),
    .S(_08752_),
    .Z(_00299_)
  );
  MUX2_X1 _16753_ (
    .A(alu_io_out[27]),
    .B(mem_reg_wdata[27]),
    .S(_08752_),
    .Z(_00300_)
  );
  MUX2_X1 _16754_ (
    .A(alu_io_out[28]),
    .B(mem_reg_wdata[28]),
    .S(_08752_),
    .Z(_00301_)
  );
  MUX2_X1 _16755_ (
    .A(alu_io_out[29]),
    .B(mem_reg_wdata[29]),
    .S(_08752_),
    .Z(_00302_)
  );
  MUX2_X1 _16756_ (
    .A(alu_io_out[30]),
    .B(mem_reg_wdata[30]),
    .S(_08752_),
    .Z(_00303_)
  );
  MUX2_X1 _16757_ (
    .A(alu_io_out[31]),
    .B(mem_reg_wdata[31]),
    .S(_08752_),
    .Z(_00304_)
  );
  MUX2_X1 _16758_ (
    .A(ex_reg_raw_inst[0]),
    .B(mem_reg_raw_inst[0]),
    .S(_08752_),
    .Z(_00305_)
  );
  MUX2_X1 _16759_ (
    .A(ex_reg_raw_inst[1]),
    .B(mem_reg_raw_inst[1]),
    .S(_08752_),
    .Z(_00306_)
  );
  MUX2_X1 _16760_ (
    .A(ex_reg_raw_inst[2]),
    .B(mem_reg_raw_inst[2]),
    .S(_08752_),
    .Z(_00307_)
  );
  MUX2_X1 _16761_ (
    .A(ex_reg_raw_inst[3]),
    .B(mem_reg_raw_inst[3]),
    .S(_08752_),
    .Z(_00308_)
  );
  MUX2_X1 _16762_ (
    .A(ex_reg_raw_inst[4]),
    .B(mem_reg_raw_inst[4]),
    .S(_08752_),
    .Z(_00309_)
  );
  MUX2_X1 _16763_ (
    .A(ex_reg_raw_inst[5]),
    .B(mem_reg_raw_inst[5]),
    .S(_08752_),
    .Z(_00310_)
  );
  MUX2_X1 _16764_ (
    .A(ex_reg_raw_inst[6]),
    .B(mem_reg_raw_inst[6]),
    .S(_08752_),
    .Z(_00311_)
  );
  MUX2_X1 _16765_ (
    .A(ex_reg_raw_inst[7]),
    .B(mem_reg_raw_inst[7]),
    .S(_08752_),
    .Z(_00312_)
  );
  MUX2_X1 _16766_ (
    .A(ex_reg_raw_inst[8]),
    .B(mem_reg_raw_inst[8]),
    .S(_08752_),
    .Z(_00313_)
  );
  MUX2_X1 _16767_ (
    .A(ex_reg_raw_inst[9]),
    .B(mem_reg_raw_inst[9]),
    .S(_08752_),
    .Z(_00314_)
  );
  MUX2_X1 _16768_ (
    .A(ex_reg_raw_inst[10]),
    .B(mem_reg_raw_inst[10]),
    .S(_08752_),
    .Z(_00315_)
  );
  MUX2_X1 _16769_ (
    .A(ex_reg_raw_inst[11]),
    .B(mem_reg_raw_inst[11]),
    .S(_08752_),
    .Z(_00316_)
  );
  MUX2_X1 _16770_ (
    .A(ex_reg_raw_inst[12]),
    .B(mem_reg_raw_inst[12]),
    .S(_08752_),
    .Z(_00317_)
  );
  MUX2_X1 _16771_ (
    .A(ex_reg_raw_inst[13]),
    .B(mem_reg_raw_inst[13]),
    .S(_08752_),
    .Z(_00318_)
  );
  MUX2_X1 _16772_ (
    .A(ex_reg_raw_inst[14]),
    .B(mem_reg_raw_inst[14]),
    .S(_08752_),
    .Z(_00319_)
  );
  MUX2_X1 _16773_ (
    .A(ex_reg_raw_inst[15]),
    .B(mem_reg_raw_inst[15]),
    .S(_08752_),
    .Z(_00320_)
  );
  MUX2_X1 _16774_ (
    .A(ex_reg_inst[7]),
    .B(mem_reg_inst[7]),
    .S(_08752_),
    .Z(_00321_)
  );
  MUX2_X1 _16775_ (
    .A(ex_reg_inst[8]),
    .B(mem_reg_inst[8]),
    .S(_08752_),
    .Z(_00322_)
  );
  MUX2_X1 _16776_ (
    .A(ex_reg_inst[9]),
    .B(mem_reg_inst[9]),
    .S(_08752_),
    .Z(_00323_)
  );
  MUX2_X1 _16777_ (
    .A(ex_reg_inst[10]),
    .B(mem_reg_inst[10]),
    .S(_08752_),
    .Z(_00324_)
  );
  MUX2_X1 _16778_ (
    .A(ex_reg_inst[11]),
    .B(mem_reg_inst[11]),
    .S(_08752_),
    .Z(_00325_)
  );
  MUX2_X1 _16779_ (
    .A(ex_reg_inst[12]),
    .B(mem_reg_inst[12]),
    .S(_08752_),
    .Z(_00326_)
  );
  MUX2_X1 _16780_ (
    .A(ex_reg_inst[13]),
    .B(mem_reg_inst[13]),
    .S(_08752_),
    .Z(_00327_)
  );
  MUX2_X1 _16781_ (
    .A(ex_reg_inst[14]),
    .B(mem_reg_inst[14]),
    .S(_08752_),
    .Z(_00328_)
  );
  MUX2_X1 _16782_ (
    .A(ex_reg_inst[15]),
    .B(mem_reg_inst[15]),
    .S(_08752_),
    .Z(_00329_)
  );
  MUX2_X1 _16783_ (
    .A(ex_reg_inst[16]),
    .B(mem_reg_inst[16]),
    .S(_08752_),
    .Z(_00330_)
  );
  MUX2_X1 _16784_ (
    .A(ex_reg_inst[17]),
    .B(mem_reg_inst[17]),
    .S(_08752_),
    .Z(_00331_)
  );
  MUX2_X1 _16785_ (
    .A(ex_reg_inst[18]),
    .B(mem_reg_inst[18]),
    .S(_08752_),
    .Z(_00332_)
  );
  MUX2_X1 _16786_ (
    .A(ex_reg_inst[19]),
    .B(mem_reg_inst[19]),
    .S(_08752_),
    .Z(_00333_)
  );
  MUX2_X1 _16787_ (
    .A(ex_reg_inst[20]),
    .B(mem_reg_inst[20]),
    .S(_08752_),
    .Z(_00334_)
  );
  MUX2_X1 _16788_ (
    .A(ex_reg_inst[21]),
    .B(mem_reg_inst[21]),
    .S(_08752_),
    .Z(_00335_)
  );
  MUX2_X1 _16789_ (
    .A(ex_reg_inst[22]),
    .B(mem_reg_inst[22]),
    .S(_08752_),
    .Z(_00336_)
  );
  MUX2_X1 _16790_ (
    .A(ex_reg_inst[23]),
    .B(mem_reg_inst[23]),
    .S(_08752_),
    .Z(_00337_)
  );
  MUX2_X1 _16791_ (
    .A(ex_reg_inst[24]),
    .B(mem_reg_inst[24]),
    .S(_08752_),
    .Z(_00338_)
  );
  MUX2_X1 _16792_ (
    .A(ex_reg_inst[25]),
    .B(mem_reg_inst[25]),
    .S(_08752_),
    .Z(_00339_)
  );
  MUX2_X1 _16793_ (
    .A(ex_reg_inst[26]),
    .B(mem_reg_inst[26]),
    .S(_08752_),
    .Z(_00340_)
  );
  MUX2_X1 _16794_ (
    .A(ex_reg_inst[27]),
    .B(mem_reg_inst[27]),
    .S(_08752_),
    .Z(_00341_)
  );
  MUX2_X1 _16795_ (
    .A(ex_reg_inst[28]),
    .B(mem_reg_inst[28]),
    .S(_08752_),
    .Z(_00342_)
  );
  MUX2_X1 _16796_ (
    .A(ex_reg_inst[29]),
    .B(mem_reg_inst[29]),
    .S(_08752_),
    .Z(_00343_)
  );
  MUX2_X1 _16797_ (
    .A(ex_reg_inst[30]),
    .B(mem_reg_inst[30]),
    .S(_08752_),
    .Z(_00344_)
  );
  MUX2_X1 _16798_ (
    .A(ex_reg_inst[31]),
    .B(mem_reg_inst[31]),
    .S(_08752_),
    .Z(_00345_)
  );
  MUX2_X1 _16799_ (
    .A(ex_reg_pc[0]),
    .B(mem_reg_pc[0]),
    .S(_08752_),
    .Z(_00346_)
  );
  MUX2_X1 _16800_ (
    .A(ex_reg_pc[1]),
    .B(mem_reg_pc[1]),
    .S(_08752_),
    .Z(_00347_)
  );
  MUX2_X1 _16801_ (
    .A(ex_reg_pc[2]),
    .B(mem_reg_pc[2]),
    .S(_08752_),
    .Z(_00348_)
  );
  MUX2_X1 _16802_ (
    .A(ex_reg_pc[3]),
    .B(mem_reg_pc[3]),
    .S(_08752_),
    .Z(_00349_)
  );
  MUX2_X1 _16803_ (
    .A(ex_reg_pc[4]),
    .B(mem_reg_pc[4]),
    .S(_08752_),
    .Z(_00350_)
  );
  MUX2_X1 _16804_ (
    .A(ex_reg_pc[5]),
    .B(mem_reg_pc[5]),
    .S(_08752_),
    .Z(_00351_)
  );
  MUX2_X1 _16805_ (
    .A(ex_reg_pc[6]),
    .B(mem_reg_pc[6]),
    .S(_08752_),
    .Z(_00352_)
  );
  MUX2_X1 _16806_ (
    .A(ex_reg_pc[7]),
    .B(mem_reg_pc[7]),
    .S(_08752_),
    .Z(_00353_)
  );
  MUX2_X1 _16807_ (
    .A(ex_reg_pc[8]),
    .B(mem_reg_pc[8]),
    .S(_08752_),
    .Z(_00354_)
  );
  MUX2_X1 _16808_ (
    .A(ex_reg_pc[9]),
    .B(mem_reg_pc[9]),
    .S(_08752_),
    .Z(_00355_)
  );
  MUX2_X1 _16809_ (
    .A(ex_reg_pc[10]),
    .B(mem_reg_pc[10]),
    .S(_08752_),
    .Z(_00356_)
  );
  MUX2_X1 _16810_ (
    .A(ex_reg_pc[11]),
    .B(mem_reg_pc[11]),
    .S(_08752_),
    .Z(_00357_)
  );
  MUX2_X1 _16811_ (
    .A(ex_reg_pc[12]),
    .B(mem_reg_pc[12]),
    .S(_08752_),
    .Z(_00358_)
  );
  MUX2_X1 _16812_ (
    .A(ex_reg_pc[13]),
    .B(mem_reg_pc[13]),
    .S(_08752_),
    .Z(_00359_)
  );
  MUX2_X1 _16813_ (
    .A(ex_reg_pc[14]),
    .B(mem_reg_pc[14]),
    .S(_08752_),
    .Z(_00360_)
  );
  MUX2_X1 _16814_ (
    .A(ex_reg_pc[15]),
    .B(mem_reg_pc[15]),
    .S(_08752_),
    .Z(_00361_)
  );
  MUX2_X1 _16815_ (
    .A(ex_reg_pc[16]),
    .B(mem_reg_pc[16]),
    .S(_08752_),
    .Z(_00362_)
  );
  MUX2_X1 _16816_ (
    .A(ex_reg_pc[17]),
    .B(mem_reg_pc[17]),
    .S(_08752_),
    .Z(_00363_)
  );
  MUX2_X1 _16817_ (
    .A(ex_reg_pc[18]),
    .B(mem_reg_pc[18]),
    .S(_08752_),
    .Z(_00364_)
  );
  MUX2_X1 _16818_ (
    .A(ex_reg_pc[19]),
    .B(mem_reg_pc[19]),
    .S(_08752_),
    .Z(_00365_)
  );
  MUX2_X1 _16819_ (
    .A(ex_reg_pc[20]),
    .B(mem_reg_pc[20]),
    .S(_08752_),
    .Z(_00366_)
  );
  MUX2_X1 _16820_ (
    .A(ex_reg_pc[21]),
    .B(mem_reg_pc[21]),
    .S(_08752_),
    .Z(_00367_)
  );
  MUX2_X1 _16821_ (
    .A(ex_reg_pc[22]),
    .B(mem_reg_pc[22]),
    .S(_08752_),
    .Z(_00368_)
  );
  MUX2_X1 _16822_ (
    .A(ex_reg_pc[23]),
    .B(mem_reg_pc[23]),
    .S(_08752_),
    .Z(_00369_)
  );
  MUX2_X1 _16823_ (
    .A(ex_reg_pc[24]),
    .B(mem_reg_pc[24]),
    .S(_08752_),
    .Z(_00370_)
  );
  MUX2_X1 _16824_ (
    .A(ex_reg_pc[25]),
    .B(mem_reg_pc[25]),
    .S(_08752_),
    .Z(_00371_)
  );
  MUX2_X1 _16825_ (
    .A(ex_reg_pc[26]),
    .B(mem_reg_pc[26]),
    .S(_08752_),
    .Z(_00372_)
  );
  MUX2_X1 _16826_ (
    .A(ex_reg_pc[27]),
    .B(mem_reg_pc[27]),
    .S(_08752_),
    .Z(_00373_)
  );
  MUX2_X1 _16827_ (
    .A(ex_reg_pc[28]),
    .B(mem_reg_pc[28]),
    .S(_08752_),
    .Z(_00374_)
  );
  MUX2_X1 _16828_ (
    .A(ex_reg_pc[29]),
    .B(mem_reg_pc[29]),
    .S(_08752_),
    .Z(_00375_)
  );
  MUX2_X1 _16829_ (
    .A(ex_reg_pc[30]),
    .B(mem_reg_pc[30]),
    .S(_08752_),
    .Z(_00376_)
  );
  MUX2_X1 _16830_ (
    .A(ex_reg_pc[31]),
    .B(mem_reg_pc[31]),
    .S(_08752_),
    .Z(_00377_)
  );
  AND2_X1 _16831_ (
    .A1(mem_reg_store),
    .A2(_08752_),
    .ZN(_01667_)
  );
  AND2_X1 _16832_ (
    .A1(ex_ctrl_mem_cmd[2]),
    .A2(_00025_),
    .ZN(_01668_)
  );
  OR2_X1 _16833_ (
    .A1(_00024_),
    .A2(_01668_),
    .ZN(_01669_)
  );
  OR2_X1 _16834_ (
    .A1(ex_ctrl_mem_cmd[3]),
    .A2(_00025_),
    .ZN(_01670_)
  );
  INV_X1 _16835_ (
    .A(_01670_),
    .ZN(_01671_)
  );
  OR2_X1 _16836_ (
    .A1(ex_ctrl_mem_cmd[0]),
    .A2(ex_ctrl_mem_cmd[1]),
    .ZN(_01672_)
  );
  OR2_X1 _16837_ (
    .A1(_01670_),
    .A2(_01672_),
    .ZN(_01673_)
  );
  AND2_X1 _16838_ (
    .A1(_01669_),
    .A2(_01673_),
    .ZN(_01674_)
  );
  AND2_X1 _16839_ (
    .A1(ex_ctrl_mem_cmd[0]),
    .A2(_00027_),
    .ZN(_01675_)
  );
  INV_X1 _16840_ (
    .A(_01675_),
    .ZN(_01676_)
  );
  AND2_X1 _16841_ (
    .A1(ex_ctrl_mem_cmd[1]),
    .A2(_00026_),
    .ZN(_01677_)
  );
  OR2_X1 _16842_ (
    .A1(_01674_),
    .A2(_01677_),
    .ZN(_01678_)
  );
  INV_X1 _16843_ (
    .A(_01678_),
    .ZN(_01679_)
  );
  AND2_X1 _16844_ (
    .A1(_01676_),
    .A2(_01679_),
    .ZN(_01680_)
  );
  AND2_X1 _16845_ (
    .A1(_03057_),
    .A2(_01671_),
    .ZN(_01681_)
  );
  OR2_X1 _16846_ (
    .A1(ex_ctrl_mem_cmd[2]),
    .A2(ex_ctrl_mem_cmd[3]),
    .ZN(_01682_)
  );
  OR2_X1 _16847_ (
    .A1(ex_ctrl_mem_cmd[1]),
    .A2(_01682_),
    .ZN(_01683_)
  );
  INV_X1 _16848_ (
    .A(_01683_),
    .ZN(_01684_)
  );
  OR2_X1 _16849_ (
    .A1(_01681_),
    .A2(_01684_),
    .ZN(_01685_)
  );
  AND2_X1 _16850_ (
    .A1(_03056_),
    .A2(_01685_),
    .ZN(_01686_)
  );
  OR2_X1 _16851_ (
    .A1(_01680_),
    .A2(_01686_),
    .ZN(_01687_)
  );
  AND2_X1 _16852_ (
    .A1(_08764_),
    .A2(_01687_),
    .ZN(_01688_)
  );
  OR2_X1 _16853_ (
    .A1(_01667_),
    .A2(_01688_),
    .ZN(_00378_)
  );
  AND2_X1 _16854_ (
    .A1(mem_reg_load),
    .A2(_08752_),
    .ZN(_01689_)
  );
  AND2_X1 _16855_ (
    .A1(_03032_),
    .A2(_01685_),
    .ZN(_01690_)
  );
  AND2_X1 _16856_ (
    .A1(_03056_),
    .A2(_01681_),
    .ZN(_01691_)
  );
  OR2_X1 _16857_ (
    .A1(_01690_),
    .A2(_01691_),
    .ZN(_01692_)
  );
  OR2_X1 _16858_ (
    .A1(_01680_),
    .A2(_01692_),
    .ZN(_01693_)
  );
  AND2_X1 _16859_ (
    .A1(_08764_),
    .A2(_01693_),
    .ZN(_01694_)
  );
  OR2_X1 _16860_ (
    .A1(_01689_),
    .A2(_01694_),
    .ZN(_00379_)
  );
  OR2_X1 _16861_ (
    .A1(_10442_[1]),
    .A2(_01691_),
    .ZN(_01695_)
  );
  MUX2_X1 _16862_ (
    .A(mem_reg_slow_bypass),
    .B(_01695_),
    .S(_08753_),
    .Z(_00380_)
  );
  MUX2_X1 _16863_ (
    .A(ex_reg_cause[0]),
    .B(mem_reg_cause[0]),
    .S(_08752_),
    .Z(_00381_)
  );
  MUX2_X1 _16864_ (
    .A(ex_reg_cause[1]),
    .B(mem_reg_cause[1]),
    .S(_08752_),
    .Z(_00382_)
  );
  MUX2_X1 _16865_ (
    .A(ex_reg_cause[2]),
    .B(mem_reg_cause[2]),
    .S(_08752_),
    .Z(_00383_)
  );
  MUX2_X1 _16866_ (
    .A(ex_reg_cause[3]),
    .B(mem_reg_cause[3]),
    .S(_08752_),
    .Z(_00384_)
  );
  MUX2_X1 _16867_ (
    .A(ex_reg_cause[4]),
    .B(mem_reg_cause[4]),
    .S(_08752_),
    .Z(_00385_)
  );
  MUX2_X1 _16868_ (
    .A(ex_reg_cause[5]),
    .B(mem_reg_cause[5]),
    .S(_08752_),
    .Z(_00386_)
  );
  MUX2_X1 _16869_ (
    .A(ex_reg_cause[6]),
    .B(mem_reg_cause[6]),
    .S(_08752_),
    .Z(_00387_)
  );
  MUX2_X1 _16870_ (
    .A(ex_reg_cause[7]),
    .B(mem_reg_cause[7]),
    .S(_08752_),
    .Z(_00388_)
  );
  MUX2_X1 _16871_ (
    .A(ex_reg_cause[8]),
    .B(mem_reg_cause[8]),
    .S(_08752_),
    .Z(_00389_)
  );
  MUX2_X1 _16872_ (
    .A(ex_reg_cause[9]),
    .B(mem_reg_cause[9]),
    .S(_08752_),
    .Z(_00390_)
  );
  MUX2_X1 _16873_ (
    .A(ex_reg_cause[10]),
    .B(mem_reg_cause[10]),
    .S(_08752_),
    .Z(_00391_)
  );
  MUX2_X1 _16874_ (
    .A(ex_reg_cause[11]),
    .B(mem_reg_cause[11]),
    .S(_08752_),
    .Z(_00392_)
  );
  MUX2_X1 _16875_ (
    .A(ex_reg_cause[12]),
    .B(mem_reg_cause[12]),
    .S(_08752_),
    .Z(_00393_)
  );
  MUX2_X1 _16876_ (
    .A(ex_reg_cause[13]),
    .B(mem_reg_cause[13]),
    .S(_08752_),
    .Z(_00394_)
  );
  MUX2_X1 _16877_ (
    .A(ex_reg_cause[14]),
    .B(mem_reg_cause[14]),
    .S(_08752_),
    .Z(_00395_)
  );
  MUX2_X1 _16878_ (
    .A(ex_reg_cause[15]),
    .B(mem_reg_cause[15]),
    .S(_08752_),
    .Z(_00396_)
  );
  MUX2_X1 _16879_ (
    .A(ex_reg_cause[16]),
    .B(mem_reg_cause[16]),
    .S(_08752_),
    .Z(_00397_)
  );
  MUX2_X1 _16880_ (
    .A(ex_reg_cause[17]),
    .B(mem_reg_cause[17]),
    .S(_08752_),
    .Z(_00398_)
  );
  MUX2_X1 _16881_ (
    .A(ex_reg_cause[18]),
    .B(mem_reg_cause[18]),
    .S(_08752_),
    .Z(_00399_)
  );
  MUX2_X1 _16882_ (
    .A(ex_reg_cause[19]),
    .B(mem_reg_cause[19]),
    .S(_08752_),
    .Z(_00400_)
  );
  MUX2_X1 _16883_ (
    .A(ex_reg_cause[20]),
    .B(mem_reg_cause[20]),
    .S(_08752_),
    .Z(_00401_)
  );
  MUX2_X1 _16884_ (
    .A(ex_reg_cause[21]),
    .B(mem_reg_cause[21]),
    .S(_08752_),
    .Z(_00402_)
  );
  MUX2_X1 _16885_ (
    .A(ex_reg_cause[22]),
    .B(mem_reg_cause[22]),
    .S(_08752_),
    .Z(_00403_)
  );
  MUX2_X1 _16886_ (
    .A(ex_reg_cause[23]),
    .B(mem_reg_cause[23]),
    .S(_08752_),
    .Z(_00404_)
  );
  MUX2_X1 _16887_ (
    .A(ex_reg_cause[24]),
    .B(mem_reg_cause[24]),
    .S(_08752_),
    .Z(_00405_)
  );
  MUX2_X1 _16888_ (
    .A(ex_reg_cause[25]),
    .B(mem_reg_cause[25]),
    .S(_08752_),
    .Z(_00406_)
  );
  MUX2_X1 _16889_ (
    .A(ex_reg_cause[26]),
    .B(mem_reg_cause[26]),
    .S(_08752_),
    .Z(_00407_)
  );
  MUX2_X1 _16890_ (
    .A(ex_reg_cause[27]),
    .B(mem_reg_cause[27]),
    .S(_08752_),
    .Z(_00408_)
  );
  MUX2_X1 _16891_ (
    .A(ex_reg_cause[28]),
    .B(mem_reg_cause[28]),
    .S(_08752_),
    .Z(_00409_)
  );
  MUX2_X1 _16892_ (
    .A(ex_reg_cause[29]),
    .B(mem_reg_cause[29]),
    .S(_08752_),
    .Z(_00410_)
  );
  MUX2_X1 _16893_ (
    .A(ex_reg_cause[30]),
    .B(mem_reg_cause[30]),
    .S(_08752_),
    .Z(_00411_)
  );
  MUX2_X1 _16894_ (
    .A(ex_reg_cause[31]),
    .B(mem_reg_cause[31]),
    .S(_08752_),
    .Z(_00412_)
  );
  AND2_X1 _16895_ (
    .A1(ex_ctrl_jalr),
    .A2(bpu_io_status_debug),
    .ZN(_01696_)
  );
  OR2_X1 _16896_ (
    .A1(ex_reg_flush_pipe),
    .A2(_01696_),
    .ZN(_01697_)
  );
  MUX2_X1 _16897_ (
    .A(_01697_),
    .B(mem_reg_flush_pipe),
    .S(_08752_),
    .Z(_00413_)
  );
  MUX2_X1 _16898_ (
    .A(ex_reg_rvc),
    .B(mem_reg_rvc),
    .S(_08752_),
    .Z(_00414_)
  );
  OR2_X1 _16899_ (
    .A1(_03586_),
    .A2(_04039_),
    .ZN(_01698_)
  );
  INV_X1 _16900_ (
    .A(_01698_),
    .ZN(_01699_)
  );
  MUX2_X1 _16901_ (
    .A(ex_reg_raw_inst[0]),
    .B(ibuf_io_inst_0_bits_raw[0]),
    .S(_01698_),
    .Z(_00415_)
  );
  MUX2_X1 _16902_ (
    .A(ex_reg_raw_inst[1]),
    .B(ibuf_io_inst_0_bits_raw[1]),
    .S(_01698_),
    .Z(_00416_)
  );
  MUX2_X1 _16903_ (
    .A(ex_reg_raw_inst[2]),
    .B(ibuf_io_inst_0_bits_raw[2]),
    .S(_01698_),
    .Z(_00417_)
  );
  MUX2_X1 _16904_ (
    .A(ex_reg_raw_inst[3]),
    .B(ibuf_io_inst_0_bits_raw[3]),
    .S(_01698_),
    .Z(_00418_)
  );
  MUX2_X1 _16905_ (
    .A(ex_reg_raw_inst[4]),
    .B(ibuf_io_inst_0_bits_raw[4]),
    .S(_01698_),
    .Z(_00419_)
  );
  MUX2_X1 _16906_ (
    .A(ex_reg_raw_inst[5]),
    .B(ibuf_io_inst_0_bits_raw[5]),
    .S(_01698_),
    .Z(_00420_)
  );
  MUX2_X1 _16907_ (
    .A(ex_reg_raw_inst[6]),
    .B(ibuf_io_inst_0_bits_raw[6]),
    .S(_01698_),
    .Z(_00421_)
  );
  MUX2_X1 _16908_ (
    .A(ex_reg_raw_inst[7]),
    .B(ibuf_io_inst_0_bits_raw[7]),
    .S(_01698_),
    .Z(_00422_)
  );
  MUX2_X1 _16909_ (
    .A(ex_reg_raw_inst[8]),
    .B(ibuf_io_inst_0_bits_raw[8]),
    .S(_01698_),
    .Z(_00423_)
  );
  MUX2_X1 _16910_ (
    .A(ex_reg_raw_inst[9]),
    .B(ibuf_io_inst_0_bits_raw[9]),
    .S(_01698_),
    .Z(_00424_)
  );
  MUX2_X1 _16911_ (
    .A(ex_reg_raw_inst[10]),
    .B(ibuf_io_inst_0_bits_raw[10]),
    .S(_01698_),
    .Z(_00425_)
  );
  MUX2_X1 _16912_ (
    .A(ex_reg_raw_inst[11]),
    .B(ibuf_io_inst_0_bits_raw[11]),
    .S(_01698_),
    .Z(_00426_)
  );
  MUX2_X1 _16913_ (
    .A(ex_reg_raw_inst[12]),
    .B(ibuf_io_inst_0_bits_raw[12]),
    .S(_01698_),
    .Z(_00427_)
  );
  MUX2_X1 _16914_ (
    .A(ex_reg_raw_inst[13]),
    .B(ibuf_io_inst_0_bits_raw[13]),
    .S(_01698_),
    .Z(_00428_)
  );
  MUX2_X1 _16915_ (
    .A(ex_reg_raw_inst[14]),
    .B(ibuf_io_inst_0_bits_raw[14]),
    .S(_01698_),
    .Z(_00429_)
  );
  MUX2_X1 _16916_ (
    .A(ex_reg_raw_inst[15]),
    .B(ibuf_io_inst_0_bits_raw[15]),
    .S(_01698_),
    .Z(_00430_)
  );
  MUX2_X1 _16917_ (
    .A(ex_reg_inst[7]),
    .B(csr_io_decode_0_inst[7]),
    .S(_01698_),
    .Z(_00431_)
  );
  MUX2_X1 _16918_ (
    .A(ex_reg_inst[8]),
    .B(csr_io_decode_0_inst[8]),
    .S(_01698_),
    .Z(_00432_)
  );
  MUX2_X1 _16919_ (
    .A(ex_reg_inst[9]),
    .B(csr_io_decode_0_inst[9]),
    .S(_01698_),
    .Z(_00433_)
  );
  MUX2_X1 _16920_ (
    .A(ex_reg_inst[10]),
    .B(csr_io_decode_0_inst[10]),
    .S(_01698_),
    .Z(_00434_)
  );
  MUX2_X1 _16921_ (
    .A(ex_reg_inst[11]),
    .B(csr_io_decode_0_inst[11]),
    .S(_01698_),
    .Z(_00435_)
  );
  MUX2_X1 _16922_ (
    .A(ex_reg_inst[12]),
    .B(csr_io_decode_0_inst[12]),
    .S(_01698_),
    .Z(_00436_)
  );
  MUX2_X1 _16923_ (
    .A(ex_reg_inst[13]),
    .B(csr_io_decode_0_inst[13]),
    .S(_01698_),
    .Z(_00437_)
  );
  MUX2_X1 _16924_ (
    .A(ex_reg_inst[14]),
    .B(csr_io_decode_0_inst[14]),
    .S(_01698_),
    .Z(_00438_)
  );
  MUX2_X1 _16925_ (
    .A(ex_reg_inst[15]),
    .B(csr_io_decode_0_inst[15]),
    .S(_01698_),
    .Z(_00439_)
  );
  MUX2_X1 _16926_ (
    .A(ex_reg_inst[16]),
    .B(csr_io_decode_0_inst[16]),
    .S(_01698_),
    .Z(_00440_)
  );
  MUX2_X1 _16927_ (
    .A(ex_reg_inst[17]),
    .B(csr_io_decode_0_inst[17]),
    .S(_01698_),
    .Z(_00441_)
  );
  MUX2_X1 _16928_ (
    .A(ex_reg_inst[18]),
    .B(csr_io_decode_0_inst[18]),
    .S(_01698_),
    .Z(_00442_)
  );
  MUX2_X1 _16929_ (
    .A(ex_reg_inst[19]),
    .B(csr_io_decode_0_inst[19]),
    .S(_01698_),
    .Z(_00443_)
  );
  MUX2_X1 _16930_ (
    .A(ex_reg_inst[20]),
    .B(csr_io_decode_0_inst[20]),
    .S(_01698_),
    .Z(_00444_)
  );
  MUX2_X1 _16931_ (
    .A(ex_reg_inst[21]),
    .B(csr_io_decode_0_inst[21]),
    .S(_01698_),
    .Z(_00445_)
  );
  MUX2_X1 _16932_ (
    .A(ex_reg_inst[22]),
    .B(csr_io_decode_0_inst[22]),
    .S(_01698_),
    .Z(_00446_)
  );
  MUX2_X1 _16933_ (
    .A(ex_reg_inst[23]),
    .B(csr_io_decode_0_inst[23]),
    .S(_01698_),
    .Z(_00447_)
  );
  MUX2_X1 _16934_ (
    .A(ex_reg_inst[24]),
    .B(csr_io_decode_0_inst[24]),
    .S(_01698_),
    .Z(_00448_)
  );
  MUX2_X1 _16935_ (
    .A(ex_reg_inst[25]),
    .B(csr_io_decode_0_inst[25]),
    .S(_01698_),
    .Z(_00449_)
  );
  MUX2_X1 _16936_ (
    .A(ex_reg_inst[26]),
    .B(csr_io_decode_0_inst[26]),
    .S(_01698_),
    .Z(_00450_)
  );
  MUX2_X1 _16937_ (
    .A(ex_reg_inst[27]),
    .B(csr_io_decode_0_inst[27]),
    .S(_01698_),
    .Z(_00451_)
  );
  MUX2_X1 _16938_ (
    .A(ex_reg_inst[28]),
    .B(csr_io_decode_0_inst[28]),
    .S(_01698_),
    .Z(_00452_)
  );
  MUX2_X1 _16939_ (
    .A(ex_reg_inst[29]),
    .B(csr_io_decode_0_inst[29]),
    .S(_01698_),
    .Z(_00453_)
  );
  MUX2_X1 _16940_ (
    .A(ex_reg_inst[30]),
    .B(csr_io_decode_0_inst[30]),
    .S(_01698_),
    .Z(_00454_)
  );
  MUX2_X1 _16941_ (
    .A(ex_reg_inst[31]),
    .B(csr_io_decode_0_inst[31]),
    .S(_01698_),
    .Z(_00455_)
  );
  MUX2_X1 _16942_ (
    .A(csr_io_decode_0_inst[12]),
    .B(ex_reg_mem_size[0]),
    .S(_04146_),
    .Z(_00456_)
  );
  MUX2_X1 _16943_ (
    .A(csr_io_decode_0_inst[13]),
    .B(ex_reg_mem_size[1]),
    .S(_04146_),
    .Z(_00457_)
  );
  AND2_X1 _16944_ (
    .A1(ex_reg_cause[5]),
    .A2(_01699_),
    .ZN(_01700_)
  );
  AND2_X1 _16945_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[5]),
    .ZN(_01701_)
  );
  OR2_X1 _16946_ (
    .A1(_01700_),
    .A2(_01701_),
    .ZN(_00458_)
  );
  AND2_X1 _16947_ (
    .A1(ex_reg_cause[6]),
    .A2(_01699_),
    .ZN(_01702_)
  );
  AND2_X1 _16948_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[6]),
    .ZN(_01703_)
  );
  OR2_X1 _16949_ (
    .A1(_01702_),
    .A2(_01703_),
    .ZN(_00459_)
  );
  AND2_X1 _16950_ (
    .A1(ex_reg_cause[7]),
    .A2(_01699_),
    .ZN(_01704_)
  );
  AND2_X1 _16951_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[7]),
    .ZN(_01705_)
  );
  OR2_X1 _16952_ (
    .A1(_01704_),
    .A2(_01705_),
    .ZN(_00460_)
  );
  AND2_X1 _16953_ (
    .A1(ex_reg_cause[8]),
    .A2(_01699_),
    .ZN(_01706_)
  );
  AND2_X1 _16954_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[8]),
    .ZN(_01707_)
  );
  OR2_X1 _16955_ (
    .A1(_01706_),
    .A2(_01707_),
    .ZN(_00461_)
  );
  AND2_X1 _16956_ (
    .A1(ex_reg_cause[9]),
    .A2(_01699_),
    .ZN(_01708_)
  );
  AND2_X1 _16957_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[9]),
    .ZN(_01709_)
  );
  OR2_X1 _16958_ (
    .A1(_01708_),
    .A2(_01709_),
    .ZN(_00462_)
  );
  AND2_X1 _16959_ (
    .A1(ex_reg_cause[10]),
    .A2(_01699_),
    .ZN(_01710_)
  );
  AND2_X1 _16960_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[10]),
    .ZN(_01711_)
  );
  OR2_X1 _16961_ (
    .A1(_01710_),
    .A2(_01711_),
    .ZN(_00463_)
  );
  AND2_X1 _16962_ (
    .A1(ex_reg_cause[11]),
    .A2(_01699_),
    .ZN(_01712_)
  );
  AND2_X1 _16963_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[11]),
    .ZN(_01713_)
  );
  OR2_X1 _16964_ (
    .A1(_01712_),
    .A2(_01713_),
    .ZN(_00464_)
  );
  AND2_X1 _16965_ (
    .A1(ex_reg_cause[12]),
    .A2(_01699_),
    .ZN(_01714_)
  );
  AND2_X1 _16966_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[12]),
    .ZN(_01715_)
  );
  OR2_X1 _16967_ (
    .A1(_01714_),
    .A2(_01715_),
    .ZN(_00465_)
  );
  AND2_X1 _16968_ (
    .A1(ex_reg_cause[13]),
    .A2(_01699_),
    .ZN(_01716_)
  );
  AND2_X1 _16969_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[13]),
    .ZN(_01717_)
  );
  OR2_X1 _16970_ (
    .A1(_01716_),
    .A2(_01717_),
    .ZN(_00466_)
  );
  AND2_X1 _16971_ (
    .A1(ex_reg_cause[14]),
    .A2(_01699_),
    .ZN(_01718_)
  );
  AND2_X1 _16972_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[14]),
    .ZN(_01719_)
  );
  OR2_X1 _16973_ (
    .A1(_01718_),
    .A2(_01719_),
    .ZN(_00467_)
  );
  AND2_X1 _16974_ (
    .A1(ex_reg_cause[15]),
    .A2(_01699_),
    .ZN(_01720_)
  );
  AND2_X1 _16975_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[15]),
    .ZN(_01721_)
  );
  OR2_X1 _16976_ (
    .A1(_01720_),
    .A2(_01721_),
    .ZN(_00468_)
  );
  AND2_X1 _16977_ (
    .A1(ex_reg_cause[16]),
    .A2(_01699_),
    .ZN(_01722_)
  );
  AND2_X1 _16978_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[16]),
    .ZN(_01723_)
  );
  OR2_X1 _16979_ (
    .A1(_01722_),
    .A2(_01723_),
    .ZN(_00469_)
  );
  AND2_X1 _16980_ (
    .A1(ex_reg_cause[17]),
    .A2(_01699_),
    .ZN(_01724_)
  );
  AND2_X1 _16981_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[17]),
    .ZN(_01725_)
  );
  OR2_X1 _16982_ (
    .A1(_01724_),
    .A2(_01725_),
    .ZN(_00470_)
  );
  AND2_X1 _16983_ (
    .A1(ex_reg_cause[18]),
    .A2(_01699_),
    .ZN(_01726_)
  );
  AND2_X1 _16984_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[18]),
    .ZN(_01727_)
  );
  OR2_X1 _16985_ (
    .A1(_01726_),
    .A2(_01727_),
    .ZN(_00471_)
  );
  AND2_X1 _16986_ (
    .A1(ex_reg_cause[19]),
    .A2(_01699_),
    .ZN(_01728_)
  );
  AND2_X1 _16987_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[19]),
    .ZN(_01729_)
  );
  OR2_X1 _16988_ (
    .A1(_01728_),
    .A2(_01729_),
    .ZN(_00472_)
  );
  AND2_X1 _16989_ (
    .A1(ex_reg_cause[20]),
    .A2(_01699_),
    .ZN(_01730_)
  );
  AND2_X1 _16990_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[20]),
    .ZN(_01731_)
  );
  OR2_X1 _16991_ (
    .A1(_01730_),
    .A2(_01731_),
    .ZN(_00473_)
  );
  AND2_X1 _16992_ (
    .A1(ex_reg_cause[21]),
    .A2(_01699_),
    .ZN(_01732_)
  );
  AND2_X1 _16993_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[21]),
    .ZN(_01733_)
  );
  OR2_X1 _16994_ (
    .A1(_01732_),
    .A2(_01733_),
    .ZN(_00474_)
  );
  AND2_X1 _16995_ (
    .A1(ex_reg_cause[22]),
    .A2(_01699_),
    .ZN(_01734_)
  );
  AND2_X1 _16996_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[22]),
    .ZN(_01735_)
  );
  OR2_X1 _16997_ (
    .A1(_01734_),
    .A2(_01735_),
    .ZN(_00475_)
  );
  AND2_X1 _16998_ (
    .A1(ex_reg_cause[23]),
    .A2(_01699_),
    .ZN(_01736_)
  );
  AND2_X1 _16999_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[23]),
    .ZN(_01737_)
  );
  OR2_X1 _17000_ (
    .A1(_01736_),
    .A2(_01737_),
    .ZN(_00476_)
  );
  AND2_X1 _17001_ (
    .A1(ex_reg_cause[24]),
    .A2(_01699_),
    .ZN(_01738_)
  );
  AND2_X1 _17002_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[24]),
    .ZN(_01739_)
  );
  OR2_X1 _17003_ (
    .A1(_01738_),
    .A2(_01739_),
    .ZN(_00477_)
  );
  AND2_X1 _17004_ (
    .A1(ex_reg_cause[25]),
    .A2(_01699_),
    .ZN(_01740_)
  );
  AND2_X1 _17005_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[25]),
    .ZN(_01741_)
  );
  OR2_X1 _17006_ (
    .A1(_01740_),
    .A2(_01741_),
    .ZN(_00478_)
  );
  AND2_X1 _17007_ (
    .A1(ex_reg_cause[26]),
    .A2(_01699_),
    .ZN(_01742_)
  );
  AND2_X1 _17008_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[26]),
    .ZN(_01743_)
  );
  OR2_X1 _17009_ (
    .A1(_01742_),
    .A2(_01743_),
    .ZN(_00479_)
  );
  AND2_X1 _17010_ (
    .A1(ex_reg_cause[27]),
    .A2(_01699_),
    .ZN(_01744_)
  );
  AND2_X1 _17011_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[27]),
    .ZN(_01745_)
  );
  OR2_X1 _17012_ (
    .A1(_01744_),
    .A2(_01745_),
    .ZN(_00480_)
  );
  AND2_X1 _17013_ (
    .A1(ex_reg_cause[28]),
    .A2(_01699_),
    .ZN(_01746_)
  );
  AND2_X1 _17014_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[28]),
    .ZN(_01747_)
  );
  OR2_X1 _17015_ (
    .A1(_01746_),
    .A2(_01747_),
    .ZN(_00481_)
  );
  AND2_X1 _17016_ (
    .A1(ex_reg_cause[29]),
    .A2(_01699_),
    .ZN(_01748_)
  );
  AND2_X1 _17017_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[29]),
    .ZN(_01749_)
  );
  OR2_X1 _17018_ (
    .A1(_01748_),
    .A2(_01749_),
    .ZN(_00482_)
  );
  AND2_X1 _17019_ (
    .A1(ex_reg_cause[30]),
    .A2(_01699_),
    .ZN(_01750_)
  );
  AND2_X1 _17020_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[30]),
    .ZN(_01751_)
  );
  OR2_X1 _17021_ (
    .A1(_01750_),
    .A2(_01751_),
    .ZN(_00483_)
  );
  AND2_X1 _17022_ (
    .A1(ex_reg_cause[31]),
    .A2(_01699_),
    .ZN(_01752_)
  );
  AND2_X1 _17023_ (
    .A1(csr_io_interrupt_cause[31]),
    .A2(csr_io_interrupt),
    .ZN(_01753_)
  );
  OR2_X1 _17024_ (
    .A1(_01752_),
    .A2(_01753_),
    .ZN(_00484_)
  );
  MUX2_X1 _17025_ (
    .A(ex_reg_pc[0]),
    .B(bpu_io_pc[0]),
    .S(_01698_),
    .Z(_00485_)
  );
  MUX2_X1 _17026_ (
    .A(ex_reg_pc[1]),
    .B(bpu_io_pc[1]),
    .S(_01698_),
    .Z(_00486_)
  );
  MUX2_X1 _17027_ (
    .A(ex_reg_pc[2]),
    .B(bpu_io_pc[2]),
    .S(_01698_),
    .Z(_00487_)
  );
  MUX2_X1 _17028_ (
    .A(ex_reg_pc[3]),
    .B(bpu_io_pc[3]),
    .S(_01698_),
    .Z(_00488_)
  );
  MUX2_X1 _17029_ (
    .A(ex_reg_pc[4]),
    .B(bpu_io_pc[4]),
    .S(_01698_),
    .Z(_00489_)
  );
  MUX2_X1 _17030_ (
    .A(ex_reg_pc[5]),
    .B(bpu_io_pc[5]),
    .S(_01698_),
    .Z(_00490_)
  );
  MUX2_X1 _17031_ (
    .A(ex_reg_pc[6]),
    .B(bpu_io_pc[6]),
    .S(_01698_),
    .Z(_00491_)
  );
  MUX2_X1 _17032_ (
    .A(ex_reg_pc[7]),
    .B(bpu_io_pc[7]),
    .S(_01698_),
    .Z(_00492_)
  );
  MUX2_X1 _17033_ (
    .A(ex_reg_pc[8]),
    .B(bpu_io_pc[8]),
    .S(_01698_),
    .Z(_00493_)
  );
  MUX2_X1 _17034_ (
    .A(ex_reg_pc[9]),
    .B(bpu_io_pc[9]),
    .S(_01698_),
    .Z(_00494_)
  );
  MUX2_X1 _17035_ (
    .A(ex_reg_pc[10]),
    .B(bpu_io_pc[10]),
    .S(_01698_),
    .Z(_00495_)
  );
  MUX2_X1 _17036_ (
    .A(ex_reg_pc[11]),
    .B(bpu_io_pc[11]),
    .S(_01698_),
    .Z(_00496_)
  );
  MUX2_X1 _17037_ (
    .A(ex_reg_pc[12]),
    .B(bpu_io_pc[12]),
    .S(_01698_),
    .Z(_00497_)
  );
  MUX2_X1 _17038_ (
    .A(ex_reg_pc[13]),
    .B(bpu_io_pc[13]),
    .S(_01698_),
    .Z(_00498_)
  );
  MUX2_X1 _17039_ (
    .A(ex_reg_pc[14]),
    .B(bpu_io_pc[14]),
    .S(_01698_),
    .Z(_00499_)
  );
  MUX2_X1 _17040_ (
    .A(ex_reg_pc[15]),
    .B(bpu_io_pc[15]),
    .S(_01698_),
    .Z(_00500_)
  );
  MUX2_X1 _17041_ (
    .A(ex_reg_pc[16]),
    .B(bpu_io_pc[16]),
    .S(_01698_),
    .Z(_00501_)
  );
  MUX2_X1 _17042_ (
    .A(ex_reg_pc[17]),
    .B(bpu_io_pc[17]),
    .S(_01698_),
    .Z(_00502_)
  );
  MUX2_X1 _17043_ (
    .A(ex_reg_pc[18]),
    .B(bpu_io_pc[18]),
    .S(_01698_),
    .Z(_00503_)
  );
  MUX2_X1 _17044_ (
    .A(ex_reg_pc[19]),
    .B(bpu_io_pc[19]),
    .S(_01698_),
    .Z(_00504_)
  );
  MUX2_X1 _17045_ (
    .A(ex_reg_pc[20]),
    .B(bpu_io_pc[20]),
    .S(_01698_),
    .Z(_00505_)
  );
  MUX2_X1 _17046_ (
    .A(ex_reg_pc[21]),
    .B(bpu_io_pc[21]),
    .S(_01698_),
    .Z(_00506_)
  );
  MUX2_X1 _17047_ (
    .A(ex_reg_pc[22]),
    .B(bpu_io_pc[22]),
    .S(_01698_),
    .Z(_00507_)
  );
  MUX2_X1 _17048_ (
    .A(ex_reg_pc[23]),
    .B(bpu_io_pc[23]),
    .S(_01698_),
    .Z(_00508_)
  );
  MUX2_X1 _17049_ (
    .A(ex_reg_pc[24]),
    .B(bpu_io_pc[24]),
    .S(_01698_),
    .Z(_00509_)
  );
  MUX2_X1 _17050_ (
    .A(ex_reg_pc[25]),
    .B(bpu_io_pc[25]),
    .S(_01698_),
    .Z(_00510_)
  );
  MUX2_X1 _17051_ (
    .A(ex_reg_pc[26]),
    .B(bpu_io_pc[26]),
    .S(_01698_),
    .Z(_00511_)
  );
  MUX2_X1 _17052_ (
    .A(ex_reg_pc[27]),
    .B(bpu_io_pc[27]),
    .S(_01698_),
    .Z(_00512_)
  );
  MUX2_X1 _17053_ (
    .A(ex_reg_pc[28]),
    .B(bpu_io_pc[28]),
    .S(_01698_),
    .Z(_00513_)
  );
  MUX2_X1 _17054_ (
    .A(ex_reg_pc[29]),
    .B(bpu_io_pc[29]),
    .S(_01698_),
    .Z(_00514_)
  );
  MUX2_X1 _17055_ (
    .A(ex_reg_pc[30]),
    .B(bpu_io_pc[30]),
    .S(_01698_),
    .Z(_00515_)
  );
  MUX2_X1 _17056_ (
    .A(ex_reg_pc[31]),
    .B(bpu_io_pc[31]),
    .S(_01698_),
    .Z(_00516_)
  );
  AND2_X1 _17057_ (
    .A1(mem_ctrl_mem),
    .A2(_03933_),
    .ZN(_01754_)
  );
  MUX2_X1 _17058_ (
    .A(_01754_),
    .B(ex_reg_load_use),
    .S(_04041_),
    .Z(_00517_)
  );
  OR2_X1 _17059_ (
    .A1(ex_reg_flush_pipe),
    .A2(_ex_reg_valid_T),
    .ZN(_01755_)
  );
  AND2_X1 _17060_ (
    .A1(csr_io_decode_0_write_flush),
    .A2(_03562_),
    .ZN(_01756_)
  );
  AND2_X1 _17061_ (
    .A1(_03569_),
    .A2(_01756_),
    .ZN(_01757_)
  );
  OR2_X1 _17062_ (
    .A1(_03566_),
    .A2(_01757_),
    .ZN(_01758_)
  );
  OR2_X1 _17063_ (
    .A1(_03882_),
    .A2(_04041_),
    .ZN(_01759_)
  );
  OR2_X1 _17064_ (
    .A1(_01758_),
    .A2(_01759_),
    .ZN(_01760_)
  );
  AND2_X1 _17065_ (
    .A1(_01755_),
    .A2(_01760_),
    .ZN(_00518_)
  );
  MUX2_X1 _17066_ (
    .A(wb_ctrl_fence_i),
    .B(mem_ctrl_fence_i),
    .S(_06433_),
    .Z(_00519_)
  );
  MUX2_X1 _17067_ (
    .A(wb_ctrl_csr[0]),
    .B(mem_ctrl_csr[0]),
    .S(_06433_),
    .Z(_00520_)
  );
  MUX2_X1 _17068_ (
    .A(wb_ctrl_csr[1]),
    .B(mem_ctrl_csr[1]),
    .S(_06433_),
    .Z(_00521_)
  );
  MUX2_X1 _17069_ (
    .A(wb_ctrl_csr[2]),
    .B(mem_ctrl_csr[2]),
    .S(_06433_),
    .Z(_00522_)
  );
  MUX2_X1 _17070_ (
    .A(wb_ctrl_wxd),
    .B(mem_ctrl_wxd),
    .S(_06433_),
    .Z(_00523_)
  );
  MUX2_X1 _17071_ (
    .A(wb_ctrl_div),
    .B(mem_ctrl_div),
    .S(_06433_),
    .Z(_00524_)
  );
  MUX2_X1 _17072_ (
    .A(wb_ctrl_mem),
    .B(mem_ctrl_mem),
    .S(_06433_),
    .Z(_00525_)
  );
  MUX2_X1 _17073_ (
    .A(wb_reg_inst[7]),
    .B(mem_reg_inst[7]),
    .S(_06433_),
    .Z(_00526_)
  );
  MUX2_X1 _17074_ (
    .A(wb_reg_inst[8]),
    .B(mem_reg_inst[8]),
    .S(_06433_),
    .Z(_00527_)
  );
  MUX2_X1 _17075_ (
    .A(wb_reg_inst[9]),
    .B(mem_reg_inst[9]),
    .S(_06433_),
    .Z(_00528_)
  );
  MUX2_X1 _17076_ (
    .A(wb_reg_inst[10]),
    .B(mem_reg_inst[10]),
    .S(_06433_),
    .Z(_00529_)
  );
  MUX2_X1 _17077_ (
    .A(wb_reg_inst[11]),
    .B(mem_reg_inst[11]),
    .S(_06433_),
    .Z(_00530_)
  );
  MUX2_X1 _17078_ (
    .A(wb_reg_inst[16]),
    .B(mem_reg_inst[16]),
    .S(_06433_),
    .Z(_00531_)
  );
  MUX2_X1 _17079_ (
    .A(wb_reg_inst[17]),
    .B(mem_reg_inst[17]),
    .S(_06433_),
    .Z(_00532_)
  );
  MUX2_X1 _17080_ (
    .A(wb_reg_inst[18]),
    .B(mem_reg_inst[18]),
    .S(_06433_),
    .Z(_00533_)
  );
  MUX2_X1 _17081_ (
    .A(wb_reg_inst[19]),
    .B(mem_reg_inst[19]),
    .S(_06433_),
    .Z(_00534_)
  );
  MUX2_X1 _17082_ (
    .A(wb_reg_inst[20]),
    .B(mem_reg_inst[20]),
    .S(_06433_),
    .Z(_00535_)
  );
  MUX2_X1 _17083_ (
    .A(wb_reg_inst[21]),
    .B(mem_reg_inst[21]),
    .S(_06433_),
    .Z(_00536_)
  );
  MUX2_X1 _17084_ (
    .A(wb_reg_inst[22]),
    .B(mem_reg_inst[22]),
    .S(_06433_),
    .Z(_00537_)
  );
  MUX2_X1 _17085_ (
    .A(wb_reg_inst[23]),
    .B(mem_reg_inst[23]),
    .S(_06433_),
    .Z(_00538_)
  );
  MUX2_X1 _17086_ (
    .A(wb_reg_inst[24]),
    .B(mem_reg_inst[24]),
    .S(_06433_),
    .Z(_00539_)
  );
  MUX2_X1 _17087_ (
    .A(wb_reg_inst[25]),
    .B(mem_reg_inst[25]),
    .S(_06433_),
    .Z(_00540_)
  );
  MUX2_X1 _17088_ (
    .A(wb_reg_inst[26]),
    .B(mem_reg_inst[26]),
    .S(_06433_),
    .Z(_00541_)
  );
  MUX2_X1 _17089_ (
    .A(wb_reg_inst[27]),
    .B(mem_reg_inst[27]),
    .S(_06433_),
    .Z(_00542_)
  );
  MUX2_X1 _17090_ (
    .A(wb_reg_inst[28]),
    .B(mem_reg_inst[28]),
    .S(_06433_),
    .Z(_00543_)
  );
  MUX2_X1 _17091_ (
    .A(wb_reg_inst[29]),
    .B(mem_reg_inst[29]),
    .S(_06433_),
    .Z(_00544_)
  );
  MUX2_X1 _17092_ (
    .A(wb_reg_inst[30]),
    .B(mem_reg_inst[30]),
    .S(_06433_),
    .Z(_00545_)
  );
  MUX2_X1 _17093_ (
    .A(wb_reg_inst[31]),
    .B(mem_reg_inst[31]),
    .S(_06433_),
    .Z(_00546_)
  );
  OR2_X1 _17094_ (
    .A1(ex_ctrl_fence_i),
    .A2(_01696_),
    .ZN(_01761_)
  );
  MUX2_X1 _17095_ (
    .A(_01761_),
    .B(mem_ctrl_fence_i),
    .S(_08752_),
    .Z(_00547_)
  );
  MUX2_X1 _17096_ (
    .A(ex_ctrl_csr[0]),
    .B(mem_ctrl_csr[0]),
    .S(_08752_),
    .Z(_00548_)
  );
  MUX2_X1 _17097_ (
    .A(ex_ctrl_csr[1]),
    .B(mem_ctrl_csr[1]),
    .S(_08752_),
    .Z(_00549_)
  );
  MUX2_X1 _17098_ (
    .A(ex_ctrl_csr[2]),
    .B(mem_ctrl_csr[2]),
    .S(_08752_),
    .Z(_00550_)
  );
  MUX2_X1 _17099_ (
    .A(ex_ctrl_wxd),
    .B(mem_ctrl_wxd),
    .S(_08752_),
    .Z(_00551_)
  );
  MUX2_X1 _17100_ (
    .A(ex_ctrl_div),
    .B(mem_ctrl_div),
    .S(_08752_),
    .Z(_00552_)
  );
  MUX2_X1 _17101_ (
    .A(ex_ctrl_mem),
    .B(mem_ctrl_mem),
    .S(_08752_),
    .Z(_00553_)
  );
  MUX2_X1 _17102_ (
    .A(ex_ctrl_jalr),
    .B(mem_ctrl_jalr),
    .S(_08752_),
    .Z(_00554_)
  );
  MUX2_X1 _17103_ (
    .A(ex_ctrl_jal),
    .B(mem_ctrl_jal),
    .S(_08752_),
    .Z(_00555_)
  );
  MUX2_X1 _17104_ (
    .A(ex_ctrl_branch),
    .B(mem_ctrl_branch),
    .S(_08752_),
    .Z(_00556_)
  );
  MUX2_X1 _17105_ (
    .A(_03541_),
    .B(ex_ctrl_csr[1]),
    .S(_04146_),
    .Z(_00557_)
  );
  MUX2_X1 _17106_ (
    .A(_03882_),
    .B(ex_ctrl_fence_i),
    .S(_04041_),
    .Z(_00558_)
  );
  MUX2_X1 _17107_ (
    .A(_03601_),
    .B(ex_ctrl_wxd),
    .S(_04146_),
    .Z(_00559_)
  );
  MUX2_X1 _17108_ (
    .A(_03574_),
    .B(ex_ctrl_div),
    .S(_04146_),
    .Z(_00560_)
  );
  AND2_X1 _17109_ (
    .A1(_03414_),
    .A2(_03426_),
    .ZN(_01762_)
  );
  AND2_X1 _17110_ (
    .A1(csr_io_decode_0_inst[29]),
    .A2(_03386_),
    .ZN(_01763_)
  );
  AND2_X1 _17111_ (
    .A1(_03036_),
    .A2(_03800_),
    .ZN(_01764_)
  );
  OR2_X1 _17112_ (
    .A1(_01763_),
    .A2(_01764_),
    .ZN(_01765_)
  );
  OR2_X1 _17113_ (
    .A1(_01762_),
    .A2(_01765_),
    .ZN(_01766_)
  );
  MUX2_X1 _17114_ (
    .A(_01766_),
    .B(ex_ctrl_mem_cmd[0]),
    .S(_04041_),
    .Z(_00561_)
  );
  AND2_X1 _17115_ (
    .A1(csr_io_decode_0_inst[30]),
    .A2(_03386_),
    .ZN(_01767_)
  );
  OR2_X1 _17116_ (
    .A1(_03425_),
    .A2(_01762_),
    .ZN(_01768_)
  );
  OR2_X1 _17117_ (
    .A1(_01767_),
    .A2(_01768_),
    .ZN(_01769_)
  );
  MUX2_X1 _17118_ (
    .A(_01769_),
    .B(ex_ctrl_mem_cmd[1]),
    .S(_04041_),
    .Z(_00562_)
  );
  AND2_X1 _17119_ (
    .A1(csr_io_decode_0_inst[31]),
    .A2(_03386_),
    .ZN(_01770_)
  );
  OR2_X1 _17120_ (
    .A1(_03428_),
    .A2(_01770_),
    .ZN(_01771_)
  );
  MUX2_X1 _17121_ (
    .A(_01771_),
    .B(ex_ctrl_mem_cmd[2]),
    .S(_04041_),
    .Z(_00563_)
  );
  MUX2_X1 _17122_ (
    .A(_03386_),
    .B(ex_ctrl_mem_cmd[3]),
    .S(_04041_),
    .Z(_00564_)
  );
  OR2_X1 _17123_ (
    .A1(csr_io_decode_0_inst[14]),
    .A2(csr_io_decode_0_inst[25]),
    .ZN(_01772_)
  );
  INV_X1 _17124_ (
    .A(_01772_),
    .ZN(_01773_)
  );
  AND2_X1 _17125_ (
    .A1(_03432_),
    .A2(_01772_),
    .ZN(_01774_)
  );
  OR2_X1 _17126_ (
    .A1(_03368_),
    .A2(_01774_),
    .ZN(_01775_)
  );
  AND2_X1 _17127_ (
    .A1(csr_io_decode_0_inst[12]),
    .A2(_01775_),
    .ZN(_01776_)
  );
  AND2_X1 _17128_ (
    .A1(_03365_),
    .A2(_03524_),
    .ZN(_01777_)
  );
  OR2_X1 _17129_ (
    .A1(_03599_),
    .A2(_01777_),
    .ZN(_01778_)
  );
  OR2_X1 _17130_ (
    .A1(_01776_),
    .A2(_01778_),
    .ZN(_01779_)
  );
  AND2_X1 _17131_ (
    .A1(_03038_),
    .A2(_03349_),
    .ZN(_01780_)
  );
  AND2_X1 _17132_ (
    .A1(_03591_),
    .A2(_01780_),
    .ZN(_01781_)
  );
  OR2_X1 _17133_ (
    .A1(_01779_),
    .A2(_01781_),
    .ZN(_01782_)
  );
  AND2_X1 _17134_ (
    .A1(_03066_),
    .A2(_03067_),
    .ZN(_01783_)
  );
  OR2_X1 _17135_ (
    .A1(ibuf_io_inst_0_bits_xcpt0_ae_inst),
    .A2(bpu_io_xcpt_if),
    .ZN(_01784_)
  );
  AND2_X1 _17136_ (
    .A1(_08716_),
    .A2(_01783_),
    .ZN(_01785_)
  );
  INV_X1 _17137_ (
    .A(_01785_),
    .ZN(_01786_)
  );
  OR2_X1 _17138_ (
    .A1(csr_io_interrupt),
    .A2(bpu_io_debug_if),
    .ZN(_01787_)
  );
  OR2_X1 _17139_ (
    .A1(_03582_),
    .A2(_01787_),
    .ZN(_01788_)
  );
  INV_X1 _17140_ (
    .A(_01788_),
    .ZN(_01789_)
  );
  AND2_X1 _17141_ (
    .A1(_01785_),
    .A2(_01789_),
    .ZN(_01790_)
  );
  AND2_X1 _17142_ (
    .A1(_01782_),
    .A2(_01790_),
    .ZN(_01791_)
  );
  MUX2_X1 _17143_ (
    .A(_01791_),
    .B(ex_ctrl_alu_fn[0]),
    .S(_04041_),
    .Z(_00565_)
  );
  OR2_X1 _17144_ (
    .A1(csr_io_decode_0_inst[25]),
    .A2(_03331_),
    .ZN(_01792_)
  );
  AND2_X1 _17145_ (
    .A1(csr_io_decode_0_inst[13]),
    .A2(_01792_),
    .ZN(_01793_)
  );
  AND2_X1 _17146_ (
    .A1(csr_io_decode_0_inst[4]),
    .A2(_03321_),
    .ZN(_01794_)
  );
  AND2_X1 _17147_ (
    .A1(_03592_),
    .A2(_01794_),
    .ZN(_01795_)
  );
  OR2_X1 _17148_ (
    .A1(_03432_),
    .A2(_01795_),
    .ZN(_01796_)
  );
  AND2_X1 _17149_ (
    .A1(_01793_),
    .A2(_01796_),
    .ZN(_01797_)
  );
  OR2_X1 _17150_ (
    .A1(_03327_),
    .A2(_03591_),
    .ZN(_01798_)
  );
  AND2_X1 _17151_ (
    .A1(_03366_),
    .A2(_01798_),
    .ZN(_01799_)
  );
  AND2_X1 _17152_ (
    .A1(_03352_),
    .A2(_01773_),
    .ZN(_01800_)
  );
  AND2_X1 _17153_ (
    .A1(_03322_),
    .A2(_01800_),
    .ZN(_01801_)
  );
  AND2_X1 _17154_ (
    .A1(_03431_),
    .A2(_01801_),
    .ZN(_01802_)
  );
  OR2_X1 _17155_ (
    .A1(_03370_),
    .A2(_01802_),
    .ZN(_01803_)
  );
  AND2_X1 _17156_ (
    .A1(csr_io_decode_0_inst[30]),
    .A2(_03359_),
    .ZN(_01804_)
  );
  AND2_X1 _17157_ (
    .A1(_01803_),
    .A2(_01804_),
    .ZN(_01805_)
  );
  OR2_X1 _17158_ (
    .A1(_01799_),
    .A2(_01805_),
    .ZN(_01806_)
  );
  OR2_X1 _17159_ (
    .A1(_01797_),
    .A2(_01806_),
    .ZN(_01807_)
  );
  AND2_X1 _17160_ (
    .A1(_01790_),
    .A2(_01807_),
    .ZN(_01808_)
  );
  MUX2_X1 _17161_ (
    .A(_01808_),
    .B(ex_ctrl_alu_fn[1]),
    .S(_04041_),
    .Z(_00566_)
  );
  AND2_X1 _17162_ (
    .A1(_03378_),
    .A2(_03401_),
    .ZN(_01809_)
  );
  OR2_X1 _17163_ (
    .A1(_03362_),
    .A2(_01809_),
    .ZN(_01810_)
  );
  AND2_X1 _17164_ (
    .A1(csr_io_decode_0_inst[14]),
    .A2(_01810_),
    .ZN(_01811_)
  );
  AND2_X1 _17165_ (
    .A1(csr_io_decode_0_inst[13]),
    .A2(_03004_),
    .ZN(_01812_)
  );
  OR2_X1 _17166_ (
    .A1(csr_io_decode_0_inst[14]),
    .A2(_01812_),
    .ZN(_01813_)
  );
  AND2_X1 _17167_ (
    .A1(_03432_),
    .A2(_01813_),
    .ZN(_01814_)
  );
  OR2_X1 _17168_ (
    .A1(_03368_),
    .A2(_03379_),
    .ZN(_01815_)
  );
  OR2_X1 _17169_ (
    .A1(_01814_),
    .A2(_01815_),
    .ZN(_01816_)
  );
  OR2_X1 _17170_ (
    .A1(_01811_),
    .A2(_01816_),
    .ZN(_01817_)
  );
  AND2_X1 _17171_ (
    .A1(_01790_),
    .A2(_01817_),
    .ZN(_01818_)
  );
  MUX2_X1 _17172_ (
    .A(_01818_),
    .B(ex_ctrl_alu_fn[2]),
    .S(_04041_),
    .Z(_00567_)
  );
  AND2_X1 _17173_ (
    .A1(_03388_),
    .A2(_01794_),
    .ZN(_01819_)
  );
  AND2_X1 _17174_ (
    .A1(_03377_),
    .A2(_01800_),
    .ZN(_01820_)
  );
  AND2_X1 _17175_ (
    .A1(_03430_),
    .A2(_01820_),
    .ZN(_01821_)
  );
  AND2_X1 _17176_ (
    .A1(_03360_),
    .A2(_01821_),
    .ZN(_01822_)
  );
  OR2_X1 _17177_ (
    .A1(_03368_),
    .A2(_01822_),
    .ZN(_01823_)
  );
  OR2_X1 _17178_ (
    .A1(_01819_),
    .A2(_01823_),
    .ZN(_01824_)
  );
  OR2_X1 _17179_ (
    .A1(_01805_),
    .A2(_01824_),
    .ZN(_01825_)
  );
  AND2_X1 _17180_ (
    .A1(_01790_),
    .A2(_01825_),
    .ZN(_01826_)
  );
  MUX2_X1 _17181_ (
    .A(_01826_),
    .B(ex_ctrl_alu_fn[3]),
    .S(_04041_),
    .Z(_00568_)
  );
  MUX2_X1 _17182_ (
    .A(_03888_),
    .B(ex_ctrl_mem),
    .S(_04041_),
    .Z(_00569_)
  );
  AND2_X1 _17183_ (
    .A1(_03323_),
    .A2(_03367_),
    .ZN(_01827_)
  );
  OR2_X1 _17184_ (
    .A1(_03343_),
    .A2(_01827_),
    .ZN(_01828_)
  );
  AND2_X1 _17185_ (
    .A1(_03319_),
    .A2(_01828_),
    .ZN(_01829_)
  );
  OR2_X1 _17186_ (
    .A1(_03544_),
    .A2(_01829_),
    .ZN(_01830_)
  );
  MUX2_X1 _17187_ (
    .A(_01830_),
    .B(ex_ctrl_sel_imm[0]),
    .S(_04146_),
    .Z(_00570_)
  );
  OR2_X1 _17188_ (
    .A1(_03493_),
    .A2(_03544_),
    .ZN(_01831_)
  );
  MUX2_X1 _17189_ (
    .A(_01831_),
    .B(ex_ctrl_sel_imm[1]),
    .S(_04146_),
    .Z(_00571_)
  );
  AND2_X1 _17190_ (
    .A1(_03347_),
    .A2(_01827_),
    .ZN(_01832_)
  );
  OR2_X1 _17191_ (
    .A1(_03590_),
    .A2(_01832_),
    .ZN(_01833_)
  );
  AND2_X1 _17192_ (
    .A1(_03038_),
    .A2(_03599_),
    .ZN(_01834_)
  );
  OR2_X1 _17193_ (
    .A1(_01833_),
    .A2(_01834_),
    .ZN(_01835_)
  );
  OR2_X1 _17194_ (
    .A1(_03379_),
    .A2(_01835_),
    .ZN(_01836_)
  );
  OR2_X1 _17195_ (
    .A1(_03595_),
    .A2(_01836_),
    .ZN(_01837_)
  );
  MUX2_X1 _17196_ (
    .A(_01837_),
    .B(ex_ctrl_sel_imm[2]),
    .S(_04146_),
    .Z(_00572_)
  );
  OR2_X1 _17197_ (
    .A1(_03447_),
    .A2(_01788_),
    .ZN(_01838_)
  );
  AND2_X1 _17198_ (
    .A1(_01785_),
    .A2(_01838_),
    .ZN(_01839_)
  );
  MUX2_X1 _17199_ (
    .A(_01839_),
    .B(ex_ctrl_sel_alu1[0]),
    .S(_04146_),
    .Z(_00573_)
  );
  AND2_X1 _17200_ (
    .A1(_03038_),
    .A2(_03493_),
    .ZN(_01840_)
  );
  OR2_X1 _17201_ (
    .A1(_03543_),
    .A2(_01840_),
    .ZN(_01841_)
  );
  AND2_X1 _17202_ (
    .A1(_01789_),
    .A2(_01841_),
    .ZN(_01842_)
  );
  OR2_X1 _17203_ (
    .A1(_01786_),
    .A2(_01842_),
    .ZN(_01843_)
  );
  MUX2_X1 _17204_ (
    .A(_01843_),
    .B(ex_ctrl_sel_alu1[1]),
    .S(_04146_),
    .Z(_00574_)
  );
  OR2_X1 _17205_ (
    .A1(_03340_),
    .A2(_01831_),
    .ZN(_01844_)
  );
  OR2_X1 _17206_ (
    .A1(_01836_),
    .A2(_01844_),
    .ZN(_01845_)
  );
  AND2_X1 _17207_ (
    .A1(_01789_),
    .A2(_01845_),
    .ZN(_01846_)
  );
  OR2_X1 _17208_ (
    .A1(_08715_),
    .A2(_01846_),
    .ZN(_01847_)
  );
  AND2_X1 _17209_ (
    .A1(_01783_),
    .A2(_01847_),
    .ZN(_01848_)
  );
  MUX2_X1 _17210_ (
    .A(_01848_),
    .B(ex_ctrl_sel_alu2[0]),
    .S(_04146_),
    .Z(_00575_)
  );
  MUX2_X1 _17211_ (
    .A(_03806_),
    .B(ex_ctrl_rxs2),
    .S(_04146_),
    .Z(_00576_)
  );
  MUX2_X1 _17212_ (
    .A(_03590_),
    .B(ex_ctrl_jalr),
    .S(_04146_),
    .Z(_00577_)
  );
  MUX2_X1 _17213_ (
    .A(_03544_),
    .B(ex_ctrl_jal),
    .S(_04146_),
    .Z(_00578_)
  );
  AND2_X1 _17214_ (
    .A1(_03366_),
    .A2(_03389_),
    .ZN(_01849_)
  );
  MUX2_X1 _17215_ (
    .A(_01849_),
    .B(ex_ctrl_branch),
    .S(_04146_),
    .Z(_00579_)
  );
  OR2_X1 _17216_ (
    .A1(_03910_),
    .A2(_06338_),
    .ZN(_01850_)
  );
  OR2_X1 _17217_ (
    .A1(_06424_),
    .A2(_01850_),
    .ZN(_01851_)
  );
  AND2_X1 _17218_ (
    .A1(_03811_),
    .A2(_01851_),
    .ZN(_01852_)
  );
  OR2_X1 _17219_ (
    .A1(\rf[26] [0]),
    .A2(_03050_),
    .ZN(_01853_)
  );
  OR2_X1 _17220_ (
    .A1(\rf[30] [0]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_01854_)
  );
  AND2_X1 _17221_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_01854_),
    .ZN(_01855_)
  );
  AND2_X1 _17222_ (
    .A1(_01853_),
    .A2(_01855_),
    .ZN(_01856_)
  );
  AND2_X1 _17223_ (
    .A1(\rf[27] [0]),
    .A2(_03817_),
    .ZN(_01857_)
  );
  OR2_X1 _17224_ (
    .A1(_01856_),
    .A2(_01857_),
    .ZN(_01858_)
  );
  MUX2_X1 _17225_ (
    .A(\rf[13] [0]),
    .B(\rf[9] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_01859_)
  );
  OR2_X1 _17226_ (
    .A1(\rf[8] [0]),
    .A2(_03050_),
    .ZN(_01860_)
  );
  OR2_X1 _17227_ (
    .A1(\rf[12] [0]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_01861_)
  );
  MUX2_X1 _17228_ (
    .A(\rf[15] [0]),
    .B(\rf[11] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_01862_)
  );
  OR2_X1 _17229_ (
    .A1(\rf[14] [0]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_01863_)
  );
  OR2_X1 _17230_ (
    .A1(\rf[10] [0]),
    .A2(_03050_),
    .ZN(_01864_)
  );
  MUX2_X1 _17231_ (
    .A(\rf[29] [0]),
    .B(\rf[25] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_01865_)
  );
  AND2_X1 _17232_ (
    .A1(_03048_),
    .A2(_01865_),
    .ZN(_01866_)
  );
  OR2_X1 _17233_ (
    .A1(\rf[28] [0]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_01867_)
  );
  OR2_X1 _17234_ (
    .A1(\rf[24] [0]),
    .A2(_03050_),
    .ZN(_01868_)
  );
  AND2_X1 _17235_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_01868_),
    .ZN(_01869_)
  );
  AND2_X1 _17236_ (
    .A1(_01867_),
    .A2(_01869_),
    .ZN(_01870_)
  );
  OR2_X1 _17237_ (
    .A1(_03049_),
    .A2(_01870_),
    .ZN(_01871_)
  );
  OR2_X1 _17238_ (
    .A1(_01866_),
    .A2(_01871_),
    .ZN(_01872_)
  );
  OR2_X1 _17239_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_01858_),
    .ZN(_01873_)
  );
  AND2_X1 _17240_ (
    .A1(_03051_),
    .A2(_01873_),
    .ZN(_01874_)
  );
  AND2_X1 _17241_ (
    .A1(_01872_),
    .A2(_01874_),
    .ZN(_01875_)
  );
  MUX2_X1 _17242_ (
    .A(\rf[21] [0]),
    .B(\rf[17] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_01876_)
  );
  AND2_X1 _17243_ (
    .A1(_03048_),
    .A2(_01876_),
    .ZN(_01877_)
  );
  OR2_X1 _17244_ (
    .A1(\rf[20] [0]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_01878_)
  );
  OR2_X1 _17245_ (
    .A1(\rf[16] [0]),
    .A2(_03050_),
    .ZN(_01879_)
  );
  AND2_X1 _17246_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_01878_),
    .ZN(_01880_)
  );
  AND2_X1 _17247_ (
    .A1(_01879_),
    .A2(_01880_),
    .ZN(_01881_)
  );
  OR2_X1 _17248_ (
    .A1(_03049_),
    .A2(_01877_),
    .ZN(_01882_)
  );
  OR2_X1 _17249_ (
    .A1(_01881_),
    .A2(_01882_),
    .ZN(_01883_)
  );
  OR2_X1 _17250_ (
    .A1(\rf[18] [0]),
    .A2(_03050_),
    .ZN(_01884_)
  );
  OR2_X1 _17251_ (
    .A1(\rf[22] [0]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_01885_)
  );
  AND2_X1 _17252_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_01885_),
    .ZN(_01886_)
  );
  AND2_X1 _17253_ (
    .A1(_01884_),
    .A2(_01886_),
    .ZN(_01887_)
  );
  MUX2_X1 _17254_ (
    .A(\rf[23] [0]),
    .B(\rf[19] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_01888_)
  );
  AND2_X1 _17255_ (
    .A1(_03048_),
    .A2(_01888_),
    .ZN(_01889_)
  );
  OR2_X1 _17256_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_01889_),
    .ZN(_01890_)
  );
  OR2_X1 _17257_ (
    .A1(_01887_),
    .A2(_01890_),
    .ZN(_01891_)
  );
  AND2_X1 _17258_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_01891_),
    .ZN(_01892_)
  );
  AND2_X1 _17259_ (
    .A1(_01883_),
    .A2(_01892_),
    .ZN(_01893_)
  );
  OR2_X1 _17260_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[4]),
    .A2(_01893_),
    .ZN(_01894_)
  );
  OR2_X1 _17261_ (
    .A1(_01875_),
    .A2(_01894_),
    .ZN(_01895_)
  );
  AND2_X1 _17262_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_01863_),
    .ZN(_01896_)
  );
  AND2_X1 _17263_ (
    .A1(_01864_),
    .A2(_01896_),
    .ZN(_01897_)
  );
  AND2_X1 _17264_ (
    .A1(_03048_),
    .A2(_01862_),
    .ZN(_01898_)
  );
  OR2_X1 _17265_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_01898_),
    .ZN(_01899_)
  );
  OR2_X1 _17266_ (
    .A1(_01897_),
    .A2(_01899_),
    .ZN(_01900_)
  );
  AND2_X1 _17267_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_01861_),
    .ZN(_01901_)
  );
  AND2_X1 _17268_ (
    .A1(_01860_),
    .A2(_01901_),
    .ZN(_01902_)
  );
  AND2_X1 _17269_ (
    .A1(_03048_),
    .A2(_01859_),
    .ZN(_01903_)
  );
  OR2_X1 _17270_ (
    .A1(_03049_),
    .A2(_01903_),
    .ZN(_01904_)
  );
  OR2_X1 _17271_ (
    .A1(_01902_),
    .A2(_01904_),
    .ZN(_01905_)
  );
  AND2_X1 _17272_ (
    .A1(_03051_),
    .A2(_01905_),
    .ZN(_01906_)
  );
  AND2_X1 _17273_ (
    .A1(_01900_),
    .A2(_01906_),
    .ZN(_01907_)
  );
  OR2_X1 _17274_ (
    .A1(\rf[0] [0]),
    .A2(_03050_),
    .ZN(_01908_)
  );
  OR2_X1 _17275_ (
    .A1(\rf[4] [0]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_01909_)
  );
  AND2_X1 _17276_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_01909_),
    .ZN(_01910_)
  );
  AND2_X1 _17277_ (
    .A1(_01908_),
    .A2(_01910_),
    .ZN(_01911_)
  );
  MUX2_X1 _17278_ (
    .A(\rf[5] [0]),
    .B(\rf[1] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_01912_)
  );
  AND2_X1 _17279_ (
    .A1(_03048_),
    .A2(_01912_),
    .ZN(_01913_)
  );
  OR2_X1 _17280_ (
    .A1(_03049_),
    .A2(_01913_),
    .ZN(_01914_)
  );
  OR2_X1 _17281_ (
    .A1(_01911_),
    .A2(_01914_),
    .ZN(_01915_)
  );
  MUX2_X1 _17282_ (
    .A(\rf[7] [0]),
    .B(\rf[3] [0]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_01916_)
  );
  AND2_X1 _17283_ (
    .A1(_03048_),
    .A2(_01916_),
    .ZN(_01917_)
  );
  OR2_X1 _17284_ (
    .A1(\rf[2] [0]),
    .A2(_03050_),
    .ZN(_01918_)
  );
  OR2_X1 _17285_ (
    .A1(\rf[6] [0]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_01919_)
  );
  AND2_X1 _17286_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_01919_),
    .ZN(_01920_)
  );
  AND2_X1 _17287_ (
    .A1(_01918_),
    .A2(_01920_),
    .ZN(_01921_)
  );
  OR2_X1 _17288_ (
    .A1(_01917_),
    .A2(_01921_),
    .ZN(_01922_)
  );
  OR2_X1 _17289_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_01922_),
    .ZN(_01923_)
  );
  AND2_X1 _17290_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_01915_),
    .ZN(_01924_)
  );
  AND2_X1 _17291_ (
    .A1(_01923_),
    .A2(_01924_),
    .ZN(_01925_)
  );
  OR2_X1 _17292_ (
    .A1(_03064_),
    .A2(_01907_),
    .ZN(_01926_)
  );
  OR2_X1 _17293_ (
    .A1(_01925_),
    .A2(_01926_),
    .ZN(_01927_)
  );
  AND2_X1 _17294_ (
    .A1(_01895_),
    .A2(_01927_),
    .ZN(_01928_)
  );
  AND2_X1 _17295_ (
    .A1(_06266_),
    .A2(_06791_),
    .ZN(_01929_)
  );
  AND2_X1 _17296_ (
    .A1(_06792_),
    .A2(_01928_),
    .ZN(_01930_)
  );
  OR2_X1 _17297_ (
    .A1(_06779_),
    .A2(_01929_),
    .ZN(_01931_)
  );
  OR2_X1 _17298_ (
    .A1(_01930_),
    .A2(_01931_),
    .ZN(_01932_)
  );
  AND2_X1 _17299_ (
    .A1(_01852_),
    .A2(_01932_),
    .ZN(_01933_)
  );
  MUX2_X1 _17300_ (
    .A(_01933_),
    .B(ex_reg_rs_lsb_1[0]),
    .S(_04146_),
    .Z(_00580_)
  );
  OR2_X1 _17301_ (
    .A1(\rf[26] [1]),
    .A2(_03050_),
    .ZN(_01934_)
  );
  OR2_X1 _17302_ (
    .A1(\rf[30] [1]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_01935_)
  );
  AND2_X1 _17303_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_01935_),
    .ZN(_01936_)
  );
  AND2_X1 _17304_ (
    .A1(_01934_),
    .A2(_01936_),
    .ZN(_01937_)
  );
  AND2_X1 _17305_ (
    .A1(\rf[27] [1]),
    .A2(_03817_),
    .ZN(_01938_)
  );
  OR2_X1 _17306_ (
    .A1(_01937_),
    .A2(_01938_),
    .ZN(_01939_)
  );
  MUX2_X1 _17307_ (
    .A(\rf[13] [1]),
    .B(\rf[9] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_01940_)
  );
  OR2_X1 _17308_ (
    .A1(\rf[8] [1]),
    .A2(_03050_),
    .ZN(_01941_)
  );
  OR2_X1 _17309_ (
    .A1(\rf[12] [1]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_01942_)
  );
  MUX2_X1 _17310_ (
    .A(\rf[15] [1]),
    .B(\rf[11] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_01943_)
  );
  OR2_X1 _17311_ (
    .A1(\rf[14] [1]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_01944_)
  );
  OR2_X1 _17312_ (
    .A1(\rf[10] [1]),
    .A2(_03050_),
    .ZN(_01945_)
  );
  MUX2_X1 _17313_ (
    .A(\rf[29] [1]),
    .B(\rf[25] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_01946_)
  );
  AND2_X1 _17314_ (
    .A1(_03048_),
    .A2(_01946_),
    .ZN(_01947_)
  );
  OR2_X1 _17315_ (
    .A1(\rf[28] [1]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_01948_)
  );
  OR2_X1 _17316_ (
    .A1(\rf[24] [1]),
    .A2(_03050_),
    .ZN(_01949_)
  );
  AND2_X1 _17317_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_01949_),
    .ZN(_01950_)
  );
  AND2_X1 _17318_ (
    .A1(_01948_),
    .A2(_01950_),
    .ZN(_01951_)
  );
  OR2_X1 _17319_ (
    .A1(_03049_),
    .A2(_01951_),
    .ZN(_01952_)
  );
  OR2_X1 _17320_ (
    .A1(_01947_),
    .A2(_01952_),
    .ZN(_01953_)
  );
  OR2_X1 _17321_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_01939_),
    .ZN(_01954_)
  );
  AND2_X1 _17322_ (
    .A1(_03051_),
    .A2(_01954_),
    .ZN(_01955_)
  );
  AND2_X1 _17323_ (
    .A1(_01953_),
    .A2(_01955_),
    .ZN(_01956_)
  );
  MUX2_X1 _17324_ (
    .A(\rf[21] [1]),
    .B(\rf[17] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_01957_)
  );
  AND2_X1 _17325_ (
    .A1(_03048_),
    .A2(_01957_),
    .ZN(_01958_)
  );
  OR2_X1 _17326_ (
    .A1(\rf[20] [1]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_01959_)
  );
  OR2_X1 _17327_ (
    .A1(\rf[16] [1]),
    .A2(_03050_),
    .ZN(_01960_)
  );
  AND2_X1 _17328_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_01959_),
    .ZN(_01961_)
  );
  AND2_X1 _17329_ (
    .A1(_01960_),
    .A2(_01961_),
    .ZN(_01962_)
  );
  OR2_X1 _17330_ (
    .A1(_03049_),
    .A2(_01958_),
    .ZN(_01963_)
  );
  OR2_X1 _17331_ (
    .A1(_01962_),
    .A2(_01963_),
    .ZN(_01964_)
  );
  OR2_X1 _17332_ (
    .A1(\rf[18] [1]),
    .A2(_03050_),
    .ZN(_01965_)
  );
  OR2_X1 _17333_ (
    .A1(\rf[22] [1]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_01966_)
  );
  AND2_X1 _17334_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_01966_),
    .ZN(_01967_)
  );
  AND2_X1 _17335_ (
    .A1(_01965_),
    .A2(_01967_),
    .ZN(_01968_)
  );
  MUX2_X1 _17336_ (
    .A(\rf[23] [1]),
    .B(\rf[19] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_01969_)
  );
  AND2_X1 _17337_ (
    .A1(_03048_),
    .A2(_01969_),
    .ZN(_01970_)
  );
  OR2_X1 _17338_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_01970_),
    .ZN(_01971_)
  );
  OR2_X1 _17339_ (
    .A1(_01968_),
    .A2(_01971_),
    .ZN(_01972_)
  );
  AND2_X1 _17340_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_01972_),
    .ZN(_01973_)
  );
  AND2_X1 _17341_ (
    .A1(_01964_),
    .A2(_01973_),
    .ZN(_01974_)
  );
  OR2_X1 _17342_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[4]),
    .A2(_01974_),
    .ZN(_01975_)
  );
  OR2_X1 _17343_ (
    .A1(_01956_),
    .A2(_01975_),
    .ZN(_01976_)
  );
  AND2_X1 _17344_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_01944_),
    .ZN(_01977_)
  );
  AND2_X1 _17345_ (
    .A1(_01945_),
    .A2(_01977_),
    .ZN(_01978_)
  );
  AND2_X1 _17346_ (
    .A1(_03048_),
    .A2(_01943_),
    .ZN(_01979_)
  );
  OR2_X1 _17347_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_01979_),
    .ZN(_01980_)
  );
  OR2_X1 _17348_ (
    .A1(_01978_),
    .A2(_01980_),
    .ZN(_01981_)
  );
  AND2_X1 _17349_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_01942_),
    .ZN(_01982_)
  );
  AND2_X1 _17350_ (
    .A1(_01941_),
    .A2(_01982_),
    .ZN(_01983_)
  );
  AND2_X1 _17351_ (
    .A1(_03048_),
    .A2(_01940_),
    .ZN(_01984_)
  );
  OR2_X1 _17352_ (
    .A1(_03049_),
    .A2(_01984_),
    .ZN(_01985_)
  );
  OR2_X1 _17353_ (
    .A1(_01983_),
    .A2(_01985_),
    .ZN(_01986_)
  );
  AND2_X1 _17354_ (
    .A1(_03051_),
    .A2(_01986_),
    .ZN(_01987_)
  );
  AND2_X1 _17355_ (
    .A1(_01981_),
    .A2(_01987_),
    .ZN(_01988_)
  );
  OR2_X1 _17356_ (
    .A1(\rf[0] [1]),
    .A2(_03050_),
    .ZN(_01989_)
  );
  OR2_X1 _17357_ (
    .A1(\rf[4] [1]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_01990_)
  );
  AND2_X1 _17358_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_01990_),
    .ZN(_01991_)
  );
  AND2_X1 _17359_ (
    .A1(_01989_),
    .A2(_01991_),
    .ZN(_01992_)
  );
  MUX2_X1 _17360_ (
    .A(\rf[5] [1]),
    .B(\rf[1] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_01993_)
  );
  AND2_X1 _17361_ (
    .A1(_03048_),
    .A2(_01993_),
    .ZN(_01994_)
  );
  OR2_X1 _17362_ (
    .A1(_03049_),
    .A2(_01994_),
    .ZN(_01995_)
  );
  OR2_X1 _17363_ (
    .A1(_01992_),
    .A2(_01995_),
    .ZN(_01996_)
  );
  MUX2_X1 _17364_ (
    .A(\rf[7] [1]),
    .B(\rf[3] [1]),
    .S(ibuf_io_inst_0_bits_inst_rs2[2]),
    .Z(_01997_)
  );
  AND2_X1 _17365_ (
    .A1(_03048_),
    .A2(_01997_),
    .ZN(_01998_)
  );
  OR2_X1 _17366_ (
    .A1(\rf[2] [1]),
    .A2(_03050_),
    .ZN(_01999_)
  );
  OR2_X1 _17367_ (
    .A1(\rf[6] [1]),
    .A2(ibuf_io_inst_0_bits_inst_rs2[2]),
    .ZN(_02000_)
  );
  AND2_X1 _17368_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[0]),
    .A2(_02000_),
    .ZN(_02001_)
  );
  AND2_X1 _17369_ (
    .A1(_01999_),
    .A2(_02001_),
    .ZN(_02002_)
  );
  OR2_X1 _17370_ (
    .A1(_01998_),
    .A2(_02002_),
    .ZN(_02003_)
  );
  OR2_X1 _17371_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[1]),
    .A2(_02003_),
    .ZN(_02004_)
  );
  AND2_X1 _17372_ (
    .A1(ibuf_io_inst_0_bits_inst_rs2[3]),
    .A2(_01996_),
    .ZN(_02005_)
  );
  AND2_X1 _17373_ (
    .A1(_02004_),
    .A2(_02005_),
    .ZN(_02006_)
  );
  OR2_X1 _17374_ (
    .A1(_03064_),
    .A2(_01988_),
    .ZN(_02007_)
  );
  OR2_X1 _17375_ (
    .A1(_02006_),
    .A2(_02007_),
    .ZN(_02008_)
  );
  AND2_X1 _17376_ (
    .A1(_01976_),
    .A2(_02008_),
    .ZN(_02009_)
  );
  MUX2_X1 _17377_ (
    .A(_02009_),
    .B(_06420_),
    .S(_06791_),
    .Z(_02010_)
  );
  OR2_X1 _17378_ (
    .A1(_06779_),
    .A2(_02010_),
    .ZN(_02011_)
  );
  AND2_X1 _17379_ (
    .A1(_06426_),
    .A2(_02011_),
    .ZN(_02012_)
  );
  MUX2_X1 _17380_ (
    .A(_02012_),
    .B(ex_reg_rs_lsb_1[1]),
    .S(_04146_),
    .Z(_00581_)
  );
  AND2_X1 _17381_ (
    .A1(_03421_),
    .A2(_03558_),
    .ZN(_02013_)
  );
  AND2_X1 _17382_ (
    .A1(_ex_reg_valid_T),
    .A2(_02013_),
    .ZN(_02014_)
  );
  OR2_X1 _17383_ (
    .A1(id_reg_pause),
    .A2(_02014_),
    .ZN(_02015_)
  );
  OR2_X1 _17384_ (
    .A1(csr_io_time[0]),
    .A2(csr_io_time[1]),
    .ZN(_02016_)
  );
  OR2_X1 _17385_ (
    .A1(csr_io_time[2]),
    .A2(csr_io_time[4]),
    .ZN(_02017_)
  );
  OR2_X1 _17386_ (
    .A1(_02016_),
    .A2(_02017_),
    .ZN(_02018_)
  );
  OR2_X1 _17387_ (
    .A1(csr_io_time[3]),
    .A2(_02018_),
    .ZN(_02019_)
  );
  AND2_X1 _17388_ (
    .A1(_03095_),
    .A2(_02019_),
    .ZN(_02020_)
  );
  AND2_X1 _17389_ (
    .A1(_04036_),
    .A2(_02020_),
    .ZN(_02021_)
  );
  AND2_X1 _17390_ (
    .A1(_02015_),
    .A2(_02021_),
    .ZN(_00582_)
  );
  AND2_X1 _17391_ (
    .A1(csr_io_decode_0_inst[26]),
    .A2(_03578_),
    .ZN(_02022_)
  );
  OR2_X1 _17392_ (
    .A1(_03558_),
    .A2(_02022_),
    .ZN(_02023_)
  );
  AND2_X1 _17393_ (
    .A1(_ex_reg_valid_T),
    .A2(_02023_),
    .ZN(_02024_)
  );
  OR2_X1 _17394_ (
    .A1(_03701_),
    .A2(_02024_),
    .ZN(_02025_)
  );
  AND2_X1 _17395_ (
    .A1(_02979_),
    .A2(_02025_),
    .ZN(_00583_)
  );
  AND2_X1 _17396_ (
    .A1(ibuf_io_inst_0_bits_xcpt1_pf_inst),
    .A2(_01783_),
    .ZN(_02026_)
  );
  OR2_X1 _17397_ (
    .A1(bpu_io_debug_if),
    .A2(_02026_),
    .ZN(_02027_)
  );
  INV_X1 _17398_ (
    .A(_02027_),
    .ZN(_02028_)
  );
  OR2_X1 _17399_ (
    .A1(csr_io_interrupt),
    .A2(_02028_),
    .ZN(_02029_)
  );
  AND2_X1 _17400_ (
    .A1(ibuf_io_inst_0_bits_xcpt1_ae_inst),
    .A2(_03060_),
    .ZN(_02030_)
  );
  OR2_X1 _17401_ (
    .A1(_01784_),
    .A2(_02030_),
    .ZN(_02031_)
  );
  MUX2_X1 _17402_ (
    .A(csr_io_interrupt_cause[0]),
    .B(_02031_),
    .S(_02978_),
    .Z(_02032_)
  );
  AND2_X1 _17403_ (
    .A1(_02029_),
    .A2(_02032_),
    .ZN(_02033_)
  );
  MUX2_X1 _17404_ (
    .A(ex_reg_cause[0]),
    .B(_02033_),
    .S(_01698_),
    .Z(_00584_)
  );
  OR2_X1 _17405_ (
    .A1(_02978_),
    .A2(csr_io_interrupt_cause[1]),
    .ZN(_02034_)
  );
  OR2_X1 _17406_ (
    .A1(bpu_io_xcpt_if),
    .A2(_01787_),
    .ZN(_02035_)
  );
  OR2_X1 _17407_ (
    .A1(_01785_),
    .A2(_02035_),
    .ZN(_02036_)
  );
  AND2_X1 _17408_ (
    .A1(_02034_),
    .A2(_02036_),
    .ZN(_02037_)
  );
  MUX2_X1 _17409_ (
    .A(ex_reg_cause[1]),
    .B(_02037_),
    .S(_01698_),
    .Z(_00585_)
  );
  AND2_X1 _17410_ (
    .A1(ibuf_io_inst_0_bits_xcpt1_gf_inst),
    .A2(_01783_),
    .ZN(_02038_)
  );
  OR2_X1 _17411_ (
    .A1(ibuf_io_inst_0_bits_xcpt1_pf_inst),
    .A2(_01787_),
    .ZN(_02039_)
  );
  INV_X1 _17412_ (
    .A(_02039_),
    .ZN(_02040_)
  );
  AND2_X1 _17413_ (
    .A1(_02038_),
    .A2(_02040_),
    .ZN(_02041_)
  );
  MUX2_X1 _17414_ (
    .A(csr_io_interrupt_cause[2]),
    .B(_02027_),
    .S(_02978_),
    .Z(_02042_)
  );
  OR2_X1 _17415_ (
    .A1(_02041_),
    .A2(_02042_),
    .ZN(_02043_)
  );
  MUX2_X1 _17416_ (
    .A(ex_reg_cause[2]),
    .B(_02043_),
    .S(_01698_),
    .Z(_00586_)
  );
  MUX2_X1 _17417_ (
    .A(csr_io_interrupt_cause[3]),
    .B(_02027_),
    .S(_02978_),
    .Z(_02044_)
  );
  MUX2_X1 _17418_ (
    .A(ex_reg_cause[3]),
    .B(_02044_),
    .S(_01698_),
    .Z(_00587_)
  );
  AND2_X1 _17419_ (
    .A1(csr_io_interrupt),
    .A2(csr_io_interrupt_cause[4]),
    .ZN(_02045_)
  );
  OR2_X1 _17420_ (
    .A1(_02041_),
    .A2(_02045_),
    .ZN(_02046_)
  );
  MUX2_X1 _17421_ (
    .A(ex_reg_cause[4]),
    .B(_02046_),
    .S(_01698_),
    .Z(_00588_)
  );
  AND2_X1 _17422_ (
    .A1(_03561_),
    .A2(_03569_),
    .ZN(_02047_)
  );
  MUX2_X1 _17423_ (
    .A(_02047_),
    .B(ex_ctrl_csr[0]),
    .S(_04146_),
    .Z(_00589_)
  );
  AND2_X1 _17424_ (
    .A1(_03565_),
    .A2(_03569_),
    .ZN(_02048_)
  );
  MUX2_X1 _17425_ (
    .A(_02048_),
    .B(ex_ctrl_csr[2]),
    .S(_04146_),
    .Z(_00590_)
  );
  OR2_X1 _17426_ (
    .A1(wb_reg_cause[0]),
    .A2(_06433_),
    .ZN(_02049_)
  );
  AND2_X1 _17427_ (
    .A1(mem_reg_load),
    .A2(bpu_io_debug_ld),
    .ZN(_02050_)
  );
  AND2_X1 _17428_ (
    .A1(mem_reg_store),
    .A2(bpu_io_debug_st),
    .ZN(_02051_)
  );
  OR2_X1 _17429_ (
    .A1(_02050_),
    .A2(_02051_),
    .ZN(_02052_)
  );
  INV_X1 _17430_ (
    .A(_02052_),
    .ZN(_02053_)
  );
  AND2_X1 _17431_ (
    .A1(mem_reg_valid),
    .A2(_06439_),
    .ZN(_02054_)
  );
  INV_X1 _17432_ (
    .A(_02054_),
    .ZN(_02055_)
  );
  AND2_X1 _17433_ (
    .A1(_08719_),
    .A2(_02055_),
    .ZN(_02056_)
  );
  INV_X1 _17434_ (
    .A(_02056_),
    .ZN(_02057_)
  );
  AND2_X1 _17435_ (
    .A1(_02053_),
    .A2(_02056_),
    .ZN(_02058_)
  );
  AND2_X1 _17436_ (
    .A1(mem_reg_cause[0]),
    .A2(_08718_),
    .ZN(_02059_)
  );
  OR2_X1 _17437_ (
    .A1(_06432_),
    .A2(_02059_),
    .ZN(_02060_)
  );
  OR2_X1 _17438_ (
    .A1(_02058_),
    .A2(_02060_),
    .ZN(_02061_)
  );
  AND2_X1 _17439_ (
    .A1(_02049_),
    .A2(_02061_),
    .ZN(_00591_)
  );
  OR2_X1 _17440_ (
    .A1(wb_reg_cause[1]),
    .A2(_06433_),
    .ZN(_02062_)
  );
  AND2_X1 _17441_ (
    .A1(mem_reg_cause[1]),
    .A2(_08718_),
    .ZN(_02063_)
  );
  OR2_X1 _17442_ (
    .A1(_06432_),
    .A2(_02063_),
    .ZN(_02064_)
  );
  OR2_X1 _17443_ (
    .A1(_02056_),
    .A2(_02064_),
    .ZN(_02065_)
  );
  AND2_X1 _17444_ (
    .A1(_02062_),
    .A2(_02065_),
    .ZN(_00592_)
  );
  OR2_X1 _17445_ (
    .A1(wb_reg_cause[2]),
    .A2(_06433_),
    .ZN(_02066_)
  );
  AND2_X1 _17446_ (
    .A1(_02052_),
    .A2(_02056_),
    .ZN(_02067_)
  );
  AND2_X1 _17447_ (
    .A1(mem_reg_cause[2]),
    .A2(_08718_),
    .ZN(_02068_)
  );
  OR2_X1 _17448_ (
    .A1(_06432_),
    .A2(_02068_),
    .ZN(_02069_)
  );
  OR2_X1 _17449_ (
    .A1(_02067_),
    .A2(_02069_),
    .ZN(_02070_)
  );
  AND2_X1 _17450_ (
    .A1(_02066_),
    .A2(_02070_),
    .ZN(_00593_)
  );
  OR2_X1 _17451_ (
    .A1(wb_reg_cause[3]),
    .A2(_06433_),
    .ZN(_02071_)
  );
  AND2_X1 _17452_ (
    .A1(mem_reg_cause[3]),
    .A2(_08718_),
    .ZN(_02072_)
  );
  OR2_X1 _17453_ (
    .A1(_06432_),
    .A2(_02072_),
    .ZN(_02073_)
  );
  OR2_X1 _17454_ (
    .A1(_02067_),
    .A2(_02073_),
    .ZN(_02074_)
  );
  AND2_X1 _17455_ (
    .A1(_02071_),
    .A2(_02074_),
    .ZN(_00594_)
  );
  AND2_X1 _17456_ (
    .A1(_04050_),
    .A2(_04062_),
    .ZN(_02075_)
  );
  INV_X1 _17457_ (
    .A(_02075_),
    .ZN(_02076_)
  );
  AND2_X1 _17458_ (
    .A1(_04047_),
    .A2(_02075_),
    .ZN(_02077_)
  );
  AND2_X1 _17459_ (
    .A1(_04057_),
    .A2(_04062_),
    .ZN(_02078_)
  );
  OR2_X1 _17460_ (
    .A1(_04056_),
    .A2(_04063_),
    .ZN(_02079_)
  );
  AND2_X1 _17461_ (
    .A1(_04054_),
    .A2(_02078_),
    .ZN(_02080_)
  );
  AND2_X1 _17462_ (
    .A1(_04053_),
    .A2(_02080_),
    .ZN(_02081_)
  );
  AND2_X1 _17463_ (
    .A1(_02077_),
    .A2(_02081_),
    .ZN(_02082_)
  );
  AND2_X1 _17464_ (
    .A1(_04062_),
    .A2(_06192_),
    .ZN(_02083_)
  );
  MUX2_X1 _17465_ (
    .A(\rf[9] [31]),
    .B(_02083_),
    .S(_02082_),
    .Z(_00595_)
  );
  AND2_X1 _17466_ (
    .A1(_04048_),
    .A2(_04062_),
    .ZN(_02084_)
  );
  OR2_X1 _17467_ (
    .A1(_04047_),
    .A2(_04063_),
    .ZN(_02085_)
  );
  AND2_X1 _17468_ (
    .A1(_02076_),
    .A2(_02085_),
    .ZN(_02086_)
  );
  AND2_X1 _17469_ (
    .A1(_02081_),
    .A2(_02086_),
    .ZN(_02087_)
  );
  MUX2_X1 _17470_ (
    .A(\rf[8] [31]),
    .B(_02083_),
    .S(_02087_),
    .Z(_00596_)
  );
  AND2_X1 _17471_ (
    .A1(_04048_),
    .A2(_02075_),
    .ZN(_02088_)
  );
  AND2_X1 _17472_ (
    .A1(_04052_),
    .A2(_04062_),
    .ZN(_02089_)
  );
  OR2_X1 _17473_ (
    .A1(_04053_),
    .A2(_04063_),
    .ZN(_02090_)
  );
  AND2_X1 _17474_ (
    .A1(_04055_),
    .A2(_04062_),
    .ZN(_02091_)
  );
  OR2_X1 _17475_ (
    .A1(_04054_),
    .A2(_04063_),
    .ZN(_02092_)
  );
  AND2_X1 _17476_ (
    .A1(_02079_),
    .A2(_02092_),
    .ZN(_02093_)
  );
  AND2_X1 _17477_ (
    .A1(_02089_),
    .A2(_02093_),
    .ZN(_02094_)
  );
  AND2_X1 _17478_ (
    .A1(_02088_),
    .A2(_02094_),
    .ZN(_02095_)
  );
  MUX2_X1 _17479_ (
    .A(\rf[7] [31]),
    .B(_06192_),
    .S(_02095_),
    .Z(_00597_)
  );
  AND2_X1 _17480_ (
    .A1(_04049_),
    .A2(_02084_),
    .ZN(_02096_)
  );
  AND2_X1 _17481_ (
    .A1(_02094_),
    .A2(_02096_),
    .ZN(_02097_)
  );
  MUX2_X1 _17482_ (
    .A(\rf[6] [31]),
    .B(_02083_),
    .S(_02097_),
    .Z(_00598_)
  );
  AND2_X1 _17483_ (
    .A1(_02077_),
    .A2(_02094_),
    .ZN(_02098_)
  );
  MUX2_X1 _17484_ (
    .A(\rf[5] [31]),
    .B(_02083_),
    .S(_02098_),
    .Z(_00599_)
  );
  AND2_X1 _17485_ (
    .A1(_02086_),
    .A2(_02094_),
    .ZN(_02099_)
  );
  MUX2_X1 _17486_ (
    .A(\rf[4] [31]),
    .B(_02083_),
    .S(_02099_),
    .Z(_00600_)
  );
  AND2_X1 _17487_ (
    .A1(_02090_),
    .A2(_02093_),
    .ZN(_02100_)
  );
  AND2_X1 _17488_ (
    .A1(_02088_),
    .A2(_02100_),
    .ZN(_02101_)
  );
  MUX2_X1 _17489_ (
    .A(\rf[3] [31]),
    .B(_02083_),
    .S(_02101_),
    .Z(_00601_)
  );
  AND2_X1 _17490_ (
    .A1(_04059_),
    .A2(_02096_),
    .ZN(_02102_)
  );
  MUX2_X1 _17491_ (
    .A(\rf[30] [31]),
    .B(_02083_),
    .S(_02102_),
    .Z(_00602_)
  );
  AND2_X1 _17492_ (
    .A1(_02096_),
    .A2(_02100_),
    .ZN(_02103_)
  );
  MUX2_X1 _17493_ (
    .A(\rf[2] [31]),
    .B(_02083_),
    .S(_02103_),
    .Z(_00603_)
  );
  AND2_X1 _17494_ (
    .A1(_04059_),
    .A2(_02077_),
    .ZN(_02104_)
  );
  MUX2_X1 _17495_ (
    .A(\rf[29] [31]),
    .B(_02083_),
    .S(_02104_),
    .Z(_00604_)
  );
  AND2_X1 _17496_ (
    .A1(_04062_),
    .A2(_02086_),
    .ZN(_02105_)
  );
  AND2_X1 _17497_ (
    .A1(_04059_),
    .A2(_02105_),
    .ZN(_02106_)
  );
  MUX2_X1 _17498_ (
    .A(\rf[28] [31]),
    .B(_02083_),
    .S(_02106_),
    .Z(_00605_)
  );
  AND2_X1 _17499_ (
    .A1(_04053_),
    .A2(_04058_),
    .ZN(_02107_)
  );
  AND2_X1 _17500_ (
    .A1(_02088_),
    .A2(_02107_),
    .ZN(_02108_)
  );
  MUX2_X1 _17501_ (
    .A(\rf[27] [31]),
    .B(_02083_),
    .S(_02108_),
    .Z(_00606_)
  );
  AND2_X1 _17502_ (
    .A1(_02096_),
    .A2(_02107_),
    .ZN(_02109_)
  );
  MUX2_X1 _17503_ (
    .A(\rf[26] [31]),
    .B(_02083_),
    .S(_02109_),
    .Z(_00607_)
  );
  AND2_X1 _17504_ (
    .A1(_02077_),
    .A2(_02107_),
    .ZN(_02110_)
  );
  MUX2_X1 _17505_ (
    .A(\rf[25] [31]),
    .B(_02083_),
    .S(_02110_),
    .Z(_00608_)
  );
  AND2_X1 _17506_ (
    .A1(_02105_),
    .A2(_02107_),
    .ZN(_02111_)
  );
  MUX2_X1 _17507_ (
    .A(\rf[24] [31]),
    .B(_06192_),
    .S(_02111_),
    .Z(_00609_)
  );
  AND2_X1 _17508_ (
    .A1(_04056_),
    .A2(_02091_),
    .ZN(_02112_)
  );
  AND2_X1 _17509_ (
    .A1(_04052_),
    .A2(_02112_),
    .ZN(_02113_)
  );
  AND2_X1 _17510_ (
    .A1(_02088_),
    .A2(_02113_),
    .ZN(_02114_)
  );
  MUX2_X1 _17511_ (
    .A(\rf[23] [31]),
    .B(_02083_),
    .S(_02114_),
    .Z(_00610_)
  );
  AND2_X1 _17512_ (
    .A1(_02096_),
    .A2(_02113_),
    .ZN(_02115_)
  );
  MUX2_X1 _17513_ (
    .A(\rf[22] [31]),
    .B(_02083_),
    .S(_02115_),
    .Z(_00611_)
  );
  AND2_X1 _17514_ (
    .A1(_02077_),
    .A2(_02113_),
    .ZN(_02116_)
  );
  MUX2_X1 _17515_ (
    .A(\rf[21] [31]),
    .B(_02083_),
    .S(_02116_),
    .Z(_00612_)
  );
  AND2_X1 _17516_ (
    .A1(_02086_),
    .A2(_02113_),
    .ZN(_02117_)
  );
  MUX2_X1 _17517_ (
    .A(\rf[20] [31]),
    .B(_02083_),
    .S(_02117_),
    .Z(_00613_)
  );
  AND2_X1 _17518_ (
    .A1(_02077_),
    .A2(_02100_),
    .ZN(_02118_)
  );
  MUX2_X1 _17519_ (
    .A(\rf[1] [31]),
    .B(_02083_),
    .S(_02118_),
    .Z(_00614_)
  );
  AND2_X1 _17520_ (
    .A1(_04053_),
    .A2(_02112_),
    .ZN(_02119_)
  );
  AND2_X1 _17521_ (
    .A1(_02088_),
    .A2(_02119_),
    .ZN(_02120_)
  );
  MUX2_X1 _17522_ (
    .A(\rf[19] [31]),
    .B(_06192_),
    .S(_02120_),
    .Z(_00615_)
  );
  AND2_X1 _17523_ (
    .A1(_02096_),
    .A2(_02119_),
    .ZN(_02121_)
  );
  MUX2_X1 _17524_ (
    .A(\rf[18] [31]),
    .B(_02083_),
    .S(_02121_),
    .Z(_00616_)
  );
  AND2_X1 _17525_ (
    .A1(_02077_),
    .A2(_02119_),
    .ZN(_02122_)
  );
  MUX2_X1 _17526_ (
    .A(\rf[17] [31]),
    .B(_02083_),
    .S(_02122_),
    .Z(_00617_)
  );
  AND2_X1 _17527_ (
    .A1(_02086_),
    .A2(_02119_),
    .ZN(_02123_)
  );
  MUX2_X1 _17528_ (
    .A(\rf[16] [31]),
    .B(_02083_),
    .S(_02123_),
    .Z(_00618_)
  );
  AND2_X1 _17529_ (
    .A1(_04052_),
    .A2(_02080_),
    .ZN(_02124_)
  );
  AND2_X1 _17530_ (
    .A1(_02088_),
    .A2(_02124_),
    .ZN(_02125_)
  );
  MUX2_X1 _17531_ (
    .A(\rf[15] [31]),
    .B(_02083_),
    .S(_02125_),
    .Z(_00619_)
  );
  AND2_X1 _17532_ (
    .A1(_02096_),
    .A2(_02124_),
    .ZN(_02126_)
  );
  MUX2_X1 _17533_ (
    .A(\rf[14] [31]),
    .B(_02083_),
    .S(_02126_),
    .Z(_00620_)
  );
  AND2_X1 _17534_ (
    .A1(_02077_),
    .A2(_02124_),
    .ZN(_02127_)
  );
  MUX2_X1 _17535_ (
    .A(\rf[13] [31]),
    .B(_02083_),
    .S(_02127_),
    .Z(_00621_)
  );
  AND2_X1 _17536_ (
    .A1(_02086_),
    .A2(_02124_),
    .ZN(_02128_)
  );
  MUX2_X1 _17537_ (
    .A(\rf[12] [31]),
    .B(_02083_),
    .S(_02128_),
    .Z(_00622_)
  );
  AND2_X1 _17538_ (
    .A1(_02081_),
    .A2(_02088_),
    .ZN(_02129_)
  );
  MUX2_X1 _17539_ (
    .A(\rf[11] [31]),
    .B(_06192_),
    .S(_02129_),
    .Z(_00623_)
  );
  AND2_X1 _17540_ (
    .A1(_02081_),
    .A2(_02096_),
    .ZN(_02130_)
  );
  MUX2_X1 _17541_ (
    .A(\rf[10] [31]),
    .B(_02083_),
    .S(_02130_),
    .Z(_00624_)
  );
  AND2_X1 _17542_ (
    .A1(_02100_),
    .A2(_02105_),
    .ZN(_02131_)
  );
  MUX2_X1 _17543_ (
    .A(\rf[0] [31]),
    .B(_06192_),
    .S(_02131_),
    .Z(_00625_)
  );
  AND2_X1 _17544_ (
    .A1(_04062_),
    .A2(_06266_),
    .ZN(_02132_)
  );
  MUX2_X1 _17545_ (
    .A(\rf[25] [0]),
    .B(_02132_),
    .S(_02110_),
    .Z(_00626_)
  );
  AND2_X1 _17546_ (
    .A1(_04062_),
    .A2(_06420_),
    .ZN(_02133_)
  );
  MUX2_X1 _17547_ (
    .A(\rf[25] [1]),
    .B(_02133_),
    .S(_02110_),
    .Z(_00627_)
  );
  AND2_X1 _17548_ (
    .A1(_04062_),
    .A2(_04080_),
    .ZN(_02134_)
  );
  MUX2_X1 _17549_ (
    .A(\rf[25] [2]),
    .B(_02134_),
    .S(_02110_),
    .Z(_00628_)
  );
  AND2_X1 _17550_ (
    .A1(_04062_),
    .A2(_04150_),
    .ZN(_02135_)
  );
  MUX2_X1 _17551_ (
    .A(\rf[25] [3]),
    .B(_02135_),
    .S(_02110_),
    .Z(_00629_)
  );
  AND2_X1 _17552_ (
    .A1(_04062_),
    .A2(_04233_),
    .ZN(_02136_)
  );
  MUX2_X1 _17553_ (
    .A(\rf[25] [4]),
    .B(_02136_),
    .S(_02110_),
    .Z(_00630_)
  );
  AND2_X1 _17554_ (
    .A1(_04062_),
    .A2(_04305_),
    .ZN(_02137_)
  );
  MUX2_X1 _17555_ (
    .A(\rf[25] [5]),
    .B(_02137_),
    .S(_02110_),
    .Z(_00631_)
  );
  AND2_X1 _17556_ (
    .A1(_04062_),
    .A2(_04379_),
    .ZN(_02138_)
  );
  MUX2_X1 _17557_ (
    .A(\rf[25] [6]),
    .B(_02138_),
    .S(_02110_),
    .Z(_00632_)
  );
  AND2_X1 _17558_ (
    .A1(_04062_),
    .A2(_04450_),
    .ZN(_02139_)
  );
  MUX2_X1 _17559_ (
    .A(\rf[25] [7]),
    .B(_02139_),
    .S(_02110_),
    .Z(_00633_)
  );
  AND2_X1 _17560_ (
    .A1(_04062_),
    .A2(_04521_),
    .ZN(_02140_)
  );
  MUX2_X1 _17561_ (
    .A(\rf[25] [8]),
    .B(_02140_),
    .S(_02110_),
    .Z(_00634_)
  );
  AND2_X1 _17562_ (
    .A1(_04062_),
    .A2(_04590_),
    .ZN(_02141_)
  );
  MUX2_X1 _17563_ (
    .A(\rf[25] [9]),
    .B(_02141_),
    .S(_02110_),
    .Z(_00635_)
  );
  AND2_X1 _17564_ (
    .A1(_04062_),
    .A2(_04659_),
    .ZN(_02142_)
  );
  MUX2_X1 _17565_ (
    .A(\rf[25] [10]),
    .B(_02142_),
    .S(_02110_),
    .Z(_00636_)
  );
  AND2_X1 _17566_ (
    .A1(_04062_),
    .A2(_04742_),
    .ZN(_02143_)
  );
  MUX2_X1 _17567_ (
    .A(\rf[25] [11]),
    .B(_02143_),
    .S(_02110_),
    .Z(_00637_)
  );
  AND2_X1 _17568_ (
    .A1(_04062_),
    .A2(_04811_),
    .ZN(_02144_)
  );
  MUX2_X1 _17569_ (
    .A(\rf[25] [12]),
    .B(_02144_),
    .S(_02110_),
    .Z(_00638_)
  );
  AND2_X1 _17570_ (
    .A1(_04062_),
    .A2(_04882_),
    .ZN(_02145_)
  );
  MUX2_X1 _17571_ (
    .A(\rf[25] [13]),
    .B(_02145_),
    .S(_02110_),
    .Z(_00639_)
  );
  AND2_X1 _17572_ (
    .A1(_04062_),
    .A2(_04953_),
    .ZN(_02146_)
  );
  MUX2_X1 _17573_ (
    .A(\rf[25] [14]),
    .B(_02146_),
    .S(_02110_),
    .Z(_00640_)
  );
  AND2_X1 _17574_ (
    .A1(_04062_),
    .A2(_05027_),
    .ZN(_02147_)
  );
  MUX2_X1 _17575_ (
    .A(\rf[25] [15]),
    .B(_02147_),
    .S(_02110_),
    .Z(_00641_)
  );
  AND2_X1 _17576_ (
    .A1(_04062_),
    .A2(_05095_),
    .ZN(_02148_)
  );
  MUX2_X1 _17577_ (
    .A(\rf[25] [16]),
    .B(_02148_),
    .S(_02110_),
    .Z(_00642_)
  );
  AND2_X1 _17578_ (
    .A1(_04062_),
    .A2(_05170_),
    .ZN(_02149_)
  );
  MUX2_X1 _17579_ (
    .A(\rf[25] [17]),
    .B(_02149_),
    .S(_02110_),
    .Z(_00643_)
  );
  AND2_X1 _17580_ (
    .A1(_04062_),
    .A2(_05302_),
    .ZN(_02150_)
  );
  MUX2_X1 _17581_ (
    .A(\rf[25] [18]),
    .B(_02150_),
    .S(_02110_),
    .Z(_00644_)
  );
  AND2_X1 _17582_ (
    .A1(_04062_),
    .A2(_05310_),
    .ZN(_02151_)
  );
  MUX2_X1 _17583_ (
    .A(\rf[25] [19]),
    .B(_02151_),
    .S(_02110_),
    .Z(_00645_)
  );
  AND2_X1 _17584_ (
    .A1(_04062_),
    .A2(_05442_),
    .ZN(_02152_)
  );
  MUX2_X1 _17585_ (
    .A(\rf[25] [20]),
    .B(_02152_),
    .S(_02110_),
    .Z(_00646_)
  );
  AND2_X1 _17586_ (
    .A1(_04062_),
    .A2(_05450_),
    .ZN(_02153_)
  );
  MUX2_X1 _17587_ (
    .A(\rf[25] [21]),
    .B(_02153_),
    .S(_02110_),
    .Z(_00647_)
  );
  AND2_X1 _17588_ (
    .A1(_04062_),
    .A2(_05592_),
    .ZN(_02154_)
  );
  MUX2_X1 _17589_ (
    .A(\rf[25] [22]),
    .B(_02154_),
    .S(_02110_),
    .Z(_00648_)
  );
  AND2_X1 _17590_ (
    .A1(_04062_),
    .A2(_05657_),
    .ZN(_02155_)
  );
  MUX2_X1 _17591_ (
    .A(\rf[25] [23]),
    .B(_02155_),
    .S(_02110_),
    .Z(_00649_)
  );
  AND2_X1 _17592_ (
    .A1(_04062_),
    .A2(_05665_),
    .ZN(_02156_)
  );
  MUX2_X1 _17593_ (
    .A(\rf[25] [24]),
    .B(_02156_),
    .S(_02110_),
    .Z(_00650_)
  );
  AND2_X1 _17594_ (
    .A1(_04062_),
    .A2(_05740_),
    .ZN(_02157_)
  );
  MUX2_X1 _17595_ (
    .A(\rf[25] [25]),
    .B(_02157_),
    .S(_02110_),
    .Z(_00651_)
  );
  AND2_X1 _17596_ (
    .A1(_04062_),
    .A2(_05882_),
    .ZN(_02158_)
  );
  MUX2_X1 _17597_ (
    .A(\rf[25] [26]),
    .B(_02158_),
    .S(_02110_),
    .Z(_00652_)
  );
  AND2_X1 _17598_ (
    .A1(_04062_),
    .A2(_05957_),
    .ZN(_02159_)
  );
  MUX2_X1 _17599_ (
    .A(\rf[25] [27]),
    .B(_02159_),
    .S(_02110_),
    .Z(_00653_)
  );
  AND2_X1 _17600_ (
    .A1(_04062_),
    .A2(_06032_),
    .ZN(_02160_)
  );
  MUX2_X1 _17601_ (
    .A(\rf[25] [28]),
    .B(_02160_),
    .S(_02110_),
    .Z(_00654_)
  );
  AND2_X1 _17602_ (
    .A1(_04062_),
    .A2(_06109_),
    .ZN(_02161_)
  );
  MUX2_X1 _17603_ (
    .A(\rf[25] [29]),
    .B(_02161_),
    .S(_02110_),
    .Z(_00655_)
  );
  AND2_X1 _17604_ (
    .A1(_04062_),
    .A2(_06117_),
    .ZN(_02162_)
  );
  MUX2_X1 _17605_ (
    .A(\rf[25] [30]),
    .B(_02162_),
    .S(_02110_),
    .Z(_00656_)
  );
  MUX2_X1 _17606_ (
    .A(\rf[23] [0]),
    .B(_06266_),
    .S(_02114_),
    .Z(_00657_)
  );
  MUX2_X1 _17607_ (
    .A(\rf[23] [1]),
    .B(_02133_),
    .S(_02114_),
    .Z(_00658_)
  );
  MUX2_X1 _17608_ (
    .A(\rf[23] [2]),
    .B(_04080_),
    .S(_02114_),
    .Z(_00659_)
  );
  MUX2_X1 _17609_ (
    .A(\rf[23] [3]),
    .B(_04150_),
    .S(_02114_),
    .Z(_00660_)
  );
  MUX2_X1 _17610_ (
    .A(\rf[23] [4]),
    .B(_04233_),
    .S(_02114_),
    .Z(_00661_)
  );
  MUX2_X1 _17611_ (
    .A(\rf[23] [5]),
    .B(_04305_),
    .S(_02114_),
    .Z(_00662_)
  );
  MUX2_X1 _17612_ (
    .A(\rf[23] [6]),
    .B(_04379_),
    .S(_02114_),
    .Z(_00663_)
  );
  MUX2_X1 _17613_ (
    .A(\rf[23] [7]),
    .B(_02139_),
    .S(_02114_),
    .Z(_00664_)
  );
  MUX2_X1 _17614_ (
    .A(\rf[23] [8]),
    .B(_04521_),
    .S(_02114_),
    .Z(_00665_)
  );
  MUX2_X1 _17615_ (
    .A(\rf[23] [9]),
    .B(_04590_),
    .S(_02114_),
    .Z(_00666_)
  );
  MUX2_X1 _17616_ (
    .A(\rf[23] [10]),
    .B(_02142_),
    .S(_02114_),
    .Z(_00667_)
  );
  MUX2_X1 _17617_ (
    .A(\rf[23] [11]),
    .B(_04742_),
    .S(_02114_),
    .Z(_00668_)
  );
  MUX2_X1 _17618_ (
    .A(\rf[23] [12]),
    .B(_04811_),
    .S(_02114_),
    .Z(_00669_)
  );
  MUX2_X1 _17619_ (
    .A(\rf[23] [13]),
    .B(_04882_),
    .S(_02114_),
    .Z(_00670_)
  );
  MUX2_X1 _17620_ (
    .A(\rf[23] [14]),
    .B(_04953_),
    .S(_02114_),
    .Z(_00671_)
  );
  MUX2_X1 _17621_ (
    .A(\rf[23] [15]),
    .B(_05027_),
    .S(_02114_),
    .Z(_00672_)
  );
  MUX2_X1 _17622_ (
    .A(\rf[23] [16]),
    .B(_02148_),
    .S(_02114_),
    .Z(_00673_)
  );
  MUX2_X1 _17623_ (
    .A(\rf[23] [17]),
    .B(_05170_),
    .S(_02114_),
    .Z(_00674_)
  );
  MUX2_X1 _17624_ (
    .A(\rf[23] [18]),
    .B(_05302_),
    .S(_02114_),
    .Z(_00675_)
  );
  MUX2_X1 _17625_ (
    .A(\rf[23] [19]),
    .B(_02151_),
    .S(_02114_),
    .Z(_00676_)
  );
  MUX2_X1 _17626_ (
    .A(\rf[23] [20]),
    .B(_05442_),
    .S(_02114_),
    .Z(_00677_)
  );
  MUX2_X1 _17627_ (
    .A(\rf[23] [21]),
    .B(_02153_),
    .S(_02114_),
    .Z(_00678_)
  );
  MUX2_X1 _17628_ (
    .A(\rf[23] [22]),
    .B(_05592_),
    .S(_02114_),
    .Z(_00679_)
  );
  MUX2_X1 _17629_ (
    .A(\rf[23] [23]),
    .B(_05657_),
    .S(_02114_),
    .Z(_00680_)
  );
  MUX2_X1 _17630_ (
    .A(\rf[23] [24]),
    .B(_05665_),
    .S(_02114_),
    .Z(_00681_)
  );
  MUX2_X1 _17631_ (
    .A(\rf[23] [25]),
    .B(_05740_),
    .S(_02114_),
    .Z(_00682_)
  );
  MUX2_X1 _17632_ (
    .A(\rf[23] [26]),
    .B(_05882_),
    .S(_02114_),
    .Z(_00683_)
  );
  MUX2_X1 _17633_ (
    .A(\rf[23] [27]),
    .B(_05957_),
    .S(_02114_),
    .Z(_00684_)
  );
  MUX2_X1 _17634_ (
    .A(\rf[23] [28]),
    .B(_06032_),
    .S(_02114_),
    .Z(_00685_)
  );
  MUX2_X1 _17635_ (
    .A(\rf[23] [29]),
    .B(_06109_),
    .S(_02114_),
    .Z(_00686_)
  );
  MUX2_X1 _17636_ (
    .A(\rf[23] [30]),
    .B(_06117_),
    .S(_02114_),
    .Z(_00687_)
  );
  MUX2_X1 _17637_ (
    .A(\rf[4] [26]),
    .B(_02158_),
    .S(_02099_),
    .Z(_00688_)
  );
  MUX2_X1 _17638_ (
    .A(\rf[4] [28]),
    .B(_02160_),
    .S(_02099_),
    .Z(_00689_)
  );
  MUX2_X1 _17639_ (
    .A(\rf[4] [30]),
    .B(_02162_),
    .S(_02099_),
    .Z(_00690_)
  );
  MUX2_X1 _17640_ (
    .A(\rf[6] [0]),
    .B(_02132_),
    .S(_02097_),
    .Z(_00691_)
  );
  MUX2_X1 _17641_ (
    .A(\rf[6] [1]),
    .B(_02133_),
    .S(_02097_),
    .Z(_00692_)
  );
  MUX2_X1 _17642_ (
    .A(\rf[6] [2]),
    .B(_02134_),
    .S(_02097_),
    .Z(_00693_)
  );
  MUX2_X1 _17643_ (
    .A(\rf[6] [3]),
    .B(_02135_),
    .S(_02097_),
    .Z(_00694_)
  );
  MUX2_X1 _17644_ (
    .A(\rf[6] [4]),
    .B(_02136_),
    .S(_02097_),
    .Z(_00695_)
  );
  MUX2_X1 _17645_ (
    .A(\rf[6] [5]),
    .B(_02137_),
    .S(_02097_),
    .Z(_00696_)
  );
  MUX2_X1 _17646_ (
    .A(\rf[6] [6]),
    .B(_02138_),
    .S(_02097_),
    .Z(_00697_)
  );
  MUX2_X1 _17647_ (
    .A(\rf[6] [7]),
    .B(_02139_),
    .S(_02097_),
    .Z(_00698_)
  );
  MUX2_X1 _17648_ (
    .A(\rf[6] [8]),
    .B(_02140_),
    .S(_02097_),
    .Z(_00699_)
  );
  MUX2_X1 _17649_ (
    .A(\rf[6] [9]),
    .B(_02141_),
    .S(_02097_),
    .Z(_00700_)
  );
  MUX2_X1 _17650_ (
    .A(\rf[6] [10]),
    .B(_02142_),
    .S(_02097_),
    .Z(_00701_)
  );
  MUX2_X1 _17651_ (
    .A(\rf[6] [11]),
    .B(_02143_),
    .S(_02097_),
    .Z(_00702_)
  );
  MUX2_X1 _17652_ (
    .A(\rf[6] [12]),
    .B(_02144_),
    .S(_02097_),
    .Z(_00703_)
  );
  MUX2_X1 _17653_ (
    .A(\rf[6] [13]),
    .B(_02145_),
    .S(_02097_),
    .Z(_00704_)
  );
  MUX2_X1 _17654_ (
    .A(\rf[6] [14]),
    .B(_02146_),
    .S(_02097_),
    .Z(_00705_)
  );
  MUX2_X1 _17655_ (
    .A(\rf[6] [15]),
    .B(_02147_),
    .S(_02097_),
    .Z(_00706_)
  );
  MUX2_X1 _17656_ (
    .A(\rf[6] [16]),
    .B(_02148_),
    .S(_02097_),
    .Z(_00707_)
  );
  MUX2_X1 _17657_ (
    .A(\rf[6] [17]),
    .B(_02149_),
    .S(_02097_),
    .Z(_00708_)
  );
  MUX2_X1 _17658_ (
    .A(\rf[6] [18]),
    .B(_02150_),
    .S(_02097_),
    .Z(_00709_)
  );
  MUX2_X1 _17659_ (
    .A(\rf[6] [19]),
    .B(_02151_),
    .S(_02097_),
    .Z(_00710_)
  );
  MUX2_X1 _17660_ (
    .A(\rf[6] [20]),
    .B(_02152_),
    .S(_02097_),
    .Z(_00711_)
  );
  MUX2_X1 _17661_ (
    .A(\rf[6] [21]),
    .B(_02153_),
    .S(_02097_),
    .Z(_00712_)
  );
  MUX2_X1 _17662_ (
    .A(\rf[6] [22]),
    .B(_02154_),
    .S(_02097_),
    .Z(_00713_)
  );
  MUX2_X1 _17663_ (
    .A(\rf[6] [23]),
    .B(_02155_),
    .S(_02097_),
    .Z(_00714_)
  );
  MUX2_X1 _17664_ (
    .A(\rf[6] [24]),
    .B(_02156_),
    .S(_02097_),
    .Z(_00715_)
  );
  MUX2_X1 _17665_ (
    .A(\rf[6] [25]),
    .B(_02157_),
    .S(_02097_),
    .Z(_00716_)
  );
  MUX2_X1 _17666_ (
    .A(\rf[6] [26]),
    .B(_02158_),
    .S(_02097_),
    .Z(_00717_)
  );
  MUX2_X1 _17667_ (
    .A(\rf[6] [27]),
    .B(_02159_),
    .S(_02097_),
    .Z(_00718_)
  );
  MUX2_X1 _17668_ (
    .A(\rf[6] [28]),
    .B(_02160_),
    .S(_02097_),
    .Z(_00719_)
  );
  MUX2_X1 _17669_ (
    .A(\rf[6] [29]),
    .B(_02161_),
    .S(_02097_),
    .Z(_00720_)
  );
  MUX2_X1 _17670_ (
    .A(\rf[6] [30]),
    .B(_02162_),
    .S(_02097_),
    .Z(_00721_)
  );
  MUX2_X1 _17671_ (
    .A(\rf[4] [0]),
    .B(_02132_),
    .S(_02099_),
    .Z(_00722_)
  );
  MUX2_X1 _17672_ (
    .A(\rf[4] [1]),
    .B(_02133_),
    .S(_02099_),
    .Z(_00723_)
  );
  MUX2_X1 _17673_ (
    .A(\rf[4] [2]),
    .B(_02134_),
    .S(_02099_),
    .Z(_00724_)
  );
  MUX2_X1 _17674_ (
    .A(\rf[4] [3]),
    .B(_02135_),
    .S(_02099_),
    .Z(_00725_)
  );
  MUX2_X1 _17675_ (
    .A(\rf[4] [4]),
    .B(_02136_),
    .S(_02099_),
    .Z(_00726_)
  );
  MUX2_X1 _17676_ (
    .A(\rf[4] [5]),
    .B(_02137_),
    .S(_02099_),
    .Z(_00727_)
  );
  MUX2_X1 _17677_ (
    .A(\rf[4] [6]),
    .B(_02138_),
    .S(_02099_),
    .Z(_00728_)
  );
  MUX2_X1 _17678_ (
    .A(\rf[4] [7]),
    .B(_02139_),
    .S(_02099_),
    .Z(_00729_)
  );
  MUX2_X1 _17679_ (
    .A(\rf[4] [8]),
    .B(_02140_),
    .S(_02099_),
    .Z(_00730_)
  );
  MUX2_X1 _17680_ (
    .A(\rf[4] [9]),
    .B(_02141_),
    .S(_02099_),
    .Z(_00731_)
  );
  MUX2_X1 _17681_ (
    .A(\rf[4] [10]),
    .B(_02142_),
    .S(_02099_),
    .Z(_00732_)
  );
  MUX2_X1 _17682_ (
    .A(\rf[4] [11]),
    .B(_02143_),
    .S(_02099_),
    .Z(_00733_)
  );
  MUX2_X1 _17683_ (
    .A(\rf[4] [12]),
    .B(_02144_),
    .S(_02099_),
    .Z(_00734_)
  );
  MUX2_X1 _17684_ (
    .A(\rf[4] [13]),
    .B(_02145_),
    .S(_02099_),
    .Z(_00735_)
  );
  MUX2_X1 _17685_ (
    .A(\rf[4] [14]),
    .B(_02146_),
    .S(_02099_),
    .Z(_00736_)
  );
  MUX2_X1 _17686_ (
    .A(\rf[4] [15]),
    .B(_02147_),
    .S(_02099_),
    .Z(_00737_)
  );
  MUX2_X1 _17687_ (
    .A(\rf[4] [16]),
    .B(_02148_),
    .S(_02099_),
    .Z(_00738_)
  );
  MUX2_X1 _17688_ (
    .A(\rf[4] [17]),
    .B(_02149_),
    .S(_02099_),
    .Z(_00739_)
  );
  MUX2_X1 _17689_ (
    .A(\rf[4] [18]),
    .B(_02150_),
    .S(_02099_),
    .Z(_00740_)
  );
  MUX2_X1 _17690_ (
    .A(\rf[4] [19]),
    .B(_02151_),
    .S(_02099_),
    .Z(_00741_)
  );
  MUX2_X1 _17691_ (
    .A(\rf[4] [20]),
    .B(_02152_),
    .S(_02099_),
    .Z(_00742_)
  );
  MUX2_X1 _17692_ (
    .A(\rf[4] [21]),
    .B(_02153_),
    .S(_02099_),
    .Z(_00743_)
  );
  MUX2_X1 _17693_ (
    .A(\rf[4] [23]),
    .B(_02155_),
    .S(_02099_),
    .Z(_00744_)
  );
  MUX2_X1 _17694_ (
    .A(\rf[4] [24]),
    .B(_02156_),
    .S(_02099_),
    .Z(_00745_)
  );
  MUX2_X1 _17695_ (
    .A(\rf[4] [22]),
    .B(_02154_),
    .S(_02099_),
    .Z(_00746_)
  );
  OR2_X1 _17696_ (
    .A1(_03379_),
    .A2(_01829_),
    .ZN(_02163_)
  );
  OR2_X1 _17697_ (
    .A1(_03371_),
    .A2(_02163_),
    .ZN(_02164_)
  );
  OR2_X1 _17698_ (
    .A1(_03364_),
    .A2(_02164_),
    .ZN(_02165_)
  );
  OR2_X1 _17699_ (
    .A1(_03494_),
    .A2(_02165_),
    .ZN(_02166_)
  );
  AND2_X1 _17700_ (
    .A1(_01790_),
    .A2(_02166_),
    .ZN(_02167_)
  );
  MUX2_X1 _17701_ (
    .A(_02167_),
    .B(ex_ctrl_sel_alu2[1]),
    .S(_04041_),
    .Z(_00747_)
  );
  MUX2_X1 _17702_ (
    .A(\rf[4] [25]),
    .B(_02157_),
    .S(_02099_),
    .Z(_00748_)
  );
  MUX2_X1 _17703_ (
    .A(\rf[4] [27]),
    .B(_02159_),
    .S(_02099_),
    .Z(_00749_)
  );
  MUX2_X1 _17704_ (
    .A(\rf[4] [29]),
    .B(_02161_),
    .S(_02099_),
    .Z(_00750_)
  );
  MUX2_X1 _17705_ (
    .A(\rf[0] [0]),
    .B(_06266_),
    .S(_02131_),
    .Z(_00751_)
  );
  MUX2_X1 _17706_ (
    .A(\rf[0] [1]),
    .B(_06420_),
    .S(_02131_),
    .Z(_00752_)
  );
  MUX2_X1 _17707_ (
    .A(\rf[0] [2]),
    .B(_04080_),
    .S(_02131_),
    .Z(_00753_)
  );
  MUX2_X1 _17708_ (
    .A(\rf[0] [3]),
    .B(_04150_),
    .S(_02131_),
    .Z(_00754_)
  );
  MUX2_X1 _17709_ (
    .A(\rf[0] [4]),
    .B(_04233_),
    .S(_02131_),
    .Z(_00755_)
  );
  MUX2_X1 _17710_ (
    .A(\rf[0] [5]),
    .B(_04305_),
    .S(_02131_),
    .Z(_00756_)
  );
  MUX2_X1 _17711_ (
    .A(\rf[0] [6]),
    .B(_04379_),
    .S(_02131_),
    .Z(_00757_)
  );
  MUX2_X1 _17712_ (
    .A(\rf[0] [7]),
    .B(_04450_),
    .S(_02131_),
    .Z(_00758_)
  );
  MUX2_X1 _17713_ (
    .A(\rf[0] [8]),
    .B(_04521_),
    .S(_02131_),
    .Z(_00759_)
  );
  MUX2_X1 _17714_ (
    .A(\rf[0] [9]),
    .B(_04590_),
    .S(_02131_),
    .Z(_00760_)
  );
  MUX2_X1 _17715_ (
    .A(\rf[0] [10]),
    .B(_04659_),
    .S(_02131_),
    .Z(_00761_)
  );
  MUX2_X1 _17716_ (
    .A(\rf[0] [11]),
    .B(_04742_),
    .S(_02131_),
    .Z(_00762_)
  );
  MUX2_X1 _17717_ (
    .A(\rf[0] [12]),
    .B(_04811_),
    .S(_02131_),
    .Z(_00763_)
  );
  MUX2_X1 _17718_ (
    .A(\rf[0] [13]),
    .B(_04882_),
    .S(_02131_),
    .Z(_00764_)
  );
  MUX2_X1 _17719_ (
    .A(\rf[0] [14]),
    .B(_04953_),
    .S(_02131_),
    .Z(_00765_)
  );
  MUX2_X1 _17720_ (
    .A(\rf[0] [15]),
    .B(_05027_),
    .S(_02131_),
    .Z(_00766_)
  );
  MUX2_X1 _17721_ (
    .A(\rf[0] [16]),
    .B(_05095_),
    .S(_02131_),
    .Z(_00767_)
  );
  MUX2_X1 _17722_ (
    .A(\rf[0] [17]),
    .B(_05170_),
    .S(_02131_),
    .Z(_00768_)
  );
  MUX2_X1 _17723_ (
    .A(\rf[0] [18]),
    .B(_05302_),
    .S(_02131_),
    .Z(_00769_)
  );
  MUX2_X1 _17724_ (
    .A(\rf[0] [19]),
    .B(_05310_),
    .S(_02131_),
    .Z(_00770_)
  );
  MUX2_X1 _17725_ (
    .A(\rf[0] [20]),
    .B(_05442_),
    .S(_02131_),
    .Z(_00771_)
  );
  MUX2_X1 _17726_ (
    .A(\rf[0] [21]),
    .B(_05450_),
    .S(_02131_),
    .Z(_00772_)
  );
  MUX2_X1 _17727_ (
    .A(\rf[0] [22]),
    .B(_05592_),
    .S(_02131_),
    .Z(_00773_)
  );
  MUX2_X1 _17728_ (
    .A(\rf[0] [23]),
    .B(_05657_),
    .S(_02131_),
    .Z(_00774_)
  );
  MUX2_X1 _17729_ (
    .A(\rf[0] [24]),
    .B(_05665_),
    .S(_02131_),
    .Z(_00775_)
  );
  MUX2_X1 _17730_ (
    .A(\rf[0] [25]),
    .B(_05740_),
    .S(_02131_),
    .Z(_00776_)
  );
  MUX2_X1 _17731_ (
    .A(\rf[0] [26]),
    .B(_05882_),
    .S(_02131_),
    .Z(_00777_)
  );
  MUX2_X1 _17732_ (
    .A(\rf[0] [27]),
    .B(_05957_),
    .S(_02131_),
    .Z(_00778_)
  );
  MUX2_X1 _17733_ (
    .A(\rf[0] [28]),
    .B(_06032_),
    .S(_02131_),
    .Z(_00779_)
  );
  MUX2_X1 _17734_ (
    .A(\rf[0] [29]),
    .B(_06109_),
    .S(_02131_),
    .Z(_00780_)
  );
  MUX2_X1 _17735_ (
    .A(\rf[0] [30]),
    .B(_06117_),
    .S(_02131_),
    .Z(_00781_)
  );
  MUX2_X1 _17736_ (
    .A(\rf[15] [0]),
    .B(_02132_),
    .S(_02125_),
    .Z(_00782_)
  );
  MUX2_X1 _17737_ (
    .A(\rf[15] [1]),
    .B(_02133_),
    .S(_02125_),
    .Z(_00783_)
  );
  MUX2_X1 _17738_ (
    .A(\rf[15] [2]),
    .B(_04080_),
    .S(_02125_),
    .Z(_00784_)
  );
  MUX2_X1 _17739_ (
    .A(\rf[15] [3]),
    .B(_04150_),
    .S(_02125_),
    .Z(_00785_)
  );
  MUX2_X1 _17740_ (
    .A(\rf[15] [4]),
    .B(_04233_),
    .S(_02125_),
    .Z(_00786_)
  );
  MUX2_X1 _17741_ (
    .A(\rf[15] [5]),
    .B(_04305_),
    .S(_02125_),
    .Z(_00787_)
  );
  MUX2_X1 _17742_ (
    .A(\rf[15] [6]),
    .B(_02138_),
    .S(_02125_),
    .Z(_00788_)
  );
  MUX2_X1 _17743_ (
    .A(\rf[15] [7]),
    .B(_02139_),
    .S(_02125_),
    .Z(_00789_)
  );
  MUX2_X1 _17744_ (
    .A(\rf[15] [8]),
    .B(_04521_),
    .S(_02125_),
    .Z(_00790_)
  );
  MUX2_X1 _17745_ (
    .A(\rf[15] [9]),
    .B(_04590_),
    .S(_02125_),
    .Z(_00791_)
  );
  MUX2_X1 _17746_ (
    .A(\rf[15] [10]),
    .B(_04659_),
    .S(_02125_),
    .Z(_00792_)
  );
  MUX2_X1 _17747_ (
    .A(\rf[15] [11]),
    .B(_04742_),
    .S(_02125_),
    .Z(_00793_)
  );
  MUX2_X1 _17748_ (
    .A(\rf[15] [12]),
    .B(_04811_),
    .S(_02125_),
    .Z(_00794_)
  );
  MUX2_X1 _17749_ (
    .A(\rf[15] [13]),
    .B(_04882_),
    .S(_02125_),
    .Z(_00795_)
  );
  MUX2_X1 _17750_ (
    .A(\rf[15] [14]),
    .B(_04953_),
    .S(_02125_),
    .Z(_00796_)
  );
  MUX2_X1 _17751_ (
    .A(\rf[15] [15]),
    .B(_05027_),
    .S(_02125_),
    .Z(_00797_)
  );
  MUX2_X1 _17752_ (
    .A(\rf[15] [16]),
    .B(_02148_),
    .S(_02125_),
    .Z(_00798_)
  );
  MUX2_X1 _17753_ (
    .A(\rf[15] [17]),
    .B(_05170_),
    .S(_02125_),
    .Z(_00799_)
  );
  MUX2_X1 _17754_ (
    .A(\rf[15] [18]),
    .B(_02150_),
    .S(_02125_),
    .Z(_00800_)
  );
  MUX2_X1 _17755_ (
    .A(\rf[15] [19]),
    .B(_02151_),
    .S(_02125_),
    .Z(_00801_)
  );
  MUX2_X1 _17756_ (
    .A(\rf[15] [20]),
    .B(_05442_),
    .S(_02125_),
    .Z(_00802_)
  );
  MUX2_X1 _17757_ (
    .A(\rf[15] [21]),
    .B(_05450_),
    .S(_02125_),
    .Z(_00803_)
  );
  MUX2_X1 _17758_ (
    .A(\rf[15] [22]),
    .B(_05592_),
    .S(_02125_),
    .Z(_00804_)
  );
  MUX2_X1 _17759_ (
    .A(\rf[15] [23]),
    .B(_05657_),
    .S(_02125_),
    .Z(_00805_)
  );
  MUX2_X1 _17760_ (
    .A(\rf[15] [24]),
    .B(_05665_),
    .S(_02125_),
    .Z(_00806_)
  );
  MUX2_X1 _17761_ (
    .A(\rf[15] [25]),
    .B(_05740_),
    .S(_02125_),
    .Z(_00807_)
  );
  MUX2_X1 _17762_ (
    .A(\rf[15] [26]),
    .B(_05882_),
    .S(_02125_),
    .Z(_00808_)
  );
  MUX2_X1 _17763_ (
    .A(\rf[15] [27]),
    .B(_05957_),
    .S(_02125_),
    .Z(_00809_)
  );
  MUX2_X1 _17764_ (
    .A(\rf[15] [28]),
    .B(_02160_),
    .S(_02125_),
    .Z(_00810_)
  );
  MUX2_X1 _17765_ (
    .A(\rf[15] [29]),
    .B(_06109_),
    .S(_02125_),
    .Z(_00811_)
  );
  MUX2_X1 _17766_ (
    .A(\rf[15] [30]),
    .B(_06117_),
    .S(_02125_),
    .Z(_00812_)
  );
  MUX2_X1 _17767_ (
    .A(\rf[8] [0]),
    .B(_02132_),
    .S(_02087_),
    .Z(_00813_)
  );
  MUX2_X1 _17768_ (
    .A(\rf[8] [1]),
    .B(_02133_),
    .S(_02087_),
    .Z(_00814_)
  );
  MUX2_X1 _17769_ (
    .A(\rf[8] [2]),
    .B(_02134_),
    .S(_02087_),
    .Z(_00815_)
  );
  MUX2_X1 _17770_ (
    .A(\rf[8] [3]),
    .B(_02135_),
    .S(_02087_),
    .Z(_00816_)
  );
  MUX2_X1 _17771_ (
    .A(\rf[8] [4]),
    .B(_02136_),
    .S(_02087_),
    .Z(_00817_)
  );
  MUX2_X1 _17772_ (
    .A(\rf[8] [5]),
    .B(_02137_),
    .S(_02087_),
    .Z(_00818_)
  );
  MUX2_X1 _17773_ (
    .A(\rf[8] [6]),
    .B(_02138_),
    .S(_02087_),
    .Z(_00819_)
  );
  MUX2_X1 _17774_ (
    .A(\rf[8] [7]),
    .B(_02139_),
    .S(_02087_),
    .Z(_00820_)
  );
  MUX2_X1 _17775_ (
    .A(\rf[8] [8]),
    .B(_02140_),
    .S(_02087_),
    .Z(_00821_)
  );
  MUX2_X1 _17776_ (
    .A(\rf[8] [9]),
    .B(_02141_),
    .S(_02087_),
    .Z(_00822_)
  );
  MUX2_X1 _17777_ (
    .A(\rf[8] [10]),
    .B(_02142_),
    .S(_02087_),
    .Z(_00823_)
  );
  MUX2_X1 _17778_ (
    .A(\rf[8] [11]),
    .B(_02143_),
    .S(_02087_),
    .Z(_00824_)
  );
  MUX2_X1 _17779_ (
    .A(\rf[8] [12]),
    .B(_02144_),
    .S(_02087_),
    .Z(_00825_)
  );
  MUX2_X1 _17780_ (
    .A(\rf[8] [13]),
    .B(_02145_),
    .S(_02087_),
    .Z(_00826_)
  );
  MUX2_X1 _17781_ (
    .A(\rf[8] [14]),
    .B(_02146_),
    .S(_02087_),
    .Z(_00827_)
  );
  MUX2_X1 _17782_ (
    .A(\rf[8] [15]),
    .B(_02147_),
    .S(_02087_),
    .Z(_00828_)
  );
  MUX2_X1 _17783_ (
    .A(\rf[8] [16]),
    .B(_02148_),
    .S(_02087_),
    .Z(_00829_)
  );
  MUX2_X1 _17784_ (
    .A(\rf[8] [17]),
    .B(_02149_),
    .S(_02087_),
    .Z(_00830_)
  );
  MUX2_X1 _17785_ (
    .A(\rf[8] [18]),
    .B(_02150_),
    .S(_02087_),
    .Z(_00831_)
  );
  MUX2_X1 _17786_ (
    .A(\rf[8] [19]),
    .B(_02151_),
    .S(_02087_),
    .Z(_00832_)
  );
  MUX2_X1 _17787_ (
    .A(\rf[8] [20]),
    .B(_02152_),
    .S(_02087_),
    .Z(_00833_)
  );
  MUX2_X1 _17788_ (
    .A(\rf[8] [21]),
    .B(_02153_),
    .S(_02087_),
    .Z(_00834_)
  );
  MUX2_X1 _17789_ (
    .A(\rf[8] [22]),
    .B(_02154_),
    .S(_02087_),
    .Z(_00835_)
  );
  MUX2_X1 _17790_ (
    .A(\rf[8] [23]),
    .B(_02155_),
    .S(_02087_),
    .Z(_00836_)
  );
  MUX2_X1 _17791_ (
    .A(\rf[8] [24]),
    .B(_02156_),
    .S(_02087_),
    .Z(_00837_)
  );
  MUX2_X1 _17792_ (
    .A(\rf[8] [25]),
    .B(_02157_),
    .S(_02087_),
    .Z(_00838_)
  );
  MUX2_X1 _17793_ (
    .A(\rf[8] [26]),
    .B(_02158_),
    .S(_02087_),
    .Z(_00839_)
  );
  MUX2_X1 _17794_ (
    .A(\rf[8] [27]),
    .B(_02159_),
    .S(_02087_),
    .Z(_00840_)
  );
  MUX2_X1 _17795_ (
    .A(\rf[8] [28]),
    .B(_02160_),
    .S(_02087_),
    .Z(_00841_)
  );
  MUX2_X1 _17796_ (
    .A(\rf[8] [29]),
    .B(_02161_),
    .S(_02087_),
    .Z(_00842_)
  );
  MUX2_X1 _17797_ (
    .A(\rf[8] [30]),
    .B(_02162_),
    .S(_02087_),
    .Z(_00843_)
  );
  MUX2_X1 _17798_ (
    .A(\rf[16] [0]),
    .B(_02132_),
    .S(_02123_),
    .Z(_00844_)
  );
  MUX2_X1 _17799_ (
    .A(\rf[16] [1]),
    .B(_02133_),
    .S(_02123_),
    .Z(_00845_)
  );
  MUX2_X1 _17800_ (
    .A(\rf[16] [2]),
    .B(_02134_),
    .S(_02123_),
    .Z(_00846_)
  );
  MUX2_X1 _17801_ (
    .A(\rf[16] [3]),
    .B(_02135_),
    .S(_02123_),
    .Z(_00847_)
  );
  MUX2_X1 _17802_ (
    .A(\rf[16] [4]),
    .B(_02136_),
    .S(_02123_),
    .Z(_00848_)
  );
  MUX2_X1 _17803_ (
    .A(\rf[16] [5]),
    .B(_02137_),
    .S(_02123_),
    .Z(_00849_)
  );
  MUX2_X1 _17804_ (
    .A(\rf[16] [6]),
    .B(_02138_),
    .S(_02123_),
    .Z(_00850_)
  );
  MUX2_X1 _17805_ (
    .A(\rf[16] [7]),
    .B(_02139_),
    .S(_02123_),
    .Z(_00851_)
  );
  MUX2_X1 _17806_ (
    .A(\rf[16] [8]),
    .B(_02140_),
    .S(_02123_),
    .Z(_00852_)
  );
  MUX2_X1 _17807_ (
    .A(\rf[16] [9]),
    .B(_02141_),
    .S(_02123_),
    .Z(_00853_)
  );
  MUX2_X1 _17808_ (
    .A(\rf[16] [10]),
    .B(_02142_),
    .S(_02123_),
    .Z(_00854_)
  );
  MUX2_X1 _17809_ (
    .A(\rf[16] [11]),
    .B(_02143_),
    .S(_02123_),
    .Z(_00855_)
  );
  MUX2_X1 _17810_ (
    .A(\rf[16] [12]),
    .B(_02144_),
    .S(_02123_),
    .Z(_00856_)
  );
  MUX2_X1 _17811_ (
    .A(\rf[16] [13]),
    .B(_02145_),
    .S(_02123_),
    .Z(_00857_)
  );
  MUX2_X1 _17812_ (
    .A(\rf[16] [14]),
    .B(_02146_),
    .S(_02123_),
    .Z(_00858_)
  );
  MUX2_X1 _17813_ (
    .A(\rf[16] [15]),
    .B(_02147_),
    .S(_02123_),
    .Z(_00859_)
  );
  MUX2_X1 _17814_ (
    .A(\rf[16] [16]),
    .B(_02148_),
    .S(_02123_),
    .Z(_00860_)
  );
  MUX2_X1 _17815_ (
    .A(\rf[16] [17]),
    .B(_02149_),
    .S(_02123_),
    .Z(_00861_)
  );
  MUX2_X1 _17816_ (
    .A(\rf[16] [18]),
    .B(_02150_),
    .S(_02123_),
    .Z(_00862_)
  );
  MUX2_X1 _17817_ (
    .A(\rf[16] [19]),
    .B(_02151_),
    .S(_02123_),
    .Z(_00863_)
  );
  MUX2_X1 _17818_ (
    .A(\rf[16] [20]),
    .B(_02152_),
    .S(_02123_),
    .Z(_00864_)
  );
  MUX2_X1 _17819_ (
    .A(\rf[16] [21]),
    .B(_02153_),
    .S(_02123_),
    .Z(_00865_)
  );
  MUX2_X1 _17820_ (
    .A(\rf[16] [22]),
    .B(_02154_),
    .S(_02123_),
    .Z(_00866_)
  );
  MUX2_X1 _17821_ (
    .A(\rf[16] [23]),
    .B(_02155_),
    .S(_02123_),
    .Z(_00867_)
  );
  MUX2_X1 _17822_ (
    .A(\rf[16] [24]),
    .B(_02156_),
    .S(_02123_),
    .Z(_00868_)
  );
  MUX2_X1 _17823_ (
    .A(\rf[16] [25]),
    .B(_02157_),
    .S(_02123_),
    .Z(_00869_)
  );
  MUX2_X1 _17824_ (
    .A(\rf[16] [26]),
    .B(_02158_),
    .S(_02123_),
    .Z(_00870_)
  );
  MUX2_X1 _17825_ (
    .A(\rf[16] [27]),
    .B(_02159_),
    .S(_02123_),
    .Z(_00871_)
  );
  MUX2_X1 _17826_ (
    .A(\rf[16] [28]),
    .B(_02160_),
    .S(_02123_),
    .Z(_00872_)
  );
  MUX2_X1 _17827_ (
    .A(\rf[16] [29]),
    .B(_02161_),
    .S(_02123_),
    .Z(_00873_)
  );
  MUX2_X1 _17828_ (
    .A(\rf[16] [30]),
    .B(_02162_),
    .S(_02123_),
    .Z(_00874_)
  );
  MUX2_X1 _17829_ (
    .A(\rf[17] [0]),
    .B(_02132_),
    .S(_02122_),
    .Z(_00875_)
  );
  MUX2_X1 _17830_ (
    .A(\rf[17] [1]),
    .B(_02133_),
    .S(_02122_),
    .Z(_00876_)
  );
  MUX2_X1 _17831_ (
    .A(\rf[17] [2]),
    .B(_02134_),
    .S(_02122_),
    .Z(_00877_)
  );
  MUX2_X1 _17832_ (
    .A(\rf[17] [3]),
    .B(_02135_),
    .S(_02122_),
    .Z(_00878_)
  );
  MUX2_X1 _17833_ (
    .A(\rf[17] [4]),
    .B(_02136_),
    .S(_02122_),
    .Z(_00879_)
  );
  MUX2_X1 _17834_ (
    .A(\rf[17] [5]),
    .B(_02137_),
    .S(_02122_),
    .Z(_00880_)
  );
  MUX2_X1 _17835_ (
    .A(\rf[17] [6]),
    .B(_02138_),
    .S(_02122_),
    .Z(_00881_)
  );
  MUX2_X1 _17836_ (
    .A(\rf[17] [7]),
    .B(_02139_),
    .S(_02122_),
    .Z(_00882_)
  );
  MUX2_X1 _17837_ (
    .A(\rf[17] [8]),
    .B(_02140_),
    .S(_02122_),
    .Z(_00883_)
  );
  MUX2_X1 _17838_ (
    .A(\rf[17] [9]),
    .B(_02141_),
    .S(_02122_),
    .Z(_00884_)
  );
  MUX2_X1 _17839_ (
    .A(\rf[17] [10]),
    .B(_02142_),
    .S(_02122_),
    .Z(_00885_)
  );
  MUX2_X1 _17840_ (
    .A(\rf[17] [11]),
    .B(_02143_),
    .S(_02122_),
    .Z(_00886_)
  );
  MUX2_X1 _17841_ (
    .A(\rf[17] [12]),
    .B(_02144_),
    .S(_02122_),
    .Z(_00887_)
  );
  MUX2_X1 _17842_ (
    .A(\rf[17] [13]),
    .B(_02145_),
    .S(_02122_),
    .Z(_00888_)
  );
  MUX2_X1 _17843_ (
    .A(\rf[17] [14]),
    .B(_02146_),
    .S(_02122_),
    .Z(_00889_)
  );
  MUX2_X1 _17844_ (
    .A(\rf[17] [15]),
    .B(_02147_),
    .S(_02122_),
    .Z(_00890_)
  );
  MUX2_X1 _17845_ (
    .A(\rf[17] [16]),
    .B(_02148_),
    .S(_02122_),
    .Z(_00891_)
  );
  MUX2_X1 _17846_ (
    .A(\rf[17] [17]),
    .B(_02149_),
    .S(_02122_),
    .Z(_00892_)
  );
  MUX2_X1 _17847_ (
    .A(\rf[17] [18]),
    .B(_02150_),
    .S(_02122_),
    .Z(_00893_)
  );
  MUX2_X1 _17848_ (
    .A(\rf[17] [19]),
    .B(_02151_),
    .S(_02122_),
    .Z(_00894_)
  );
  MUX2_X1 _17849_ (
    .A(\rf[17] [20]),
    .B(_02152_),
    .S(_02122_),
    .Z(_00895_)
  );
  MUX2_X1 _17850_ (
    .A(\rf[17] [21]),
    .B(_02153_),
    .S(_02122_),
    .Z(_00896_)
  );
  MUX2_X1 _17851_ (
    .A(\rf[17] [22]),
    .B(_02154_),
    .S(_02122_),
    .Z(_00897_)
  );
  MUX2_X1 _17852_ (
    .A(\rf[17] [23]),
    .B(_02155_),
    .S(_02122_),
    .Z(_00898_)
  );
  MUX2_X1 _17853_ (
    .A(\rf[17] [24]),
    .B(_02156_),
    .S(_02122_),
    .Z(_00899_)
  );
  MUX2_X1 _17854_ (
    .A(\rf[17] [25]),
    .B(_02157_),
    .S(_02122_),
    .Z(_00900_)
  );
  MUX2_X1 _17855_ (
    .A(\rf[17] [26]),
    .B(_02158_),
    .S(_02122_),
    .Z(_00901_)
  );
  MUX2_X1 _17856_ (
    .A(\rf[17] [27]),
    .B(_02159_),
    .S(_02122_),
    .Z(_00902_)
  );
  MUX2_X1 _17857_ (
    .A(\rf[17] [28]),
    .B(_02160_),
    .S(_02122_),
    .Z(_00903_)
  );
  MUX2_X1 _17858_ (
    .A(\rf[17] [29]),
    .B(_02161_),
    .S(_02122_),
    .Z(_00904_)
  );
  MUX2_X1 _17859_ (
    .A(\rf[17] [30]),
    .B(_02162_),
    .S(_02122_),
    .Z(_00905_)
  );
  MUX2_X1 _17860_ (
    .A(\rf[10] [0]),
    .B(_02132_),
    .S(_02130_),
    .Z(_00906_)
  );
  MUX2_X1 _17861_ (
    .A(\rf[10] [1]),
    .B(_02133_),
    .S(_02130_),
    .Z(_00907_)
  );
  MUX2_X1 _17862_ (
    .A(\rf[10] [2]),
    .B(_02134_),
    .S(_02130_),
    .Z(_00908_)
  );
  MUX2_X1 _17863_ (
    .A(\rf[10] [3]),
    .B(_02135_),
    .S(_02130_),
    .Z(_00909_)
  );
  MUX2_X1 _17864_ (
    .A(\rf[10] [4]),
    .B(_02136_),
    .S(_02130_),
    .Z(_00910_)
  );
  MUX2_X1 _17865_ (
    .A(\rf[10] [5]),
    .B(_02137_),
    .S(_02130_),
    .Z(_00911_)
  );
  MUX2_X1 _17866_ (
    .A(\rf[10] [6]),
    .B(_02138_),
    .S(_02130_),
    .Z(_00912_)
  );
  MUX2_X1 _17867_ (
    .A(\rf[10] [7]),
    .B(_02139_),
    .S(_02130_),
    .Z(_00913_)
  );
  MUX2_X1 _17868_ (
    .A(\rf[10] [8]),
    .B(_02140_),
    .S(_02130_),
    .Z(_00914_)
  );
  MUX2_X1 _17869_ (
    .A(\rf[10] [9]),
    .B(_02141_),
    .S(_02130_),
    .Z(_00915_)
  );
  MUX2_X1 _17870_ (
    .A(\rf[10] [10]),
    .B(_02142_),
    .S(_02130_),
    .Z(_00916_)
  );
  MUX2_X1 _17871_ (
    .A(\rf[10] [11]),
    .B(_02143_),
    .S(_02130_),
    .Z(_00917_)
  );
  MUX2_X1 _17872_ (
    .A(\rf[10] [12]),
    .B(_02144_),
    .S(_02130_),
    .Z(_00918_)
  );
  MUX2_X1 _17873_ (
    .A(\rf[10] [13]),
    .B(_02145_),
    .S(_02130_),
    .Z(_00919_)
  );
  MUX2_X1 _17874_ (
    .A(\rf[10] [14]),
    .B(_02146_),
    .S(_02130_),
    .Z(_00920_)
  );
  MUX2_X1 _17875_ (
    .A(\rf[10] [15]),
    .B(_02147_),
    .S(_02130_),
    .Z(_00921_)
  );
  MUX2_X1 _17876_ (
    .A(\rf[10] [16]),
    .B(_02148_),
    .S(_02130_),
    .Z(_00922_)
  );
  MUX2_X1 _17877_ (
    .A(\rf[10] [17]),
    .B(_02149_),
    .S(_02130_),
    .Z(_00923_)
  );
  MUX2_X1 _17878_ (
    .A(\rf[10] [18]),
    .B(_02150_),
    .S(_02130_),
    .Z(_00924_)
  );
  MUX2_X1 _17879_ (
    .A(\rf[10] [19]),
    .B(_02151_),
    .S(_02130_),
    .Z(_00925_)
  );
  MUX2_X1 _17880_ (
    .A(\rf[10] [20]),
    .B(_02152_),
    .S(_02130_),
    .Z(_00926_)
  );
  MUX2_X1 _17881_ (
    .A(\rf[10] [21]),
    .B(_02153_),
    .S(_02130_),
    .Z(_00927_)
  );
  MUX2_X1 _17882_ (
    .A(\rf[10] [22]),
    .B(_02154_),
    .S(_02130_),
    .Z(_00928_)
  );
  MUX2_X1 _17883_ (
    .A(\rf[10] [23]),
    .B(_02155_),
    .S(_02130_),
    .Z(_00929_)
  );
  MUX2_X1 _17884_ (
    .A(\rf[10] [24]),
    .B(_02156_),
    .S(_02130_),
    .Z(_00930_)
  );
  MUX2_X1 _17885_ (
    .A(\rf[10] [25]),
    .B(_02157_),
    .S(_02130_),
    .Z(_00931_)
  );
  MUX2_X1 _17886_ (
    .A(\rf[10] [26]),
    .B(_02158_),
    .S(_02130_),
    .Z(_00932_)
  );
  MUX2_X1 _17887_ (
    .A(\rf[10] [27]),
    .B(_02159_),
    .S(_02130_),
    .Z(_00933_)
  );
  MUX2_X1 _17888_ (
    .A(\rf[10] [28]),
    .B(_02160_),
    .S(_02130_),
    .Z(_00934_)
  );
  MUX2_X1 _17889_ (
    .A(\rf[10] [29]),
    .B(_02161_),
    .S(_02130_),
    .Z(_00935_)
  );
  MUX2_X1 _17890_ (
    .A(\rf[10] [30]),
    .B(_02162_),
    .S(_02130_),
    .Z(_00936_)
  );
  MUX2_X1 _17891_ (
    .A(\rf[18] [0]),
    .B(_02132_),
    .S(_02121_),
    .Z(_00937_)
  );
  MUX2_X1 _17892_ (
    .A(\rf[18] [1]),
    .B(_02133_),
    .S(_02121_),
    .Z(_00938_)
  );
  MUX2_X1 _17893_ (
    .A(\rf[18] [2]),
    .B(_02134_),
    .S(_02121_),
    .Z(_00939_)
  );
  MUX2_X1 _17894_ (
    .A(\rf[18] [3]),
    .B(_02135_),
    .S(_02121_),
    .Z(_00940_)
  );
  MUX2_X1 _17895_ (
    .A(\rf[18] [4]),
    .B(_02136_),
    .S(_02121_),
    .Z(_00941_)
  );
  MUX2_X1 _17896_ (
    .A(\rf[18] [5]),
    .B(_02137_),
    .S(_02121_),
    .Z(_00942_)
  );
  MUX2_X1 _17897_ (
    .A(\rf[18] [6]),
    .B(_02138_),
    .S(_02121_),
    .Z(_00943_)
  );
  MUX2_X1 _17898_ (
    .A(\rf[18] [7]),
    .B(_02139_),
    .S(_02121_),
    .Z(_00944_)
  );
  MUX2_X1 _17899_ (
    .A(\rf[18] [8]),
    .B(_02140_),
    .S(_02121_),
    .Z(_00945_)
  );
  MUX2_X1 _17900_ (
    .A(\rf[18] [9]),
    .B(_02141_),
    .S(_02121_),
    .Z(_00946_)
  );
  MUX2_X1 _17901_ (
    .A(\rf[18] [10]),
    .B(_02142_),
    .S(_02121_),
    .Z(_00947_)
  );
  MUX2_X1 _17902_ (
    .A(\rf[18] [11]),
    .B(_02143_),
    .S(_02121_),
    .Z(_00948_)
  );
  MUX2_X1 _17903_ (
    .A(\rf[18] [12]),
    .B(_02144_),
    .S(_02121_),
    .Z(_00949_)
  );
  MUX2_X1 _17904_ (
    .A(\rf[18] [13]),
    .B(_02145_),
    .S(_02121_),
    .Z(_00950_)
  );
  MUX2_X1 _17905_ (
    .A(\rf[18] [14]),
    .B(_02146_),
    .S(_02121_),
    .Z(_00951_)
  );
  MUX2_X1 _17906_ (
    .A(\rf[18] [15]),
    .B(_02147_),
    .S(_02121_),
    .Z(_00952_)
  );
  MUX2_X1 _17907_ (
    .A(\rf[18] [16]),
    .B(_02148_),
    .S(_02121_),
    .Z(_00953_)
  );
  MUX2_X1 _17908_ (
    .A(\rf[18] [17]),
    .B(_02149_),
    .S(_02121_),
    .Z(_00954_)
  );
  MUX2_X1 _17909_ (
    .A(\rf[18] [18]),
    .B(_02150_),
    .S(_02121_),
    .Z(_00955_)
  );
  MUX2_X1 _17910_ (
    .A(\rf[18] [19]),
    .B(_02151_),
    .S(_02121_),
    .Z(_00956_)
  );
  MUX2_X1 _17911_ (
    .A(\rf[18] [20]),
    .B(_02152_),
    .S(_02121_),
    .Z(_00957_)
  );
  MUX2_X1 _17912_ (
    .A(\rf[18] [21]),
    .B(_02153_),
    .S(_02121_),
    .Z(_00958_)
  );
  MUX2_X1 _17913_ (
    .A(\rf[18] [22]),
    .B(_02154_),
    .S(_02121_),
    .Z(_00959_)
  );
  MUX2_X1 _17914_ (
    .A(\rf[18] [23]),
    .B(_02155_),
    .S(_02121_),
    .Z(_00960_)
  );
  MUX2_X1 _17915_ (
    .A(\rf[18] [24]),
    .B(_02156_),
    .S(_02121_),
    .Z(_00961_)
  );
  MUX2_X1 _17916_ (
    .A(\rf[18] [25]),
    .B(_02157_),
    .S(_02121_),
    .Z(_00962_)
  );
  MUX2_X1 _17917_ (
    .A(\rf[18] [26]),
    .B(_02158_),
    .S(_02121_),
    .Z(_00963_)
  );
  MUX2_X1 _17918_ (
    .A(\rf[18] [27]),
    .B(_02159_),
    .S(_02121_),
    .Z(_00964_)
  );
  MUX2_X1 _17919_ (
    .A(\rf[18] [28]),
    .B(_02160_),
    .S(_02121_),
    .Z(_00965_)
  );
  MUX2_X1 _17920_ (
    .A(\rf[18] [29]),
    .B(_02161_),
    .S(_02121_),
    .Z(_00966_)
  );
  MUX2_X1 _17921_ (
    .A(\rf[18] [30]),
    .B(_02162_),
    .S(_02121_),
    .Z(_00967_)
  );
  MUX2_X1 _17922_ (
    .A(\rf[11] [0]),
    .B(_02132_),
    .S(_02129_),
    .Z(_00968_)
  );
  MUX2_X1 _17923_ (
    .A(\rf[11] [1]),
    .B(_02133_),
    .S(_02129_),
    .Z(_00969_)
  );
  MUX2_X1 _17924_ (
    .A(\rf[11] [2]),
    .B(_04080_),
    .S(_02129_),
    .Z(_00970_)
  );
  MUX2_X1 _17925_ (
    .A(\rf[11] [3]),
    .B(_04150_),
    .S(_02129_),
    .Z(_00971_)
  );
  MUX2_X1 _17926_ (
    .A(\rf[11] [4]),
    .B(_04233_),
    .S(_02129_),
    .Z(_00972_)
  );
  MUX2_X1 _17927_ (
    .A(\rf[11] [5]),
    .B(_04305_),
    .S(_02129_),
    .Z(_00973_)
  );
  MUX2_X1 _17928_ (
    .A(\rf[11] [6]),
    .B(_02138_),
    .S(_02129_),
    .Z(_00974_)
  );
  MUX2_X1 _17929_ (
    .A(\rf[11] [7]),
    .B(_02139_),
    .S(_02129_),
    .Z(_00975_)
  );
  MUX2_X1 _17930_ (
    .A(\rf[11] [8]),
    .B(_02140_),
    .S(_02129_),
    .Z(_00976_)
  );
  MUX2_X1 _17931_ (
    .A(\rf[11] [9]),
    .B(_02141_),
    .S(_02129_),
    .Z(_00977_)
  );
  MUX2_X1 _17932_ (
    .A(\rf[11] [10]),
    .B(_02142_),
    .S(_02129_),
    .Z(_00978_)
  );
  MUX2_X1 _17933_ (
    .A(\rf[11] [11]),
    .B(_04742_),
    .S(_02129_),
    .Z(_00979_)
  );
  MUX2_X1 _17934_ (
    .A(\rf[11] [12]),
    .B(_04811_),
    .S(_02129_),
    .Z(_00980_)
  );
  MUX2_X1 _17935_ (
    .A(\rf[11] [13]),
    .B(_04882_),
    .S(_02129_),
    .Z(_00981_)
  );
  MUX2_X1 _17936_ (
    .A(\rf[11] [14]),
    .B(_02146_),
    .S(_02129_),
    .Z(_00982_)
  );
  MUX2_X1 _17937_ (
    .A(\rf[11] [15]),
    .B(_05027_),
    .S(_02129_),
    .Z(_00983_)
  );
  MUX2_X1 _17938_ (
    .A(\rf[11] [16]),
    .B(_02148_),
    .S(_02129_),
    .Z(_00984_)
  );
  MUX2_X1 _17939_ (
    .A(\rf[11] [17]),
    .B(_05170_),
    .S(_02129_),
    .Z(_00985_)
  );
  MUX2_X1 _17940_ (
    .A(\rf[11] [18]),
    .B(_02150_),
    .S(_02129_),
    .Z(_00986_)
  );
  MUX2_X1 _17941_ (
    .A(\rf[11] [19]),
    .B(_02151_),
    .S(_02129_),
    .Z(_00987_)
  );
  MUX2_X1 _17942_ (
    .A(\rf[11] [20]),
    .B(_05442_),
    .S(_02129_),
    .Z(_00988_)
  );
  MUX2_X1 _17943_ (
    .A(\rf[11] [21]),
    .B(_02153_),
    .S(_02129_),
    .Z(_00989_)
  );
  MUX2_X1 _17944_ (
    .A(\rf[11] [22]),
    .B(_05592_),
    .S(_02129_),
    .Z(_00990_)
  );
  MUX2_X1 _17945_ (
    .A(\rf[11] [23]),
    .B(_05657_),
    .S(_02129_),
    .Z(_00991_)
  );
  MUX2_X1 _17946_ (
    .A(\rf[11] [24]),
    .B(_05665_),
    .S(_02129_),
    .Z(_00992_)
  );
  MUX2_X1 _17947_ (
    .A(\rf[11] [25]),
    .B(_02157_),
    .S(_02129_),
    .Z(_00993_)
  );
  MUX2_X1 _17948_ (
    .A(\rf[11] [26]),
    .B(_05882_),
    .S(_02129_),
    .Z(_00994_)
  );
  MUX2_X1 _17949_ (
    .A(\rf[11] [27]),
    .B(_02159_),
    .S(_02129_),
    .Z(_00995_)
  );
  MUX2_X1 _17950_ (
    .A(\rf[11] [28]),
    .B(_02160_),
    .S(_02129_),
    .Z(_00996_)
  );
  MUX2_X1 _17951_ (
    .A(\rf[11] [29]),
    .B(_02161_),
    .S(_02129_),
    .Z(_00997_)
  );
  MUX2_X1 _17952_ (
    .A(\rf[11] [30]),
    .B(_06117_),
    .S(_02129_),
    .Z(_00998_)
  );
  MUX2_X1 _17953_ (
    .A(\rf[19] [0]),
    .B(_06266_),
    .S(_02120_),
    .Z(_00999_)
  );
  MUX2_X1 _17954_ (
    .A(\rf[19] [1]),
    .B(_02133_),
    .S(_02120_),
    .Z(_01000_)
  );
  MUX2_X1 _17955_ (
    .A(\rf[19] [2]),
    .B(_04080_),
    .S(_02120_),
    .Z(_01001_)
  );
  MUX2_X1 _17956_ (
    .A(\rf[19] [3]),
    .B(_04150_),
    .S(_02120_),
    .Z(_01002_)
  );
  MUX2_X1 _17957_ (
    .A(\rf[19] [4]),
    .B(_04233_),
    .S(_02120_),
    .Z(_01003_)
  );
  MUX2_X1 _17958_ (
    .A(\rf[19] [5]),
    .B(_04305_),
    .S(_02120_),
    .Z(_01004_)
  );
  MUX2_X1 _17959_ (
    .A(\rf[19] [6]),
    .B(_04379_),
    .S(_02120_),
    .Z(_01005_)
  );
  MUX2_X1 _17960_ (
    .A(\rf[19] [7]),
    .B(_02139_),
    .S(_02120_),
    .Z(_01006_)
  );
  MUX2_X1 _17961_ (
    .A(\rf[19] [8]),
    .B(_04521_),
    .S(_02120_),
    .Z(_01007_)
  );
  MUX2_X1 _17962_ (
    .A(\rf[19] [9]),
    .B(_04590_),
    .S(_02120_),
    .Z(_01008_)
  );
  MUX2_X1 _17963_ (
    .A(\rf[19] [10]),
    .B(_04659_),
    .S(_02120_),
    .Z(_01009_)
  );
  MUX2_X1 _17964_ (
    .A(\rf[19] [11]),
    .B(_04742_),
    .S(_02120_),
    .Z(_01010_)
  );
  MUX2_X1 _17965_ (
    .A(\rf[19] [12]),
    .B(_04811_),
    .S(_02120_),
    .Z(_01011_)
  );
  MUX2_X1 _17966_ (
    .A(\rf[19] [13]),
    .B(_04882_),
    .S(_02120_),
    .Z(_01012_)
  );
  MUX2_X1 _17967_ (
    .A(\rf[19] [14]),
    .B(_04953_),
    .S(_02120_),
    .Z(_01013_)
  );
  MUX2_X1 _17968_ (
    .A(\rf[19] [15]),
    .B(_05027_),
    .S(_02120_),
    .Z(_01014_)
  );
  MUX2_X1 _17969_ (
    .A(\rf[19] [16]),
    .B(_02148_),
    .S(_02120_),
    .Z(_01015_)
  );
  MUX2_X1 _17970_ (
    .A(\rf[19] [17]),
    .B(_05170_),
    .S(_02120_),
    .Z(_01016_)
  );
  MUX2_X1 _17971_ (
    .A(\rf[19] [18]),
    .B(_05302_),
    .S(_02120_),
    .Z(_01017_)
  );
  MUX2_X1 _17972_ (
    .A(\rf[19] [19]),
    .B(_02151_),
    .S(_02120_),
    .Z(_01018_)
  );
  MUX2_X1 _17973_ (
    .A(\rf[19] [20]),
    .B(_05442_),
    .S(_02120_),
    .Z(_01019_)
  );
  MUX2_X1 _17974_ (
    .A(\rf[19] [21]),
    .B(_02153_),
    .S(_02120_),
    .Z(_01020_)
  );
  MUX2_X1 _17975_ (
    .A(\rf[19] [22]),
    .B(_05592_),
    .S(_02120_),
    .Z(_01021_)
  );
  MUX2_X1 _17976_ (
    .A(\rf[19] [23]),
    .B(_05657_),
    .S(_02120_),
    .Z(_01022_)
  );
  MUX2_X1 _17977_ (
    .A(\rf[19] [24]),
    .B(_05665_),
    .S(_02120_),
    .Z(_01023_)
  );
  MUX2_X1 _17978_ (
    .A(\rf[19] [25]),
    .B(_02157_),
    .S(_02120_),
    .Z(_01024_)
  );
  MUX2_X1 _17979_ (
    .A(\rf[19] [26]),
    .B(_05882_),
    .S(_02120_),
    .Z(_01025_)
  );
  MUX2_X1 _17980_ (
    .A(\rf[19] [27]),
    .B(_05957_),
    .S(_02120_),
    .Z(_01026_)
  );
  MUX2_X1 _17981_ (
    .A(\rf[19] [28]),
    .B(_06032_),
    .S(_02120_),
    .Z(_01027_)
  );
  MUX2_X1 _17982_ (
    .A(\rf[19] [29]),
    .B(_06109_),
    .S(_02120_),
    .Z(_01028_)
  );
  MUX2_X1 _17983_ (
    .A(\rf[19] [30]),
    .B(_06117_),
    .S(_02120_),
    .Z(_01029_)
  );
  MUX2_X1 _17984_ (
    .A(\rf[12] [0]),
    .B(_02132_),
    .S(_02128_),
    .Z(_01030_)
  );
  MUX2_X1 _17985_ (
    .A(\rf[12] [1]),
    .B(_02133_),
    .S(_02128_),
    .Z(_01031_)
  );
  MUX2_X1 _17986_ (
    .A(\rf[12] [2]),
    .B(_02134_),
    .S(_02128_),
    .Z(_01032_)
  );
  MUX2_X1 _17987_ (
    .A(\rf[12] [3]),
    .B(_02135_),
    .S(_02128_),
    .Z(_01033_)
  );
  MUX2_X1 _17988_ (
    .A(\rf[12] [4]),
    .B(_02136_),
    .S(_02128_),
    .Z(_01034_)
  );
  MUX2_X1 _17989_ (
    .A(\rf[12] [5]),
    .B(_02137_),
    .S(_02128_),
    .Z(_01035_)
  );
  MUX2_X1 _17990_ (
    .A(\rf[12] [6]),
    .B(_02138_),
    .S(_02128_),
    .Z(_01036_)
  );
  MUX2_X1 _17991_ (
    .A(\rf[12] [7]),
    .B(_02139_),
    .S(_02128_),
    .Z(_01037_)
  );
  MUX2_X1 _17992_ (
    .A(\rf[12] [8]),
    .B(_02140_),
    .S(_02128_),
    .Z(_01038_)
  );
  MUX2_X1 _17993_ (
    .A(\rf[12] [9]),
    .B(_02141_),
    .S(_02128_),
    .Z(_01039_)
  );
  MUX2_X1 _17994_ (
    .A(\rf[12] [10]),
    .B(_02142_),
    .S(_02128_),
    .Z(_01040_)
  );
  MUX2_X1 _17995_ (
    .A(\rf[12] [11]),
    .B(_02143_),
    .S(_02128_),
    .Z(_01041_)
  );
  MUX2_X1 _17996_ (
    .A(\rf[12] [12]),
    .B(_02144_),
    .S(_02128_),
    .Z(_01042_)
  );
  MUX2_X1 _17997_ (
    .A(\rf[12] [13]),
    .B(_02145_),
    .S(_02128_),
    .Z(_01043_)
  );
  MUX2_X1 _17998_ (
    .A(\rf[12] [14]),
    .B(_02146_),
    .S(_02128_),
    .Z(_01044_)
  );
  MUX2_X1 _17999_ (
    .A(\rf[12] [15]),
    .B(_02147_),
    .S(_02128_),
    .Z(_01045_)
  );
  MUX2_X1 _18000_ (
    .A(\rf[12] [16]),
    .B(_02148_),
    .S(_02128_),
    .Z(_01046_)
  );
  MUX2_X1 _18001_ (
    .A(\rf[12] [17]),
    .B(_02149_),
    .S(_02128_),
    .Z(_01047_)
  );
  MUX2_X1 _18002_ (
    .A(\rf[12] [18]),
    .B(_02150_),
    .S(_02128_),
    .Z(_01048_)
  );
  MUX2_X1 _18003_ (
    .A(\rf[12] [19]),
    .B(_02151_),
    .S(_02128_),
    .Z(_01049_)
  );
  MUX2_X1 _18004_ (
    .A(\rf[12] [20]),
    .B(_02152_),
    .S(_02128_),
    .Z(_01050_)
  );
  MUX2_X1 _18005_ (
    .A(\rf[12] [21]),
    .B(_02153_),
    .S(_02128_),
    .Z(_01051_)
  );
  MUX2_X1 _18006_ (
    .A(\rf[12] [22]),
    .B(_02154_),
    .S(_02128_),
    .Z(_01052_)
  );
  MUX2_X1 _18007_ (
    .A(\rf[12] [23]),
    .B(_02155_),
    .S(_02128_),
    .Z(_01053_)
  );
  MUX2_X1 _18008_ (
    .A(\rf[12] [24]),
    .B(_02156_),
    .S(_02128_),
    .Z(_01054_)
  );
  MUX2_X1 _18009_ (
    .A(\rf[12] [25]),
    .B(_02157_),
    .S(_02128_),
    .Z(_01055_)
  );
  MUX2_X1 _18010_ (
    .A(\rf[12] [26]),
    .B(_02158_),
    .S(_02128_),
    .Z(_01056_)
  );
  MUX2_X1 _18011_ (
    .A(\rf[12] [27]),
    .B(_02159_),
    .S(_02128_),
    .Z(_01057_)
  );
  MUX2_X1 _18012_ (
    .A(\rf[12] [28]),
    .B(_02160_),
    .S(_02128_),
    .Z(_01058_)
  );
  MUX2_X1 _18013_ (
    .A(\rf[12] [29]),
    .B(_02161_),
    .S(_02128_),
    .Z(_01059_)
  );
  MUX2_X1 _18014_ (
    .A(\rf[12] [30]),
    .B(_02162_),
    .S(_02128_),
    .Z(_01060_)
  );
  MUX2_X1 _18015_ (
    .A(\rf[20] [0]),
    .B(_02132_),
    .S(_02117_),
    .Z(_01061_)
  );
  MUX2_X1 _18016_ (
    .A(\rf[20] [1]),
    .B(_02133_),
    .S(_02117_),
    .Z(_01062_)
  );
  MUX2_X1 _18017_ (
    .A(\rf[20] [2]),
    .B(_02134_),
    .S(_02117_),
    .Z(_01063_)
  );
  MUX2_X1 _18018_ (
    .A(\rf[20] [3]),
    .B(_02135_),
    .S(_02117_),
    .Z(_01064_)
  );
  MUX2_X1 _18019_ (
    .A(\rf[20] [4]),
    .B(_02136_),
    .S(_02117_),
    .Z(_01065_)
  );
  MUX2_X1 _18020_ (
    .A(\rf[20] [5]),
    .B(_02137_),
    .S(_02117_),
    .Z(_01066_)
  );
  MUX2_X1 _18021_ (
    .A(\rf[20] [6]),
    .B(_02138_),
    .S(_02117_),
    .Z(_01067_)
  );
  MUX2_X1 _18022_ (
    .A(\rf[20] [7]),
    .B(_02139_),
    .S(_02117_),
    .Z(_01068_)
  );
  MUX2_X1 _18023_ (
    .A(\rf[20] [8]),
    .B(_02140_),
    .S(_02117_),
    .Z(_01069_)
  );
  MUX2_X1 _18024_ (
    .A(\rf[20] [9]),
    .B(_02141_),
    .S(_02117_),
    .Z(_01070_)
  );
  MUX2_X1 _18025_ (
    .A(\rf[20] [10]),
    .B(_02142_),
    .S(_02117_),
    .Z(_01071_)
  );
  MUX2_X1 _18026_ (
    .A(\rf[20] [11]),
    .B(_02143_),
    .S(_02117_),
    .Z(_01072_)
  );
  MUX2_X1 _18027_ (
    .A(\rf[20] [12]),
    .B(_02144_),
    .S(_02117_),
    .Z(_01073_)
  );
  MUX2_X1 _18028_ (
    .A(\rf[20] [13]),
    .B(_02145_),
    .S(_02117_),
    .Z(_01074_)
  );
  MUX2_X1 _18029_ (
    .A(\rf[20] [14]),
    .B(_02146_),
    .S(_02117_),
    .Z(_01075_)
  );
  MUX2_X1 _18030_ (
    .A(\rf[20] [15]),
    .B(_02147_),
    .S(_02117_),
    .Z(_01076_)
  );
  MUX2_X1 _18031_ (
    .A(\rf[20] [16]),
    .B(_02148_),
    .S(_02117_),
    .Z(_01077_)
  );
  MUX2_X1 _18032_ (
    .A(\rf[20] [17]),
    .B(_02149_),
    .S(_02117_),
    .Z(_01078_)
  );
  MUX2_X1 _18033_ (
    .A(\rf[20] [18]),
    .B(_02150_),
    .S(_02117_),
    .Z(_01079_)
  );
  MUX2_X1 _18034_ (
    .A(\rf[20] [19]),
    .B(_02151_),
    .S(_02117_),
    .Z(_01080_)
  );
  MUX2_X1 _18035_ (
    .A(\rf[20] [20]),
    .B(_02152_),
    .S(_02117_),
    .Z(_01081_)
  );
  MUX2_X1 _18036_ (
    .A(\rf[20] [21]),
    .B(_02153_),
    .S(_02117_),
    .Z(_01082_)
  );
  MUX2_X1 _18037_ (
    .A(\rf[20] [22]),
    .B(_02154_),
    .S(_02117_),
    .Z(_01083_)
  );
  MUX2_X1 _18038_ (
    .A(\rf[20] [23]),
    .B(_02155_),
    .S(_02117_),
    .Z(_01084_)
  );
  MUX2_X1 _18039_ (
    .A(\rf[20] [24]),
    .B(_02156_),
    .S(_02117_),
    .Z(_01085_)
  );
  MUX2_X1 _18040_ (
    .A(\rf[20] [25]),
    .B(_02157_),
    .S(_02117_),
    .Z(_01086_)
  );
  MUX2_X1 _18041_ (
    .A(\rf[20] [26]),
    .B(_02158_),
    .S(_02117_),
    .Z(_01087_)
  );
  MUX2_X1 _18042_ (
    .A(\rf[20] [27]),
    .B(_02159_),
    .S(_02117_),
    .Z(_01088_)
  );
  MUX2_X1 _18043_ (
    .A(\rf[20] [28]),
    .B(_02160_),
    .S(_02117_),
    .Z(_01089_)
  );
  MUX2_X1 _18044_ (
    .A(\rf[20] [29]),
    .B(_02161_),
    .S(_02117_),
    .Z(_01090_)
  );
  MUX2_X1 _18045_ (
    .A(\rf[20] [30]),
    .B(_02162_),
    .S(_02117_),
    .Z(_01091_)
  );
  MUX2_X1 _18046_ (
    .A(\rf[9] [0]),
    .B(_02132_),
    .S(_02082_),
    .Z(_01092_)
  );
  MUX2_X1 _18047_ (
    .A(\rf[9] [1]),
    .B(_02133_),
    .S(_02082_),
    .Z(_01093_)
  );
  MUX2_X1 _18048_ (
    .A(\rf[9] [2]),
    .B(_02134_),
    .S(_02082_),
    .Z(_01094_)
  );
  MUX2_X1 _18049_ (
    .A(\rf[9] [3]),
    .B(_02135_),
    .S(_02082_),
    .Z(_01095_)
  );
  MUX2_X1 _18050_ (
    .A(\rf[9] [4]),
    .B(_02136_),
    .S(_02082_),
    .Z(_01096_)
  );
  MUX2_X1 _18051_ (
    .A(\rf[9] [5]),
    .B(_02137_),
    .S(_02082_),
    .Z(_01097_)
  );
  MUX2_X1 _18052_ (
    .A(\rf[9] [6]),
    .B(_02138_),
    .S(_02082_),
    .Z(_01098_)
  );
  MUX2_X1 _18053_ (
    .A(\rf[9] [7]),
    .B(_02139_),
    .S(_02082_),
    .Z(_01099_)
  );
  MUX2_X1 _18054_ (
    .A(\rf[9] [8]),
    .B(_02140_),
    .S(_02082_),
    .Z(_01100_)
  );
  MUX2_X1 _18055_ (
    .A(\rf[9] [9]),
    .B(_02141_),
    .S(_02082_),
    .Z(_01101_)
  );
  MUX2_X1 _18056_ (
    .A(\rf[9] [10]),
    .B(_02142_),
    .S(_02082_),
    .Z(_01102_)
  );
  MUX2_X1 _18057_ (
    .A(\rf[9] [11]),
    .B(_02143_),
    .S(_02082_),
    .Z(_01103_)
  );
  MUX2_X1 _18058_ (
    .A(\rf[9] [12]),
    .B(_02144_),
    .S(_02082_),
    .Z(_01104_)
  );
  MUX2_X1 _18059_ (
    .A(\rf[9] [13]),
    .B(_02145_),
    .S(_02082_),
    .Z(_01105_)
  );
  MUX2_X1 _18060_ (
    .A(\rf[9] [14]),
    .B(_02146_),
    .S(_02082_),
    .Z(_01106_)
  );
  MUX2_X1 _18061_ (
    .A(\rf[9] [15]),
    .B(_02147_),
    .S(_02082_),
    .Z(_01107_)
  );
  MUX2_X1 _18062_ (
    .A(\rf[9] [16]),
    .B(_02148_),
    .S(_02082_),
    .Z(_01108_)
  );
  MUX2_X1 _18063_ (
    .A(\rf[9] [17]),
    .B(_02149_),
    .S(_02082_),
    .Z(_01109_)
  );
  MUX2_X1 _18064_ (
    .A(\rf[9] [18]),
    .B(_02150_),
    .S(_02082_),
    .Z(_01110_)
  );
  MUX2_X1 _18065_ (
    .A(\rf[9] [19]),
    .B(_02151_),
    .S(_02082_),
    .Z(_01111_)
  );
  MUX2_X1 _18066_ (
    .A(\rf[9] [20]),
    .B(_02152_),
    .S(_02082_),
    .Z(_01112_)
  );
  MUX2_X1 _18067_ (
    .A(\rf[9] [21]),
    .B(_02153_),
    .S(_02082_),
    .Z(_01113_)
  );
  MUX2_X1 _18068_ (
    .A(\rf[9] [22]),
    .B(_02154_),
    .S(_02082_),
    .Z(_01114_)
  );
  MUX2_X1 _18069_ (
    .A(\rf[9] [23]),
    .B(_02155_),
    .S(_02082_),
    .Z(_01115_)
  );
  MUX2_X1 _18070_ (
    .A(\rf[9] [24]),
    .B(_02156_),
    .S(_02082_),
    .Z(_01116_)
  );
  MUX2_X1 _18071_ (
    .A(\rf[9] [25]),
    .B(_02157_),
    .S(_02082_),
    .Z(_01117_)
  );
  MUX2_X1 _18072_ (
    .A(\rf[9] [26]),
    .B(_02158_),
    .S(_02082_),
    .Z(_01118_)
  );
  MUX2_X1 _18073_ (
    .A(\rf[9] [27]),
    .B(_02159_),
    .S(_02082_),
    .Z(_01119_)
  );
  MUX2_X1 _18074_ (
    .A(\rf[9] [28]),
    .B(_02160_),
    .S(_02082_),
    .Z(_01120_)
  );
  MUX2_X1 _18075_ (
    .A(\rf[9] [29]),
    .B(_02161_),
    .S(_02082_),
    .Z(_01121_)
  );
  MUX2_X1 _18076_ (
    .A(\rf[9] [30]),
    .B(_02162_),
    .S(_02082_),
    .Z(_01122_)
  );
  MUX2_X1 _18077_ (
    .A(\rf[21] [0]),
    .B(_02132_),
    .S(_02116_),
    .Z(_01123_)
  );
  MUX2_X1 _18078_ (
    .A(\rf[21] [1]),
    .B(_02133_),
    .S(_02116_),
    .Z(_01124_)
  );
  MUX2_X1 _18079_ (
    .A(\rf[21] [2]),
    .B(_02134_),
    .S(_02116_),
    .Z(_01125_)
  );
  MUX2_X1 _18080_ (
    .A(\rf[21] [3]),
    .B(_02135_),
    .S(_02116_),
    .Z(_01126_)
  );
  MUX2_X1 _18081_ (
    .A(\rf[21] [4]),
    .B(_02136_),
    .S(_02116_),
    .Z(_01127_)
  );
  MUX2_X1 _18082_ (
    .A(\rf[21] [5]),
    .B(_02137_),
    .S(_02116_),
    .Z(_01128_)
  );
  MUX2_X1 _18083_ (
    .A(\rf[21] [6]),
    .B(_02138_),
    .S(_02116_),
    .Z(_01129_)
  );
  MUX2_X1 _18084_ (
    .A(\rf[21] [7]),
    .B(_02139_),
    .S(_02116_),
    .Z(_01130_)
  );
  MUX2_X1 _18085_ (
    .A(\rf[21] [8]),
    .B(_02140_),
    .S(_02116_),
    .Z(_01131_)
  );
  MUX2_X1 _18086_ (
    .A(\rf[21] [9]),
    .B(_02141_),
    .S(_02116_),
    .Z(_01132_)
  );
  MUX2_X1 _18087_ (
    .A(\rf[21] [10]),
    .B(_02142_),
    .S(_02116_),
    .Z(_01133_)
  );
  MUX2_X1 _18088_ (
    .A(\rf[21] [11]),
    .B(_02143_),
    .S(_02116_),
    .Z(_01134_)
  );
  MUX2_X1 _18089_ (
    .A(\rf[21] [12]),
    .B(_02144_),
    .S(_02116_),
    .Z(_01135_)
  );
  MUX2_X1 _18090_ (
    .A(\rf[21] [13]),
    .B(_02145_),
    .S(_02116_),
    .Z(_01136_)
  );
  MUX2_X1 _18091_ (
    .A(\rf[21] [14]),
    .B(_02146_),
    .S(_02116_),
    .Z(_01137_)
  );
  MUX2_X1 _18092_ (
    .A(\rf[21] [15]),
    .B(_02147_),
    .S(_02116_),
    .Z(_01138_)
  );
  MUX2_X1 _18093_ (
    .A(\rf[21] [16]),
    .B(_02148_),
    .S(_02116_),
    .Z(_01139_)
  );
  MUX2_X1 _18094_ (
    .A(\rf[21] [17]),
    .B(_02149_),
    .S(_02116_),
    .Z(_01140_)
  );
  MUX2_X1 _18095_ (
    .A(\rf[21] [18]),
    .B(_02150_),
    .S(_02116_),
    .Z(_01141_)
  );
  MUX2_X1 _18096_ (
    .A(\rf[21] [19]),
    .B(_02151_),
    .S(_02116_),
    .Z(_01142_)
  );
  MUX2_X1 _18097_ (
    .A(\rf[21] [20]),
    .B(_02152_),
    .S(_02116_),
    .Z(_01143_)
  );
  MUX2_X1 _18098_ (
    .A(\rf[21] [21]),
    .B(_02153_),
    .S(_02116_),
    .Z(_01144_)
  );
  MUX2_X1 _18099_ (
    .A(\rf[21] [22]),
    .B(_02154_),
    .S(_02116_),
    .Z(_01145_)
  );
  MUX2_X1 _18100_ (
    .A(\rf[21] [23]),
    .B(_02155_),
    .S(_02116_),
    .Z(_01146_)
  );
  MUX2_X1 _18101_ (
    .A(\rf[21] [24]),
    .B(_02156_),
    .S(_02116_),
    .Z(_01147_)
  );
  MUX2_X1 _18102_ (
    .A(\rf[21] [25]),
    .B(_02157_),
    .S(_02116_),
    .Z(_01148_)
  );
  MUX2_X1 _18103_ (
    .A(\rf[21] [26]),
    .B(_02158_),
    .S(_02116_),
    .Z(_01149_)
  );
  MUX2_X1 _18104_ (
    .A(\rf[21] [27]),
    .B(_02159_),
    .S(_02116_),
    .Z(_01150_)
  );
  MUX2_X1 _18105_ (
    .A(\rf[21] [28]),
    .B(_02160_),
    .S(_02116_),
    .Z(_01151_)
  );
  MUX2_X1 _18106_ (
    .A(\rf[21] [29]),
    .B(_02161_),
    .S(_02116_),
    .Z(_01152_)
  );
  MUX2_X1 _18107_ (
    .A(\rf[21] [30]),
    .B(_02162_),
    .S(_02116_),
    .Z(_01153_)
  );
  MUX2_X1 _18108_ (
    .A(\rf[13] [0]),
    .B(_02132_),
    .S(_02127_),
    .Z(_01154_)
  );
  MUX2_X1 _18109_ (
    .A(\rf[13] [1]),
    .B(_02133_),
    .S(_02127_),
    .Z(_01155_)
  );
  MUX2_X1 _18110_ (
    .A(\rf[13] [2]),
    .B(_02134_),
    .S(_02127_),
    .Z(_01156_)
  );
  MUX2_X1 _18111_ (
    .A(\rf[13] [3]),
    .B(_02135_),
    .S(_02127_),
    .Z(_01157_)
  );
  MUX2_X1 _18112_ (
    .A(\rf[13] [4]),
    .B(_02136_),
    .S(_02127_),
    .Z(_01158_)
  );
  MUX2_X1 _18113_ (
    .A(\rf[13] [5]),
    .B(_02137_),
    .S(_02127_),
    .Z(_01159_)
  );
  MUX2_X1 _18114_ (
    .A(\rf[13] [6]),
    .B(_02138_),
    .S(_02127_),
    .Z(_01160_)
  );
  MUX2_X1 _18115_ (
    .A(\rf[13] [7]),
    .B(_02139_),
    .S(_02127_),
    .Z(_01161_)
  );
  MUX2_X1 _18116_ (
    .A(\rf[13] [8]),
    .B(_02140_),
    .S(_02127_),
    .Z(_01162_)
  );
  MUX2_X1 _18117_ (
    .A(\rf[13] [9]),
    .B(_02141_),
    .S(_02127_),
    .Z(_01163_)
  );
  MUX2_X1 _18118_ (
    .A(\rf[13] [10]),
    .B(_02142_),
    .S(_02127_),
    .Z(_01164_)
  );
  MUX2_X1 _18119_ (
    .A(\rf[13] [11]),
    .B(_02143_),
    .S(_02127_),
    .Z(_01165_)
  );
  MUX2_X1 _18120_ (
    .A(\rf[13] [12]),
    .B(_02144_),
    .S(_02127_),
    .Z(_01166_)
  );
  MUX2_X1 _18121_ (
    .A(\rf[13] [13]),
    .B(_02145_),
    .S(_02127_),
    .Z(_01167_)
  );
  MUX2_X1 _18122_ (
    .A(\rf[13] [14]),
    .B(_02146_),
    .S(_02127_),
    .Z(_01168_)
  );
  MUX2_X1 _18123_ (
    .A(\rf[13] [15]),
    .B(_02147_),
    .S(_02127_),
    .Z(_01169_)
  );
  MUX2_X1 _18124_ (
    .A(\rf[13] [16]),
    .B(_02148_),
    .S(_02127_),
    .Z(_01170_)
  );
  MUX2_X1 _18125_ (
    .A(\rf[13] [17]),
    .B(_02149_),
    .S(_02127_),
    .Z(_01171_)
  );
  MUX2_X1 _18126_ (
    .A(\rf[13] [18]),
    .B(_02150_),
    .S(_02127_),
    .Z(_01172_)
  );
  MUX2_X1 _18127_ (
    .A(\rf[13] [19]),
    .B(_02151_),
    .S(_02127_),
    .Z(_01173_)
  );
  MUX2_X1 _18128_ (
    .A(\rf[13] [20]),
    .B(_02152_),
    .S(_02127_),
    .Z(_01174_)
  );
  MUX2_X1 _18129_ (
    .A(\rf[13] [21]),
    .B(_02153_),
    .S(_02127_),
    .Z(_01175_)
  );
  MUX2_X1 _18130_ (
    .A(\rf[13] [22]),
    .B(_02154_),
    .S(_02127_),
    .Z(_01176_)
  );
  MUX2_X1 _18131_ (
    .A(\rf[13] [23]),
    .B(_02155_),
    .S(_02127_),
    .Z(_01177_)
  );
  MUX2_X1 _18132_ (
    .A(\rf[13] [24]),
    .B(_02156_),
    .S(_02127_),
    .Z(_01178_)
  );
  MUX2_X1 _18133_ (
    .A(\rf[13] [25]),
    .B(_02157_),
    .S(_02127_),
    .Z(_01179_)
  );
  MUX2_X1 _18134_ (
    .A(\rf[13] [26]),
    .B(_02158_),
    .S(_02127_),
    .Z(_01180_)
  );
  MUX2_X1 _18135_ (
    .A(\rf[13] [27]),
    .B(_02159_),
    .S(_02127_),
    .Z(_01181_)
  );
  MUX2_X1 _18136_ (
    .A(\rf[13] [28]),
    .B(_02160_),
    .S(_02127_),
    .Z(_01182_)
  );
  MUX2_X1 _18137_ (
    .A(\rf[13] [29]),
    .B(_02161_),
    .S(_02127_),
    .Z(_01183_)
  );
  MUX2_X1 _18138_ (
    .A(\rf[13] [30]),
    .B(_02162_),
    .S(_02127_),
    .Z(_01184_)
  );
  MUX2_X1 _18139_ (
    .A(\rf[28] [0]),
    .B(_02132_),
    .S(_02106_),
    .Z(_01185_)
  );
  MUX2_X1 _18140_ (
    .A(\rf[28] [1]),
    .B(_02133_),
    .S(_02106_),
    .Z(_01186_)
  );
  MUX2_X1 _18141_ (
    .A(\rf[28] [2]),
    .B(_02134_),
    .S(_02106_),
    .Z(_01187_)
  );
  MUX2_X1 _18142_ (
    .A(\rf[28] [3]),
    .B(_02135_),
    .S(_02106_),
    .Z(_01188_)
  );
  MUX2_X1 _18143_ (
    .A(\rf[28] [4]),
    .B(_02136_),
    .S(_02106_),
    .Z(_01189_)
  );
  MUX2_X1 _18144_ (
    .A(\rf[28] [5]),
    .B(_02137_),
    .S(_02106_),
    .Z(_01190_)
  );
  MUX2_X1 _18145_ (
    .A(\rf[28] [6]),
    .B(_02138_),
    .S(_02106_),
    .Z(_01191_)
  );
  MUX2_X1 _18146_ (
    .A(\rf[28] [7]),
    .B(_02139_),
    .S(_02106_),
    .Z(_01192_)
  );
  MUX2_X1 _18147_ (
    .A(\rf[28] [8]),
    .B(_02140_),
    .S(_02106_),
    .Z(_01193_)
  );
  MUX2_X1 _18148_ (
    .A(\rf[28] [9]),
    .B(_02141_),
    .S(_02106_),
    .Z(_01194_)
  );
  MUX2_X1 _18149_ (
    .A(\rf[28] [10]),
    .B(_02142_),
    .S(_02106_),
    .Z(_01195_)
  );
  MUX2_X1 _18150_ (
    .A(\rf[28] [11]),
    .B(_02143_),
    .S(_02106_),
    .Z(_01196_)
  );
  MUX2_X1 _18151_ (
    .A(\rf[28] [12]),
    .B(_02144_),
    .S(_02106_),
    .Z(_01197_)
  );
  MUX2_X1 _18152_ (
    .A(\rf[28] [13]),
    .B(_02145_),
    .S(_02106_),
    .Z(_01198_)
  );
  MUX2_X1 _18153_ (
    .A(\rf[28] [14]),
    .B(_02146_),
    .S(_02106_),
    .Z(_01199_)
  );
  MUX2_X1 _18154_ (
    .A(\rf[28] [15]),
    .B(_02147_),
    .S(_02106_),
    .Z(_01200_)
  );
  MUX2_X1 _18155_ (
    .A(\rf[28] [16]),
    .B(_02148_),
    .S(_02106_),
    .Z(_01201_)
  );
  MUX2_X1 _18156_ (
    .A(\rf[28] [17]),
    .B(_02149_),
    .S(_02106_),
    .Z(_01202_)
  );
  MUX2_X1 _18157_ (
    .A(\rf[28] [18]),
    .B(_02150_),
    .S(_02106_),
    .Z(_01203_)
  );
  MUX2_X1 _18158_ (
    .A(\rf[28] [19]),
    .B(_02151_),
    .S(_02106_),
    .Z(_01204_)
  );
  MUX2_X1 _18159_ (
    .A(\rf[28] [20]),
    .B(_02152_),
    .S(_02106_),
    .Z(_01205_)
  );
  MUX2_X1 _18160_ (
    .A(\rf[28] [21]),
    .B(_02153_),
    .S(_02106_),
    .Z(_01206_)
  );
  MUX2_X1 _18161_ (
    .A(\rf[28] [22]),
    .B(_02154_),
    .S(_02106_),
    .Z(_01207_)
  );
  MUX2_X1 _18162_ (
    .A(\rf[28] [23]),
    .B(_02155_),
    .S(_02106_),
    .Z(_01208_)
  );
  MUX2_X1 _18163_ (
    .A(\rf[28] [24]),
    .B(_02156_),
    .S(_02106_),
    .Z(_01209_)
  );
  MUX2_X1 _18164_ (
    .A(\rf[28] [25]),
    .B(_02157_),
    .S(_02106_),
    .Z(_01210_)
  );
  MUX2_X1 _18165_ (
    .A(\rf[28] [26]),
    .B(_02158_),
    .S(_02106_),
    .Z(_01211_)
  );
  MUX2_X1 _18166_ (
    .A(\rf[28] [27]),
    .B(_02159_),
    .S(_02106_),
    .Z(_01212_)
  );
  MUX2_X1 _18167_ (
    .A(\rf[28] [28]),
    .B(_02160_),
    .S(_02106_),
    .Z(_01213_)
  );
  MUX2_X1 _18168_ (
    .A(\rf[28] [29]),
    .B(_02161_),
    .S(_02106_),
    .Z(_01214_)
  );
  MUX2_X1 _18169_ (
    .A(\rf[28] [30]),
    .B(_02162_),
    .S(_02106_),
    .Z(_01215_)
  );
  MUX2_X1 _18170_ (
    .A(\rf[29] [0]),
    .B(_02132_),
    .S(_02104_),
    .Z(_01216_)
  );
  MUX2_X1 _18171_ (
    .A(\rf[29] [1]),
    .B(_02133_),
    .S(_02104_),
    .Z(_01217_)
  );
  MUX2_X1 _18172_ (
    .A(\rf[29] [2]),
    .B(_02134_),
    .S(_02104_),
    .Z(_01218_)
  );
  MUX2_X1 _18173_ (
    .A(\rf[29] [3]),
    .B(_02135_),
    .S(_02104_),
    .Z(_01219_)
  );
  MUX2_X1 _18174_ (
    .A(\rf[29] [4]),
    .B(_02136_),
    .S(_02104_),
    .Z(_01220_)
  );
  MUX2_X1 _18175_ (
    .A(\rf[29] [5]),
    .B(_02137_),
    .S(_02104_),
    .Z(_01221_)
  );
  MUX2_X1 _18176_ (
    .A(\rf[29] [6]),
    .B(_02138_),
    .S(_02104_),
    .Z(_01222_)
  );
  MUX2_X1 _18177_ (
    .A(\rf[29] [7]),
    .B(_02139_),
    .S(_02104_),
    .Z(_01223_)
  );
  MUX2_X1 _18178_ (
    .A(\rf[29] [8]),
    .B(_02140_),
    .S(_02104_),
    .Z(_01224_)
  );
  MUX2_X1 _18179_ (
    .A(\rf[29] [9]),
    .B(_02141_),
    .S(_02104_),
    .Z(_01225_)
  );
  MUX2_X1 _18180_ (
    .A(\rf[29] [10]),
    .B(_02142_),
    .S(_02104_),
    .Z(_01226_)
  );
  MUX2_X1 _18181_ (
    .A(\rf[29] [11]),
    .B(_02143_),
    .S(_02104_),
    .Z(_01227_)
  );
  MUX2_X1 _18182_ (
    .A(\rf[29] [12]),
    .B(_02144_),
    .S(_02104_),
    .Z(_01228_)
  );
  MUX2_X1 _18183_ (
    .A(\rf[29] [13]),
    .B(_02145_),
    .S(_02104_),
    .Z(_01229_)
  );
  MUX2_X1 _18184_ (
    .A(\rf[29] [14]),
    .B(_02146_),
    .S(_02104_),
    .Z(_01230_)
  );
  MUX2_X1 _18185_ (
    .A(\rf[29] [15]),
    .B(_02147_),
    .S(_02104_),
    .Z(_01231_)
  );
  MUX2_X1 _18186_ (
    .A(\rf[29] [16]),
    .B(_02148_),
    .S(_02104_),
    .Z(_01232_)
  );
  MUX2_X1 _18187_ (
    .A(\rf[29] [17]),
    .B(_02149_),
    .S(_02104_),
    .Z(_01233_)
  );
  MUX2_X1 _18188_ (
    .A(\rf[29] [18]),
    .B(_02150_),
    .S(_02104_),
    .Z(_01234_)
  );
  MUX2_X1 _18189_ (
    .A(\rf[29] [19]),
    .B(_02151_),
    .S(_02104_),
    .Z(_01235_)
  );
  MUX2_X1 _18190_ (
    .A(\rf[29] [20]),
    .B(_02152_),
    .S(_02104_),
    .Z(_01236_)
  );
  MUX2_X1 _18191_ (
    .A(\rf[29] [21]),
    .B(_02153_),
    .S(_02104_),
    .Z(_01237_)
  );
  MUX2_X1 _18192_ (
    .A(\rf[29] [22]),
    .B(_02154_),
    .S(_02104_),
    .Z(_01238_)
  );
  MUX2_X1 _18193_ (
    .A(\rf[29] [23]),
    .B(_02155_),
    .S(_02104_),
    .Z(_01239_)
  );
  MUX2_X1 _18194_ (
    .A(\rf[29] [24]),
    .B(_02156_),
    .S(_02104_),
    .Z(_01240_)
  );
  MUX2_X1 _18195_ (
    .A(\rf[29] [25]),
    .B(_02157_),
    .S(_02104_),
    .Z(_01241_)
  );
  MUX2_X1 _18196_ (
    .A(\rf[29] [26]),
    .B(_02158_),
    .S(_02104_),
    .Z(_01242_)
  );
  MUX2_X1 _18197_ (
    .A(\rf[29] [27]),
    .B(_02159_),
    .S(_02104_),
    .Z(_01243_)
  );
  MUX2_X1 _18198_ (
    .A(\rf[29] [28]),
    .B(_02160_),
    .S(_02104_),
    .Z(_01244_)
  );
  MUX2_X1 _18199_ (
    .A(\rf[29] [29]),
    .B(_02161_),
    .S(_02104_),
    .Z(_01245_)
  );
  MUX2_X1 _18200_ (
    .A(\rf[29] [30]),
    .B(_02162_),
    .S(_02104_),
    .Z(_01246_)
  );
  MUX2_X1 _18201_ (
    .A(\rf[30] [0]),
    .B(_02132_),
    .S(_02102_),
    .Z(_01247_)
  );
  MUX2_X1 _18202_ (
    .A(\rf[30] [1]),
    .B(_02133_),
    .S(_02102_),
    .Z(_01248_)
  );
  MUX2_X1 _18203_ (
    .A(\rf[30] [2]),
    .B(_02134_),
    .S(_02102_),
    .Z(_01249_)
  );
  MUX2_X1 _18204_ (
    .A(\rf[30] [3]),
    .B(_02135_),
    .S(_02102_),
    .Z(_01250_)
  );
  MUX2_X1 _18205_ (
    .A(\rf[30] [4]),
    .B(_02136_),
    .S(_02102_),
    .Z(_01251_)
  );
  MUX2_X1 _18206_ (
    .A(\rf[30] [5]),
    .B(_02137_),
    .S(_02102_),
    .Z(_01252_)
  );
  MUX2_X1 _18207_ (
    .A(\rf[30] [6]),
    .B(_02138_),
    .S(_02102_),
    .Z(_01253_)
  );
  MUX2_X1 _18208_ (
    .A(\rf[30] [7]),
    .B(_02139_),
    .S(_02102_),
    .Z(_01254_)
  );
  MUX2_X1 _18209_ (
    .A(\rf[30] [8]),
    .B(_02140_),
    .S(_02102_),
    .Z(_01255_)
  );
  MUX2_X1 _18210_ (
    .A(\rf[30] [9]),
    .B(_02141_),
    .S(_02102_),
    .Z(_01256_)
  );
  MUX2_X1 _18211_ (
    .A(\rf[30] [10]),
    .B(_02142_),
    .S(_02102_),
    .Z(_01257_)
  );
  MUX2_X1 _18212_ (
    .A(\rf[30] [11]),
    .B(_02143_),
    .S(_02102_),
    .Z(_01258_)
  );
  MUX2_X1 _18213_ (
    .A(\rf[30] [12]),
    .B(_02144_),
    .S(_02102_),
    .Z(_01259_)
  );
  MUX2_X1 _18214_ (
    .A(\rf[30] [13]),
    .B(_02145_),
    .S(_02102_),
    .Z(_01260_)
  );
  MUX2_X1 _18215_ (
    .A(\rf[30] [14]),
    .B(_02146_),
    .S(_02102_),
    .Z(_01261_)
  );
  MUX2_X1 _18216_ (
    .A(\rf[30] [15]),
    .B(_02147_),
    .S(_02102_),
    .Z(_01262_)
  );
  MUX2_X1 _18217_ (
    .A(\rf[30] [16]),
    .B(_02148_),
    .S(_02102_),
    .Z(_01263_)
  );
  MUX2_X1 _18218_ (
    .A(\rf[30] [17]),
    .B(_02149_),
    .S(_02102_),
    .Z(_01264_)
  );
  MUX2_X1 _18219_ (
    .A(\rf[30] [18]),
    .B(_02150_),
    .S(_02102_),
    .Z(_01265_)
  );
  MUX2_X1 _18220_ (
    .A(\rf[30] [19]),
    .B(_02151_),
    .S(_02102_),
    .Z(_01266_)
  );
  MUX2_X1 _18221_ (
    .A(\rf[30] [20]),
    .B(_02152_),
    .S(_02102_),
    .Z(_01267_)
  );
  MUX2_X1 _18222_ (
    .A(\rf[30] [21]),
    .B(_02153_),
    .S(_02102_),
    .Z(_01268_)
  );
  MUX2_X1 _18223_ (
    .A(\rf[30] [22]),
    .B(_02154_),
    .S(_02102_),
    .Z(_01269_)
  );
  MUX2_X1 _18224_ (
    .A(\rf[30] [23]),
    .B(_02155_),
    .S(_02102_),
    .Z(_01270_)
  );
  MUX2_X1 _18225_ (
    .A(\rf[30] [24]),
    .B(_02156_),
    .S(_02102_),
    .Z(_01271_)
  );
  MUX2_X1 _18226_ (
    .A(\rf[30] [25]),
    .B(_02157_),
    .S(_02102_),
    .Z(_01272_)
  );
  MUX2_X1 _18227_ (
    .A(\rf[30] [26]),
    .B(_02158_),
    .S(_02102_),
    .Z(_01273_)
  );
  MUX2_X1 _18228_ (
    .A(\rf[30] [27]),
    .B(_02159_),
    .S(_02102_),
    .Z(_01274_)
  );
  MUX2_X1 _18229_ (
    .A(\rf[30] [28]),
    .B(_02160_),
    .S(_02102_),
    .Z(_01275_)
  );
  MUX2_X1 _18230_ (
    .A(\rf[30] [29]),
    .B(_02161_),
    .S(_02102_),
    .Z(_01276_)
  );
  MUX2_X1 _18231_ (
    .A(\rf[30] [30]),
    .B(_02162_),
    .S(_02102_),
    .Z(_01277_)
  );
  MUX2_X1 _18232_ (
    .A(\rf[14] [0]),
    .B(_02132_),
    .S(_02126_),
    .Z(_01278_)
  );
  MUX2_X1 _18233_ (
    .A(\rf[14] [1]),
    .B(_02133_),
    .S(_02126_),
    .Z(_01279_)
  );
  MUX2_X1 _18234_ (
    .A(\rf[14] [2]),
    .B(_02134_),
    .S(_02126_),
    .Z(_01280_)
  );
  MUX2_X1 _18235_ (
    .A(\rf[14] [3]),
    .B(_02135_),
    .S(_02126_),
    .Z(_01281_)
  );
  MUX2_X1 _18236_ (
    .A(\rf[14] [4]),
    .B(_02136_),
    .S(_02126_),
    .Z(_01282_)
  );
  MUX2_X1 _18237_ (
    .A(\rf[14] [5]),
    .B(_02137_),
    .S(_02126_),
    .Z(_01283_)
  );
  MUX2_X1 _18238_ (
    .A(\rf[14] [6]),
    .B(_02138_),
    .S(_02126_),
    .Z(_01284_)
  );
  MUX2_X1 _18239_ (
    .A(\rf[14] [7]),
    .B(_02139_),
    .S(_02126_),
    .Z(_01285_)
  );
  MUX2_X1 _18240_ (
    .A(\rf[14] [8]),
    .B(_02140_),
    .S(_02126_),
    .Z(_01286_)
  );
  MUX2_X1 _18241_ (
    .A(\rf[14] [9]),
    .B(_02141_),
    .S(_02126_),
    .Z(_01287_)
  );
  MUX2_X1 _18242_ (
    .A(\rf[14] [10]),
    .B(_02142_),
    .S(_02126_),
    .Z(_01288_)
  );
  MUX2_X1 _18243_ (
    .A(\rf[14] [11]),
    .B(_02143_),
    .S(_02126_),
    .Z(_01289_)
  );
  MUX2_X1 _18244_ (
    .A(\rf[14] [12]),
    .B(_02144_),
    .S(_02126_),
    .Z(_01290_)
  );
  MUX2_X1 _18245_ (
    .A(\rf[14] [13]),
    .B(_02145_),
    .S(_02126_),
    .Z(_01291_)
  );
  MUX2_X1 _18246_ (
    .A(\rf[14] [14]),
    .B(_02146_),
    .S(_02126_),
    .Z(_01292_)
  );
  MUX2_X1 _18247_ (
    .A(\rf[14] [15]),
    .B(_02147_),
    .S(_02126_),
    .Z(_01293_)
  );
  MUX2_X1 _18248_ (
    .A(\rf[14] [16]),
    .B(_02148_),
    .S(_02126_),
    .Z(_01294_)
  );
  MUX2_X1 _18249_ (
    .A(\rf[14] [17]),
    .B(_02149_),
    .S(_02126_),
    .Z(_01295_)
  );
  MUX2_X1 _18250_ (
    .A(\rf[14] [18]),
    .B(_02150_),
    .S(_02126_),
    .Z(_01296_)
  );
  MUX2_X1 _18251_ (
    .A(\rf[14] [19]),
    .B(_02151_),
    .S(_02126_),
    .Z(_01297_)
  );
  MUX2_X1 _18252_ (
    .A(\rf[14] [20]),
    .B(_02152_),
    .S(_02126_),
    .Z(_01298_)
  );
  MUX2_X1 _18253_ (
    .A(\rf[14] [21]),
    .B(_02153_),
    .S(_02126_),
    .Z(_01299_)
  );
  MUX2_X1 _18254_ (
    .A(\rf[14] [22]),
    .B(_02154_),
    .S(_02126_),
    .Z(_01300_)
  );
  MUX2_X1 _18255_ (
    .A(\rf[14] [23]),
    .B(_02155_),
    .S(_02126_),
    .Z(_01301_)
  );
  MUX2_X1 _18256_ (
    .A(\rf[14] [24]),
    .B(_02156_),
    .S(_02126_),
    .Z(_01302_)
  );
  MUX2_X1 _18257_ (
    .A(\rf[14] [25]),
    .B(_02157_),
    .S(_02126_),
    .Z(_01303_)
  );
  MUX2_X1 _18258_ (
    .A(\rf[14] [26]),
    .B(_02158_),
    .S(_02126_),
    .Z(_01304_)
  );
  MUX2_X1 _18259_ (
    .A(\rf[14] [27]),
    .B(_02159_),
    .S(_02126_),
    .Z(_01305_)
  );
  MUX2_X1 _18260_ (
    .A(\rf[14] [28]),
    .B(_02160_),
    .S(_02126_),
    .Z(_01306_)
  );
  MUX2_X1 _18261_ (
    .A(\rf[14] [29]),
    .B(_02161_),
    .S(_02126_),
    .Z(_01307_)
  );
  MUX2_X1 _18262_ (
    .A(\rf[14] [30]),
    .B(_02162_),
    .S(_02126_),
    .Z(_01308_)
  );
  MUX2_X1 _18263_ (
    .A(\rf[22] [0]),
    .B(_02132_),
    .S(_02115_),
    .Z(_01309_)
  );
  MUX2_X1 _18264_ (
    .A(\rf[22] [1]),
    .B(_02133_),
    .S(_02115_),
    .Z(_01310_)
  );
  MUX2_X1 _18265_ (
    .A(\rf[22] [2]),
    .B(_02134_),
    .S(_02115_),
    .Z(_01311_)
  );
  MUX2_X1 _18266_ (
    .A(\rf[22] [3]),
    .B(_02135_),
    .S(_02115_),
    .Z(_01312_)
  );
  MUX2_X1 _18267_ (
    .A(\rf[22] [4]),
    .B(_02136_),
    .S(_02115_),
    .Z(_01313_)
  );
  MUX2_X1 _18268_ (
    .A(\rf[22] [5]),
    .B(_02137_),
    .S(_02115_),
    .Z(_01314_)
  );
  MUX2_X1 _18269_ (
    .A(\rf[22] [6]),
    .B(_02138_),
    .S(_02115_),
    .Z(_01315_)
  );
  MUX2_X1 _18270_ (
    .A(\rf[22] [7]),
    .B(_02139_),
    .S(_02115_),
    .Z(_01316_)
  );
  MUX2_X1 _18271_ (
    .A(\rf[22] [8]),
    .B(_02140_),
    .S(_02115_),
    .Z(_01317_)
  );
  MUX2_X1 _18272_ (
    .A(\rf[22] [9]),
    .B(_02141_),
    .S(_02115_),
    .Z(_01318_)
  );
  MUX2_X1 _18273_ (
    .A(\rf[22] [10]),
    .B(_02142_),
    .S(_02115_),
    .Z(_01319_)
  );
  MUX2_X1 _18274_ (
    .A(\rf[22] [11]),
    .B(_02143_),
    .S(_02115_),
    .Z(_01320_)
  );
  MUX2_X1 _18275_ (
    .A(\rf[22] [12]),
    .B(_02144_),
    .S(_02115_),
    .Z(_01321_)
  );
  MUX2_X1 _18276_ (
    .A(\rf[22] [13]),
    .B(_02145_),
    .S(_02115_),
    .Z(_01322_)
  );
  MUX2_X1 _18277_ (
    .A(\rf[22] [14]),
    .B(_02146_),
    .S(_02115_),
    .Z(_01323_)
  );
  MUX2_X1 _18278_ (
    .A(\rf[22] [15]),
    .B(_02147_),
    .S(_02115_),
    .Z(_01324_)
  );
  MUX2_X1 _18279_ (
    .A(\rf[22] [16]),
    .B(_02148_),
    .S(_02115_),
    .Z(_01325_)
  );
  MUX2_X1 _18280_ (
    .A(\rf[22] [17]),
    .B(_02149_),
    .S(_02115_),
    .Z(_01326_)
  );
  MUX2_X1 _18281_ (
    .A(\rf[22] [18]),
    .B(_02150_),
    .S(_02115_),
    .Z(_01327_)
  );
  MUX2_X1 _18282_ (
    .A(\rf[22] [19]),
    .B(_02151_),
    .S(_02115_),
    .Z(_01328_)
  );
  MUX2_X1 _18283_ (
    .A(\rf[22] [20]),
    .B(_02152_),
    .S(_02115_),
    .Z(_01329_)
  );
  MUX2_X1 _18284_ (
    .A(\rf[22] [21]),
    .B(_02153_),
    .S(_02115_),
    .Z(_01330_)
  );
  MUX2_X1 _18285_ (
    .A(\rf[22] [22]),
    .B(_02154_),
    .S(_02115_),
    .Z(_01331_)
  );
  MUX2_X1 _18286_ (
    .A(\rf[22] [23]),
    .B(_02155_),
    .S(_02115_),
    .Z(_01332_)
  );
  MUX2_X1 _18287_ (
    .A(\rf[22] [24]),
    .B(_02156_),
    .S(_02115_),
    .Z(_01333_)
  );
  MUX2_X1 _18288_ (
    .A(\rf[22] [25]),
    .B(_02157_),
    .S(_02115_),
    .Z(_01334_)
  );
  MUX2_X1 _18289_ (
    .A(\rf[22] [26]),
    .B(_02158_),
    .S(_02115_),
    .Z(_01335_)
  );
  MUX2_X1 _18290_ (
    .A(\rf[22] [27]),
    .B(_02159_),
    .S(_02115_),
    .Z(_01336_)
  );
  MUX2_X1 _18291_ (
    .A(\rf[22] [28]),
    .B(_02160_),
    .S(_02115_),
    .Z(_01337_)
  );
  MUX2_X1 _18292_ (
    .A(\rf[22] [29]),
    .B(_02161_),
    .S(_02115_),
    .Z(_01338_)
  );
  MUX2_X1 _18293_ (
    .A(\rf[22] [30]),
    .B(_02162_),
    .S(_02115_),
    .Z(_01339_)
  );
  MUX2_X1 _18294_ (
    .A(\rf[26] [0]),
    .B(_02132_),
    .S(_02109_),
    .Z(_01340_)
  );
  MUX2_X1 _18295_ (
    .A(\rf[26] [1]),
    .B(_02133_),
    .S(_02109_),
    .Z(_01341_)
  );
  MUX2_X1 _18296_ (
    .A(\rf[26] [2]),
    .B(_02134_),
    .S(_02109_),
    .Z(_01342_)
  );
  MUX2_X1 _18297_ (
    .A(\rf[26] [3]),
    .B(_02135_),
    .S(_02109_),
    .Z(_01343_)
  );
  MUX2_X1 _18298_ (
    .A(\rf[26] [4]),
    .B(_02136_),
    .S(_02109_),
    .Z(_01344_)
  );
  MUX2_X1 _18299_ (
    .A(\rf[26] [5]),
    .B(_02137_),
    .S(_02109_),
    .Z(_01345_)
  );
  MUX2_X1 _18300_ (
    .A(\rf[26] [6]),
    .B(_02138_),
    .S(_02109_),
    .Z(_01346_)
  );
  MUX2_X1 _18301_ (
    .A(\rf[26] [7]),
    .B(_02139_),
    .S(_02109_),
    .Z(_01347_)
  );
  MUX2_X1 _18302_ (
    .A(\rf[26] [8]),
    .B(_02140_),
    .S(_02109_),
    .Z(_01348_)
  );
  MUX2_X1 _18303_ (
    .A(\rf[26] [9]),
    .B(_02141_),
    .S(_02109_),
    .Z(_01349_)
  );
  MUX2_X1 _18304_ (
    .A(\rf[26] [10]),
    .B(_02142_),
    .S(_02109_),
    .Z(_01350_)
  );
  MUX2_X1 _18305_ (
    .A(\rf[26] [11]),
    .B(_02143_),
    .S(_02109_),
    .Z(_01351_)
  );
  MUX2_X1 _18306_ (
    .A(\rf[26] [12]),
    .B(_02144_),
    .S(_02109_),
    .Z(_01352_)
  );
  MUX2_X1 _18307_ (
    .A(\rf[26] [13]),
    .B(_02145_),
    .S(_02109_),
    .Z(_01353_)
  );
  MUX2_X1 _18308_ (
    .A(\rf[26] [14]),
    .B(_02146_),
    .S(_02109_),
    .Z(_01354_)
  );
  MUX2_X1 _18309_ (
    .A(\rf[26] [15]),
    .B(_02147_),
    .S(_02109_),
    .Z(_01355_)
  );
  MUX2_X1 _18310_ (
    .A(\rf[26] [16]),
    .B(_02148_),
    .S(_02109_),
    .Z(_01356_)
  );
  MUX2_X1 _18311_ (
    .A(\rf[26] [17]),
    .B(_02149_),
    .S(_02109_),
    .Z(_01357_)
  );
  MUX2_X1 _18312_ (
    .A(\rf[26] [18]),
    .B(_02150_),
    .S(_02109_),
    .Z(_01358_)
  );
  MUX2_X1 _18313_ (
    .A(\rf[26] [19]),
    .B(_02151_),
    .S(_02109_),
    .Z(_01359_)
  );
  MUX2_X1 _18314_ (
    .A(\rf[26] [20]),
    .B(_02152_),
    .S(_02109_),
    .Z(_01360_)
  );
  MUX2_X1 _18315_ (
    .A(\rf[26] [21]),
    .B(_02153_),
    .S(_02109_),
    .Z(_01361_)
  );
  MUX2_X1 _18316_ (
    .A(\rf[26] [22]),
    .B(_02154_),
    .S(_02109_),
    .Z(_01362_)
  );
  MUX2_X1 _18317_ (
    .A(\rf[26] [23]),
    .B(_02155_),
    .S(_02109_),
    .Z(_01363_)
  );
  MUX2_X1 _18318_ (
    .A(\rf[26] [24]),
    .B(_02156_),
    .S(_02109_),
    .Z(_01364_)
  );
  MUX2_X1 _18319_ (
    .A(\rf[26] [25]),
    .B(_02157_),
    .S(_02109_),
    .Z(_01365_)
  );
  MUX2_X1 _18320_ (
    .A(\rf[26] [26]),
    .B(_02158_),
    .S(_02109_),
    .Z(_01366_)
  );
  MUX2_X1 _18321_ (
    .A(\rf[26] [27]),
    .B(_02159_),
    .S(_02109_),
    .Z(_01367_)
  );
  MUX2_X1 _18322_ (
    .A(\rf[26] [28]),
    .B(_02160_),
    .S(_02109_),
    .Z(_01368_)
  );
  MUX2_X1 _18323_ (
    .A(\rf[26] [29]),
    .B(_02161_),
    .S(_02109_),
    .Z(_01369_)
  );
  MUX2_X1 _18324_ (
    .A(\rf[26] [30]),
    .B(_02162_),
    .S(_02109_),
    .Z(_01370_)
  );
  MUX2_X1 _18325_ (
    .A(\rf[2] [0]),
    .B(_02132_),
    .S(_02103_),
    .Z(_01371_)
  );
  MUX2_X1 _18326_ (
    .A(\rf[2] [1]),
    .B(_02133_),
    .S(_02103_),
    .Z(_01372_)
  );
  MUX2_X1 _18327_ (
    .A(\rf[2] [2]),
    .B(_02134_),
    .S(_02103_),
    .Z(_01373_)
  );
  MUX2_X1 _18328_ (
    .A(\rf[2] [3]),
    .B(_02135_),
    .S(_02103_),
    .Z(_01374_)
  );
  MUX2_X1 _18329_ (
    .A(\rf[2] [4]),
    .B(_02136_),
    .S(_02103_),
    .Z(_01375_)
  );
  MUX2_X1 _18330_ (
    .A(\rf[2] [5]),
    .B(_02137_),
    .S(_02103_),
    .Z(_01376_)
  );
  MUX2_X1 _18331_ (
    .A(\rf[2] [6]),
    .B(_02138_),
    .S(_02103_),
    .Z(_01377_)
  );
  MUX2_X1 _18332_ (
    .A(\rf[2] [7]),
    .B(_02139_),
    .S(_02103_),
    .Z(_01378_)
  );
  MUX2_X1 _18333_ (
    .A(\rf[2] [8]),
    .B(_02140_),
    .S(_02103_),
    .Z(_01379_)
  );
  MUX2_X1 _18334_ (
    .A(\rf[2] [9]),
    .B(_02141_),
    .S(_02103_),
    .Z(_01380_)
  );
  MUX2_X1 _18335_ (
    .A(\rf[2] [10]),
    .B(_02142_),
    .S(_02103_),
    .Z(_01381_)
  );
  MUX2_X1 _18336_ (
    .A(\rf[2] [11]),
    .B(_02143_),
    .S(_02103_),
    .Z(_01382_)
  );
  MUX2_X1 _18337_ (
    .A(\rf[2] [12]),
    .B(_02144_),
    .S(_02103_),
    .Z(_01383_)
  );
  MUX2_X1 _18338_ (
    .A(\rf[2] [13]),
    .B(_02145_),
    .S(_02103_),
    .Z(_01384_)
  );
  MUX2_X1 _18339_ (
    .A(\rf[2] [14]),
    .B(_02146_),
    .S(_02103_),
    .Z(_01385_)
  );
  MUX2_X1 _18340_ (
    .A(\rf[2] [15]),
    .B(_02147_),
    .S(_02103_),
    .Z(_01386_)
  );
  MUX2_X1 _18341_ (
    .A(\rf[2] [16]),
    .B(_02148_),
    .S(_02103_),
    .Z(_01387_)
  );
  MUX2_X1 _18342_ (
    .A(\rf[2] [17]),
    .B(_02149_),
    .S(_02103_),
    .Z(_01388_)
  );
  MUX2_X1 _18343_ (
    .A(\rf[2] [18]),
    .B(_02150_),
    .S(_02103_),
    .Z(_01389_)
  );
  MUX2_X1 _18344_ (
    .A(\rf[2] [19]),
    .B(_02151_),
    .S(_02103_),
    .Z(_01390_)
  );
  MUX2_X1 _18345_ (
    .A(\rf[2] [20]),
    .B(_02152_),
    .S(_02103_),
    .Z(_01391_)
  );
  MUX2_X1 _18346_ (
    .A(\rf[2] [21]),
    .B(_02153_),
    .S(_02103_),
    .Z(_01392_)
  );
  MUX2_X1 _18347_ (
    .A(\rf[2] [22]),
    .B(_02154_),
    .S(_02103_),
    .Z(_01393_)
  );
  MUX2_X1 _18348_ (
    .A(\rf[2] [23]),
    .B(_02155_),
    .S(_02103_),
    .Z(_01394_)
  );
  MUX2_X1 _18349_ (
    .A(\rf[2] [24]),
    .B(_02156_),
    .S(_02103_),
    .Z(_01395_)
  );
  MUX2_X1 _18350_ (
    .A(\rf[2] [25]),
    .B(_02157_),
    .S(_02103_),
    .Z(_01396_)
  );
  MUX2_X1 _18351_ (
    .A(\rf[2] [26]),
    .B(_02158_),
    .S(_02103_),
    .Z(_01397_)
  );
  MUX2_X1 _18352_ (
    .A(\rf[2] [27]),
    .B(_02159_),
    .S(_02103_),
    .Z(_01398_)
  );
  MUX2_X1 _18353_ (
    .A(\rf[2] [28]),
    .B(_02160_),
    .S(_02103_),
    .Z(_01399_)
  );
  MUX2_X1 _18354_ (
    .A(\rf[2] [29]),
    .B(_02161_),
    .S(_02103_),
    .Z(_01400_)
  );
  MUX2_X1 _18355_ (
    .A(\rf[2] [30]),
    .B(_02162_),
    .S(_02103_),
    .Z(_01401_)
  );
  MUX2_X1 _18356_ (
    .A(\rf[27] [0]),
    .B(_02132_),
    .S(_02108_),
    .Z(_01402_)
  );
  MUX2_X1 _18357_ (
    .A(\rf[27] [1]),
    .B(_02133_),
    .S(_02108_),
    .Z(_01403_)
  );
  MUX2_X1 _18358_ (
    .A(\rf[27] [2]),
    .B(_02134_),
    .S(_02108_),
    .Z(_01404_)
  );
  MUX2_X1 _18359_ (
    .A(\rf[27] [3]),
    .B(_02135_),
    .S(_02108_),
    .Z(_01405_)
  );
  MUX2_X1 _18360_ (
    .A(\rf[27] [4]),
    .B(_02136_),
    .S(_02108_),
    .Z(_01406_)
  );
  MUX2_X1 _18361_ (
    .A(\rf[27] [5]),
    .B(_02137_),
    .S(_02108_),
    .Z(_01407_)
  );
  MUX2_X1 _18362_ (
    .A(\rf[27] [6]),
    .B(_02138_),
    .S(_02108_),
    .Z(_01408_)
  );
  MUX2_X1 _18363_ (
    .A(\rf[27] [7]),
    .B(_02139_),
    .S(_02108_),
    .Z(_01409_)
  );
  MUX2_X1 _18364_ (
    .A(\rf[27] [8]),
    .B(_02140_),
    .S(_02108_),
    .Z(_01410_)
  );
  MUX2_X1 _18365_ (
    .A(\rf[27] [9]),
    .B(_02141_),
    .S(_02108_),
    .Z(_01411_)
  );
  MUX2_X1 _18366_ (
    .A(\rf[27] [10]),
    .B(_02142_),
    .S(_02108_),
    .Z(_01412_)
  );
  MUX2_X1 _18367_ (
    .A(\rf[27] [11]),
    .B(_02143_),
    .S(_02108_),
    .Z(_01413_)
  );
  MUX2_X1 _18368_ (
    .A(\rf[27] [12]),
    .B(_02144_),
    .S(_02108_),
    .Z(_01414_)
  );
  MUX2_X1 _18369_ (
    .A(\rf[27] [13]),
    .B(_02145_),
    .S(_02108_),
    .Z(_01415_)
  );
  MUX2_X1 _18370_ (
    .A(\rf[27] [14]),
    .B(_02146_),
    .S(_02108_),
    .Z(_01416_)
  );
  MUX2_X1 _18371_ (
    .A(\rf[27] [15]),
    .B(_02147_),
    .S(_02108_),
    .Z(_01417_)
  );
  MUX2_X1 _18372_ (
    .A(\rf[27] [16]),
    .B(_02148_),
    .S(_02108_),
    .Z(_01418_)
  );
  MUX2_X1 _18373_ (
    .A(\rf[27] [17]),
    .B(_02149_),
    .S(_02108_),
    .Z(_01419_)
  );
  MUX2_X1 _18374_ (
    .A(\rf[27] [18]),
    .B(_02150_),
    .S(_02108_),
    .Z(_01420_)
  );
  MUX2_X1 _18375_ (
    .A(\rf[27] [19]),
    .B(_02151_),
    .S(_02108_),
    .Z(_01421_)
  );
  MUX2_X1 _18376_ (
    .A(\rf[27] [20]),
    .B(_02152_),
    .S(_02108_),
    .Z(_01422_)
  );
  MUX2_X1 _18377_ (
    .A(\rf[27] [21]),
    .B(_02153_),
    .S(_02108_),
    .Z(_01423_)
  );
  MUX2_X1 _18378_ (
    .A(\rf[27] [22]),
    .B(_02154_),
    .S(_02108_),
    .Z(_01424_)
  );
  MUX2_X1 _18379_ (
    .A(\rf[27] [23]),
    .B(_02155_),
    .S(_02108_),
    .Z(_01425_)
  );
  MUX2_X1 _18380_ (
    .A(\rf[27] [24]),
    .B(_02156_),
    .S(_02108_),
    .Z(_01426_)
  );
  MUX2_X1 _18381_ (
    .A(\rf[27] [25]),
    .B(_02157_),
    .S(_02108_),
    .Z(_01427_)
  );
  MUX2_X1 _18382_ (
    .A(\rf[27] [26]),
    .B(_02158_),
    .S(_02108_),
    .Z(_01428_)
  );
  MUX2_X1 _18383_ (
    .A(\rf[27] [27]),
    .B(_02159_),
    .S(_02108_),
    .Z(_01429_)
  );
  MUX2_X1 _18384_ (
    .A(\rf[27] [28]),
    .B(_02160_),
    .S(_02108_),
    .Z(_01430_)
  );
  MUX2_X1 _18385_ (
    .A(\rf[27] [29]),
    .B(_02161_),
    .S(_02108_),
    .Z(_01431_)
  );
  MUX2_X1 _18386_ (
    .A(\rf[27] [30]),
    .B(_02162_),
    .S(_02108_),
    .Z(_01432_)
  );
  MUX2_X1 _18387_ (
    .A(\rf[24] [0]),
    .B(_06266_),
    .S(_02111_),
    .Z(_01433_)
  );
  MUX2_X1 _18388_ (
    .A(\rf[24] [1]),
    .B(_06420_),
    .S(_02111_),
    .Z(_01434_)
  );
  MUX2_X1 _18389_ (
    .A(\rf[24] [2]),
    .B(_04080_),
    .S(_02111_),
    .Z(_01435_)
  );
  MUX2_X1 _18390_ (
    .A(\rf[24] [3]),
    .B(_04150_),
    .S(_02111_),
    .Z(_01436_)
  );
  MUX2_X1 _18391_ (
    .A(\rf[24] [4]),
    .B(_04233_),
    .S(_02111_),
    .Z(_01437_)
  );
  MUX2_X1 _18392_ (
    .A(\rf[24] [5]),
    .B(_04305_),
    .S(_02111_),
    .Z(_01438_)
  );
  MUX2_X1 _18393_ (
    .A(\rf[24] [6]),
    .B(_04379_),
    .S(_02111_),
    .Z(_01439_)
  );
  MUX2_X1 _18394_ (
    .A(\rf[24] [7]),
    .B(_04450_),
    .S(_02111_),
    .Z(_01440_)
  );
  MUX2_X1 _18395_ (
    .A(\rf[24] [8]),
    .B(_04521_),
    .S(_02111_),
    .Z(_01441_)
  );
  MUX2_X1 _18396_ (
    .A(\rf[24] [9]),
    .B(_04590_),
    .S(_02111_),
    .Z(_01442_)
  );
  MUX2_X1 _18397_ (
    .A(\rf[24] [10]),
    .B(_04659_),
    .S(_02111_),
    .Z(_01443_)
  );
  MUX2_X1 _18398_ (
    .A(\rf[24] [11]),
    .B(_04742_),
    .S(_02111_),
    .Z(_01444_)
  );
  MUX2_X1 _18399_ (
    .A(\rf[24] [12]),
    .B(_04811_),
    .S(_02111_),
    .Z(_01445_)
  );
  MUX2_X1 _18400_ (
    .A(\rf[24] [13]),
    .B(_04882_),
    .S(_02111_),
    .Z(_01446_)
  );
  MUX2_X1 _18401_ (
    .A(\rf[24] [14]),
    .B(_04953_),
    .S(_02111_),
    .Z(_01447_)
  );
  MUX2_X1 _18402_ (
    .A(\rf[24] [15]),
    .B(_05027_),
    .S(_02111_),
    .Z(_01448_)
  );
  MUX2_X1 _18403_ (
    .A(\rf[24] [16]),
    .B(_05095_),
    .S(_02111_),
    .Z(_01449_)
  );
  MUX2_X1 _18404_ (
    .A(\rf[24] [17]),
    .B(_05170_),
    .S(_02111_),
    .Z(_01450_)
  );
  MUX2_X1 _18405_ (
    .A(\rf[24] [18]),
    .B(_05302_),
    .S(_02111_),
    .Z(_01451_)
  );
  MUX2_X1 _18406_ (
    .A(\rf[24] [19]),
    .B(_05310_),
    .S(_02111_),
    .Z(_01452_)
  );
  MUX2_X1 _18407_ (
    .A(\rf[24] [20]),
    .B(_05442_),
    .S(_02111_),
    .Z(_01453_)
  );
  MUX2_X1 _18408_ (
    .A(\rf[24] [21]),
    .B(_05450_),
    .S(_02111_),
    .Z(_01454_)
  );
  MUX2_X1 _18409_ (
    .A(\rf[24] [22]),
    .B(_05592_),
    .S(_02111_),
    .Z(_01455_)
  );
  MUX2_X1 _18410_ (
    .A(\rf[24] [23]),
    .B(_05657_),
    .S(_02111_),
    .Z(_01456_)
  );
  MUX2_X1 _18411_ (
    .A(\rf[24] [24]),
    .B(_05665_),
    .S(_02111_),
    .Z(_01457_)
  );
  MUX2_X1 _18412_ (
    .A(\rf[24] [25]),
    .B(_05740_),
    .S(_02111_),
    .Z(_01458_)
  );
  MUX2_X1 _18413_ (
    .A(\rf[24] [26]),
    .B(_05882_),
    .S(_02111_),
    .Z(_01459_)
  );
  MUX2_X1 _18414_ (
    .A(\rf[24] [27]),
    .B(_05957_),
    .S(_02111_),
    .Z(_01460_)
  );
  MUX2_X1 _18415_ (
    .A(\rf[24] [28]),
    .B(_06032_),
    .S(_02111_),
    .Z(_01461_)
  );
  MUX2_X1 _18416_ (
    .A(\rf[24] [29]),
    .B(_06109_),
    .S(_02111_),
    .Z(_01462_)
  );
  MUX2_X1 _18417_ (
    .A(\rf[24] [30]),
    .B(_06117_),
    .S(_02111_),
    .Z(_01463_)
  );
  MUX2_X1 _18418_ (
    .A(\rf[5] [0]),
    .B(_02132_),
    .S(_02098_),
    .Z(_01464_)
  );
  MUX2_X1 _18419_ (
    .A(\rf[5] [1]),
    .B(_02133_),
    .S(_02098_),
    .Z(_01465_)
  );
  MUX2_X1 _18420_ (
    .A(\rf[5] [2]),
    .B(_02134_),
    .S(_02098_),
    .Z(_01466_)
  );
  MUX2_X1 _18421_ (
    .A(\rf[5] [3]),
    .B(_02135_),
    .S(_02098_),
    .Z(_01467_)
  );
  MUX2_X1 _18422_ (
    .A(\rf[5] [4]),
    .B(_02136_),
    .S(_02098_),
    .Z(_01468_)
  );
  MUX2_X1 _18423_ (
    .A(\rf[5] [5]),
    .B(_02137_),
    .S(_02098_),
    .Z(_01469_)
  );
  MUX2_X1 _18424_ (
    .A(\rf[5] [6]),
    .B(_02138_),
    .S(_02098_),
    .Z(_01470_)
  );
  MUX2_X1 _18425_ (
    .A(\rf[5] [7]),
    .B(_02139_),
    .S(_02098_),
    .Z(_01471_)
  );
  MUX2_X1 _18426_ (
    .A(\rf[5] [8]),
    .B(_02140_),
    .S(_02098_),
    .Z(_01472_)
  );
  MUX2_X1 _18427_ (
    .A(\rf[5] [9]),
    .B(_02141_),
    .S(_02098_),
    .Z(_01473_)
  );
  MUX2_X1 _18428_ (
    .A(\rf[5] [10]),
    .B(_02142_),
    .S(_02098_),
    .Z(_01474_)
  );
  MUX2_X1 _18429_ (
    .A(\rf[5] [11]),
    .B(_02143_),
    .S(_02098_),
    .Z(_01475_)
  );
  MUX2_X1 _18430_ (
    .A(\rf[5] [12]),
    .B(_02144_),
    .S(_02098_),
    .Z(_01476_)
  );
  MUX2_X1 _18431_ (
    .A(\rf[5] [13]),
    .B(_02145_),
    .S(_02098_),
    .Z(_01477_)
  );
  MUX2_X1 _18432_ (
    .A(\rf[5] [14]),
    .B(_02146_),
    .S(_02098_),
    .Z(_01478_)
  );
  MUX2_X1 _18433_ (
    .A(\rf[5] [15]),
    .B(_02147_),
    .S(_02098_),
    .Z(_01479_)
  );
  MUX2_X1 _18434_ (
    .A(\rf[5] [16]),
    .B(_02148_),
    .S(_02098_),
    .Z(_01480_)
  );
  MUX2_X1 _18435_ (
    .A(\rf[5] [17]),
    .B(_02149_),
    .S(_02098_),
    .Z(_01481_)
  );
  MUX2_X1 _18436_ (
    .A(\rf[5] [18]),
    .B(_02150_),
    .S(_02098_),
    .Z(_01482_)
  );
  MUX2_X1 _18437_ (
    .A(\rf[5] [19]),
    .B(_02151_),
    .S(_02098_),
    .Z(_01483_)
  );
  MUX2_X1 _18438_ (
    .A(\rf[5] [20]),
    .B(_02152_),
    .S(_02098_),
    .Z(_01484_)
  );
  MUX2_X1 _18439_ (
    .A(\rf[5] [21]),
    .B(_02153_),
    .S(_02098_),
    .Z(_01485_)
  );
  MUX2_X1 _18440_ (
    .A(\rf[5] [22]),
    .B(_02154_),
    .S(_02098_),
    .Z(_01486_)
  );
  MUX2_X1 _18441_ (
    .A(\rf[5] [23]),
    .B(_02155_),
    .S(_02098_),
    .Z(_01487_)
  );
  MUX2_X1 _18442_ (
    .A(\rf[5] [24]),
    .B(_02156_),
    .S(_02098_),
    .Z(_01488_)
  );
  MUX2_X1 _18443_ (
    .A(\rf[5] [25]),
    .B(_02157_),
    .S(_02098_),
    .Z(_01489_)
  );
  MUX2_X1 _18444_ (
    .A(\rf[5] [26]),
    .B(_02158_),
    .S(_02098_),
    .Z(_01490_)
  );
  MUX2_X1 _18445_ (
    .A(\rf[5] [27]),
    .B(_02159_),
    .S(_02098_),
    .Z(_01491_)
  );
  MUX2_X1 _18446_ (
    .A(\rf[5] [28]),
    .B(_02160_),
    .S(_02098_),
    .Z(_01492_)
  );
  MUX2_X1 _18447_ (
    .A(\rf[5] [29]),
    .B(_02161_),
    .S(_02098_),
    .Z(_01493_)
  );
  MUX2_X1 _18448_ (
    .A(\rf[5] [30]),
    .B(_02162_),
    .S(_02098_),
    .Z(_01494_)
  );
  MUX2_X1 _18449_ (
    .A(\rf[7] [0]),
    .B(_06266_),
    .S(_02095_),
    .Z(_01495_)
  );
  MUX2_X1 _18450_ (
    .A(\rf[7] [1]),
    .B(_02133_),
    .S(_02095_),
    .Z(_01496_)
  );
  MUX2_X1 _18451_ (
    .A(\rf[7] [2]),
    .B(_04080_),
    .S(_02095_),
    .Z(_01497_)
  );
  MUX2_X1 _18452_ (
    .A(\rf[7] [3]),
    .B(_04150_),
    .S(_02095_),
    .Z(_01498_)
  );
  MUX2_X1 _18453_ (
    .A(\rf[7] [4]),
    .B(_04233_),
    .S(_02095_),
    .Z(_01499_)
  );
  MUX2_X1 _18454_ (
    .A(\rf[7] [5]),
    .B(_04305_),
    .S(_02095_),
    .Z(_01500_)
  );
  MUX2_X1 _18455_ (
    .A(\rf[7] [6]),
    .B(_04379_),
    .S(_02095_),
    .Z(_01501_)
  );
  MUX2_X1 _18456_ (
    .A(\rf[7] [7]),
    .B(_02139_),
    .S(_02095_),
    .Z(_01502_)
  );
  MUX2_X1 _18457_ (
    .A(\rf[7] [8]),
    .B(_04521_),
    .S(_02095_),
    .Z(_01503_)
  );
  MUX2_X1 _18458_ (
    .A(\rf[7] [9]),
    .B(_04590_),
    .S(_02095_),
    .Z(_01504_)
  );
  MUX2_X1 _18459_ (
    .A(\rf[7] [10]),
    .B(_04659_),
    .S(_02095_),
    .Z(_01505_)
  );
  MUX2_X1 _18460_ (
    .A(\rf[7] [11]),
    .B(_04742_),
    .S(_02095_),
    .Z(_01506_)
  );
  MUX2_X1 _18461_ (
    .A(\rf[7] [12]),
    .B(_04811_),
    .S(_02095_),
    .Z(_01507_)
  );
  MUX2_X1 _18462_ (
    .A(\rf[7] [13]),
    .B(_04882_),
    .S(_02095_),
    .Z(_01508_)
  );
  MUX2_X1 _18463_ (
    .A(\rf[7] [14]),
    .B(_02146_),
    .S(_02095_),
    .Z(_01509_)
  );
  MUX2_X1 _18464_ (
    .A(\rf[7] [15]),
    .B(_05027_),
    .S(_02095_),
    .Z(_01510_)
  );
  MUX2_X1 _18465_ (
    .A(\rf[7] [16]),
    .B(_02148_),
    .S(_02095_),
    .Z(_01511_)
  );
  MUX2_X1 _18466_ (
    .A(\rf[7] [17]),
    .B(_05170_),
    .S(_02095_),
    .Z(_01512_)
  );
  MUX2_X1 _18467_ (
    .A(\rf[7] [18]),
    .B(_02150_),
    .S(_02095_),
    .Z(_01513_)
  );
  MUX2_X1 _18468_ (
    .A(\rf[7] [19]),
    .B(_02151_),
    .S(_02095_),
    .Z(_01514_)
  );
  MUX2_X1 _18469_ (
    .A(\rf[7] [20]),
    .B(_05442_),
    .S(_02095_),
    .Z(_01515_)
  );
  MUX2_X1 _18470_ (
    .A(\rf[7] [21]),
    .B(_05450_),
    .S(_02095_),
    .Z(_01516_)
  );
  MUX2_X1 _18471_ (
    .A(\rf[7] [22]),
    .B(_05592_),
    .S(_02095_),
    .Z(_01517_)
  );
  MUX2_X1 _18472_ (
    .A(\rf[7] [23]),
    .B(_05657_),
    .S(_02095_),
    .Z(_01518_)
  );
  MUX2_X1 _18473_ (
    .A(\rf[7] [24]),
    .B(_05665_),
    .S(_02095_),
    .Z(_01519_)
  );
  MUX2_X1 _18474_ (
    .A(\rf[7] [25]),
    .B(_05740_),
    .S(_02095_),
    .Z(_01520_)
  );
  MUX2_X1 _18475_ (
    .A(\rf[7] [26]),
    .B(_05882_),
    .S(_02095_),
    .Z(_01521_)
  );
  MUX2_X1 _18476_ (
    .A(\rf[7] [27]),
    .B(_02159_),
    .S(_02095_),
    .Z(_01522_)
  );
  MUX2_X1 _18477_ (
    .A(\rf[7] [28]),
    .B(_02160_),
    .S(_02095_),
    .Z(_01523_)
  );
  MUX2_X1 _18478_ (
    .A(\rf[7] [29]),
    .B(_02161_),
    .S(_02095_),
    .Z(_01524_)
  );
  MUX2_X1 _18479_ (
    .A(\rf[7] [30]),
    .B(_06117_),
    .S(_02095_),
    .Z(_01525_)
  );
  MUX2_X1 _18480_ (
    .A(\rf[3] [0]),
    .B(_06266_),
    .S(_02101_),
    .Z(_01526_)
  );
  MUX2_X1 _18481_ (
    .A(\rf[3] [1]),
    .B(_06420_),
    .S(_02101_),
    .Z(_01527_)
  );
  MUX2_X1 _18482_ (
    .A(\rf[3] [2]),
    .B(_04080_),
    .S(_02101_),
    .Z(_01528_)
  );
  MUX2_X1 _18483_ (
    .A(\rf[3] [3]),
    .B(_04150_),
    .S(_02101_),
    .Z(_01529_)
  );
  MUX2_X1 _18484_ (
    .A(\rf[3] [4]),
    .B(_04233_),
    .S(_02101_),
    .Z(_01530_)
  );
  MUX2_X1 _18485_ (
    .A(\rf[3] [5]),
    .B(_04305_),
    .S(_02101_),
    .Z(_01531_)
  );
  MUX2_X1 _18486_ (
    .A(\rf[3] [6]),
    .B(_04379_),
    .S(_02101_),
    .Z(_01532_)
  );
  MUX2_X1 _18487_ (
    .A(\rf[3] [7]),
    .B(_02139_),
    .S(_02101_),
    .Z(_01533_)
  );
  MUX2_X1 _18488_ (
    .A(\rf[3] [8]),
    .B(_04521_),
    .S(_02101_),
    .Z(_01534_)
  );
  MUX2_X1 _18489_ (
    .A(\rf[3] [9]),
    .B(_04590_),
    .S(_02101_),
    .Z(_01535_)
  );
  MUX2_X1 _18490_ (
    .A(\rf[3] [10]),
    .B(_04659_),
    .S(_02101_),
    .Z(_01536_)
  );
  MUX2_X1 _18491_ (
    .A(\rf[3] [11]),
    .B(_04742_),
    .S(_02101_),
    .Z(_01537_)
  );
  MUX2_X1 _18492_ (
    .A(\rf[3] [12]),
    .B(_04811_),
    .S(_02101_),
    .Z(_01538_)
  );
  MUX2_X1 _18493_ (
    .A(\rf[3] [13]),
    .B(_04882_),
    .S(_02101_),
    .Z(_01539_)
  );
  MUX2_X1 _18494_ (
    .A(\rf[3] [14]),
    .B(_04953_),
    .S(_02101_),
    .Z(_01540_)
  );
  MUX2_X1 _18495_ (
    .A(\rf[3] [15]),
    .B(_05027_),
    .S(_02101_),
    .Z(_01541_)
  );
  MUX2_X1 _18496_ (
    .A(\rf[3] [16]),
    .B(_02148_),
    .S(_02101_),
    .Z(_01542_)
  );
  MUX2_X1 _18497_ (
    .A(\rf[3] [17]),
    .B(_05170_),
    .S(_02101_),
    .Z(_01543_)
  );
  MUX2_X1 _18498_ (
    .A(\rf[3] [18]),
    .B(_02150_),
    .S(_02101_),
    .Z(_01544_)
  );
  MUX2_X1 _18499_ (
    .A(\rf[3] [19]),
    .B(_02151_),
    .S(_02101_),
    .Z(_01545_)
  );
  MUX2_X1 _18500_ (
    .A(\rf[3] [20]),
    .B(_05442_),
    .S(_02101_),
    .Z(_01546_)
  );
  MUX2_X1 _18501_ (
    .A(\rf[3] [21]),
    .B(_05450_),
    .S(_02101_),
    .Z(_01547_)
  );
  MUX2_X1 _18502_ (
    .A(\rf[3] [22]),
    .B(_05592_),
    .S(_02101_),
    .Z(_01548_)
  );
  MUX2_X1 _18503_ (
    .A(\rf[3] [23]),
    .B(_05657_),
    .S(_02101_),
    .Z(_01549_)
  );
  MUX2_X1 _18504_ (
    .A(\rf[3] [24]),
    .B(_05665_),
    .S(_02101_),
    .Z(_01550_)
  );
  MUX2_X1 _18505_ (
    .A(\rf[3] [25]),
    .B(_05740_),
    .S(_02101_),
    .Z(_01551_)
  );
  MUX2_X1 _18506_ (
    .A(\rf[3] [26]),
    .B(_05882_),
    .S(_02101_),
    .Z(_01552_)
  );
  MUX2_X1 _18507_ (
    .A(\rf[3] [27]),
    .B(_05957_),
    .S(_02101_),
    .Z(_01553_)
  );
  MUX2_X1 _18508_ (
    .A(\rf[3] [28]),
    .B(_02160_),
    .S(_02101_),
    .Z(_01554_)
  );
  MUX2_X1 _18509_ (
    .A(\rf[3] [29]),
    .B(_02161_),
    .S(_02101_),
    .Z(_01555_)
  );
  MUX2_X1 _18510_ (
    .A(\rf[3] [30]),
    .B(_06117_),
    .S(_02101_),
    .Z(_01556_)
  );
  MUX2_X1 _18511_ (
    .A(\rf[1] [0]),
    .B(_02132_),
    .S(_02118_),
    .Z(_01557_)
  );
  MUX2_X1 _18512_ (
    .A(\rf[1] [1]),
    .B(_02133_),
    .S(_02118_),
    .Z(_01558_)
  );
  MUX2_X1 _18513_ (
    .A(\rf[1] [2]),
    .B(_02134_),
    .S(_02118_),
    .Z(_01559_)
  );
  MUX2_X1 _18514_ (
    .A(\rf[1] [3]),
    .B(_02135_),
    .S(_02118_),
    .Z(_01560_)
  );
  MUX2_X1 _18515_ (
    .A(\rf[1] [4]),
    .B(_02136_),
    .S(_02118_),
    .Z(_01561_)
  );
  MUX2_X1 _18516_ (
    .A(\rf[1] [5]),
    .B(_02137_),
    .S(_02118_),
    .Z(_01562_)
  );
  MUX2_X1 _18517_ (
    .A(\rf[1] [6]),
    .B(_02138_),
    .S(_02118_),
    .Z(_01563_)
  );
  MUX2_X1 _18518_ (
    .A(\rf[1] [7]),
    .B(_02139_),
    .S(_02118_),
    .Z(_01564_)
  );
  MUX2_X1 _18519_ (
    .A(\rf[1] [8]),
    .B(_02140_),
    .S(_02118_),
    .Z(_01565_)
  );
  MUX2_X1 _18520_ (
    .A(\rf[1] [9]),
    .B(_02141_),
    .S(_02118_),
    .Z(_01566_)
  );
  MUX2_X1 _18521_ (
    .A(\rf[1] [10]),
    .B(_02142_),
    .S(_02118_),
    .Z(_01567_)
  );
  MUX2_X1 _18522_ (
    .A(\rf[1] [11]),
    .B(_02143_),
    .S(_02118_),
    .Z(_01568_)
  );
  MUX2_X1 _18523_ (
    .A(\rf[1] [12]),
    .B(_02144_),
    .S(_02118_),
    .Z(_01569_)
  );
  MUX2_X1 _18524_ (
    .A(\rf[1] [13]),
    .B(_02145_),
    .S(_02118_),
    .Z(_01570_)
  );
  MUX2_X1 _18525_ (
    .A(\rf[1] [14]),
    .B(_02146_),
    .S(_02118_),
    .Z(_01571_)
  );
  MUX2_X1 _18526_ (
    .A(\rf[1] [15]),
    .B(_02147_),
    .S(_02118_),
    .Z(_01572_)
  );
  MUX2_X1 _18527_ (
    .A(\rf[1] [16]),
    .B(_02148_),
    .S(_02118_),
    .Z(_01573_)
  );
  MUX2_X1 _18528_ (
    .A(\rf[1] [17]),
    .B(_02149_),
    .S(_02118_),
    .Z(_01574_)
  );
  MUX2_X1 _18529_ (
    .A(\rf[1] [18]),
    .B(_02150_),
    .S(_02118_),
    .Z(_01575_)
  );
  MUX2_X1 _18530_ (
    .A(\rf[1] [19]),
    .B(_02151_),
    .S(_02118_),
    .Z(_01576_)
  );
  MUX2_X1 _18531_ (
    .A(\rf[1] [20]),
    .B(_02152_),
    .S(_02118_),
    .Z(_01577_)
  );
  MUX2_X1 _18532_ (
    .A(\rf[1] [21]),
    .B(_02153_),
    .S(_02118_),
    .Z(_01578_)
  );
  MUX2_X1 _18533_ (
    .A(\rf[1] [22]),
    .B(_02154_),
    .S(_02118_),
    .Z(_01579_)
  );
  MUX2_X1 _18534_ (
    .A(\rf[1] [23]),
    .B(_02155_),
    .S(_02118_),
    .Z(_01580_)
  );
  MUX2_X1 _18535_ (
    .A(\rf[1] [24]),
    .B(_02156_),
    .S(_02118_),
    .Z(_01581_)
  );
  MUX2_X1 _18536_ (
    .A(\rf[1] [25]),
    .B(_02157_),
    .S(_02118_),
    .Z(_01582_)
  );
  MUX2_X1 _18537_ (
    .A(\rf[1] [26]),
    .B(_02158_),
    .S(_02118_),
    .Z(_01583_)
  );
  MUX2_X1 _18538_ (
    .A(\rf[1] [27]),
    .B(_02159_),
    .S(_02118_),
    .Z(_01584_)
  );
  MUX2_X1 _18539_ (
    .A(\rf[1] [28]),
    .B(_02160_),
    .S(_02118_),
    .Z(_01585_)
  );
  MUX2_X1 _18540_ (
    .A(\rf[1] [29]),
    .B(_02161_),
    .S(_02118_),
    .Z(_01586_)
  );
  MUX2_X1 _18541_ (
    .A(\rf[1] [30]),
    .B(_02162_),
    .S(_02118_),
    .Z(_01587_)
  );
  OR2_X1 _18542_ (
    .A1(_00032_),
    .A2(_00031_),
    .ZN(_02168_)
  );
  AND2_X1 _18543_ (
    .A1(_02980_),
    .A2(_03061_),
    .ZN(_02169_)
  );
  INV_X1 _18544_ (
    .A(_02169_),
    .ZN(_02170_)
  );
  OR2_X1 _18545_ (
    .A1(ex_reg_rs_lsb_0[1]),
    .A2(_00032_),
    .ZN(_02171_)
  );
  INV_X1 _18546_ (
    .A(_02171_),
    .ZN(_02172_)
  );
  AND2_X1 _18547_ (
    .A1(_02170_),
    .A2(_02172_),
    .ZN(_02173_)
  );
  AND2_X1 _18548_ (
    .A1(mem_reg_wdata[0]),
    .A2(_02173_),
    .ZN(_02174_)
  );
  AND2_X1 _18549_ (
    .A1(wb_reg_wdata[0]),
    .A2(_02169_),
    .ZN(_02175_)
  );
  OR2_X1 _18550_ (
    .A1(_02174_),
    .A2(_02175_),
    .ZN(_02176_)
  );
  MUX2_X1 _18551_ (
    .A(io_dmem_resp_bits_data_word_bypass[0]),
    .B(_02176_),
    .S(_02168_),
    .Z(_02177_)
  );
  MUX2_X1 _18552_ (
    .A(ex_reg_rs_lsb_0[0]),
    .B(_02177_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[0])
  );
  AND2_X1 _18553_ (
    .A1(mem_reg_wdata[1]),
    .A2(_02173_),
    .ZN(_02178_)
  );
  AND2_X1 _18554_ (
    .A1(wb_reg_wdata[1]),
    .A2(_02169_),
    .ZN(_02179_)
  );
  OR2_X1 _18555_ (
    .A1(_02178_),
    .A2(_02179_),
    .ZN(_02180_)
  );
  MUX2_X1 _18556_ (
    .A(io_dmem_resp_bits_data_word_bypass[1]),
    .B(_02180_),
    .S(_02168_),
    .Z(_02181_)
  );
  MUX2_X1 _18557_ (
    .A(ex_reg_rs_lsb_0[1]),
    .B(_02181_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[1])
  );
  AND2_X1 _18558_ (
    .A1(mem_reg_wdata[2]),
    .A2(_02173_),
    .ZN(_02182_)
  );
  AND2_X1 _18559_ (
    .A1(wb_reg_wdata[2]),
    .A2(_02169_),
    .ZN(_02183_)
  );
  OR2_X1 _18560_ (
    .A1(_02182_),
    .A2(_02183_),
    .ZN(_02184_)
  );
  MUX2_X1 _18561_ (
    .A(io_dmem_resp_bits_data_word_bypass[2]),
    .B(_02184_),
    .S(_02168_),
    .Z(_02185_)
  );
  MUX2_X1 _18562_ (
    .A(ex_reg_rs_msb_0[0]),
    .B(_02185_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[2])
  );
  AND2_X1 _18563_ (
    .A1(mem_reg_wdata[3]),
    .A2(_02173_),
    .ZN(_02186_)
  );
  AND2_X1 _18564_ (
    .A1(wb_reg_wdata[3]),
    .A2(_02169_),
    .ZN(_02187_)
  );
  OR2_X1 _18565_ (
    .A1(_02186_),
    .A2(_02187_),
    .ZN(_02188_)
  );
  MUX2_X1 _18566_ (
    .A(io_dmem_resp_bits_data_word_bypass[3]),
    .B(_02188_),
    .S(_02168_),
    .Z(_02189_)
  );
  MUX2_X1 _18567_ (
    .A(ex_reg_rs_msb_0[1]),
    .B(_02189_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[3])
  );
  AND2_X1 _18568_ (
    .A1(mem_reg_wdata[4]),
    .A2(_02173_),
    .ZN(_02190_)
  );
  AND2_X1 _18569_ (
    .A1(wb_reg_wdata[4]),
    .A2(_02169_),
    .ZN(_02191_)
  );
  OR2_X1 _18570_ (
    .A1(_02190_),
    .A2(_02191_),
    .ZN(_02192_)
  );
  MUX2_X1 _18571_ (
    .A(io_dmem_resp_bits_data_word_bypass[4]),
    .B(_02192_),
    .S(_02168_),
    .Z(_02193_)
  );
  MUX2_X1 _18572_ (
    .A(ex_reg_rs_msb_0[2]),
    .B(_02193_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[4])
  );
  AND2_X1 _18573_ (
    .A1(mem_reg_wdata[5]),
    .A2(_02173_),
    .ZN(_02194_)
  );
  AND2_X1 _18574_ (
    .A1(wb_reg_wdata[5]),
    .A2(_02169_),
    .ZN(_02195_)
  );
  OR2_X1 _18575_ (
    .A1(_02194_),
    .A2(_02195_),
    .ZN(_02196_)
  );
  MUX2_X1 _18576_ (
    .A(io_dmem_resp_bits_data_word_bypass[5]),
    .B(_02196_),
    .S(_02168_),
    .Z(_02197_)
  );
  MUX2_X1 _18577_ (
    .A(ex_reg_rs_msb_0[3]),
    .B(_02197_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[5])
  );
  AND2_X1 _18578_ (
    .A1(mem_reg_wdata[6]),
    .A2(_02173_),
    .ZN(_02198_)
  );
  AND2_X1 _18579_ (
    .A1(wb_reg_wdata[6]),
    .A2(_02169_),
    .ZN(_02199_)
  );
  OR2_X1 _18580_ (
    .A1(_02198_),
    .A2(_02199_),
    .ZN(_02200_)
  );
  MUX2_X1 _18581_ (
    .A(io_dmem_resp_bits_data_word_bypass[6]),
    .B(_02200_),
    .S(_02168_),
    .Z(_02201_)
  );
  MUX2_X1 _18582_ (
    .A(ex_reg_rs_msb_0[4]),
    .B(_02201_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[6])
  );
  AND2_X1 _18583_ (
    .A1(mem_reg_wdata[7]),
    .A2(_02173_),
    .ZN(_02202_)
  );
  AND2_X1 _18584_ (
    .A1(wb_reg_wdata[7]),
    .A2(_02169_),
    .ZN(_02203_)
  );
  OR2_X1 _18585_ (
    .A1(_02202_),
    .A2(_02203_),
    .ZN(_02204_)
  );
  MUX2_X1 _18586_ (
    .A(io_dmem_resp_bits_data_word_bypass[7]),
    .B(_02204_),
    .S(_02168_),
    .Z(_02205_)
  );
  MUX2_X1 _18587_ (
    .A(ex_reg_rs_msb_0[5]),
    .B(_02205_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[7])
  );
  AND2_X1 _18588_ (
    .A1(mem_reg_wdata[8]),
    .A2(_02173_),
    .ZN(_02206_)
  );
  AND2_X1 _18589_ (
    .A1(wb_reg_wdata[8]),
    .A2(_02169_),
    .ZN(_02207_)
  );
  OR2_X1 _18590_ (
    .A1(_02206_),
    .A2(_02207_),
    .ZN(_02208_)
  );
  MUX2_X1 _18591_ (
    .A(io_dmem_resp_bits_data_word_bypass[8]),
    .B(_02208_),
    .S(_02168_),
    .Z(_02209_)
  );
  MUX2_X1 _18592_ (
    .A(ex_reg_rs_msb_0[6]),
    .B(_02209_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[8])
  );
  AND2_X1 _18593_ (
    .A1(mem_reg_wdata[9]),
    .A2(_02173_),
    .ZN(_02210_)
  );
  AND2_X1 _18594_ (
    .A1(wb_reg_wdata[9]),
    .A2(_02169_),
    .ZN(_02211_)
  );
  OR2_X1 _18595_ (
    .A1(_02210_),
    .A2(_02211_),
    .ZN(_02212_)
  );
  MUX2_X1 _18596_ (
    .A(io_dmem_resp_bits_data_word_bypass[9]),
    .B(_02212_),
    .S(_02168_),
    .Z(_02213_)
  );
  MUX2_X1 _18597_ (
    .A(ex_reg_rs_msb_0[7]),
    .B(_02213_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[9])
  );
  AND2_X1 _18598_ (
    .A1(mem_reg_wdata[10]),
    .A2(_02173_),
    .ZN(_02214_)
  );
  AND2_X1 _18599_ (
    .A1(wb_reg_wdata[10]),
    .A2(_02169_),
    .ZN(_02215_)
  );
  OR2_X1 _18600_ (
    .A1(_02214_),
    .A2(_02215_),
    .ZN(_02216_)
  );
  MUX2_X1 _18601_ (
    .A(io_dmem_resp_bits_data_word_bypass[10]),
    .B(_02216_),
    .S(_02168_),
    .Z(_02217_)
  );
  MUX2_X1 _18602_ (
    .A(ex_reg_rs_msb_0[8]),
    .B(_02217_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[10])
  );
  AND2_X1 _18603_ (
    .A1(mem_reg_wdata[11]),
    .A2(_02173_),
    .ZN(_02218_)
  );
  AND2_X1 _18604_ (
    .A1(wb_reg_wdata[11]),
    .A2(_02169_),
    .ZN(_02219_)
  );
  OR2_X1 _18605_ (
    .A1(_02218_),
    .A2(_02219_),
    .ZN(_02220_)
  );
  MUX2_X1 _18606_ (
    .A(io_dmem_resp_bits_data_word_bypass[11]),
    .B(_02220_),
    .S(_02168_),
    .Z(_02221_)
  );
  MUX2_X1 _18607_ (
    .A(ex_reg_rs_msb_0[9]),
    .B(_02221_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[11])
  );
  AND2_X1 _18608_ (
    .A1(mem_reg_wdata[12]),
    .A2(_02173_),
    .ZN(_02222_)
  );
  AND2_X1 _18609_ (
    .A1(wb_reg_wdata[12]),
    .A2(_02169_),
    .ZN(_02223_)
  );
  OR2_X1 _18610_ (
    .A1(_02222_),
    .A2(_02223_),
    .ZN(_02224_)
  );
  MUX2_X1 _18611_ (
    .A(io_dmem_resp_bits_data_word_bypass[12]),
    .B(_02224_),
    .S(_02168_),
    .Z(_02225_)
  );
  MUX2_X1 _18612_ (
    .A(ex_reg_rs_msb_0[10]),
    .B(_02225_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[12])
  );
  AND2_X1 _18613_ (
    .A1(mem_reg_wdata[13]),
    .A2(_02173_),
    .ZN(_02226_)
  );
  AND2_X1 _18614_ (
    .A1(wb_reg_wdata[13]),
    .A2(_02169_),
    .ZN(_02227_)
  );
  OR2_X1 _18615_ (
    .A1(_02226_),
    .A2(_02227_),
    .ZN(_02228_)
  );
  MUX2_X1 _18616_ (
    .A(io_dmem_resp_bits_data_word_bypass[13]),
    .B(_02228_),
    .S(_02168_),
    .Z(_02229_)
  );
  MUX2_X1 _18617_ (
    .A(ex_reg_rs_msb_0[11]),
    .B(_02229_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[13])
  );
  AND2_X1 _18618_ (
    .A1(mem_reg_wdata[14]),
    .A2(_02173_),
    .ZN(_02230_)
  );
  AND2_X1 _18619_ (
    .A1(wb_reg_wdata[14]),
    .A2(_02169_),
    .ZN(_02231_)
  );
  OR2_X1 _18620_ (
    .A1(_02230_),
    .A2(_02231_),
    .ZN(_02232_)
  );
  MUX2_X1 _18621_ (
    .A(io_dmem_resp_bits_data_word_bypass[14]),
    .B(_02232_),
    .S(_02168_),
    .Z(_02233_)
  );
  MUX2_X1 _18622_ (
    .A(ex_reg_rs_msb_0[12]),
    .B(_02233_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[14])
  );
  AND2_X1 _18623_ (
    .A1(mem_reg_wdata[15]),
    .A2(_02173_),
    .ZN(_02234_)
  );
  AND2_X1 _18624_ (
    .A1(wb_reg_wdata[15]),
    .A2(_02169_),
    .ZN(_02235_)
  );
  OR2_X1 _18625_ (
    .A1(_02234_),
    .A2(_02235_),
    .ZN(_02236_)
  );
  MUX2_X1 _18626_ (
    .A(io_dmem_resp_bits_data_word_bypass[15]),
    .B(_02236_),
    .S(_02168_),
    .Z(_02237_)
  );
  MUX2_X1 _18627_ (
    .A(ex_reg_rs_msb_0[13]),
    .B(_02237_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[15])
  );
  AND2_X1 _18628_ (
    .A1(mem_reg_wdata[16]),
    .A2(_02173_),
    .ZN(_02238_)
  );
  AND2_X1 _18629_ (
    .A1(wb_reg_wdata[16]),
    .A2(_02169_),
    .ZN(_02239_)
  );
  OR2_X1 _18630_ (
    .A1(_02238_),
    .A2(_02239_),
    .ZN(_02240_)
  );
  MUX2_X1 _18631_ (
    .A(io_dmem_resp_bits_data_word_bypass[16]),
    .B(_02240_),
    .S(_02168_),
    .Z(_02241_)
  );
  MUX2_X1 _18632_ (
    .A(ex_reg_rs_msb_0[14]),
    .B(_02241_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[16])
  );
  AND2_X1 _18633_ (
    .A1(mem_reg_wdata[17]),
    .A2(_02173_),
    .ZN(_02242_)
  );
  AND2_X1 _18634_ (
    .A1(wb_reg_wdata[17]),
    .A2(_02169_),
    .ZN(_02243_)
  );
  OR2_X1 _18635_ (
    .A1(_02242_),
    .A2(_02243_),
    .ZN(_02244_)
  );
  MUX2_X1 _18636_ (
    .A(io_dmem_resp_bits_data_word_bypass[17]),
    .B(_02244_),
    .S(_02168_),
    .Z(_02245_)
  );
  MUX2_X1 _18637_ (
    .A(ex_reg_rs_msb_0[15]),
    .B(_02245_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[17])
  );
  AND2_X1 _18638_ (
    .A1(mem_reg_wdata[18]),
    .A2(_02173_),
    .ZN(_02246_)
  );
  AND2_X1 _18639_ (
    .A1(wb_reg_wdata[18]),
    .A2(_02169_),
    .ZN(_02247_)
  );
  OR2_X1 _18640_ (
    .A1(_02246_),
    .A2(_02247_),
    .ZN(_02248_)
  );
  MUX2_X1 _18641_ (
    .A(io_dmem_resp_bits_data_word_bypass[18]),
    .B(_02248_),
    .S(_02168_),
    .Z(_02249_)
  );
  MUX2_X1 _18642_ (
    .A(ex_reg_rs_msb_0[16]),
    .B(_02249_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[18])
  );
  AND2_X1 _18643_ (
    .A1(mem_reg_wdata[19]),
    .A2(_02173_),
    .ZN(_02250_)
  );
  AND2_X1 _18644_ (
    .A1(wb_reg_wdata[19]),
    .A2(_02169_),
    .ZN(_02251_)
  );
  OR2_X1 _18645_ (
    .A1(_02250_),
    .A2(_02251_),
    .ZN(_02252_)
  );
  MUX2_X1 _18646_ (
    .A(io_dmem_resp_bits_data_word_bypass[19]),
    .B(_02252_),
    .S(_02168_),
    .Z(_02253_)
  );
  MUX2_X1 _18647_ (
    .A(ex_reg_rs_msb_0[17]),
    .B(_02253_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[19])
  );
  AND2_X1 _18648_ (
    .A1(mem_reg_wdata[20]),
    .A2(_02173_),
    .ZN(_02254_)
  );
  AND2_X1 _18649_ (
    .A1(wb_reg_wdata[20]),
    .A2(_02169_),
    .ZN(_02255_)
  );
  OR2_X1 _18650_ (
    .A1(_02254_),
    .A2(_02255_),
    .ZN(_02256_)
  );
  MUX2_X1 _18651_ (
    .A(io_dmem_resp_bits_data_word_bypass[20]),
    .B(_02256_),
    .S(_02168_),
    .Z(_02257_)
  );
  MUX2_X1 _18652_ (
    .A(ex_reg_rs_msb_0[18]),
    .B(_02257_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[20])
  );
  AND2_X1 _18653_ (
    .A1(mem_reg_wdata[21]),
    .A2(_02173_),
    .ZN(_02258_)
  );
  AND2_X1 _18654_ (
    .A1(wb_reg_wdata[21]),
    .A2(_02169_),
    .ZN(_02259_)
  );
  OR2_X1 _18655_ (
    .A1(_02258_),
    .A2(_02259_),
    .ZN(_02260_)
  );
  MUX2_X1 _18656_ (
    .A(io_dmem_resp_bits_data_word_bypass[21]),
    .B(_02260_),
    .S(_02168_),
    .Z(_02261_)
  );
  MUX2_X1 _18657_ (
    .A(ex_reg_rs_msb_0[19]),
    .B(_02261_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[21])
  );
  AND2_X1 _18658_ (
    .A1(mem_reg_wdata[22]),
    .A2(_02173_),
    .ZN(_02262_)
  );
  AND2_X1 _18659_ (
    .A1(wb_reg_wdata[22]),
    .A2(_02169_),
    .ZN(_02263_)
  );
  OR2_X1 _18660_ (
    .A1(_02262_),
    .A2(_02263_),
    .ZN(_02264_)
  );
  MUX2_X1 _18661_ (
    .A(io_dmem_resp_bits_data_word_bypass[22]),
    .B(_02264_),
    .S(_02168_),
    .Z(_02265_)
  );
  MUX2_X1 _18662_ (
    .A(ex_reg_rs_msb_0[20]),
    .B(_02265_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[22])
  );
  AND2_X1 _18663_ (
    .A1(mem_reg_wdata[23]),
    .A2(_02173_),
    .ZN(_02266_)
  );
  AND2_X1 _18664_ (
    .A1(wb_reg_wdata[23]),
    .A2(_02169_),
    .ZN(_02267_)
  );
  OR2_X1 _18665_ (
    .A1(_02266_),
    .A2(_02267_),
    .ZN(_02268_)
  );
  MUX2_X1 _18666_ (
    .A(io_dmem_resp_bits_data_word_bypass[23]),
    .B(_02268_),
    .S(_02168_),
    .Z(_02269_)
  );
  MUX2_X1 _18667_ (
    .A(ex_reg_rs_msb_0[21]),
    .B(_02269_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[23])
  );
  AND2_X1 _18668_ (
    .A1(mem_reg_wdata[24]),
    .A2(_02173_),
    .ZN(_02270_)
  );
  AND2_X1 _18669_ (
    .A1(wb_reg_wdata[24]),
    .A2(_02169_),
    .ZN(_02271_)
  );
  OR2_X1 _18670_ (
    .A1(_02270_),
    .A2(_02271_),
    .ZN(_02272_)
  );
  MUX2_X1 _18671_ (
    .A(io_dmem_resp_bits_data_word_bypass[24]),
    .B(_02272_),
    .S(_02168_),
    .Z(_02273_)
  );
  MUX2_X1 _18672_ (
    .A(ex_reg_rs_msb_0[22]),
    .B(_02273_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[24])
  );
  AND2_X1 _18673_ (
    .A1(mem_reg_wdata[25]),
    .A2(_02173_),
    .ZN(_02274_)
  );
  AND2_X1 _18674_ (
    .A1(wb_reg_wdata[25]),
    .A2(_02169_),
    .ZN(_02275_)
  );
  OR2_X1 _18675_ (
    .A1(_02274_),
    .A2(_02275_),
    .ZN(_02276_)
  );
  MUX2_X1 _18676_ (
    .A(io_dmem_resp_bits_data_word_bypass[25]),
    .B(_02276_),
    .S(_02168_),
    .Z(_02277_)
  );
  MUX2_X1 _18677_ (
    .A(ex_reg_rs_msb_0[23]),
    .B(_02277_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[25])
  );
  AND2_X1 _18678_ (
    .A1(mem_reg_wdata[26]),
    .A2(_02173_),
    .ZN(_02278_)
  );
  AND2_X1 _18679_ (
    .A1(wb_reg_wdata[26]),
    .A2(_02169_),
    .ZN(_02279_)
  );
  OR2_X1 _18680_ (
    .A1(_02278_),
    .A2(_02279_),
    .ZN(_02280_)
  );
  MUX2_X1 _18681_ (
    .A(io_dmem_resp_bits_data_word_bypass[26]),
    .B(_02280_),
    .S(_02168_),
    .Z(_02281_)
  );
  MUX2_X1 _18682_ (
    .A(ex_reg_rs_msb_0[24]),
    .B(_02281_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[26])
  );
  AND2_X1 _18683_ (
    .A1(mem_reg_wdata[27]),
    .A2(_02173_),
    .ZN(_02282_)
  );
  AND2_X1 _18684_ (
    .A1(wb_reg_wdata[27]),
    .A2(_02169_),
    .ZN(_02283_)
  );
  OR2_X1 _18685_ (
    .A1(_02282_),
    .A2(_02283_),
    .ZN(_02284_)
  );
  MUX2_X1 _18686_ (
    .A(io_dmem_resp_bits_data_word_bypass[27]),
    .B(_02284_),
    .S(_02168_),
    .Z(_02285_)
  );
  MUX2_X1 _18687_ (
    .A(ex_reg_rs_msb_0[25]),
    .B(_02285_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[27])
  );
  AND2_X1 _18688_ (
    .A1(mem_reg_wdata[28]),
    .A2(_02173_),
    .ZN(_02286_)
  );
  AND2_X1 _18689_ (
    .A1(wb_reg_wdata[28]),
    .A2(_02169_),
    .ZN(_02287_)
  );
  OR2_X1 _18690_ (
    .A1(_02286_),
    .A2(_02287_),
    .ZN(_02288_)
  );
  MUX2_X1 _18691_ (
    .A(io_dmem_resp_bits_data_word_bypass[28]),
    .B(_02288_),
    .S(_02168_),
    .Z(_02289_)
  );
  MUX2_X1 _18692_ (
    .A(ex_reg_rs_msb_0[26]),
    .B(_02289_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[28])
  );
  AND2_X1 _18693_ (
    .A1(mem_reg_wdata[29]),
    .A2(_02173_),
    .ZN(_02290_)
  );
  AND2_X1 _18694_ (
    .A1(wb_reg_wdata[29]),
    .A2(_02169_),
    .ZN(_02291_)
  );
  OR2_X1 _18695_ (
    .A1(_02290_),
    .A2(_02291_),
    .ZN(_02292_)
  );
  MUX2_X1 _18696_ (
    .A(io_dmem_resp_bits_data_word_bypass[29]),
    .B(_02292_),
    .S(_02168_),
    .Z(_02293_)
  );
  MUX2_X1 _18697_ (
    .A(ex_reg_rs_msb_0[27]),
    .B(_02293_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[29])
  );
  AND2_X1 _18698_ (
    .A1(mem_reg_wdata[30]),
    .A2(_02173_),
    .ZN(_02294_)
  );
  AND2_X1 _18699_ (
    .A1(wb_reg_wdata[30]),
    .A2(_02169_),
    .ZN(_02295_)
  );
  OR2_X1 _18700_ (
    .A1(_02294_),
    .A2(_02295_),
    .ZN(_02296_)
  );
  MUX2_X1 _18701_ (
    .A(io_dmem_resp_bits_data_word_bypass[30]),
    .B(_02296_),
    .S(_02168_),
    .Z(_02297_)
  );
  MUX2_X1 _18702_ (
    .A(ex_reg_rs_msb_0[28]),
    .B(_02297_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[30])
  );
  AND2_X1 _18703_ (
    .A1(mem_reg_wdata[31]),
    .A2(_02173_),
    .ZN(_02298_)
  );
  AND2_X1 _18704_ (
    .A1(wb_reg_wdata[31]),
    .A2(_02169_),
    .ZN(_02299_)
  );
  OR2_X1 _18705_ (
    .A1(_02298_),
    .A2(_02299_),
    .ZN(_02300_)
  );
  MUX2_X1 _18706_ (
    .A(io_dmem_resp_bits_data_word_bypass[31]),
    .B(_02300_),
    .S(_02168_),
    .Z(_02301_)
  );
  MUX2_X1 _18707_ (
    .A(ex_reg_rs_msb_0[29]),
    .B(_02301_),
    .S(ex_reg_rs_bypass_0),
    .Z(_ex_op1_T[31])
  );
  AND2_X1 _18708_ (
    .A1(wb_reg_raw_inst[0]),
    .A2(wb_reg_raw_inst[1]),
    .ZN(_02302_)
  );
  AND2_X1 _18709_ (
    .A1(wb_reg_inst[16]),
    .A2(_02302_),
    .ZN(_csr_io_inst_0_T_3[0])
  );
  AND2_X1 _18710_ (
    .A1(wb_reg_inst[17]),
    .A2(_02302_),
    .ZN(_csr_io_inst_0_T_3[1])
  );
  AND2_X1 _18711_ (
    .A1(wb_reg_inst[18]),
    .A2(_02302_),
    .ZN(_csr_io_inst_0_T_3[2])
  );
  AND2_X1 _18712_ (
    .A1(wb_reg_inst[19]),
    .A2(_02302_),
    .ZN(_csr_io_inst_0_T_3[3])
  );
  AND2_X1 _18713_ (
    .A1(wb_reg_inst[20]),
    .A2(_02302_),
    .ZN(_csr_io_inst_0_T_3[4])
  );
  AND2_X1 _18714_ (
    .A1(wb_reg_inst[21]),
    .A2(_02302_),
    .ZN(_csr_io_inst_0_T_3[5])
  );
  AND2_X1 _18715_ (
    .A1(wb_reg_inst[22]),
    .A2(_02302_),
    .ZN(_csr_io_inst_0_T_3[6])
  );
  AND2_X1 _18716_ (
    .A1(wb_reg_inst[23]),
    .A2(_02302_),
    .ZN(_csr_io_inst_0_T_3[7])
  );
  AND2_X1 _18717_ (
    .A1(wb_reg_inst[24]),
    .A2(_02302_),
    .ZN(_csr_io_inst_0_T_3[8])
  );
  AND2_X1 _18718_ (
    .A1(wb_reg_inst[25]),
    .A2(_02302_),
    .ZN(_csr_io_inst_0_T_3[9])
  );
  AND2_X1 _18719_ (
    .A1(wb_reg_inst[26]),
    .A2(_02302_),
    .ZN(_csr_io_inst_0_T_3[10])
  );
  AND2_X1 _18720_ (
    .A1(wb_reg_inst[27]),
    .A2(_02302_),
    .ZN(_csr_io_inst_0_T_3[11])
  );
  AND2_X1 _18721_ (
    .A1(wb_reg_inst[28]),
    .A2(_02302_),
    .ZN(_csr_io_inst_0_T_3[12])
  );
  AND2_X1 _18722_ (
    .A1(wb_reg_inst[29]),
    .A2(_02302_),
    .ZN(_csr_io_inst_0_T_3[13])
  );
  AND2_X1 _18723_ (
    .A1(wb_reg_inst[30]),
    .A2(_02302_),
    .ZN(_csr_io_inst_0_T_3[14])
  );
  AND2_X1 _18724_ (
    .A1(wb_reg_inst[31]),
    .A2(_02302_),
    .ZN(_csr_io_inst_0_T_3[15])
  );
  AND2_X1 _18725_ (
    .A1(wb_reg_pc[0]),
    .A2(_03142_),
    .ZN(_02303_)
  );
  MUX2_X1 _18726_ (
    .A(_02303_),
    .B(csr_io_evec[0]),
    .S(_04026_),
    .Z(io_imem_req_bits_pc[0])
  );
  AND2_X1 _18727_ (
    .A1(_03141_),
    .A2(_06438_),
    .ZN(_02304_)
  );
  AND2_X1 _18728_ (
    .A1(wb_reg_pc[1]),
    .A2(_03142_),
    .ZN(_02305_)
  );
  OR2_X1 _18729_ (
    .A1(_04026_),
    .A2(_02305_),
    .ZN(_02306_)
  );
  OR2_X1 _18730_ (
    .A1(_02304_),
    .A2(_02306_),
    .ZN(_02307_)
  );
  OR2_X1 _18731_ (
    .A1(csr_io_evec[1]),
    .A2(_04025_),
    .ZN(_02308_)
  );
  AND2_X1 _18732_ (
    .A1(_02307_),
    .A2(_02308_),
    .ZN(io_imem_req_bits_pc[1])
  );
  MUX2_X1 _18733_ (
    .A(mem_reg_wdata[2]),
    .B(_06451_),
    .S(_03030_),
    .Z(_02309_)
  );
  MUX2_X1 _18734_ (
    .A(wb_reg_pc[2]),
    .B(_02309_),
    .S(_03141_),
    .Z(_02310_)
  );
  MUX2_X1 _18735_ (
    .A(_02310_),
    .B(csr_io_evec[2]),
    .S(_04026_),
    .Z(io_imem_req_bits_pc[2])
  );
  MUX2_X1 _18736_ (
    .A(mem_reg_wdata[3]),
    .B(_06459_),
    .S(_03030_),
    .Z(_02311_)
  );
  INV_X1 _18737_ (
    .A(_02311_),
    .ZN(_02312_)
  );
  MUX2_X1 _18738_ (
    .A(wb_reg_pc[3]),
    .B(_02311_),
    .S(_03141_),
    .Z(_02313_)
  );
  MUX2_X1 _18739_ (
    .A(csr_io_evec[3]),
    .B(_02313_),
    .S(_04025_),
    .Z(io_imem_req_bits_pc[3])
  );
  MUX2_X1 _18740_ (
    .A(mem_reg_wdata[4]),
    .B(_06468_),
    .S(_03030_),
    .Z(_02314_)
  );
  INV_X1 _18741_ (
    .A(_02314_),
    .ZN(_02315_)
  );
  MUX2_X1 _18742_ (
    .A(wb_reg_pc[4]),
    .B(_02314_),
    .S(_03141_),
    .Z(_02316_)
  );
  MUX2_X1 _18743_ (
    .A(csr_io_evec[4]),
    .B(_02316_),
    .S(_04025_),
    .Z(io_imem_req_bits_pc[4])
  );
  AND2_X1 _18744_ (
    .A1(csr_io_evec[5]),
    .A2(_04026_),
    .ZN(_02317_)
  );
  MUX2_X1 _18745_ (
    .A(mem_reg_wdata[5]),
    .B(_06476_),
    .S(_03030_),
    .Z(_02318_)
  );
  INV_X1 _18746_ (
    .A(_02318_),
    .ZN(_02319_)
  );
  OR2_X1 _18747_ (
    .A1(_03142_),
    .A2(_02318_),
    .ZN(_02320_)
  );
  OR2_X1 _18748_ (
    .A1(wb_reg_pc[5]),
    .A2(_03141_),
    .ZN(_02321_)
  );
  AND2_X1 _18749_ (
    .A1(_04025_),
    .A2(_02321_),
    .ZN(_02322_)
  );
  AND2_X1 _18750_ (
    .A1(_02320_),
    .A2(_02322_),
    .ZN(_02323_)
  );
  OR2_X1 _18751_ (
    .A1(_02317_),
    .A2(_02323_),
    .ZN(io_imem_req_bits_pc[5])
  );
  AND2_X1 _18752_ (
    .A1(csr_io_evec[6]),
    .A2(_04026_),
    .ZN(_02324_)
  );
  MUX2_X1 _18753_ (
    .A(mem_reg_wdata[6]),
    .B(_06487_),
    .S(_03030_),
    .Z(_02325_)
  );
  INV_X1 _18754_ (
    .A(_02325_),
    .ZN(_02326_)
  );
  OR2_X1 _18755_ (
    .A1(_03142_),
    .A2(_02325_),
    .ZN(_02327_)
  );
  OR2_X1 _18756_ (
    .A1(wb_reg_pc[6]),
    .A2(_03141_),
    .ZN(_02328_)
  );
  AND2_X1 _18757_ (
    .A1(_04025_),
    .A2(_02328_),
    .ZN(_02329_)
  );
  AND2_X1 _18758_ (
    .A1(_02327_),
    .A2(_02329_),
    .ZN(_02330_)
  );
  OR2_X1 _18759_ (
    .A1(_02324_),
    .A2(_02330_),
    .ZN(io_imem_req_bits_pc[6])
  );
  AND2_X1 _18760_ (
    .A1(csr_io_evec[7]),
    .A2(_04026_),
    .ZN(_02331_)
  );
  MUX2_X1 _18761_ (
    .A(mem_reg_wdata[7]),
    .B(_06498_),
    .S(_03030_),
    .Z(_02332_)
  );
  INV_X1 _18762_ (
    .A(_02332_),
    .ZN(_02333_)
  );
  OR2_X1 _18763_ (
    .A1(_03142_),
    .A2(_02332_),
    .ZN(_02334_)
  );
  OR2_X1 _18764_ (
    .A1(wb_reg_pc[7]),
    .A2(_03141_),
    .ZN(_02335_)
  );
  AND2_X1 _18765_ (
    .A1(_04025_),
    .A2(_02335_),
    .ZN(_02336_)
  );
  AND2_X1 _18766_ (
    .A1(_02334_),
    .A2(_02336_),
    .ZN(_02337_)
  );
  OR2_X1 _18767_ (
    .A1(_02331_),
    .A2(_02337_),
    .ZN(io_imem_req_bits_pc[7])
  );
  AND2_X1 _18768_ (
    .A1(csr_io_evec[8]),
    .A2(_04026_),
    .ZN(_02338_)
  );
  MUX2_X1 _18769_ (
    .A(mem_reg_wdata[8]),
    .B(_06509_),
    .S(_03030_),
    .Z(_02339_)
  );
  INV_X1 _18770_ (
    .A(_02339_),
    .ZN(_02340_)
  );
  OR2_X1 _18771_ (
    .A1(_03142_),
    .A2(_02339_),
    .ZN(_02341_)
  );
  OR2_X1 _18772_ (
    .A1(wb_reg_pc[8]),
    .A2(_03141_),
    .ZN(_02342_)
  );
  AND2_X1 _18773_ (
    .A1(_04025_),
    .A2(_02342_),
    .ZN(_02343_)
  );
  AND2_X1 _18774_ (
    .A1(_02341_),
    .A2(_02343_),
    .ZN(_02344_)
  );
  OR2_X1 _18775_ (
    .A1(_02338_),
    .A2(_02344_),
    .ZN(io_imem_req_bits_pc[8])
  );
  AND2_X1 _18776_ (
    .A1(csr_io_evec[9]),
    .A2(_04026_),
    .ZN(_02345_)
  );
  MUX2_X1 _18777_ (
    .A(mem_reg_wdata[9]),
    .B(_06517_),
    .S(_03030_),
    .Z(_02346_)
  );
  INV_X1 _18778_ (
    .A(_02346_),
    .ZN(_02347_)
  );
  OR2_X1 _18779_ (
    .A1(_03142_),
    .A2(_02346_),
    .ZN(_02348_)
  );
  OR2_X1 _18780_ (
    .A1(wb_reg_pc[9]),
    .A2(_03141_),
    .ZN(_02349_)
  );
  AND2_X1 _18781_ (
    .A1(_04025_),
    .A2(_02349_),
    .ZN(_02350_)
  );
  AND2_X1 _18782_ (
    .A1(_02348_),
    .A2(_02350_),
    .ZN(_02351_)
  );
  OR2_X1 _18783_ (
    .A1(_02345_),
    .A2(_02351_),
    .ZN(io_imem_req_bits_pc[9])
  );
  AND2_X1 _18784_ (
    .A1(csr_io_evec[10]),
    .A2(_04026_),
    .ZN(_02352_)
  );
  MUX2_X1 _18785_ (
    .A(mem_reg_wdata[10]),
    .B(_06529_),
    .S(_03030_),
    .Z(_02353_)
  );
  INV_X1 _18786_ (
    .A(_02353_),
    .ZN(_02354_)
  );
  OR2_X1 _18787_ (
    .A1(_03142_),
    .A2(_02353_),
    .ZN(_02355_)
  );
  OR2_X1 _18788_ (
    .A1(wb_reg_pc[10]),
    .A2(_03141_),
    .ZN(_02356_)
  );
  AND2_X1 _18789_ (
    .A1(_04025_),
    .A2(_02356_),
    .ZN(_02357_)
  );
  AND2_X1 _18790_ (
    .A1(_02355_),
    .A2(_02357_),
    .ZN(_02358_)
  );
  OR2_X1 _18791_ (
    .A1(_02352_),
    .A2(_02358_),
    .ZN(io_imem_req_bits_pc[10])
  );
  AND2_X1 _18792_ (
    .A1(csr_io_evec[11]),
    .A2(_04026_),
    .ZN(_02359_)
  );
  MUX2_X1 _18793_ (
    .A(mem_reg_wdata[11]),
    .B(_06541_),
    .S(_03030_),
    .Z(_02360_)
  );
  INV_X1 _18794_ (
    .A(_02360_),
    .ZN(_02361_)
  );
  OR2_X1 _18795_ (
    .A1(_03142_),
    .A2(_02360_),
    .ZN(_02362_)
  );
  OR2_X1 _18796_ (
    .A1(wb_reg_pc[11]),
    .A2(_03141_),
    .ZN(_02363_)
  );
  AND2_X1 _18797_ (
    .A1(_04025_),
    .A2(_02363_),
    .ZN(_02364_)
  );
  AND2_X1 _18798_ (
    .A1(_02362_),
    .A2(_02364_),
    .ZN(_02365_)
  );
  OR2_X1 _18799_ (
    .A1(_02359_),
    .A2(_02365_),
    .ZN(io_imem_req_bits_pc[11])
  );
  AND2_X1 _18800_ (
    .A1(csr_io_evec[12]),
    .A2(_04026_),
    .ZN(_02366_)
  );
  MUX2_X1 _18801_ (
    .A(mem_reg_wdata[12]),
    .B(_06554_),
    .S(_03030_),
    .Z(_02367_)
  );
  INV_X1 _18802_ (
    .A(_02367_),
    .ZN(_02368_)
  );
  OR2_X1 _18803_ (
    .A1(_03142_),
    .A2(_02367_),
    .ZN(_02369_)
  );
  OR2_X1 _18804_ (
    .A1(wb_reg_pc[12]),
    .A2(_03141_),
    .ZN(_02370_)
  );
  AND2_X1 _18805_ (
    .A1(_04025_),
    .A2(_02370_),
    .ZN(_02371_)
  );
  AND2_X1 _18806_ (
    .A1(_02369_),
    .A2(_02371_),
    .ZN(_02372_)
  );
  OR2_X1 _18807_ (
    .A1(_02366_),
    .A2(_02372_),
    .ZN(io_imem_req_bits_pc[12])
  );
  AND2_X1 _18808_ (
    .A1(csr_io_evec[13]),
    .A2(_04026_),
    .ZN(_02373_)
  );
  MUX2_X1 _18809_ (
    .A(mem_reg_wdata[13]),
    .B(_06566_),
    .S(_03030_),
    .Z(_02374_)
  );
  INV_X1 _18810_ (
    .A(_02374_),
    .ZN(_02375_)
  );
  OR2_X1 _18811_ (
    .A1(_03142_),
    .A2(_02374_),
    .ZN(_02376_)
  );
  OR2_X1 _18812_ (
    .A1(wb_reg_pc[13]),
    .A2(_03141_),
    .ZN(_02377_)
  );
  AND2_X1 _18813_ (
    .A1(_04025_),
    .A2(_02377_),
    .ZN(_02378_)
  );
  AND2_X1 _18814_ (
    .A1(_02376_),
    .A2(_02378_),
    .ZN(_02379_)
  );
  OR2_X1 _18815_ (
    .A1(_02373_),
    .A2(_02379_),
    .ZN(io_imem_req_bits_pc[13])
  );
  AND2_X1 _18816_ (
    .A1(csr_io_evec[14]),
    .A2(_04026_),
    .ZN(_02380_)
  );
  MUX2_X1 _18817_ (
    .A(mem_reg_wdata[14]),
    .B(_06579_),
    .S(_03030_),
    .Z(_02381_)
  );
  INV_X1 _18818_ (
    .A(_02381_),
    .ZN(_02382_)
  );
  OR2_X1 _18819_ (
    .A1(_03142_),
    .A2(_02381_),
    .ZN(_02383_)
  );
  OR2_X1 _18820_ (
    .A1(wb_reg_pc[14]),
    .A2(_03141_),
    .ZN(_02384_)
  );
  AND2_X1 _18821_ (
    .A1(_04025_),
    .A2(_02384_),
    .ZN(_02385_)
  );
  AND2_X1 _18822_ (
    .A1(_02383_),
    .A2(_02385_),
    .ZN(_02386_)
  );
  OR2_X1 _18823_ (
    .A1(_02380_),
    .A2(_02386_),
    .ZN(io_imem_req_bits_pc[14])
  );
  AND2_X1 _18824_ (
    .A1(csr_io_evec[15]),
    .A2(_04026_),
    .ZN(_02387_)
  );
  MUX2_X1 _18825_ (
    .A(mem_reg_wdata[15]),
    .B(_06591_),
    .S(_03030_),
    .Z(_02388_)
  );
  INV_X1 _18826_ (
    .A(_02388_),
    .ZN(_02389_)
  );
  OR2_X1 _18827_ (
    .A1(_03142_),
    .A2(_02388_),
    .ZN(_02390_)
  );
  OR2_X1 _18828_ (
    .A1(wb_reg_pc[15]),
    .A2(_03141_),
    .ZN(_02391_)
  );
  AND2_X1 _18829_ (
    .A1(_04025_),
    .A2(_02391_),
    .ZN(_02392_)
  );
  AND2_X1 _18830_ (
    .A1(_02390_),
    .A2(_02392_),
    .ZN(_02393_)
  );
  OR2_X1 _18831_ (
    .A1(_02387_),
    .A2(_02393_),
    .ZN(io_imem_req_bits_pc[15])
  );
  AND2_X1 _18832_ (
    .A1(csr_io_evec[16]),
    .A2(_04026_),
    .ZN(_02394_)
  );
  MUX2_X1 _18833_ (
    .A(mem_reg_wdata[16]),
    .B(_06604_),
    .S(_03030_),
    .Z(_02395_)
  );
  INV_X1 _18834_ (
    .A(_02395_),
    .ZN(_02396_)
  );
  OR2_X1 _18835_ (
    .A1(_03142_),
    .A2(_02395_),
    .ZN(_02397_)
  );
  OR2_X1 _18836_ (
    .A1(wb_reg_pc[16]),
    .A2(_03141_),
    .ZN(_02398_)
  );
  AND2_X1 _18837_ (
    .A1(_04025_),
    .A2(_02398_),
    .ZN(_02399_)
  );
  AND2_X1 _18838_ (
    .A1(_02397_),
    .A2(_02399_),
    .ZN(_02400_)
  );
  OR2_X1 _18839_ (
    .A1(_02394_),
    .A2(_02400_),
    .ZN(io_imem_req_bits_pc[16])
  );
  AND2_X1 _18840_ (
    .A1(csr_io_evec[17]),
    .A2(_04026_),
    .ZN(_02401_)
  );
  MUX2_X1 _18841_ (
    .A(mem_reg_wdata[17]),
    .B(_06616_),
    .S(_03030_),
    .Z(_02402_)
  );
  INV_X1 _18842_ (
    .A(_02402_),
    .ZN(_02403_)
  );
  OR2_X1 _18843_ (
    .A1(_03142_),
    .A2(_02402_),
    .ZN(_02404_)
  );
  OR2_X1 _18844_ (
    .A1(wb_reg_pc[17]),
    .A2(_03141_),
    .ZN(_02405_)
  );
  AND2_X1 _18845_ (
    .A1(_04025_),
    .A2(_02405_),
    .ZN(_02406_)
  );
  AND2_X1 _18846_ (
    .A1(_02404_),
    .A2(_02406_),
    .ZN(_02407_)
  );
  OR2_X1 _18847_ (
    .A1(_02401_),
    .A2(_02407_),
    .ZN(io_imem_req_bits_pc[17])
  );
  AND2_X1 _18848_ (
    .A1(csr_io_evec[18]),
    .A2(_04026_),
    .ZN(_02408_)
  );
  MUX2_X1 _18849_ (
    .A(mem_reg_wdata[18]),
    .B(_06629_),
    .S(_03030_),
    .Z(_02409_)
  );
  OR2_X1 _18850_ (
    .A1(_03142_),
    .A2(_02409_),
    .ZN(_02410_)
  );
  OR2_X1 _18851_ (
    .A1(wb_reg_pc[18]),
    .A2(_03141_),
    .ZN(_02411_)
  );
  AND2_X1 _18852_ (
    .A1(_04025_),
    .A2(_02411_),
    .ZN(_02412_)
  );
  AND2_X1 _18853_ (
    .A1(_02410_),
    .A2(_02412_),
    .ZN(_02413_)
  );
  OR2_X1 _18854_ (
    .A1(_02408_),
    .A2(_02413_),
    .ZN(io_imem_req_bits_pc[18])
  );
  AND2_X1 _18855_ (
    .A1(csr_io_evec[19]),
    .A2(_04026_),
    .ZN(_02414_)
  );
  MUX2_X1 _18856_ (
    .A(mem_reg_wdata[19]),
    .B(_06641_),
    .S(_03030_),
    .Z(_02415_)
  );
  OR2_X1 _18857_ (
    .A1(_03142_),
    .A2(_02415_),
    .ZN(_02416_)
  );
  OR2_X1 _18858_ (
    .A1(wb_reg_pc[19]),
    .A2(_03141_),
    .ZN(_02417_)
  );
  AND2_X1 _18859_ (
    .A1(_04025_),
    .A2(_02417_),
    .ZN(_02418_)
  );
  AND2_X1 _18860_ (
    .A1(_02416_),
    .A2(_02418_),
    .ZN(_02419_)
  );
  OR2_X1 _18861_ (
    .A1(_02414_),
    .A2(_02419_),
    .ZN(io_imem_req_bits_pc[19])
  );
  AND2_X1 _18862_ (
    .A1(csr_io_evec[20]),
    .A2(_04026_),
    .ZN(_02420_)
  );
  MUX2_X1 _18863_ (
    .A(mem_reg_wdata[20]),
    .B(_06653_),
    .S(_03030_),
    .Z(_02421_)
  );
  OR2_X1 _18864_ (
    .A1(_03142_),
    .A2(_02421_),
    .ZN(_02422_)
  );
  OR2_X1 _18865_ (
    .A1(wb_reg_pc[20]),
    .A2(_03141_),
    .ZN(_02423_)
  );
  AND2_X1 _18866_ (
    .A1(_04025_),
    .A2(_02423_),
    .ZN(_02424_)
  );
  AND2_X1 _18867_ (
    .A1(_02422_),
    .A2(_02424_),
    .ZN(_02425_)
  );
  OR2_X1 _18868_ (
    .A1(_02420_),
    .A2(_02425_),
    .ZN(io_imem_req_bits_pc[20])
  );
  AND2_X1 _18869_ (
    .A1(csr_io_evec[21]),
    .A2(_04026_),
    .ZN(_02426_)
  );
  MUX2_X1 _18870_ (
    .A(mem_reg_wdata[21]),
    .B(_06662_),
    .S(_03030_),
    .Z(_02427_)
  );
  OR2_X1 _18871_ (
    .A1(_03142_),
    .A2(_02427_),
    .ZN(_02428_)
  );
  OR2_X1 _18872_ (
    .A1(wb_reg_pc[21]),
    .A2(_03141_),
    .ZN(_02429_)
  );
  AND2_X1 _18873_ (
    .A1(_04025_),
    .A2(_02429_),
    .ZN(_02430_)
  );
  AND2_X1 _18874_ (
    .A1(_02428_),
    .A2(_02430_),
    .ZN(_02431_)
  );
  OR2_X1 _18875_ (
    .A1(_02426_),
    .A2(_02431_),
    .ZN(io_imem_req_bits_pc[21])
  );
  AND2_X1 _18876_ (
    .A1(csr_io_evec[22]),
    .A2(_04026_),
    .ZN(_02432_)
  );
  MUX2_X1 _18877_ (
    .A(mem_reg_wdata[22]),
    .B(_06674_),
    .S(_03030_),
    .Z(_02433_)
  );
  OR2_X1 _18878_ (
    .A1(_03142_),
    .A2(_02433_),
    .ZN(_02434_)
  );
  OR2_X1 _18879_ (
    .A1(wb_reg_pc[22]),
    .A2(_03141_),
    .ZN(_02435_)
  );
  AND2_X1 _18880_ (
    .A1(_04025_),
    .A2(_02435_),
    .ZN(_02436_)
  );
  AND2_X1 _18881_ (
    .A1(_02434_),
    .A2(_02436_),
    .ZN(_02437_)
  );
  OR2_X1 _18882_ (
    .A1(_02432_),
    .A2(_02437_),
    .ZN(io_imem_req_bits_pc[22])
  );
  AND2_X1 _18883_ (
    .A1(csr_io_evec[23]),
    .A2(_04026_),
    .ZN(_02438_)
  );
  MUX2_X1 _18884_ (
    .A(mem_reg_wdata[23]),
    .B(_06683_),
    .S(_03030_),
    .Z(_02439_)
  );
  OR2_X1 _18885_ (
    .A1(_03142_),
    .A2(_02439_),
    .ZN(_02440_)
  );
  OR2_X1 _18886_ (
    .A1(wb_reg_pc[23]),
    .A2(_03141_),
    .ZN(_02441_)
  );
  AND2_X1 _18887_ (
    .A1(_04025_),
    .A2(_02441_),
    .ZN(_02442_)
  );
  AND2_X1 _18888_ (
    .A1(_02440_),
    .A2(_02442_),
    .ZN(_02443_)
  );
  OR2_X1 _18889_ (
    .A1(_02438_),
    .A2(_02443_),
    .ZN(io_imem_req_bits_pc[23])
  );
  AND2_X1 _18890_ (
    .A1(csr_io_evec[24]),
    .A2(_04026_),
    .ZN(_02444_)
  );
  MUX2_X1 _18891_ (
    .A(mem_reg_wdata[24]),
    .B(_06698_),
    .S(_03030_),
    .Z(_02445_)
  );
  OR2_X1 _18892_ (
    .A1(_03142_),
    .A2(_02445_),
    .ZN(_02446_)
  );
  OR2_X1 _18893_ (
    .A1(wb_reg_pc[24]),
    .A2(_03141_),
    .ZN(_02447_)
  );
  AND2_X1 _18894_ (
    .A1(_04025_),
    .A2(_02447_),
    .ZN(_02448_)
  );
  AND2_X1 _18895_ (
    .A1(_02446_),
    .A2(_02448_),
    .ZN(_02449_)
  );
  OR2_X1 _18896_ (
    .A1(_02444_),
    .A2(_02449_),
    .ZN(io_imem_req_bits_pc[24])
  );
  AND2_X1 _18897_ (
    .A1(csr_io_evec[25]),
    .A2(_04026_),
    .ZN(_02450_)
  );
  MUX2_X1 _18898_ (
    .A(mem_reg_wdata[25]),
    .B(_06707_),
    .S(_03030_),
    .Z(_02451_)
  );
  OR2_X1 _18899_ (
    .A1(_03142_),
    .A2(_02451_),
    .ZN(_02452_)
  );
  OR2_X1 _18900_ (
    .A1(wb_reg_pc[25]),
    .A2(_03141_),
    .ZN(_02453_)
  );
  AND2_X1 _18901_ (
    .A1(_04025_),
    .A2(_02453_),
    .ZN(_02454_)
  );
  AND2_X1 _18902_ (
    .A1(_02452_),
    .A2(_02454_),
    .ZN(_02455_)
  );
  OR2_X1 _18903_ (
    .A1(_02450_),
    .A2(_02455_),
    .ZN(io_imem_req_bits_pc[25])
  );
  AND2_X1 _18904_ (
    .A1(csr_io_evec[26]),
    .A2(_04026_),
    .ZN(_02456_)
  );
  MUX2_X1 _18905_ (
    .A(mem_reg_wdata[26]),
    .B(_06719_),
    .S(_03030_),
    .Z(_02457_)
  );
  OR2_X1 _18906_ (
    .A1(_03142_),
    .A2(_02457_),
    .ZN(_02458_)
  );
  OR2_X1 _18907_ (
    .A1(wb_reg_pc[26]),
    .A2(_03141_),
    .ZN(_02459_)
  );
  AND2_X1 _18908_ (
    .A1(_04025_),
    .A2(_02459_),
    .ZN(_02460_)
  );
  AND2_X1 _18909_ (
    .A1(_02458_),
    .A2(_02460_),
    .ZN(_02461_)
  );
  OR2_X1 _18910_ (
    .A1(_02456_),
    .A2(_02461_),
    .ZN(io_imem_req_bits_pc[26])
  );
  AND2_X1 _18911_ (
    .A1(csr_io_evec[27]),
    .A2(_04026_),
    .ZN(_02462_)
  );
  MUX2_X1 _18912_ (
    .A(mem_reg_wdata[27]),
    .B(_06728_),
    .S(_03030_),
    .Z(_02463_)
  );
  OR2_X1 _18913_ (
    .A1(_03142_),
    .A2(_02463_),
    .ZN(_02464_)
  );
  OR2_X1 _18914_ (
    .A1(wb_reg_pc[27]),
    .A2(_03141_),
    .ZN(_02465_)
  );
  AND2_X1 _18915_ (
    .A1(_04025_),
    .A2(_02465_),
    .ZN(_02466_)
  );
  AND2_X1 _18916_ (
    .A1(_02464_),
    .A2(_02466_),
    .ZN(_02467_)
  );
  OR2_X1 _18917_ (
    .A1(_02462_),
    .A2(_02467_),
    .ZN(io_imem_req_bits_pc[27])
  );
  AND2_X1 _18918_ (
    .A1(csr_io_evec[28]),
    .A2(_04026_),
    .ZN(_02468_)
  );
  MUX2_X1 _18919_ (
    .A(_02981_),
    .B(_06745_),
    .S(_03030_),
    .Z(_02469_)
  );
  MUX2_X1 _18920_ (
    .A(mem_reg_wdata[28]),
    .B(_06744_),
    .S(_03030_),
    .Z(_02470_)
  );
  OR2_X1 _18921_ (
    .A1(_03142_),
    .A2(_02470_),
    .ZN(_02471_)
  );
  OR2_X1 _18922_ (
    .A1(wb_reg_pc[28]),
    .A2(_03141_),
    .ZN(_02472_)
  );
  AND2_X1 _18923_ (
    .A1(_04025_),
    .A2(_02472_),
    .ZN(_02473_)
  );
  AND2_X1 _18924_ (
    .A1(_02471_),
    .A2(_02473_),
    .ZN(_02474_)
  );
  OR2_X1 _18925_ (
    .A1(_02468_),
    .A2(_02474_),
    .ZN(io_imem_req_bits_pc[28])
  );
  AND2_X1 _18926_ (
    .A1(csr_io_evec[29]),
    .A2(_04026_),
    .ZN(_02475_)
  );
  MUX2_X1 _18927_ (
    .A(mem_reg_wdata[29]),
    .B(_06755_),
    .S(_03030_),
    .Z(_02476_)
  );
  OR2_X1 _18928_ (
    .A1(_03142_),
    .A2(_02476_),
    .ZN(_02477_)
  );
  OR2_X1 _18929_ (
    .A1(wb_reg_pc[29]),
    .A2(_03141_),
    .ZN(_02478_)
  );
  AND2_X1 _18930_ (
    .A1(_04025_),
    .A2(_02478_),
    .ZN(_02479_)
  );
  AND2_X1 _18931_ (
    .A1(_02477_),
    .A2(_02479_),
    .ZN(_02480_)
  );
  OR2_X1 _18932_ (
    .A1(_02475_),
    .A2(_02480_),
    .ZN(io_imem_req_bits_pc[29])
  );
  AND2_X1 _18933_ (
    .A1(csr_io_evec[30]),
    .A2(_04026_),
    .ZN(_02481_)
  );
  MUX2_X1 _18934_ (
    .A(mem_reg_wdata[30]),
    .B(_06766_),
    .S(_03030_),
    .Z(_02482_)
  );
  OR2_X1 _18935_ (
    .A1(_03142_),
    .A2(_02482_),
    .ZN(_02483_)
  );
  OR2_X1 _18936_ (
    .A1(wb_reg_pc[30]),
    .A2(_03141_),
    .ZN(_02484_)
  );
  AND2_X1 _18937_ (
    .A1(_04025_),
    .A2(_02484_),
    .ZN(_02485_)
  );
  AND2_X1 _18938_ (
    .A1(_02483_),
    .A2(_02485_),
    .ZN(_02486_)
  );
  OR2_X1 _18939_ (
    .A1(_02481_),
    .A2(_02486_),
    .ZN(io_imem_req_bits_pc[30])
  );
  AND2_X1 _18940_ (
    .A1(csr_io_evec[31]),
    .A2(_04026_),
    .ZN(_02487_)
  );
  MUX2_X1 _18941_ (
    .A(mem_reg_wdata[31]),
    .B(_06774_),
    .S(_03030_),
    .Z(_02488_)
  );
  OR2_X1 _18942_ (
    .A1(_03142_),
    .A2(_02488_),
    .ZN(_02489_)
  );
  OR2_X1 _18943_ (
    .A1(wb_reg_pc[31]),
    .A2(_03141_),
    .ZN(_02490_)
  );
  AND2_X1 _18944_ (
    .A1(_04025_),
    .A2(_02490_),
    .ZN(_02491_)
  );
  AND2_X1 _18945_ (
    .A1(_02489_),
    .A2(_02491_),
    .ZN(_02492_)
  );
  OR2_X1 _18946_ (
    .A1(_02487_),
    .A2(_02492_),
    .ZN(io_imem_req_bits_pc[31])
  );
  OR2_X1 _18947_ (
    .A1(wb_reg_cause[0]),
    .A2(_03076_),
    .ZN(_02493_)
  );
  AND2_X1 _18948_ (
    .A1(_03136_),
    .A2(_02493_),
    .ZN(csr_io_cause[0])
  );
  AND2_X1 _18949_ (
    .A1(_03089_),
    .A2(_03138_),
    .ZN(_02494_)
  );
  OR2_X1 _18950_ (
    .A1(_03134_),
    .A2(_02494_),
    .ZN(_02495_)
  );
  AND2_X1 _18951_ (
    .A1(_03131_),
    .A2(_02495_),
    .ZN(_02496_)
  );
  MUX2_X1 _18952_ (
    .A(wb_reg_cause[1]),
    .B(_03128_),
    .S(_03076_),
    .Z(_02497_)
  );
  OR2_X1 _18953_ (
    .A1(_02496_),
    .A2(_02497_),
    .ZN(csr_io_cause[1])
  );
  OR2_X1 _18954_ (
    .A1(wb_reg_cause[2]),
    .A2(_03076_),
    .ZN(csr_io_cause[2])
  );
  OR2_X1 _18955_ (
    .A1(wb_reg_cause[3]),
    .A2(_03076_),
    .ZN(_02498_)
  );
  AND2_X1 _18956_ (
    .A1(_03132_),
    .A2(_02498_),
    .ZN(csr_io_cause[3])
  );
  AND2_X1 _18957_ (
    .A1(wb_reg_cause[4]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[4])
  );
  AND2_X1 _18958_ (
    .A1(wb_reg_cause[5]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[5])
  );
  AND2_X1 _18959_ (
    .A1(wb_reg_cause[6]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[6])
  );
  AND2_X1 _18960_ (
    .A1(wb_reg_cause[7]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[7])
  );
  AND2_X1 _18961_ (
    .A1(wb_reg_cause[8]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[8])
  );
  AND2_X1 _18962_ (
    .A1(wb_reg_cause[9]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[9])
  );
  AND2_X1 _18963_ (
    .A1(wb_reg_cause[10]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[10])
  );
  AND2_X1 _18964_ (
    .A1(wb_reg_cause[11]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[11])
  );
  AND2_X1 _18965_ (
    .A1(wb_reg_cause[12]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[12])
  );
  AND2_X1 _18966_ (
    .A1(wb_reg_cause[13]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[13])
  );
  AND2_X1 _18967_ (
    .A1(wb_reg_cause[14]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[14])
  );
  AND2_X1 _18968_ (
    .A1(wb_reg_cause[15]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[15])
  );
  AND2_X1 _18969_ (
    .A1(wb_reg_cause[16]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[16])
  );
  AND2_X1 _18970_ (
    .A1(wb_reg_cause[17]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[17])
  );
  AND2_X1 _18971_ (
    .A1(wb_reg_cause[18]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[18])
  );
  AND2_X1 _18972_ (
    .A1(wb_reg_cause[19]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[19])
  );
  AND2_X1 _18973_ (
    .A1(wb_reg_cause[20]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[20])
  );
  AND2_X1 _18974_ (
    .A1(wb_reg_cause[21]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[21])
  );
  AND2_X1 _18975_ (
    .A1(wb_reg_cause[22]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[22])
  );
  AND2_X1 _18976_ (
    .A1(wb_reg_cause[23]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[23])
  );
  AND2_X1 _18977_ (
    .A1(wb_reg_cause[24]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[24])
  );
  AND2_X1 _18978_ (
    .A1(wb_reg_cause[25]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[25])
  );
  AND2_X1 _18979_ (
    .A1(wb_reg_cause[26]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[26])
  );
  AND2_X1 _18980_ (
    .A1(wb_reg_cause[27]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[27])
  );
  AND2_X1 _18981_ (
    .A1(wb_reg_cause[28]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[28])
  );
  AND2_X1 _18982_ (
    .A1(wb_reg_cause[29]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[29])
  );
  AND2_X1 _18983_ (
    .A1(wb_reg_cause[30]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[30])
  );
  AND2_X1 _18984_ (
    .A1(wb_reg_cause[31]),
    .A2(wb_reg_xcpt),
    .ZN(csr_io_cause[31])
  );
  OR2_X1 _18985_ (
    .A1(wb_reg_cause[4]),
    .A2(wb_reg_cause[2]),
    .ZN(_02499_)
  );
  OR2_X1 _18986_ (
    .A1(wb_reg_cause[3]),
    .A2(_02499_),
    .ZN(_02500_)
  );
  OR2_X1 _18987_ (
    .A1(_00015_),
    .A2(_02500_),
    .ZN(_02501_)
  );
  OR2_X1 _18988_ (
    .A1(wb_reg_cause[3]),
    .A2(_00030_),
    .ZN(_02502_)
  );
  OR2_X1 _18989_ (
    .A1(wb_reg_cause[4]),
    .A2(_00013_),
    .ZN(_02503_)
  );
  AND2_X1 _18990_ (
    .A1(_02502_),
    .A2(_02503_),
    .ZN(_02504_)
  );
  OR2_X1 _18991_ (
    .A1(wb_reg_cause[1]),
    .A2(_00014_),
    .ZN(_02505_)
  );
  OR2_X1 _18992_ (
    .A1(_02504_),
    .A2(_02505_),
    .ZN(_02506_)
  );
  AND2_X1 _18993_ (
    .A1(_02501_),
    .A2(_02506_),
    .ZN(_02507_)
  );
  OR2_X1 _18994_ (
    .A1(wb_reg_cause[0]),
    .A2(_02507_),
    .ZN(_02508_)
  );
  AND2_X1 _18995_ (
    .A1(wb_reg_cause[1]),
    .A2(_00015_),
    .ZN(_02509_)
  );
  OR2_X1 _18996_ (
    .A1(_00016_),
    .A2(_02509_),
    .ZN(_02510_)
  );
  OR2_X1 _18997_ (
    .A1(_02500_),
    .A2(_02510_),
    .ZN(_02511_)
  );
  AND2_X1 _18998_ (
    .A1(_02508_),
    .A2(_02511_),
    .ZN(_02512_)
  );
  OR2_X1 _18999_ (
    .A1(wb_reg_cause[29]),
    .A2(wb_reg_cause[30]),
    .ZN(_02513_)
  );
  OR2_X1 _19000_ (
    .A1(wb_reg_cause[31]),
    .A2(_02513_),
    .ZN(_02514_)
  );
  OR2_X1 _19001_ (
    .A1(wb_reg_cause[25]),
    .A2(wb_reg_cause[26]),
    .ZN(_02515_)
  );
  OR2_X1 _19002_ (
    .A1(wb_reg_cause[27]),
    .A2(wb_reg_cause[28]),
    .ZN(_02516_)
  );
  OR2_X1 _19003_ (
    .A1(_02515_),
    .A2(_02516_),
    .ZN(_02517_)
  );
  OR2_X1 _19004_ (
    .A1(wb_reg_cause[21]),
    .A2(wb_reg_cause[22]),
    .ZN(_02518_)
  );
  OR2_X1 _19005_ (
    .A1(wb_reg_cause[23]),
    .A2(wb_reg_cause[24]),
    .ZN(_02519_)
  );
  OR2_X1 _19006_ (
    .A1(_02518_),
    .A2(_02519_),
    .ZN(_02520_)
  );
  OR2_X1 _19007_ (
    .A1(_02517_),
    .A2(_02520_),
    .ZN(_02521_)
  );
  OR2_X1 _19008_ (
    .A1(_02514_),
    .A2(_02521_),
    .ZN(_02522_)
  );
  OR2_X1 _19009_ (
    .A1(wb_reg_cause[19]),
    .A2(wb_reg_cause[20]),
    .ZN(_02523_)
  );
  OR2_X1 _19010_ (
    .A1(wb_reg_cause[17]),
    .A2(wb_reg_cause[18]),
    .ZN(_02524_)
  );
  OR2_X1 _19011_ (
    .A1(_02523_),
    .A2(_02524_),
    .ZN(_02525_)
  );
  OR2_X1 _19012_ (
    .A1(wb_reg_cause[13]),
    .A2(wb_reg_cause[14]),
    .ZN(_02526_)
  );
  OR2_X1 _19013_ (
    .A1(wb_reg_cause[15]),
    .A2(wb_reg_cause[16]),
    .ZN(_02527_)
  );
  OR2_X1 _19014_ (
    .A1(_02526_),
    .A2(_02527_),
    .ZN(_02528_)
  );
  OR2_X1 _19015_ (
    .A1(_02525_),
    .A2(_02528_),
    .ZN(_02529_)
  );
  OR2_X1 _19016_ (
    .A1(wb_reg_cause[11]),
    .A2(wb_reg_cause[12]),
    .ZN(_02530_)
  );
  OR2_X1 _19017_ (
    .A1(wb_reg_cause[9]),
    .A2(wb_reg_cause[10]),
    .ZN(_02531_)
  );
  OR2_X1 _19018_ (
    .A1(_02530_),
    .A2(_02531_),
    .ZN(_02532_)
  );
  OR2_X1 _19019_ (
    .A1(wb_reg_cause[5]),
    .A2(wb_reg_cause[6]),
    .ZN(_02533_)
  );
  OR2_X1 _19020_ (
    .A1(wb_reg_cause[7]),
    .A2(wb_reg_cause[8]),
    .ZN(_02534_)
  );
  OR2_X1 _19021_ (
    .A1(_02533_),
    .A2(_02534_),
    .ZN(_02535_)
  );
  OR2_X1 _19022_ (
    .A1(_02532_),
    .A2(_02535_),
    .ZN(_02536_)
  );
  OR2_X1 _19023_ (
    .A1(_02529_),
    .A2(_02536_),
    .ZN(_02537_)
  );
  OR2_X1 _19024_ (
    .A1(_02522_),
    .A2(_02537_),
    .ZN(_02538_)
  );
  OR2_X1 _19025_ (
    .A1(_02512_),
    .A2(_02538_),
    .ZN(_02539_)
  );
  INV_X1 _19026_ (
    .A(_02539_),
    .ZN(_02540_)
  );
  OR2_X1 _19027_ (
    .A1(tval_dmem_addr),
    .A2(_02540_),
    .ZN(_02541_)
  );
  AND2_X1 _19028_ (
    .A1(csr_io_exception),
    .A2(_02541_),
    .ZN(_02542_)
  );
  AND2_X1 _19029_ (
    .A1(wb_reg_wdata[0]),
    .A2(_02542_),
    .ZN(csr_io_tval[0])
  );
  AND2_X1 _19030_ (
    .A1(wb_reg_wdata[1]),
    .A2(_02542_),
    .ZN(csr_io_tval[1])
  );
  AND2_X1 _19031_ (
    .A1(wb_reg_wdata[2]),
    .A2(_02542_),
    .ZN(csr_io_tval[2])
  );
  AND2_X1 _19032_ (
    .A1(wb_reg_wdata[3]),
    .A2(_02542_),
    .ZN(csr_io_tval[3])
  );
  AND2_X1 _19033_ (
    .A1(wb_reg_wdata[4]),
    .A2(_02542_),
    .ZN(csr_io_tval[4])
  );
  AND2_X1 _19034_ (
    .A1(wb_reg_wdata[5]),
    .A2(_02542_),
    .ZN(csr_io_tval[5])
  );
  AND2_X1 _19035_ (
    .A1(wb_reg_wdata[6]),
    .A2(_02542_),
    .ZN(csr_io_tval[6])
  );
  AND2_X1 _19036_ (
    .A1(wb_reg_wdata[7]),
    .A2(_02542_),
    .ZN(csr_io_tval[7])
  );
  AND2_X1 _19037_ (
    .A1(wb_reg_wdata[8]),
    .A2(_02542_),
    .ZN(csr_io_tval[8])
  );
  AND2_X1 _19038_ (
    .A1(wb_reg_wdata[9]),
    .A2(_02542_),
    .ZN(csr_io_tval[9])
  );
  AND2_X1 _19039_ (
    .A1(wb_reg_wdata[10]),
    .A2(_02542_),
    .ZN(csr_io_tval[10])
  );
  AND2_X1 _19040_ (
    .A1(wb_reg_wdata[11]),
    .A2(_02542_),
    .ZN(csr_io_tval[11])
  );
  AND2_X1 _19041_ (
    .A1(wb_reg_wdata[12]),
    .A2(_02542_),
    .ZN(csr_io_tval[12])
  );
  AND2_X1 _19042_ (
    .A1(wb_reg_wdata[13]),
    .A2(_02542_),
    .ZN(csr_io_tval[13])
  );
  AND2_X1 _19043_ (
    .A1(wb_reg_wdata[14]),
    .A2(_02542_),
    .ZN(csr_io_tval[14])
  );
  AND2_X1 _19044_ (
    .A1(wb_reg_wdata[15]),
    .A2(_02542_),
    .ZN(csr_io_tval[15])
  );
  AND2_X1 _19045_ (
    .A1(wb_reg_wdata[16]),
    .A2(_02542_),
    .ZN(csr_io_tval[16])
  );
  AND2_X1 _19046_ (
    .A1(wb_reg_wdata[17]),
    .A2(_02542_),
    .ZN(csr_io_tval[17])
  );
  AND2_X1 _19047_ (
    .A1(wb_reg_wdata[18]),
    .A2(_02542_),
    .ZN(csr_io_tval[18])
  );
  AND2_X1 _19048_ (
    .A1(wb_reg_wdata[19]),
    .A2(_02542_),
    .ZN(csr_io_tval[19])
  );
  AND2_X1 _19049_ (
    .A1(wb_reg_wdata[20]),
    .A2(_02542_),
    .ZN(csr_io_tval[20])
  );
  AND2_X1 _19050_ (
    .A1(wb_reg_wdata[21]),
    .A2(_02542_),
    .ZN(csr_io_tval[21])
  );
  AND2_X1 _19051_ (
    .A1(wb_reg_wdata[22]),
    .A2(_02542_),
    .ZN(csr_io_tval[22])
  );
  AND2_X1 _19052_ (
    .A1(wb_reg_wdata[23]),
    .A2(_02542_),
    .ZN(csr_io_tval[23])
  );
  AND2_X1 _19053_ (
    .A1(wb_reg_wdata[24]),
    .A2(_02542_),
    .ZN(csr_io_tval[24])
  );
  AND2_X1 _19054_ (
    .A1(wb_reg_wdata[25]),
    .A2(_02542_),
    .ZN(csr_io_tval[25])
  );
  AND2_X1 _19055_ (
    .A1(wb_reg_wdata[26]),
    .A2(_02542_),
    .ZN(csr_io_tval[26])
  );
  AND2_X1 _19056_ (
    .A1(wb_reg_wdata[27]),
    .A2(_02542_),
    .ZN(csr_io_tval[27])
  );
  AND2_X1 _19057_ (
    .A1(wb_reg_wdata[28]),
    .A2(_02542_),
    .ZN(csr_io_tval[28])
  );
  AND2_X1 _19058_ (
    .A1(wb_reg_wdata[29]),
    .A2(_02542_),
    .ZN(csr_io_tval[29])
  );
  AND2_X1 _19059_ (
    .A1(wb_reg_wdata[30]),
    .A2(_02542_),
    .ZN(csr_io_tval[30])
  );
  AND2_X1 _19060_ (
    .A1(wb_reg_wdata[31]),
    .A2(_02542_),
    .ZN(csr_io_tval[31])
  );
  OR2_X1 _19061_ (
    .A1(ex_ctrl_sel_alu2[1]),
    .A2(_00018_),
    .ZN(_02543_)
  );
  OR2_X1 _19062_ (
    .A1(ex_ctrl_sel_alu2[0]),
    .A2(_00012_),
    .ZN(_02544_)
  );
  INV_X1 _19063_ (
    .A(_02544_),
    .ZN(_02545_)
  );
  AND2_X1 _19064_ (
    .A1(_00018_),
    .A2(_02545_),
    .ZN(_02546_)
  );
  AND2_X1 _19065_ (
    .A1(_ex_op2_T[0]),
    .A2(_02546_),
    .ZN(_02547_)
  );
  AND2_X1 _19066_ (
    .A1(_03042_),
    .A2(_03043_),
    .ZN(_02548_)
  );
  OR2_X1 _19067_ (
    .A1(ex_ctrl_sel_imm[0]),
    .A2(ex_ctrl_sel_imm[1]),
    .ZN(_02549_)
  );
  INV_X1 _19068_ (
    .A(_02549_),
    .ZN(_02550_)
  );
  OR2_X1 _19069_ (
    .A1(ex_ctrl_sel_imm[2]),
    .A2(_02549_),
    .ZN(_02551_)
  );
  OR2_X1 _19070_ (
    .A1(ex_ctrl_sel_imm[1]),
    .A2(_00023_),
    .ZN(_02552_)
  );
  OR2_X1 _19071_ (
    .A1(_00021_),
    .A2(_02552_),
    .ZN(_02553_)
  );
  INV_X1 _19072_ (
    .A(_02553_),
    .ZN(_02554_)
  );
  AND2_X1 _19073_ (
    .A1(ex_reg_inst[15]),
    .A2(_02549_),
    .ZN(_02555_)
  );
  AND2_X1 _19074_ (
    .A1(_02554_),
    .A2(_02555_),
    .ZN(_02556_)
  );
  AND2_X1 _19075_ (
    .A1(ex_reg_inst[20]),
    .A2(_03041_),
    .ZN(_02557_)
  );
  AND2_X1 _19076_ (
    .A1(_02550_),
    .A2(_02557_),
    .ZN(_02558_)
  );
  OR2_X1 _19077_ (
    .A1(_02556_),
    .A2(_02558_),
    .ZN(_02559_)
  );
  MUX2_X1 _19078_ (
    .A(ex_reg_inst[7]),
    .B(_02559_),
    .S(_02551_),
    .Z(_02560_)
  );
  AND2_X1 _19079_ (
    .A1(_02548_),
    .A2(_02560_),
    .ZN(_02561_)
  );
  OR2_X1 _19080_ (
    .A1(_02547_),
    .A2(_02561_),
    .ZN(_02562_)
  );
  AND2_X1 _19081_ (
    .A1(_02543_),
    .A2(_02562_),
    .ZN(alu_io_in2[0])
  );
  AND2_X1 _19082_ (
    .A1(_ex_op2_T[1]),
    .A2(_02546_),
    .ZN(_02563_)
  );
  OR2_X1 _19083_ (
    .A1(ex_ctrl_sel_imm[2]),
    .A2(_00022_),
    .ZN(_02564_)
  );
  OR2_X1 _19084_ (
    .A1(ex_ctrl_sel_imm[0]),
    .A2(_02564_),
    .ZN(_02565_)
  );
  AND2_X1 _19085_ (
    .A1(_02548_),
    .A2(_02565_),
    .ZN(_02566_)
  );
  OR2_X1 _19086_ (
    .A1(ex_ctrl_sel_imm[2]),
    .A2(_02552_),
    .ZN(_02567_)
  );
  AND2_X1 _19087_ (
    .A1(_02551_),
    .A2(_02567_),
    .ZN(_02568_)
  );
  INV_X1 _19088_ (
    .A(_02568_),
    .ZN(_02569_)
  );
  MUX2_X1 _19089_ (
    .A(ex_reg_inst[16]),
    .B(ex_reg_inst[21]),
    .S(_02553_),
    .Z(_02570_)
  );
  MUX2_X1 _19090_ (
    .A(ex_reg_inst[8]),
    .B(_02570_),
    .S(_02568_),
    .Z(_02571_)
  );
  AND2_X1 _19091_ (
    .A1(_02566_),
    .A2(_02571_),
    .ZN(_02572_)
  );
  OR2_X1 _19092_ (
    .A1(_02563_),
    .A2(_02572_),
    .ZN(_02573_)
  );
  MUX2_X1 _19093_ (
    .A(ex_reg_rvc),
    .B(_02573_),
    .S(_02543_),
    .Z(alu_io_in2[1])
  );
  AND2_X1 _19094_ (
    .A1(_ex_op2_T[2]),
    .A2(_02546_),
    .ZN(_02574_)
  );
  MUX2_X1 _19095_ (
    .A(ex_reg_inst[17]),
    .B(ex_reg_inst[22]),
    .S(_02553_),
    .Z(_02575_)
  );
  MUX2_X1 _19096_ (
    .A(ex_reg_inst[9]),
    .B(_02575_),
    .S(_02568_),
    .Z(_02576_)
  );
  AND2_X1 _19097_ (
    .A1(_02566_),
    .A2(_02576_),
    .ZN(_02577_)
  );
  OR2_X1 _19098_ (
    .A1(_02574_),
    .A2(_02577_),
    .ZN(_02578_)
  );
  MUX2_X1 _19099_ (
    .A(_ex_op2_T_1[2]),
    .B(_02578_),
    .S(_02543_),
    .Z(alu_io_in2[2])
  );
  AND2_X1 _19100_ (
    .A1(_ex_op2_T[3]),
    .A2(_02546_),
    .ZN(_02579_)
  );
  MUX2_X1 _19101_ (
    .A(ex_reg_inst[18]),
    .B(ex_reg_inst[23]),
    .S(_02553_),
    .Z(_02580_)
  );
  MUX2_X1 _19102_ (
    .A(ex_reg_inst[10]),
    .B(_02580_),
    .S(_02568_),
    .Z(_02581_)
  );
  AND2_X1 _19103_ (
    .A1(_02566_),
    .A2(_02581_),
    .ZN(_02582_)
  );
  OR2_X1 _19104_ (
    .A1(_02579_),
    .A2(_02582_),
    .ZN(_02583_)
  );
  AND2_X1 _19105_ (
    .A1(_02543_),
    .A2(_02583_),
    .ZN(alu_io_in2[3])
  );
  AND2_X1 _19106_ (
    .A1(_ex_op2_T[4]),
    .A2(_02546_),
    .ZN(_02584_)
  );
  MUX2_X1 _19107_ (
    .A(ex_reg_inst[19]),
    .B(ex_reg_inst[24]),
    .S(_02553_),
    .Z(_02585_)
  );
  OR2_X1 _19108_ (
    .A1(_02569_),
    .A2(_02585_),
    .ZN(_02586_)
  );
  OR2_X1 _19109_ (
    .A1(ex_reg_inst[11]),
    .A2(_02568_),
    .ZN(_02587_)
  );
  AND2_X1 _19110_ (
    .A1(_02566_),
    .A2(_02587_),
    .ZN(_02588_)
  );
  AND2_X1 _19111_ (
    .A1(_02586_),
    .A2(_02588_),
    .ZN(_02589_)
  );
  OR2_X1 _19112_ (
    .A1(_02584_),
    .A2(_02589_),
    .ZN(_02590_)
  );
  AND2_X1 _19113_ (
    .A1(_02543_),
    .A2(_02590_),
    .ZN(alu_io_in2[4])
  );
  AND2_X1 _19114_ (
    .A1(_02553_),
    .A2(_02566_),
    .ZN(_02591_)
  );
  AND2_X1 _19115_ (
    .A1(ex_reg_inst[25]),
    .A2(_02591_),
    .ZN(_02592_)
  );
  AND2_X1 _19116_ (
    .A1(_ex_op2_T[5]),
    .A2(_02546_),
    .ZN(_02593_)
  );
  OR2_X1 _19117_ (
    .A1(_02592_),
    .A2(_02593_),
    .ZN(_02594_)
  );
  AND2_X1 _19118_ (
    .A1(_02543_),
    .A2(_02594_),
    .ZN(alu_io_in2[5])
  );
  AND2_X1 _19119_ (
    .A1(ex_reg_inst[26]),
    .A2(_02591_),
    .ZN(_02595_)
  );
  AND2_X1 _19120_ (
    .A1(_ex_op2_T[6]),
    .A2(_02546_),
    .ZN(_02596_)
  );
  OR2_X1 _19121_ (
    .A1(_02595_),
    .A2(_02596_),
    .ZN(_02597_)
  );
  AND2_X1 _19122_ (
    .A1(_02543_),
    .A2(_02597_),
    .ZN(alu_io_in2[6])
  );
  AND2_X1 _19123_ (
    .A1(ex_reg_inst[27]),
    .A2(_02591_),
    .ZN(_02598_)
  );
  AND2_X1 _19124_ (
    .A1(_ex_op2_T[7]),
    .A2(_02546_),
    .ZN(_02599_)
  );
  OR2_X1 _19125_ (
    .A1(_02598_),
    .A2(_02599_),
    .ZN(_02600_)
  );
  AND2_X1 _19126_ (
    .A1(_02543_),
    .A2(_02600_),
    .ZN(alu_io_in2[7])
  );
  AND2_X1 _19127_ (
    .A1(ex_reg_inst[28]),
    .A2(_02591_),
    .ZN(_02601_)
  );
  AND2_X1 _19128_ (
    .A1(_ex_op2_T[8]),
    .A2(_02546_),
    .ZN(_02602_)
  );
  OR2_X1 _19129_ (
    .A1(_02601_),
    .A2(_02602_),
    .ZN(_02603_)
  );
  AND2_X1 _19130_ (
    .A1(_02543_),
    .A2(_02603_),
    .ZN(alu_io_in2[8])
  );
  AND2_X1 _19131_ (
    .A1(ex_reg_inst[29]),
    .A2(_02591_),
    .ZN(_02604_)
  );
  AND2_X1 _19132_ (
    .A1(_ex_op2_T[9]),
    .A2(_02546_),
    .ZN(_02605_)
  );
  OR2_X1 _19133_ (
    .A1(_02604_),
    .A2(_02605_),
    .ZN(_02606_)
  );
  AND2_X1 _19134_ (
    .A1(_02543_),
    .A2(_02606_),
    .ZN(alu_io_in2[9])
  );
  AND2_X1 _19135_ (
    .A1(ex_reg_inst[30]),
    .A2(_02591_),
    .ZN(_02607_)
  );
  AND2_X1 _19136_ (
    .A1(_ex_op2_T[10]),
    .A2(_02546_),
    .ZN(_02608_)
  );
  OR2_X1 _19137_ (
    .A1(_02607_),
    .A2(_02608_),
    .ZN(_02609_)
  );
  AND2_X1 _19138_ (
    .A1(_02543_),
    .A2(_02609_),
    .ZN(alu_io_in2[10])
  );
  AND2_X1 _19139_ (
    .A1(_ex_op2_T[11]),
    .A2(_02546_),
    .ZN(_02610_)
  );
  OR2_X1 _19140_ (
    .A1(_00023_),
    .A2(_02564_),
    .ZN(_02611_)
  );
  INV_X1 _19141_ (
    .A(_02611_),
    .ZN(_02612_)
  );
  AND2_X1 _19142_ (
    .A1(ex_reg_inst[31]),
    .A2(_02553_),
    .ZN(_02613_)
  );
  MUX2_X1 _19143_ (
    .A(ex_reg_inst[7]),
    .B(_02613_),
    .S(_02567_),
    .Z(_02614_)
  );
  OR2_X1 _19144_ (
    .A1(_02612_),
    .A2(_02614_),
    .ZN(_02615_)
  );
  OR2_X1 _19145_ (
    .A1(ex_reg_inst[20]),
    .A2(_02611_),
    .ZN(_02616_)
  );
  AND2_X1 _19146_ (
    .A1(_02591_),
    .A2(_02616_),
    .ZN(_02617_)
  );
  AND2_X1 _19147_ (
    .A1(_02615_),
    .A2(_02617_),
    .ZN(_02618_)
  );
  OR2_X1 _19148_ (
    .A1(_02610_),
    .A2(_02618_),
    .ZN(_02619_)
  );
  AND2_X1 _19149_ (
    .A1(_02543_),
    .A2(_02619_),
    .ZN(alu_io_in2[11])
  );
  AND2_X1 _19150_ (
    .A1(_02565_),
    .A2(_02611_),
    .ZN(_02620_)
  );
  MUX2_X1 _19151_ (
    .A(ex_reg_inst[12]),
    .B(_02613_),
    .S(_02620_),
    .Z(_02621_)
  );
  AND2_X1 _19152_ (
    .A1(_02548_),
    .A2(_02621_),
    .ZN(_02622_)
  );
  AND2_X1 _19153_ (
    .A1(_ex_op2_T[12]),
    .A2(_02546_),
    .ZN(_02623_)
  );
  OR2_X1 _19154_ (
    .A1(_02622_),
    .A2(_02623_),
    .ZN(_02624_)
  );
  AND2_X1 _19155_ (
    .A1(_02543_),
    .A2(_02624_),
    .ZN(alu_io_in2[12])
  );
  MUX2_X1 _19156_ (
    .A(ex_reg_inst[13]),
    .B(_02613_),
    .S(_02620_),
    .Z(_02625_)
  );
  AND2_X1 _19157_ (
    .A1(_02548_),
    .A2(_02625_),
    .ZN(_02626_)
  );
  AND2_X1 _19158_ (
    .A1(_ex_op2_T[13]),
    .A2(_02546_),
    .ZN(_02627_)
  );
  OR2_X1 _19159_ (
    .A1(_02626_),
    .A2(_02627_),
    .ZN(_02628_)
  );
  AND2_X1 _19160_ (
    .A1(_02543_),
    .A2(_02628_),
    .ZN(alu_io_in2[13])
  );
  MUX2_X1 _19161_ (
    .A(ex_reg_inst[14]),
    .B(_02613_),
    .S(_02620_),
    .Z(_02629_)
  );
  AND2_X1 _19162_ (
    .A1(_02548_),
    .A2(_02629_),
    .ZN(_02630_)
  );
  AND2_X1 _19163_ (
    .A1(_ex_op2_T[14]),
    .A2(_02546_),
    .ZN(_02631_)
  );
  OR2_X1 _19164_ (
    .A1(_02630_),
    .A2(_02631_),
    .ZN(_02632_)
  );
  AND2_X1 _19165_ (
    .A1(_02543_),
    .A2(_02632_),
    .ZN(alu_io_in2[14])
  );
  MUX2_X1 _19166_ (
    .A(ex_reg_inst[15]),
    .B(_02613_),
    .S(_02620_),
    .Z(_02633_)
  );
  AND2_X1 _19167_ (
    .A1(_02548_),
    .A2(_02633_),
    .ZN(_02634_)
  );
  AND2_X1 _19168_ (
    .A1(_ex_op2_T[15]),
    .A2(_02546_),
    .ZN(_02635_)
  );
  OR2_X1 _19169_ (
    .A1(_02634_),
    .A2(_02635_),
    .ZN(_02636_)
  );
  AND2_X1 _19170_ (
    .A1(_02543_),
    .A2(_02636_),
    .ZN(alu_io_in2[15])
  );
  MUX2_X1 _19171_ (
    .A(ex_reg_inst[16]),
    .B(_02613_),
    .S(_02620_),
    .Z(_02637_)
  );
  AND2_X1 _19172_ (
    .A1(_02548_),
    .A2(_02637_),
    .ZN(_02638_)
  );
  AND2_X1 _19173_ (
    .A1(_ex_op2_T[16]),
    .A2(_02546_),
    .ZN(_02639_)
  );
  OR2_X1 _19174_ (
    .A1(_02638_),
    .A2(_02639_),
    .ZN(_02640_)
  );
  AND2_X1 _19175_ (
    .A1(_02543_),
    .A2(_02640_),
    .ZN(alu_io_in2[16])
  );
  MUX2_X1 _19176_ (
    .A(ex_reg_inst[17]),
    .B(_02613_),
    .S(_02620_),
    .Z(_02641_)
  );
  AND2_X1 _19177_ (
    .A1(_02548_),
    .A2(_02641_),
    .ZN(_02642_)
  );
  AND2_X1 _19178_ (
    .A1(_ex_op2_T[17]),
    .A2(_02546_),
    .ZN(_02643_)
  );
  OR2_X1 _19179_ (
    .A1(_02642_),
    .A2(_02643_),
    .ZN(_02644_)
  );
  AND2_X1 _19180_ (
    .A1(_02543_),
    .A2(_02644_),
    .ZN(alu_io_in2[17])
  );
  MUX2_X1 _19181_ (
    .A(ex_reg_inst[18]),
    .B(_02613_),
    .S(_02620_),
    .Z(_02645_)
  );
  AND2_X1 _19182_ (
    .A1(_02548_),
    .A2(_02645_),
    .ZN(_02646_)
  );
  AND2_X1 _19183_ (
    .A1(_ex_op2_T[18]),
    .A2(_02546_),
    .ZN(_02647_)
  );
  OR2_X1 _19184_ (
    .A1(_02646_),
    .A2(_02647_),
    .ZN(_02648_)
  );
  AND2_X1 _19185_ (
    .A1(_02543_),
    .A2(_02648_),
    .ZN(alu_io_in2[18])
  );
  MUX2_X1 _19186_ (
    .A(ex_reg_inst[19]),
    .B(_02613_),
    .S(_02620_),
    .Z(_02649_)
  );
  AND2_X1 _19187_ (
    .A1(_02548_),
    .A2(_02649_),
    .ZN(_02650_)
  );
  AND2_X1 _19188_ (
    .A1(_ex_op2_T[19]),
    .A2(_02546_),
    .ZN(_02651_)
  );
  OR2_X1 _19189_ (
    .A1(_02650_),
    .A2(_02651_),
    .ZN(_02652_)
  );
  AND2_X1 _19190_ (
    .A1(_02543_),
    .A2(_02652_),
    .ZN(alu_io_in2[19])
  );
  MUX2_X1 _19191_ (
    .A(ex_reg_inst[20]),
    .B(_02613_),
    .S(_02565_),
    .Z(_02653_)
  );
  AND2_X1 _19192_ (
    .A1(_02548_),
    .A2(_02653_),
    .ZN(_02654_)
  );
  AND2_X1 _19193_ (
    .A1(_ex_op2_T[20]),
    .A2(_02546_),
    .ZN(_02655_)
  );
  OR2_X1 _19194_ (
    .A1(_02654_),
    .A2(_02655_),
    .ZN(_02656_)
  );
  AND2_X1 _19195_ (
    .A1(_02543_),
    .A2(_02656_),
    .ZN(alu_io_in2[20])
  );
  MUX2_X1 _19196_ (
    .A(ex_reg_inst[21]),
    .B(_02613_),
    .S(_02565_),
    .Z(_02657_)
  );
  AND2_X1 _19197_ (
    .A1(_02548_),
    .A2(_02657_),
    .ZN(_02658_)
  );
  AND2_X1 _19198_ (
    .A1(_ex_op2_T[21]),
    .A2(_02546_),
    .ZN(_02659_)
  );
  OR2_X1 _19199_ (
    .A1(_02658_),
    .A2(_02659_),
    .ZN(_02660_)
  );
  AND2_X1 _19200_ (
    .A1(_02543_),
    .A2(_02660_),
    .ZN(alu_io_in2[21])
  );
  MUX2_X1 _19201_ (
    .A(ex_reg_inst[22]),
    .B(_02613_),
    .S(_02565_),
    .Z(_02661_)
  );
  AND2_X1 _19202_ (
    .A1(_02548_),
    .A2(_02661_),
    .ZN(_02662_)
  );
  AND2_X1 _19203_ (
    .A1(_ex_op2_T[22]),
    .A2(_02546_),
    .ZN(_02663_)
  );
  OR2_X1 _19204_ (
    .A1(_02662_),
    .A2(_02663_),
    .ZN(_02664_)
  );
  AND2_X1 _19205_ (
    .A1(_02543_),
    .A2(_02664_),
    .ZN(alu_io_in2[22])
  );
  MUX2_X1 _19206_ (
    .A(ex_reg_inst[23]),
    .B(_02613_),
    .S(_02565_),
    .Z(_02665_)
  );
  AND2_X1 _19207_ (
    .A1(_02548_),
    .A2(_02665_),
    .ZN(_02666_)
  );
  AND2_X1 _19208_ (
    .A1(_ex_op2_T[23]),
    .A2(_02546_),
    .ZN(_02667_)
  );
  OR2_X1 _19209_ (
    .A1(_02666_),
    .A2(_02667_),
    .ZN(_02668_)
  );
  AND2_X1 _19210_ (
    .A1(_02543_),
    .A2(_02668_),
    .ZN(alu_io_in2[23])
  );
  MUX2_X1 _19211_ (
    .A(ex_reg_inst[24]),
    .B(_02613_),
    .S(_02565_),
    .Z(_02669_)
  );
  AND2_X1 _19212_ (
    .A1(_02548_),
    .A2(_02669_),
    .ZN(_02670_)
  );
  AND2_X1 _19213_ (
    .A1(_ex_op2_T[24]),
    .A2(_02546_),
    .ZN(_02671_)
  );
  OR2_X1 _19214_ (
    .A1(_02670_),
    .A2(_02671_),
    .ZN(_02672_)
  );
  AND2_X1 _19215_ (
    .A1(_02543_),
    .A2(_02672_),
    .ZN(alu_io_in2[24])
  );
  MUX2_X1 _19216_ (
    .A(ex_reg_inst[25]),
    .B(_02613_),
    .S(_02565_),
    .Z(_02673_)
  );
  AND2_X1 _19217_ (
    .A1(_02548_),
    .A2(_02673_),
    .ZN(_02674_)
  );
  AND2_X1 _19218_ (
    .A1(_ex_op2_T[25]),
    .A2(_02546_),
    .ZN(_02675_)
  );
  OR2_X1 _19219_ (
    .A1(_02674_),
    .A2(_02675_),
    .ZN(_02676_)
  );
  AND2_X1 _19220_ (
    .A1(_02543_),
    .A2(_02676_),
    .ZN(alu_io_in2[25])
  );
  MUX2_X1 _19221_ (
    .A(ex_reg_inst[26]),
    .B(_02613_),
    .S(_02565_),
    .Z(_02677_)
  );
  AND2_X1 _19222_ (
    .A1(_02548_),
    .A2(_02677_),
    .ZN(_02678_)
  );
  AND2_X1 _19223_ (
    .A1(_ex_op2_T[26]),
    .A2(_02546_),
    .ZN(_02679_)
  );
  OR2_X1 _19224_ (
    .A1(_02678_),
    .A2(_02679_),
    .ZN(_02680_)
  );
  AND2_X1 _19225_ (
    .A1(_02543_),
    .A2(_02680_),
    .ZN(alu_io_in2[26])
  );
  MUX2_X1 _19226_ (
    .A(ex_reg_inst[27]),
    .B(_02613_),
    .S(_02565_),
    .Z(_02681_)
  );
  AND2_X1 _19227_ (
    .A1(_02548_),
    .A2(_02681_),
    .ZN(_02682_)
  );
  AND2_X1 _19228_ (
    .A1(_ex_op2_T[27]),
    .A2(_02546_),
    .ZN(_02683_)
  );
  OR2_X1 _19229_ (
    .A1(_02682_),
    .A2(_02683_),
    .ZN(_02684_)
  );
  AND2_X1 _19230_ (
    .A1(_02543_),
    .A2(_02684_),
    .ZN(alu_io_in2[27])
  );
  MUX2_X1 _19231_ (
    .A(ex_reg_inst[28]),
    .B(_02613_),
    .S(_02565_),
    .Z(_02685_)
  );
  AND2_X1 _19232_ (
    .A1(_02548_),
    .A2(_02685_),
    .ZN(_02686_)
  );
  AND2_X1 _19233_ (
    .A1(_ex_op2_T[28]),
    .A2(_02546_),
    .ZN(_02687_)
  );
  OR2_X1 _19234_ (
    .A1(_02686_),
    .A2(_02687_),
    .ZN(_02688_)
  );
  AND2_X1 _19235_ (
    .A1(_02543_),
    .A2(_02688_),
    .ZN(alu_io_in2[28])
  );
  MUX2_X1 _19236_ (
    .A(ex_reg_inst[29]),
    .B(_02613_),
    .S(_02565_),
    .Z(_02689_)
  );
  AND2_X1 _19237_ (
    .A1(_02548_),
    .A2(_02689_),
    .ZN(_02690_)
  );
  AND2_X1 _19238_ (
    .A1(_ex_op2_T[29]),
    .A2(_02546_),
    .ZN(_02691_)
  );
  OR2_X1 _19239_ (
    .A1(_02690_),
    .A2(_02691_),
    .ZN(_02692_)
  );
  AND2_X1 _19240_ (
    .A1(_02543_),
    .A2(_02692_),
    .ZN(alu_io_in2[29])
  );
  MUX2_X1 _19241_ (
    .A(ex_reg_inst[30]),
    .B(_02613_),
    .S(_02565_),
    .Z(_02693_)
  );
  AND2_X1 _19242_ (
    .A1(_02548_),
    .A2(_02693_),
    .ZN(_02694_)
  );
  AND2_X1 _19243_ (
    .A1(_ex_op2_T[30]),
    .A2(_02546_),
    .ZN(_02695_)
  );
  OR2_X1 _19244_ (
    .A1(_02694_),
    .A2(_02695_),
    .ZN(_02696_)
  );
  AND2_X1 _19245_ (
    .A1(_02543_),
    .A2(_02696_),
    .ZN(alu_io_in2[30])
  );
  AND2_X1 _19246_ (
    .A1(_02548_),
    .A2(_02613_),
    .ZN(_02697_)
  );
  AND2_X1 _19247_ (
    .A1(_ex_op2_T[31]),
    .A2(_02546_),
    .ZN(_02698_)
  );
  OR2_X1 _19248_ (
    .A1(_02697_),
    .A2(_02698_),
    .ZN(_02699_)
  );
  AND2_X1 _19249_ (
    .A1(_02543_),
    .A2(_02699_),
    .ZN(alu_io_in2[31])
  );
  AND2_X1 _19250_ (
    .A1(_03033_),
    .A2(_03059_),
    .ZN(_02700_)
  );
  INV_X1 _19251_ (
    .A(_02700_),
    .ZN(_02701_)
  );
  AND2_X1 _19252_ (
    .A1(ex_reg_pc[0]),
    .A2(_02700_),
    .ZN(_02702_)
  );
  OR2_X1 _19253_ (
    .A1(ex_ctrl_sel_alu1[1]),
    .A2(_00020_),
    .ZN(_02703_)
  );
  INV_X1 _19254_ (
    .A(_02703_),
    .ZN(_02704_)
  );
  AND2_X1 _19255_ (
    .A1(_02701_),
    .A2(_02704_),
    .ZN(_02705_)
  );
  AND2_X1 _19256_ (
    .A1(_ex_op1_T[0]),
    .A2(_02705_),
    .ZN(_02706_)
  );
  OR2_X1 _19257_ (
    .A1(_02702_),
    .A2(_02706_),
    .ZN(alu_io_in1[0])
  );
  AND2_X1 _19258_ (
    .A1(ex_reg_pc[1]),
    .A2(_02700_),
    .ZN(_02707_)
  );
  AND2_X1 _19259_ (
    .A1(_ex_op1_T[1]),
    .A2(_02705_),
    .ZN(_02708_)
  );
  OR2_X1 _19260_ (
    .A1(_02707_),
    .A2(_02708_),
    .ZN(alu_io_in1[1])
  );
  AND2_X1 _19261_ (
    .A1(ex_reg_pc[2]),
    .A2(_02700_),
    .ZN(_02709_)
  );
  AND2_X1 _19262_ (
    .A1(_ex_op1_T[2]),
    .A2(_02705_),
    .ZN(_02710_)
  );
  OR2_X1 _19263_ (
    .A1(_02709_),
    .A2(_02710_),
    .ZN(alu_io_in1[2])
  );
  AND2_X1 _19264_ (
    .A1(ex_reg_pc[3]),
    .A2(_02700_),
    .ZN(_02711_)
  );
  AND2_X1 _19265_ (
    .A1(_ex_op1_T[3]),
    .A2(_02705_),
    .ZN(_02712_)
  );
  OR2_X1 _19266_ (
    .A1(_02711_),
    .A2(_02712_),
    .ZN(alu_io_in1[3])
  );
  AND2_X1 _19267_ (
    .A1(ex_reg_pc[4]),
    .A2(_02700_),
    .ZN(_02713_)
  );
  AND2_X1 _19268_ (
    .A1(_ex_op1_T[4]),
    .A2(_02705_),
    .ZN(_02714_)
  );
  OR2_X1 _19269_ (
    .A1(_02713_),
    .A2(_02714_),
    .ZN(alu_io_in1[4])
  );
  AND2_X1 _19270_ (
    .A1(ex_reg_pc[5]),
    .A2(_02700_),
    .ZN(_02715_)
  );
  AND2_X1 _19271_ (
    .A1(_ex_op1_T[5]),
    .A2(_02705_),
    .ZN(_02716_)
  );
  OR2_X1 _19272_ (
    .A1(_02715_),
    .A2(_02716_),
    .ZN(alu_io_in1[5])
  );
  AND2_X1 _19273_ (
    .A1(ex_reg_pc[6]),
    .A2(_02700_),
    .ZN(_02717_)
  );
  AND2_X1 _19274_ (
    .A1(_ex_op1_T[6]),
    .A2(_02705_),
    .ZN(_02718_)
  );
  OR2_X1 _19275_ (
    .A1(_02717_),
    .A2(_02718_),
    .ZN(alu_io_in1[6])
  );
  AND2_X1 _19276_ (
    .A1(ex_reg_pc[7]),
    .A2(_02700_),
    .ZN(_02719_)
  );
  AND2_X1 _19277_ (
    .A1(_ex_op1_T[7]),
    .A2(_02705_),
    .ZN(_02720_)
  );
  OR2_X1 _19278_ (
    .A1(_02719_),
    .A2(_02720_),
    .ZN(alu_io_in1[7])
  );
  AND2_X1 _19279_ (
    .A1(ex_reg_pc[8]),
    .A2(_02700_),
    .ZN(_02721_)
  );
  AND2_X1 _19280_ (
    .A1(_ex_op1_T[8]),
    .A2(_02705_),
    .ZN(_02722_)
  );
  OR2_X1 _19281_ (
    .A1(_02721_),
    .A2(_02722_),
    .ZN(alu_io_in1[8])
  );
  AND2_X1 _19282_ (
    .A1(ex_reg_pc[9]),
    .A2(_02700_),
    .ZN(_02723_)
  );
  AND2_X1 _19283_ (
    .A1(_ex_op1_T[9]),
    .A2(_02705_),
    .ZN(_02724_)
  );
  OR2_X1 _19284_ (
    .A1(_02723_),
    .A2(_02724_),
    .ZN(alu_io_in1[9])
  );
  AND2_X1 _19285_ (
    .A1(ex_reg_pc[10]),
    .A2(_02700_),
    .ZN(_02725_)
  );
  AND2_X1 _19286_ (
    .A1(_ex_op1_T[10]),
    .A2(_02705_),
    .ZN(_02726_)
  );
  OR2_X1 _19287_ (
    .A1(_02725_),
    .A2(_02726_),
    .ZN(alu_io_in1[10])
  );
  AND2_X1 _19288_ (
    .A1(ex_reg_pc[11]),
    .A2(_02700_),
    .ZN(_02727_)
  );
  AND2_X1 _19289_ (
    .A1(_ex_op1_T[11]),
    .A2(_02705_),
    .ZN(_02728_)
  );
  OR2_X1 _19290_ (
    .A1(_02727_),
    .A2(_02728_),
    .ZN(alu_io_in1[11])
  );
  AND2_X1 _19291_ (
    .A1(ex_reg_pc[12]),
    .A2(_02700_),
    .ZN(_02729_)
  );
  AND2_X1 _19292_ (
    .A1(_ex_op1_T[12]),
    .A2(_02705_),
    .ZN(_02730_)
  );
  OR2_X1 _19293_ (
    .A1(_02729_),
    .A2(_02730_),
    .ZN(alu_io_in1[12])
  );
  AND2_X1 _19294_ (
    .A1(ex_reg_pc[13]),
    .A2(_02700_),
    .ZN(_02731_)
  );
  AND2_X1 _19295_ (
    .A1(_ex_op1_T[13]),
    .A2(_02705_),
    .ZN(_02732_)
  );
  OR2_X1 _19296_ (
    .A1(_02731_),
    .A2(_02732_),
    .ZN(alu_io_in1[13])
  );
  AND2_X1 _19297_ (
    .A1(ex_reg_pc[14]),
    .A2(_02700_),
    .ZN(_02733_)
  );
  AND2_X1 _19298_ (
    .A1(_ex_op1_T[14]),
    .A2(_02705_),
    .ZN(_02734_)
  );
  OR2_X1 _19299_ (
    .A1(_02733_),
    .A2(_02734_),
    .ZN(alu_io_in1[14])
  );
  AND2_X1 _19300_ (
    .A1(ex_reg_pc[15]),
    .A2(_02700_),
    .ZN(_02735_)
  );
  AND2_X1 _19301_ (
    .A1(_ex_op1_T[15]),
    .A2(_02705_),
    .ZN(_02736_)
  );
  OR2_X1 _19302_ (
    .A1(_02735_),
    .A2(_02736_),
    .ZN(alu_io_in1[15])
  );
  AND2_X1 _19303_ (
    .A1(ex_reg_pc[16]),
    .A2(_02700_),
    .ZN(_02737_)
  );
  AND2_X1 _19304_ (
    .A1(_ex_op1_T[16]),
    .A2(_02705_),
    .ZN(_02738_)
  );
  OR2_X1 _19305_ (
    .A1(_02737_),
    .A2(_02738_),
    .ZN(alu_io_in1[16])
  );
  AND2_X1 _19306_ (
    .A1(ex_reg_pc[17]),
    .A2(_02700_),
    .ZN(_02739_)
  );
  AND2_X1 _19307_ (
    .A1(_ex_op1_T[17]),
    .A2(_02705_),
    .ZN(_02740_)
  );
  OR2_X1 _19308_ (
    .A1(_02739_),
    .A2(_02740_),
    .ZN(alu_io_in1[17])
  );
  AND2_X1 _19309_ (
    .A1(ex_reg_pc[18]),
    .A2(_02700_),
    .ZN(_02741_)
  );
  AND2_X1 _19310_ (
    .A1(_ex_op1_T[18]),
    .A2(_02705_),
    .ZN(_02742_)
  );
  OR2_X1 _19311_ (
    .A1(_02741_),
    .A2(_02742_),
    .ZN(alu_io_in1[18])
  );
  AND2_X1 _19312_ (
    .A1(ex_reg_pc[19]),
    .A2(_02700_),
    .ZN(_02743_)
  );
  AND2_X1 _19313_ (
    .A1(_ex_op1_T[19]),
    .A2(_02705_),
    .ZN(_02744_)
  );
  OR2_X1 _19314_ (
    .A1(_02743_),
    .A2(_02744_),
    .ZN(alu_io_in1[19])
  );
  AND2_X1 _19315_ (
    .A1(ex_reg_pc[20]),
    .A2(_02700_),
    .ZN(_02745_)
  );
  AND2_X1 _19316_ (
    .A1(_ex_op1_T[20]),
    .A2(_02705_),
    .ZN(_02746_)
  );
  OR2_X1 _19317_ (
    .A1(_02745_),
    .A2(_02746_),
    .ZN(alu_io_in1[20])
  );
  AND2_X1 _19318_ (
    .A1(ex_reg_pc[21]),
    .A2(_02700_),
    .ZN(_02747_)
  );
  AND2_X1 _19319_ (
    .A1(_ex_op1_T[21]),
    .A2(_02705_),
    .ZN(_02748_)
  );
  OR2_X1 _19320_ (
    .A1(_02747_),
    .A2(_02748_),
    .ZN(alu_io_in1[21])
  );
  AND2_X1 _19321_ (
    .A1(ex_reg_pc[22]),
    .A2(_02700_),
    .ZN(_02749_)
  );
  AND2_X1 _19322_ (
    .A1(_ex_op1_T[22]),
    .A2(_02705_),
    .ZN(_02750_)
  );
  OR2_X1 _19323_ (
    .A1(_02749_),
    .A2(_02750_),
    .ZN(alu_io_in1[22])
  );
  AND2_X1 _19324_ (
    .A1(ex_reg_pc[23]),
    .A2(_02700_),
    .ZN(_02751_)
  );
  AND2_X1 _19325_ (
    .A1(_ex_op1_T[23]),
    .A2(_02705_),
    .ZN(_02752_)
  );
  OR2_X1 _19326_ (
    .A1(_02751_),
    .A2(_02752_),
    .ZN(alu_io_in1[23])
  );
  AND2_X1 _19327_ (
    .A1(ex_reg_pc[24]),
    .A2(_02700_),
    .ZN(_02753_)
  );
  AND2_X1 _19328_ (
    .A1(_ex_op1_T[24]),
    .A2(_02705_),
    .ZN(_02754_)
  );
  OR2_X1 _19329_ (
    .A1(_02753_),
    .A2(_02754_),
    .ZN(alu_io_in1[24])
  );
  AND2_X1 _19330_ (
    .A1(ex_reg_pc[25]),
    .A2(_02700_),
    .ZN(_02755_)
  );
  AND2_X1 _19331_ (
    .A1(_ex_op1_T[25]),
    .A2(_02705_),
    .ZN(_02756_)
  );
  OR2_X1 _19332_ (
    .A1(_02755_),
    .A2(_02756_),
    .ZN(alu_io_in1[25])
  );
  AND2_X1 _19333_ (
    .A1(ex_reg_pc[26]),
    .A2(_02700_),
    .ZN(_02757_)
  );
  AND2_X1 _19334_ (
    .A1(_ex_op1_T[26]),
    .A2(_02705_),
    .ZN(_02758_)
  );
  OR2_X1 _19335_ (
    .A1(_02757_),
    .A2(_02758_),
    .ZN(alu_io_in1[26])
  );
  AND2_X1 _19336_ (
    .A1(ex_reg_pc[27]),
    .A2(_02700_),
    .ZN(_02759_)
  );
  AND2_X1 _19337_ (
    .A1(_ex_op1_T[27]),
    .A2(_02705_),
    .ZN(_02760_)
  );
  OR2_X1 _19338_ (
    .A1(_02759_),
    .A2(_02760_),
    .ZN(alu_io_in1[27])
  );
  AND2_X1 _19339_ (
    .A1(ex_reg_pc[28]),
    .A2(_02700_),
    .ZN(_02761_)
  );
  AND2_X1 _19340_ (
    .A1(_ex_op1_T[28]),
    .A2(_02705_),
    .ZN(_02762_)
  );
  OR2_X1 _19341_ (
    .A1(_02761_),
    .A2(_02762_),
    .ZN(alu_io_in1[28])
  );
  AND2_X1 _19342_ (
    .A1(ex_reg_pc[29]),
    .A2(_02700_),
    .ZN(_02763_)
  );
  AND2_X1 _19343_ (
    .A1(_ex_op1_T[29]),
    .A2(_02705_),
    .ZN(_02764_)
  );
  OR2_X1 _19344_ (
    .A1(_02763_),
    .A2(_02764_),
    .ZN(alu_io_in1[29])
  );
  AND2_X1 _19345_ (
    .A1(ex_reg_pc[30]),
    .A2(_02700_),
    .ZN(_02765_)
  );
  AND2_X1 _19346_ (
    .A1(_ex_op1_T[30]),
    .A2(_02705_),
    .ZN(_02766_)
  );
  OR2_X1 _19347_ (
    .A1(_02765_),
    .A2(_02766_),
    .ZN(alu_io_in1[30])
  );
  AND2_X1 _19348_ (
    .A1(ex_reg_pc[31]),
    .A2(_02700_),
    .ZN(_02767_)
  );
  AND2_X1 _19349_ (
    .A1(_ex_op1_T[31]),
    .A2(_02705_),
    .ZN(_02768_)
  );
  OR2_X1 _19350_ (
    .A1(_02767_),
    .A2(_02768_),
    .ZN(alu_io_in1[31])
  );
  AND2_X1 _19351_ (
    .A1(_03099_),
    .A2(_03113_),
    .ZN(div_io_resp_ready)
  );
  AND2_X1 _19352_ (
    .A1(ex_reg_load_use),
    .A2(_03125_),
    .ZN(_02769_)
  );
  AND2_X1 _19353_ (
    .A1(ex_ctrl_mem),
    .A2(_03085_),
    .ZN(_02770_)
  );
  AND2_X1 _19354_ (
    .A1(ex_ctrl_div),
    .A2(_03084_),
    .ZN(_02771_)
  );
  OR2_X1 _19355_ (
    .A1(_02770_),
    .A2(_02771_),
    .ZN(_02772_)
  );
  OR2_X1 _19356_ (
    .A1(_02769_),
    .A2(_02772_),
    .ZN(_02773_)
  );
  AND2_X1 _19357_ (
    .A1(ex_reg_valid),
    .A2(_02773_),
    .ZN(_02774_)
  );
  OR2_X1 _19358_ (
    .A1(ex_reg_replay),
    .A2(_02774_),
    .ZN(_02775_)
  );
  OR2_X1 _19359_ (
    .A1(_00034_),
    .A2(_02775_),
    .ZN(_02776_)
  );
  INV_X1 _19360_ (
    .A(_02776_),
    .ZN(_02777_)
  );
  AND2_X1 _19361_ (
    .A1(_04036_),
    .A2(_02777_),
    .ZN(_mem_reg_valid_T)
  );
  AND2_X1 _19362_ (
    .A1(io_dmem_replay_next),
    .A2(_03471_),
    .ZN(_02778_)
  );
  OR2_X1 _19363_ (
    .A1(mem_reg_xcpt),
    .A2(_00033_),
    .ZN(_02779_)
  );
  OR2_X1 _19364_ (
    .A1(_02778_),
    .A2(_02779_),
    .ZN(_02780_)
  );
  OR2_X1 _19365_ (
    .A1(_04029_),
    .A2(_02780_),
    .ZN(_02781_)
  );
  INV_X1 _19366_ (
    .A(_02781_),
    .ZN(_02782_)
  );
  AND2_X1 _19367_ (
    .A1(mem_reg_load),
    .A2(bpu_io_xcpt_ld),
    .ZN(_02783_)
  );
  AND2_X1 _19368_ (
    .A1(mem_reg_store),
    .A2(bpu_io_xcpt_st),
    .ZN(_02784_)
  );
  OR2_X1 _19369_ (
    .A1(_02783_),
    .A2(_02784_),
    .ZN(_02785_)
  );
  OR2_X1 _19370_ (
    .A1(_02052_),
    .A2(_02785_),
    .ZN(_02786_)
  );
  AND2_X1 _19371_ (
    .A1(mem_reg_valid),
    .A2(_02786_),
    .ZN(_02787_)
  );
  INV_X1 _19372_ (
    .A(_02787_),
    .ZN(_02788_)
  );
  AND2_X1 _19373_ (
    .A1(_02056_),
    .A2(_02788_),
    .ZN(_02789_)
  );
  OR2_X1 _19374_ (
    .A1(_02057_),
    .A2(_02787_),
    .ZN(_02790_)
  );
  AND2_X1 _19375_ (
    .A1(_02782_),
    .A2(_02789_),
    .ZN(_wb_reg_valid_T)
  );
  AND2_X1 _19376_ (
    .A1(mem_reg_valid),
    .A2(io_imem_req_bits_speculative),
    .ZN(io_imem_bht_update_valid)
  );
  XOR2_X1 _19377_ (
    .A(bpu_io_pc[29]),
    .B(_02476_),
    .Z(_02791_)
  );
  XOR2_X1 _19378_ (
    .A(bpu_io_pc[27]),
    .B(_02463_),
    .Z(_02792_)
  );
  XOR2_X1 _19379_ (
    .A(bpu_io_pc[26]),
    .B(_02457_),
    .Z(_02793_)
  );
  XOR2_X1 _19380_ (
    .A(bpu_io_pc[24]),
    .B(_02445_),
    .Z(_02794_)
  );
  XOR2_X1 _19381_ (
    .A(bpu_io_pc[22]),
    .B(_02433_),
    .Z(_02795_)
  );
  AND2_X1 _19382_ (
    .A1(bpu_io_pc[17]),
    .A2(_02403_),
    .ZN(_02796_)
  );
  AND2_X1 _19383_ (
    .A1(_03023_),
    .A2(_02402_),
    .ZN(_02797_)
  );
  AND2_X1 _19384_ (
    .A1(_03022_),
    .A2(_02381_),
    .ZN(_02798_)
  );
  AND2_X1 _19385_ (
    .A1(bpu_io_pc[14]),
    .A2(_02382_),
    .ZN(_02799_)
  );
  AND2_X1 _19386_ (
    .A1(_03021_),
    .A2(_02374_),
    .ZN(_02800_)
  );
  AND2_X1 _19387_ (
    .A1(bpu_io_pc[13]),
    .A2(_02375_),
    .ZN(_02801_)
  );
  AND2_X1 _19388_ (
    .A1(bpu_io_pc[12]),
    .A2(_02368_),
    .ZN(_02802_)
  );
  AND2_X1 _19389_ (
    .A1(_03020_),
    .A2(_02367_),
    .ZN(_02803_)
  );
  AND2_X1 _19390_ (
    .A1(_03019_),
    .A2(_02360_),
    .ZN(_02804_)
  );
  AND2_X1 _19391_ (
    .A1(bpu_io_pc[11]),
    .A2(_02361_),
    .ZN(_02805_)
  );
  AND2_X1 _19392_ (
    .A1(_03018_),
    .A2(_02353_),
    .ZN(_02806_)
  );
  AND2_X1 _19393_ (
    .A1(bpu_io_pc[10]),
    .A2(_02354_),
    .ZN(_02807_)
  );
  AND2_X1 _19394_ (
    .A1(_03017_),
    .A2(_02346_),
    .ZN(_02808_)
  );
  AND2_X1 _19395_ (
    .A1(bpu_io_pc[9]),
    .A2(_02347_),
    .ZN(_02809_)
  );
  AND2_X1 _19396_ (
    .A1(_03016_),
    .A2(_02339_),
    .ZN(_02810_)
  );
  AND2_X1 _19397_ (
    .A1(bpu_io_pc[8]),
    .A2(_02340_),
    .ZN(_02811_)
  );
  AND2_X1 _19398_ (
    .A1(bpu_io_pc[7]),
    .A2(_02333_),
    .ZN(_02812_)
  );
  AND2_X1 _19399_ (
    .A1(_03015_),
    .A2(_02332_),
    .ZN(_02813_)
  );
  AND2_X1 _19400_ (
    .A1(bpu_io_pc[6]),
    .A2(_02326_),
    .ZN(_02814_)
  );
  AND2_X1 _19401_ (
    .A1(_03014_),
    .A2(_02325_),
    .ZN(_02815_)
  );
  AND2_X1 _19402_ (
    .A1(_03013_),
    .A2(_02318_),
    .ZN(_02816_)
  );
  AND2_X1 _19403_ (
    .A1(bpu_io_pc[5]),
    .A2(_02319_),
    .ZN(_02817_)
  );
  AND2_X1 _19404_ (
    .A1(_03012_),
    .A2(_02314_),
    .ZN(_02818_)
  );
  AND2_X1 _19405_ (
    .A1(bpu_io_pc[4]),
    .A2(_02315_),
    .ZN(_02819_)
  );
  AND2_X1 _19406_ (
    .A1(bpu_io_pc[3]),
    .A2(_02312_),
    .ZN(_02820_)
  );
  AND2_X1 _19407_ (
    .A1(_03011_),
    .A2(_02311_),
    .ZN(_02821_)
  );
  XOR2_X1 _19408_ (
    .A(bpu_io_pc[1]),
    .B(_06438_),
    .Z(_02822_)
  );
  OR2_X1 _19409_ (
    .A1(ibuf_io_inst_0_valid),
    .A2(io_imem_resp_valid),
    .ZN(_02823_)
  );
  INV_X1 _19410_ (
    .A(_02823_),
    .ZN(_02824_)
  );
  OR2_X1 _19411_ (
    .A1(bpu_io_pc[0]),
    .A2(_02824_),
    .ZN(_02825_)
  );
  OR2_X1 _19412_ (
    .A1(_08749_),
    .A2(_02825_),
    .ZN(_02826_)
  );
  OR2_X1 _19413_ (
    .A1(_02822_),
    .A2(_02826_),
    .ZN(_02827_)
  );
  XOR2_X1 _19414_ (
    .A(bpu_io_pc[23]),
    .B(_02439_),
    .Z(_02828_)
  );
  AND2_X1 _19415_ (
    .A1(_03024_),
    .A2(_02470_),
    .ZN(_02829_)
  );
  AND2_X1 _19416_ (
    .A1(bpu_io_pc[28]),
    .A2(_02469_),
    .ZN(_02830_)
  );
  OR2_X1 _19417_ (
    .A1(_03031_),
    .A2(_04032_),
    .ZN(_02831_)
  );
  AND2_X1 _19418_ (
    .A1(io_imem_bht_update_valid),
    .A2(_02831_),
    .ZN(_02832_)
  );
  XOR2_X1 _19419_ (
    .A(ex_reg_pc[31]),
    .B(_02488_),
    .Z(_02833_)
  );
  XOR2_X1 _19420_ (
    .A(ex_reg_pc[29]),
    .B(_02476_),
    .Z(_02834_)
  );
  XOR2_X1 _19421_ (
    .A(ex_reg_pc[27]),
    .B(_02463_),
    .Z(_02835_)
  );
  XOR2_X1 _19422_ (
    .A(ex_reg_pc[28]),
    .B(_02470_),
    .Z(_02836_)
  );
  XOR2_X1 _19423_ (
    .A(ex_reg_pc[26]),
    .B(_02457_),
    .Z(_02837_)
  );
  XOR2_X1 _19424_ (
    .A(ex_reg_pc[25]),
    .B(_02451_),
    .Z(_02838_)
  );
  XOR2_X1 _19425_ (
    .A(ex_reg_pc[23]),
    .B(_02439_),
    .Z(_02839_)
  );
  XOR2_X1 _19426_ (
    .A(ex_reg_pc[24]),
    .B(_02445_),
    .Z(_02840_)
  );
  XOR2_X1 _19427_ (
    .A(ex_reg_pc[22]),
    .B(_02433_),
    .Z(_02841_)
  );
  AND2_X1 _19428_ (
    .A1(ex_reg_pc[17]),
    .A2(_02403_),
    .ZN(_02842_)
  );
  AND2_X1 _19429_ (
    .A1(_02999_),
    .A2(_02402_),
    .ZN(_02843_)
  );
  AND2_X1 _19430_ (
    .A1(_02998_),
    .A2(_02395_),
    .ZN(_02844_)
  );
  AND2_X1 _19431_ (
    .A1(ex_reg_pc[16]),
    .A2(_02396_),
    .ZN(_02845_)
  );
  AND2_X1 _19432_ (
    .A1(ex_reg_pc[15]),
    .A2(_02389_),
    .ZN(_02846_)
  );
  AND2_X1 _19433_ (
    .A1(_02997_),
    .A2(_02388_),
    .ZN(_02847_)
  );
  AND2_X1 _19434_ (
    .A1(_02996_),
    .A2(_02381_),
    .ZN(_02848_)
  );
  AND2_X1 _19435_ (
    .A1(ex_reg_pc[14]),
    .A2(_02382_),
    .ZN(_02849_)
  );
  AND2_X1 _19436_ (
    .A1(ex_reg_pc[13]),
    .A2(_02375_),
    .ZN(_02850_)
  );
  AND2_X1 _19437_ (
    .A1(_02995_),
    .A2(_02374_),
    .ZN(_02851_)
  );
  AND2_X1 _19438_ (
    .A1(_02994_),
    .A2(_02367_),
    .ZN(_02852_)
  );
  AND2_X1 _19439_ (
    .A1(ex_reg_pc[12]),
    .A2(_02368_),
    .ZN(_02853_)
  );
  AND2_X1 _19440_ (
    .A1(_02993_),
    .A2(_02360_),
    .ZN(_02854_)
  );
  AND2_X1 _19441_ (
    .A1(ex_reg_pc[11]),
    .A2(_02361_),
    .ZN(_02855_)
  );
  AND2_X1 _19442_ (
    .A1(_02992_),
    .A2(_02353_),
    .ZN(_02856_)
  );
  AND2_X1 _19443_ (
    .A1(ex_reg_pc[10]),
    .A2(_02354_),
    .ZN(_02857_)
  );
  XOR2_X1 _19444_ (
    .A(ex_reg_pc[6]),
    .B(_02325_),
    .Z(_02858_)
  );
  AND2_X1 _19445_ (
    .A1(ex_reg_pc[4]),
    .A2(_02315_),
    .ZN(_02859_)
  );
  AND2_X1 _19446_ (
    .A1(_02991_),
    .A2(_02314_),
    .ZN(_02860_)
  );
  OR2_X1 _19447_ (
    .A1(ex_reg_pc[0]),
    .A2(_08750_),
    .ZN(_02861_)
  );
  XOR2_X1 _19448_ (
    .A(ex_reg_pc[1]),
    .B(_06438_),
    .Z(_02862_)
  );
  OR2_X1 _19449_ (
    .A1(_02861_),
    .A2(_02862_),
    .ZN(_02863_)
  );
  XOR2_X1 _19450_ (
    .A(ex_reg_pc[2]),
    .B(_02309_),
    .Z(_02864_)
  );
  OR2_X1 _19451_ (
    .A1(_02863_),
    .A2(_02864_),
    .ZN(_02865_)
  );
  XOR2_X1 _19452_ (
    .A(ex_reg_pc[3]),
    .B(_02311_),
    .Z(_02866_)
  );
  OR2_X1 _19453_ (
    .A1(_02865_),
    .A2(_02866_),
    .ZN(_02867_)
  );
  OR2_X1 _19454_ (
    .A1(_02860_),
    .A2(_02867_),
    .ZN(_02868_)
  );
  OR2_X1 _19455_ (
    .A1(_02859_),
    .A2(_02868_),
    .ZN(_02869_)
  );
  XOR2_X1 _19456_ (
    .A(ex_reg_pc[5]),
    .B(_02318_),
    .Z(_02870_)
  );
  OR2_X1 _19457_ (
    .A1(_02869_),
    .A2(_02870_),
    .ZN(_02871_)
  );
  OR2_X1 _19458_ (
    .A1(_02858_),
    .A2(_02871_),
    .ZN(_02872_)
  );
  XOR2_X1 _19459_ (
    .A(bpu_io_pc[30]),
    .B(_02482_),
    .Z(_02873_)
  );
  XOR2_X1 _19460_ (
    .A(bpu_io_pc[25]),
    .B(_02451_),
    .Z(_02874_)
  );
  OR2_X1 _19461_ (
    .A1(_02793_),
    .A2(_02830_),
    .ZN(_02875_)
  );
  XOR2_X1 _19462_ (
    .A(bpu_io_pc[19]),
    .B(_02415_),
    .Z(_02876_)
  );
  XOR2_X1 _19463_ (
    .A(bpu_io_pc[18]),
    .B(_02409_),
    .Z(_02877_)
  );
  XOR2_X1 _19464_ (
    .A(bpu_io_pc[15]),
    .B(_02388_),
    .Z(_02878_)
  );
  OR2_X1 _19465_ (
    .A1(_02821_),
    .A2(_02827_),
    .ZN(_02879_)
  );
  OR2_X1 _19466_ (
    .A1(_02819_),
    .A2(_02879_),
    .ZN(_02880_)
  );
  OR2_X1 _19467_ (
    .A1(_02817_),
    .A2(_02880_),
    .ZN(_02881_)
  );
  OR2_X1 _19468_ (
    .A1(_02815_),
    .A2(_02881_),
    .ZN(_02882_)
  );
  OR2_X1 _19469_ (
    .A1(_02813_),
    .A2(_02882_),
    .ZN(_02883_)
  );
  OR2_X1 _19470_ (
    .A1(_02811_),
    .A2(_02883_),
    .ZN(_02884_)
  );
  OR2_X1 _19471_ (
    .A1(_02809_),
    .A2(_02884_),
    .ZN(_02885_)
  );
  OR2_X1 _19472_ (
    .A1(_02807_),
    .A2(_02885_),
    .ZN(_02886_)
  );
  OR2_X1 _19473_ (
    .A1(_02805_),
    .A2(_02886_),
    .ZN(_02887_)
  );
  OR2_X1 _19474_ (
    .A1(_02803_),
    .A2(_02887_),
    .ZN(_02888_)
  );
  OR2_X1 _19475_ (
    .A1(_02801_),
    .A2(_02888_),
    .ZN(_02889_)
  );
  OR2_X1 _19476_ (
    .A1(_02799_),
    .A2(_02889_),
    .ZN(_02890_)
  );
  XOR2_X1 _19477_ (
    .A(bpu_io_pc[2]),
    .B(_02309_),
    .Z(_02891_)
  );
  OR2_X1 _19478_ (
    .A1(_02820_),
    .A2(_02891_),
    .ZN(_02892_)
  );
  OR2_X1 _19479_ (
    .A1(_02818_),
    .A2(_02892_),
    .ZN(_02893_)
  );
  OR2_X1 _19480_ (
    .A1(_02816_),
    .A2(_02893_),
    .ZN(_02894_)
  );
  OR2_X1 _19481_ (
    .A1(_02814_),
    .A2(_02894_),
    .ZN(_02895_)
  );
  OR2_X1 _19482_ (
    .A1(_02812_),
    .A2(_02895_),
    .ZN(_02896_)
  );
  OR2_X1 _19483_ (
    .A1(_02810_),
    .A2(_02896_),
    .ZN(_02897_)
  );
  OR2_X1 _19484_ (
    .A1(_02808_),
    .A2(_02897_),
    .ZN(_02898_)
  );
  OR2_X1 _19485_ (
    .A1(_02806_),
    .A2(_02898_),
    .ZN(_02899_)
  );
  OR2_X1 _19486_ (
    .A1(_02804_),
    .A2(_02899_),
    .ZN(_02900_)
  );
  OR2_X1 _19487_ (
    .A1(_02802_),
    .A2(_02900_),
    .ZN(_02901_)
  );
  OR2_X1 _19488_ (
    .A1(_02800_),
    .A2(_02901_),
    .ZN(_02902_)
  );
  OR2_X1 _19489_ (
    .A1(_02798_),
    .A2(_02902_),
    .ZN(_02903_)
  );
  OR2_X1 _19490_ (
    .A1(_02890_),
    .A2(_02903_),
    .ZN(_02904_)
  );
  OR2_X1 _19491_ (
    .A1(_02878_),
    .A2(_02904_),
    .ZN(_02905_)
  );
  XOR2_X1 _19492_ (
    .A(bpu_io_pc[16]),
    .B(_02395_),
    .Z(_02906_)
  );
  OR2_X1 _19493_ (
    .A1(_02905_),
    .A2(_02906_),
    .ZN(_02907_)
  );
  OR2_X1 _19494_ (
    .A1(_02796_),
    .A2(_02907_),
    .ZN(_02908_)
  );
  OR2_X1 _19495_ (
    .A1(_02797_),
    .A2(_02908_),
    .ZN(_02909_)
  );
  OR2_X1 _19496_ (
    .A1(_02877_),
    .A2(_02909_),
    .ZN(_02910_)
  );
  OR2_X1 _19497_ (
    .A1(_02876_),
    .A2(_02910_),
    .ZN(_02911_)
  );
  XOR2_X1 _19498_ (
    .A(bpu_io_pc[20]),
    .B(_02421_),
    .Z(_02912_)
  );
  OR2_X1 _19499_ (
    .A1(_02911_),
    .A2(_02912_),
    .ZN(_02913_)
  );
  XOR2_X1 _19500_ (
    .A(bpu_io_pc[21]),
    .B(_02427_),
    .Z(_02914_)
  );
  OR2_X1 _19501_ (
    .A1(_02913_),
    .A2(_02914_),
    .ZN(_02915_)
  );
  OR2_X1 _19502_ (
    .A1(_02795_),
    .A2(_02915_),
    .ZN(_02916_)
  );
  OR2_X1 _19503_ (
    .A1(_02794_),
    .A2(_02916_),
    .ZN(_02917_)
  );
  OR2_X1 _19504_ (
    .A1(_02828_),
    .A2(_02917_),
    .ZN(_02918_)
  );
  OR2_X1 _19505_ (
    .A1(_02829_),
    .A2(_02918_),
    .ZN(_02919_)
  );
  OR2_X1 _19506_ (
    .A1(_02875_),
    .A2(_02919_),
    .ZN(_02920_)
  );
  OR2_X1 _19507_ (
    .A1(_02792_),
    .A2(_02920_),
    .ZN(_02921_)
  );
  OR2_X1 _19508_ (
    .A1(_02874_),
    .A2(_02921_),
    .ZN(_02922_)
  );
  OR2_X1 _19509_ (
    .A1(_02791_),
    .A2(_02922_),
    .ZN(_02923_)
  );
  OR2_X1 _19510_ (
    .A1(_02873_),
    .A2(_02923_),
    .ZN(_02924_)
  );
  XOR2_X1 _19511_ (
    .A(bpu_io_pc[31]),
    .B(_02488_),
    .Z(_02925_)
  );
  OR2_X1 _19512_ (
    .A1(_02924_),
    .A2(_02925_),
    .ZN(_02926_)
  );
  AND2_X1 _19513_ (
    .A1(_02832_),
    .A2(_02926_),
    .ZN(_02927_)
  );
  XOR2_X1 _19514_ (
    .A(ex_reg_pc[30]),
    .B(_02482_),
    .Z(_02928_)
  );
  XOR2_X1 _19515_ (
    .A(ex_reg_pc[19]),
    .B(_02415_),
    .Z(_02929_)
  );
  XOR2_X1 _19516_ (
    .A(ex_reg_pc[18]),
    .B(_02409_),
    .Z(_02930_)
  );
  XOR2_X1 _19517_ (
    .A(ex_reg_pc[7]),
    .B(_02332_),
    .Z(_02931_)
  );
  OR2_X1 _19518_ (
    .A1(_02872_),
    .A2(_02931_),
    .ZN(_02932_)
  );
  XOR2_X1 _19519_ (
    .A(ex_reg_pc[8]),
    .B(_02339_),
    .Z(_02933_)
  );
  OR2_X1 _19520_ (
    .A1(_02932_),
    .A2(_02933_),
    .ZN(_02934_)
  );
  OR2_X1 _19521_ (
    .A1(_02857_),
    .A2(_02934_),
    .ZN(_02935_)
  );
  OR2_X1 _19522_ (
    .A1(_02855_),
    .A2(_02935_),
    .ZN(_02936_)
  );
  OR2_X1 _19523_ (
    .A1(_02853_),
    .A2(_02936_),
    .ZN(_02937_)
  );
  OR2_X1 _19524_ (
    .A1(_02851_),
    .A2(_02937_),
    .ZN(_02938_)
  );
  OR2_X1 _19525_ (
    .A1(_02849_),
    .A2(_02938_),
    .ZN(_02939_)
  );
  OR2_X1 _19526_ (
    .A1(_02846_),
    .A2(_02939_),
    .ZN(_02940_)
  );
  OR2_X1 _19527_ (
    .A1(_02845_),
    .A2(_02940_),
    .ZN(_02941_)
  );
  OR2_X1 _19528_ (
    .A1(_02843_),
    .A2(_02941_),
    .ZN(_02942_)
  );
  XOR2_X1 _19529_ (
    .A(ex_reg_pc[9]),
    .B(_02346_),
    .Z(_02943_)
  );
  OR2_X1 _19530_ (
    .A1(_02856_),
    .A2(_02943_),
    .ZN(_02944_)
  );
  OR2_X1 _19531_ (
    .A1(_02854_),
    .A2(_02944_),
    .ZN(_02945_)
  );
  OR2_X1 _19532_ (
    .A1(_02852_),
    .A2(_02945_),
    .ZN(_02946_)
  );
  OR2_X1 _19533_ (
    .A1(_02850_),
    .A2(_02946_),
    .ZN(_02947_)
  );
  OR2_X1 _19534_ (
    .A1(_02848_),
    .A2(_02947_),
    .ZN(_02948_)
  );
  OR2_X1 _19535_ (
    .A1(_02847_),
    .A2(_02948_),
    .ZN(_02949_)
  );
  OR2_X1 _19536_ (
    .A1(_02844_),
    .A2(_02949_),
    .ZN(_02950_)
  );
  OR2_X1 _19537_ (
    .A1(_02842_),
    .A2(_02950_),
    .ZN(_02951_)
  );
  OR2_X1 _19538_ (
    .A1(_02942_),
    .A2(_02951_),
    .ZN(_02952_)
  );
  OR2_X1 _19539_ (
    .A1(_02930_),
    .A2(_02952_),
    .ZN(_02953_)
  );
  OR2_X1 _19540_ (
    .A1(_02929_),
    .A2(_02953_),
    .ZN(_02954_)
  );
  XOR2_X1 _19541_ (
    .A(ex_reg_pc[20]),
    .B(_02421_),
    .Z(_02955_)
  );
  OR2_X1 _19542_ (
    .A1(_02954_),
    .A2(_02955_),
    .ZN(_02956_)
  );
  XOR2_X1 _19543_ (
    .A(ex_reg_pc[21]),
    .B(_02427_),
    .Z(_02957_)
  );
  OR2_X1 _19544_ (
    .A1(_02956_),
    .A2(_02957_),
    .ZN(_02958_)
  );
  OR2_X1 _19545_ (
    .A1(_02841_),
    .A2(_02958_),
    .ZN(_02959_)
  );
  OR2_X1 _19546_ (
    .A1(_02840_),
    .A2(_02959_),
    .ZN(_02960_)
  );
  OR2_X1 _19547_ (
    .A1(_02839_),
    .A2(_02960_),
    .ZN(_02961_)
  );
  OR2_X1 _19548_ (
    .A1(_02838_),
    .A2(_02961_),
    .ZN(_02962_)
  );
  OR2_X1 _19549_ (
    .A1(_02837_),
    .A2(_02962_),
    .ZN(_02963_)
  );
  OR2_X1 _19550_ (
    .A1(_02836_),
    .A2(_02963_),
    .ZN(_02964_)
  );
  OR2_X1 _19551_ (
    .A1(_02835_),
    .A2(_02964_),
    .ZN(_02965_)
  );
  OR2_X1 _19552_ (
    .A1(_02834_),
    .A2(_02965_),
    .ZN(_02966_)
  );
  OR2_X1 _19553_ (
    .A1(_02928_),
    .A2(_02966_),
    .ZN(_02967_)
  );
  OR2_X1 _19554_ (
    .A1(_02833_),
    .A2(_02967_),
    .ZN(_02968_)
  );
  AND2_X1 _19555_ (
    .A1(_02927_),
    .A2(_02968_),
    .ZN(io_imem_btb_update_valid)
  );
  AND2_X1 _19556_ (
    .A1(wb_ctrl_fence_i),
    .A2(wb_reg_valid),
    .ZN(_02969_)
  );
  AND2_X1 _19557_ (
    .A1(_03086_),
    .A2(_02969_),
    .ZN(io_imem_flush_icache)
  );
  OR2_X1 _19558_ (
    .A1(_02781_),
    .A2(_02786_),
    .ZN(io_dmem_s1_kill)
  );
  AND2_X1 _19559_ (
    .A1(wb_ctrl_csr[2]),
    .A2(wb_reg_valid),
    .ZN(csr_io_rw_cmd[2])
  );
  AND2_X1 _19560_ (
    .A1(div_io_kill_REG),
    .A2(_02781_),
    .ZN(div_io_kill)
  );
  OR2_X1 _19561_ (
    .A1(_06433_),
    .A2(_08749_),
    .ZN(_02970_)
  );
  OR2_X1 _19562_ (
    .A1(io_ptw_customCSRs_csrs_0_value[1]),
    .A2(_02970_),
    .ZN(_00005_)
  );
  AND2_X1 _19563_ (
    .A1(csr_io_interrupt),
    .A2(_04037_),
    .ZN(_00004_)
  );
  OR2_X1 _19564_ (
    .A1(_04041_),
    .A2(_01790_),
    .ZN(_02971_)
  );
  INV_X1 _19565_ (
    .A(_02971_),
    .ZN(_00003_)
  );
  AND2_X1 _19566_ (
    .A1(ibuf_io_inst_0_bits_replay),
    .A2(_04037_),
    .ZN(_00002_)
  );
  AND2_X1 _19567_ (
    .A1(ex_reg_xcpt_interrupt),
    .A2(_04036_),
    .ZN(_00008_)
  );
  OR2_X1 _19568_ (
    .A1(ex_reg_xcpt_interrupt),
    .A2(ex_reg_xcpt),
    .ZN(_02972_)
  );
  AND2_X1 _19569_ (
    .A1(_mem_reg_valid_T),
    .A2(_02972_),
    .ZN(_00007_)
  );
  AND2_X1 _19570_ (
    .A1(_04036_),
    .A2(_02775_),
    .ZN(_00006_)
  );
  AND2_X1 _19571_ (
    .A1(io_imem_req_bits_speculative),
    .A2(_02790_),
    .ZN(_00011_)
  );
  OR2_X1 _19572_ (
    .A1(mem_reg_replay),
    .A2(_02778_),
    .ZN(_02973_)
  );
  AND2_X1 _19573_ (
    .A1(io_imem_req_bits_speculative),
    .A2(_02973_),
    .ZN(_00010_)
  );
  AND2_X1 _19574_ (
    .A1(mem_reg_flush_pipe),
    .A2(_wb_reg_valid_T),
    .ZN(_00009_)
  );
  OR2_X1 _19575_ (
    .A1(io_dmem_s2_nack),
    .A2(blocked),
    .ZN(_02974_)
  );
  OR2_X1 _19576_ (
    .A1(io_dmem_req_valid),
    .A2(_02974_),
    .ZN(_02975_)
  );
  OR2_X1 _19577_ (
    .A1(io_dmem_perf_grant),
    .A2(io_dmem_req_ready),
    .ZN(_02976_)
  );
  INV_X1 _19578_ (
    .A(_02976_),
    .ZN(_02977_)
  );
  AND2_X1 _19579_ (
    .A1(_02975_),
    .A2(_02977_),
    .ZN(_00000_)
  );
  AND2_X1 _19580_ (
    .A1(div_io_req_ready),
    .A2(div_io_req_valid),
    .ZN(_00001_)
  );
  DFF_X1 \_r[10]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00045_),
    .Q(_r[10]),
    .QN(_10421_)
  );
  DFF_X1 \_r[11]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00046_),
    .Q(_r[11]),
    .QN(_10420_)
  );
  DFF_X1 \_r[12]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00047_),
    .Q(_r[12]),
    .QN(_10419_)
  );
  DFF_X1 \_r[13]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00048_),
    .Q(_r[13]),
    .QN(_10418_)
  );
  DFF_X1 \_r[14]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00049_),
    .Q(_r[14]),
    .QN(_10417_)
  );
  DFF_X1 \_r[15]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00050_),
    .Q(_r[15]),
    .QN(_10416_)
  );
  DFF_X1 \_r[16]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00051_),
    .Q(_r[16]),
    .QN(_10415_)
  );
  DFF_X1 \_r[17]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00052_),
    .Q(_r[17]),
    .QN(_10414_)
  );
  DFF_X1 \_r[18]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00053_),
    .Q(_r[18]),
    .QN(_10413_)
  );
  DFF_X1 \_r[19]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00054_),
    .Q(_r[19]),
    .QN(_10412_)
  );
  DFF_X1 \_r[1]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00036_),
    .Q(_r[1]),
    .QN(_10430_)
  );
  DFF_X1 \_r[20]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00055_),
    .Q(_r[20]),
    .QN(_10411_)
  );
  DFF_X1 \_r[21]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00056_),
    .Q(_r[21]),
    .QN(_10410_)
  );
  DFF_X1 \_r[22]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00057_),
    .Q(_r[22]),
    .QN(_10409_)
  );
  DFF_X1 \_r[23]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00058_),
    .Q(_r[23]),
    .QN(_10408_)
  );
  DFF_X1 \_r[24]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00059_),
    .Q(_r[24]),
    .QN(_10407_)
  );
  DFF_X1 \_r[25]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00060_),
    .Q(_r[25]),
    .QN(_10406_)
  );
  DFF_X1 \_r[26]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00061_),
    .Q(_r[26]),
    .QN(_10405_)
  );
  DFF_X1 \_r[27]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00062_),
    .Q(_r[27]),
    .QN(_10404_)
  );
  DFF_X1 \_r[28]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00063_),
    .Q(_r[28]),
    .QN(_10403_)
  );
  DFF_X1 \_r[29]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00064_),
    .Q(_r[29]),
    .QN(_10402_)
  );
  DFF_X1 \_r[2]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00037_),
    .Q(_r[2]),
    .QN(_10429_)
  );
  DFF_X1 \_r[30]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00065_),
    .Q(_r[30]),
    .QN(_10401_)
  );
  DFF_X1 \_r[31]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00066_),
    .Q(_r[31]),
    .QN(_10400_)
  );
  DFF_X1 \_r[3]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00038_),
    .Q(_r[3]),
    .QN(_10428_)
  );
  DFF_X1 \_r[4]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00039_),
    .Q(_r[4]),
    .QN(_10427_)
  );
  DFF_X1 \_r[5]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00040_),
    .Q(_r[5]),
    .QN(_10426_)
  );
  DFF_X1 \_r[6]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00041_),
    .Q(_r[6]),
    .QN(_10425_)
  );
  DFF_X1 \_r[7]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00042_),
    .Q(_r[7]),
    .QN(_10424_)
  );
  DFF_X1 \_r[8]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00043_),
    .Q(_r[8]),
    .QN(_10423_)
  );
  DFF_X1 \_r[9]$_SDFFE_PP0P_  (
    .CK(clock),
    .D(_00044_),
    .Q(_r[9]),
    .QN(_10422_)
  );
  ALU alu (
    .io_adder_out(alu_io_adder_out),
    .io_cmp_out(alu_io_cmp_out),
    .io_fn(ex_ctrl_alu_fn),
    .io_in1(alu_io_in1),
    .io_in2(alu_io_in2),
    .io_out(alu_io_out)
  );
  DFF_X1 \blocked$_DFF_P_  (
    .CK(clock),
    .D(_00000_),
    .Q(blocked),
    .QN(_08905_)
  );
  BreakpointUnit bpu (
    .io_bp_0_address(bpu_io_bp_0_address),
    .io_bp_0_control_action(bpu_io_bp_0_control_action),
    .io_bp_0_control_r(bpu_io_bp_0_control_r),
    .io_bp_0_control_tmatch(bpu_io_bp_0_control_tmatch),
    .io_bp_0_control_w(bpu_io_bp_0_control_w),
    .io_bp_0_control_x(bpu_io_bp_0_control_x),
    .io_debug_if(bpu_io_debug_if),
    .io_debug_ld(bpu_io_debug_ld),
    .io_debug_st(bpu_io_debug_st),
    .io_ea(mem_reg_wdata),
    .io_pc(bpu_io_pc),
    .io_status_debug(bpu_io_status_debug),
    .io_xcpt_if(bpu_io_xcpt_if),
    .io_xcpt_ld(bpu_io_xcpt_ld),
    .io_xcpt_st(bpu_io_xcpt_st)
  );
  CSRFile csr (
    .clock(clock),
    .io_bp_0_address(bpu_io_bp_0_address),
    .io_bp_0_control_action(bpu_io_bp_0_control_action),
    .io_bp_0_control_r(bpu_io_bp_0_control_r),
    .io_bp_0_control_tmatch(bpu_io_bp_0_control_tmatch),
    .io_bp_0_control_w(bpu_io_bp_0_control_w),
    .io_bp_0_control_x(bpu_io_bp_0_control_x),
    .io_cause(csr_io_cause),
    .io_csr_stall(csr_io_csr_stall),
    .io_customCSRs_0_value({ csr_io_customCSRs_0_value[31:2], io_ptw_customCSRs_csrs_0_value[1], csr_io_customCSRs_0_value[0] }),
    .io_decode_0_fp_csr(csr_io_decode_0_fp_csr),
    .io_decode_0_fp_illegal(csr_io_decode_0_fp_illegal),
    .io_decode_0_inst(csr_io_decode_0_inst),
    .io_decode_0_read_illegal(csr_io_decode_0_read_illegal),
    .io_decode_0_rocc_illegal(csr_io_decode_0_rocc_illegal),
    .io_decode_0_system_illegal(csr_io_decode_0_system_illegal),
    .io_decode_0_write_flush(csr_io_decode_0_write_flush),
    .io_decode_0_write_illegal(csr_io_decode_0_write_illegal),
    .io_eret(csr_io_eret),
    .io_evec(csr_io_evec),
    .io_exception(csr_io_exception),
    .io_gva(1'h0),
    .io_hartid(io_hartid),
    .io_inhibit_cycle(csr_io_inhibit_cycle),
    .io_inst_0({ _csr_io_inst_0_T_3, wb_reg_raw_inst[15:0] }),
    .io_interrupt(csr_io_interrupt),
    .io_interrupt_cause(csr_io_interrupt_cause),
    .io_interrupts_debug(io_interrupts_debug),
    .io_interrupts_meip(io_interrupts_meip),
    .io_interrupts_msip(io_interrupts_msip),
    .io_interrupts_mtip(io_interrupts_mtip),
    .io_pc(wb_reg_pc),
    .io_pmp_0_addr(csr_io_pmp_0_addr),
    .io_pmp_0_cfg_a(csr_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_l(csr_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_r(csr_io_pmp_0_cfg_r),
    .io_pmp_0_cfg_w(csr_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_x(csr_io_pmp_0_cfg_x),
    .io_pmp_0_mask(csr_io_pmp_0_mask),
    .io_pmp_1_addr(csr_io_pmp_1_addr),
    .io_pmp_1_cfg_a(csr_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_l(csr_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_r(csr_io_pmp_1_cfg_r),
    .io_pmp_1_cfg_w(csr_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_x(csr_io_pmp_1_cfg_x),
    .io_pmp_1_mask(csr_io_pmp_1_mask),
    .io_pmp_2_addr(csr_io_pmp_2_addr),
    .io_pmp_2_cfg_a(csr_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_l(csr_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_r(csr_io_pmp_2_cfg_r),
    .io_pmp_2_cfg_w(csr_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_x(csr_io_pmp_2_cfg_x),
    .io_pmp_2_mask(csr_io_pmp_2_mask),
    .io_pmp_3_addr(csr_io_pmp_3_addr),
    .io_pmp_3_cfg_a(csr_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_l(csr_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_r(csr_io_pmp_3_cfg_r),
    .io_pmp_3_cfg_w(csr_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_x(csr_io_pmp_3_cfg_x),
    .io_pmp_3_mask(csr_io_pmp_3_mask),
    .io_pmp_4_addr(csr_io_pmp_4_addr),
    .io_pmp_4_cfg_a(csr_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_l(csr_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_r(csr_io_pmp_4_cfg_r),
    .io_pmp_4_cfg_w(csr_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_x(csr_io_pmp_4_cfg_x),
    .io_pmp_4_mask(csr_io_pmp_4_mask),
    .io_pmp_5_addr(csr_io_pmp_5_addr),
    .io_pmp_5_cfg_a(csr_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_l(csr_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_r(csr_io_pmp_5_cfg_r),
    .io_pmp_5_cfg_w(csr_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_x(csr_io_pmp_5_cfg_x),
    .io_pmp_5_mask(csr_io_pmp_5_mask),
    .io_pmp_6_addr(csr_io_pmp_6_addr),
    .io_pmp_6_cfg_a(csr_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_l(csr_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_r(csr_io_pmp_6_cfg_r),
    .io_pmp_6_cfg_w(csr_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_x(csr_io_pmp_6_cfg_x),
    .io_pmp_6_mask(csr_io_pmp_6_mask),
    .io_pmp_7_addr(csr_io_pmp_7_addr),
    .io_pmp_7_cfg_a(csr_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_l(csr_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_r(csr_io_pmp_7_cfg_r),
    .io_pmp_7_cfg_w(csr_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_x(csr_io_pmp_7_cfg_x),
    .io_pmp_7_mask(csr_io_pmp_7_mask),
    .io_retire(csr_io_retire),
    .io_rw_addr(wb_reg_inst[31:20]),
    .io_rw_cmd({ csr_io_rw_cmd[2], wb_ctrl_csr[1:0] }),
    .io_rw_rdata(csr_io_rw_rdata),
    .io_rw_wdata(wb_reg_wdata),
    .io_singleStep(csr_io_singleStep),
    .io_status_cease(csr_io_status_cease),
    .io_status_debug(bpu_io_status_debug),
    .io_status_dprv(csr_io_status_dprv),
    .io_status_dv(csr_io_status_dv),
    .io_status_fs(csr_io_status_fs),
    .io_status_gva(csr_io_status_gva),
    .io_status_hie(csr_io_status_hie),
    .io_status_isa(csr_io_status_isa),
    .io_status_mbe(csr_io_status_mbe),
    .io_status_mie(csr_io_status_mie),
    .io_status_mpie(csr_io_status_mpie),
    .io_status_mpp(csr_io_status_mpp),
    .io_status_mprv(csr_io_status_mprv),
    .io_status_mpv(csr_io_status_mpv),
    .io_status_mxr(csr_io_status_mxr),
    .io_status_prv(csr_io_status_prv),
    .io_status_sbe(csr_io_status_sbe),
    .io_status_sd(csr_io_status_sd),
    .io_status_sd_rv32(csr_io_status_sd_rv32),
    .io_status_sie(csr_io_status_sie),
    .io_status_spie(csr_io_status_spie),
    .io_status_spp(csr_io_status_spp),
    .io_status_sum(csr_io_status_sum),
    .io_status_sxl(csr_io_status_sxl),
    .io_status_tsr(csr_io_status_tsr),
    .io_status_tvm(csr_io_status_tvm),
    .io_status_tw(csr_io_status_tw),
    .io_status_ube(csr_io_status_ube),
    .io_status_uie(csr_io_status_uie),
    .io_status_upie(csr_io_status_upie),
    .io_status_uxl(csr_io_status_uxl),
    .io_status_v(csr_io_status_v),
    .io_status_vs(csr_io_status_vs),
    .io_status_wfi(csr_io_status_wfi),
    .io_status_xs(csr_io_status_xs),
    .io_status_zero1(csr_io_status_zero1),
    .io_status_zero2(csr_io_status_zero2),
    .io_time(csr_io_time),
    .io_trace_0_exception(csr_io_trace_0_exception),
    .io_trace_0_iaddr(csr_io_trace_0_iaddr),
    .io_trace_0_insn(csr_io_trace_0_insn),
    .io_trace_0_valid(csr_io_trace_0_valid),
    .io_tval(csr_io_tval),
    .io_ungated_clock(clock),
    .reset(reset)
  );
  MulDiv div (
    .clock(clock),
    .io_kill(div_io_kill),
    .io_req_bits_fn(ex_ctrl_alu_fn),
    .io_req_bits_in1(_ex_op1_T),
    .io_req_bits_in2(_ex_op2_T),
    .io_req_bits_tag(ex_reg_inst[11:7]),
    .io_req_ready(div_io_req_ready),
    .io_req_valid(div_io_req_valid),
    .io_resp_bits_data(div_io_resp_bits_data),
    .io_resp_bits_tag(div_io_resp_bits_tag),
    .io_resp_ready(div_io_resp_ready),
    .io_resp_valid(div_io_resp_valid),
    .reset(reset)
  );
  DFF_X1 \div_io_kill_REG$_DFF_P_  (
    .CK(clock),
    .D(_00001_),
    .Q(div_io_kill_REG),
    .QN(_10431_)
  );
  DFF_X1 \ex_ctrl_alu_fn[0]$_SDFFCE_PP0N_  (
    .CK(clock),
    .D(_00565_),
    .Q(ex_ctrl_alu_fn[0]),
    .QN(_09915_)
  );
  DFF_X1 \ex_ctrl_alu_fn[1]$_SDFFCE_PP0N_  (
    .CK(clock),
    .D(_00566_),
    .Q(ex_ctrl_alu_fn[1]),
    .QN(_09914_)
  );
  DFF_X1 \ex_ctrl_alu_fn[2]$_SDFFCE_PP0N_  (
    .CK(clock),
    .D(_00567_),
    .Q(ex_ctrl_alu_fn[2]),
    .QN(_09913_)
  );
  DFF_X1 \ex_ctrl_alu_fn[3]$_SDFFCE_PP0N_  (
    .CK(clock),
    .D(_00568_),
    .Q(ex_ctrl_alu_fn[3]),
    .QN(_09912_)
  );
  DFF_X1 \ex_ctrl_branch$_DFFE_PN_  (
    .CK(clock),
    .D(_00579_),
    .Q(ex_ctrl_branch),
    .QN(_09907_)
  );
  DFF_X1 \ex_ctrl_csr[0]$_SDFFCE_PP0N_  (
    .CK(clock),
    .D(_00589_),
    .Q(ex_ctrl_csr[0]),
    .QN(_09898_)
  );
  DFF_X1 \ex_ctrl_csr[1]$_SDFFCE_PP0N_  (
    .CK(clock),
    .D(_00557_),
    .Q(ex_ctrl_csr[1]),
    .QN(_09919_)
  );
  DFF_X1 \ex_ctrl_csr[2]$_SDFFCE_PP0N_  (
    .CK(clock),
    .D(_00590_),
    .Q(ex_ctrl_csr[2]),
    .QN(_09897_)
  );
  DFF_X1 \ex_ctrl_div$_DFFE_PN_  (
    .CK(clock),
    .D(_00560_),
    .Q(ex_ctrl_div),
    .QN(_09916_)
  );
  DFF_X1 \ex_ctrl_fence_i$_DFFE_PN_  (
    .CK(clock),
    .D(_00558_),
    .Q(ex_ctrl_fence_i),
    .QN(_09918_)
  );
  DFF_X1 \ex_ctrl_jal$_DFFE_PN_  (
    .CK(clock),
    .D(_00578_),
    .Q(ex_ctrl_jal),
    .QN(_09908_)
  );
  DFF_X1 \ex_ctrl_jalr$_DFFE_PN_  (
    .CK(clock),
    .D(_00577_),
    .Q(ex_ctrl_jalr),
    .QN(_09909_)
  );
  DFF_X1 \ex_ctrl_mem$_DFFE_PN_  (
    .CK(clock),
    .D(_00569_),
    .Q(ex_ctrl_mem),
    .QN(_09911_)
  );
  DFF_X1 \ex_ctrl_mem_cmd[0]$_DFFE_PN_  (
    .CK(clock),
    .D(_00561_),
    .Q(ex_ctrl_mem_cmd[0]),
    .QN(_00027_)
  );
  DFF_X1 \ex_ctrl_mem_cmd[1]$_DFFE_PN_  (
    .CK(clock),
    .D(_00562_),
    .Q(ex_ctrl_mem_cmd[1]),
    .QN(_00026_)
  );
  DFF_X1 \ex_ctrl_mem_cmd[2]$_DFFE_PN_  (
    .CK(clock),
    .D(_00563_),
    .Q(ex_ctrl_mem_cmd[2]),
    .QN(_00025_)
  );
  DFF_X1 \ex_ctrl_mem_cmd[3]$_DFFE_PN_  (
    .CK(clock),
    .D(_00564_),
    .Q(ex_ctrl_mem_cmd[3]),
    .QN(_00024_)
  );
  DFF_X1 \ex_ctrl_rxs2$_DFFE_PN_  (
    .CK(clock),
    .D(_00576_),
    .Q(ex_ctrl_rxs2),
    .QN(_09910_)
  );
  DFF_X1 \ex_ctrl_sel_alu1[0]$_DFFE_PN_  (
    .CK(clock),
    .D(_00573_),
    .Q(ex_ctrl_sel_alu1[0]),
    .QN(_00020_)
  );
  DFF_X1 \ex_ctrl_sel_alu1[1]$_DFFE_PN_  (
    .CK(clock),
    .D(_00574_),
    .Q(ex_ctrl_sel_alu1[1]),
    .QN(_00019_)
  );
  DFF_X1 \ex_ctrl_sel_alu2[0]$_DFFE_PN_  (
    .CK(clock),
    .D(_00575_),
    .Q(ex_ctrl_sel_alu2[0]),
    .QN(_00018_)
  );
  DFF_X1 \ex_ctrl_sel_alu2[1]$_SDFFCE_PP0N_  (
    .CK(clock),
    .D(_00747_),
    .Q(ex_ctrl_sel_alu2[1]),
    .QN(_00012_)
  );
  DFF_X1 \ex_ctrl_sel_imm[0]$_DFFE_PN_  (
    .CK(clock),
    .D(_00570_),
    .Q(ex_ctrl_sel_imm[0]),
    .QN(_00023_)
  );
  DFF_X1 \ex_ctrl_sel_imm[1]$_DFFE_PN_  (
    .CK(clock),
    .D(_00571_),
    .Q(ex_ctrl_sel_imm[1]),
    .QN(_00022_)
  );
  DFF_X1 \ex_ctrl_sel_imm[2]$_DFFE_PN_  (
    .CK(clock),
    .D(_00572_),
    .Q(ex_ctrl_sel_imm[2]),
    .QN(_00021_)
  );
  DFF_X1 \ex_ctrl_wxd$_DFFE_PN_  (
    .CK(clock),
    .D(_00559_),
    .Q(ex_ctrl_wxd),
    .QN(_09917_)
  );
  DFF_X1 \ex_reg_cause[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00584_),
    .Q(ex_reg_cause[0]),
    .QN(_09903_)
  );
  DFF_X1 \ex_reg_cause[10]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00463_),
    .Q(ex_reg_cause[10]),
    .QN(_10011_)
  );
  DFF_X1 \ex_reg_cause[11]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00464_),
    .Q(ex_reg_cause[11]),
    .QN(_10010_)
  );
  DFF_X1 \ex_reg_cause[12]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00465_),
    .Q(ex_reg_cause[12]),
    .QN(_10009_)
  );
  DFF_X1 \ex_reg_cause[13]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00466_),
    .Q(ex_reg_cause[13]),
    .QN(_10008_)
  );
  DFF_X1 \ex_reg_cause[14]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00467_),
    .Q(ex_reg_cause[14]),
    .QN(_10007_)
  );
  DFF_X1 \ex_reg_cause[15]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00468_),
    .Q(ex_reg_cause[15]),
    .QN(_10006_)
  );
  DFF_X1 \ex_reg_cause[16]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00469_),
    .Q(ex_reg_cause[16]),
    .QN(_10005_)
  );
  DFF_X1 \ex_reg_cause[17]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00470_),
    .Q(ex_reg_cause[17]),
    .QN(_10004_)
  );
  DFF_X1 \ex_reg_cause[18]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00471_),
    .Q(ex_reg_cause[18]),
    .QN(_10003_)
  );
  DFF_X1 \ex_reg_cause[19]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00472_),
    .Q(ex_reg_cause[19]),
    .QN(_10002_)
  );
  DFF_X1 \ex_reg_cause[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00585_),
    .Q(ex_reg_cause[1]),
    .QN(_09902_)
  );
  DFF_X1 \ex_reg_cause[20]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00473_),
    .Q(ex_reg_cause[20]),
    .QN(_10001_)
  );
  DFF_X1 \ex_reg_cause[21]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00474_),
    .Q(ex_reg_cause[21]),
    .QN(_10000_)
  );
  DFF_X1 \ex_reg_cause[22]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00475_),
    .Q(ex_reg_cause[22]),
    .QN(_09999_)
  );
  DFF_X1 \ex_reg_cause[23]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00476_),
    .Q(ex_reg_cause[23]),
    .QN(_09998_)
  );
  DFF_X1 \ex_reg_cause[24]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00477_),
    .Q(ex_reg_cause[24]),
    .QN(_09997_)
  );
  DFF_X1 \ex_reg_cause[25]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00478_),
    .Q(ex_reg_cause[25]),
    .QN(_09996_)
  );
  DFF_X1 \ex_reg_cause[26]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00479_),
    .Q(ex_reg_cause[26]),
    .QN(_09995_)
  );
  DFF_X1 \ex_reg_cause[27]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00480_),
    .Q(ex_reg_cause[27]),
    .QN(_09994_)
  );
  DFF_X1 \ex_reg_cause[28]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00481_),
    .Q(ex_reg_cause[28]),
    .QN(_09993_)
  );
  DFF_X1 \ex_reg_cause[29]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00482_),
    .Q(ex_reg_cause[29]),
    .QN(_09992_)
  );
  DFF_X1 \ex_reg_cause[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00586_),
    .Q(ex_reg_cause[2]),
    .QN(_09901_)
  );
  DFF_X1 \ex_reg_cause[30]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00483_),
    .Q(ex_reg_cause[30]),
    .QN(_09991_)
  );
  DFF_X1 \ex_reg_cause[31]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00484_),
    .Q(ex_reg_cause[31]),
    .QN(_09990_)
  );
  DFF_X1 \ex_reg_cause[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00587_),
    .Q(ex_reg_cause[3]),
    .QN(_09900_)
  );
  DFF_X1 \ex_reg_cause[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00588_),
    .Q(ex_reg_cause[4]),
    .QN(_09899_)
  );
  DFF_X1 \ex_reg_cause[5]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00458_),
    .Q(ex_reg_cause[5]),
    .QN(_10016_)
  );
  DFF_X1 \ex_reg_cause[6]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00459_),
    .Q(ex_reg_cause[6]),
    .QN(_10015_)
  );
  DFF_X1 \ex_reg_cause[7]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00460_),
    .Q(ex_reg_cause[7]),
    .QN(_10014_)
  );
  DFF_X1 \ex_reg_cause[8]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00461_),
    .Q(ex_reg_cause[8]),
    .QN(_10013_)
  );
  DFF_X1 \ex_reg_cause[9]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00462_),
    .Q(ex_reg_cause[9]),
    .QN(_10012_)
  );
  DFF_X1 \ex_reg_flush_pipe$_DFFE_PN_  (
    .CK(clock),
    .D(_00518_),
    .Q(ex_reg_flush_pipe),
    .QN(_10439_)
  );
  DFF_X1 \ex_reg_inst[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00434_),
    .Q(ex_reg_inst[10]),
    .QN(_10038_)
  );
  DFF_X1 \ex_reg_inst[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00435_),
    .Q(ex_reg_inst[11]),
    .QN(_10037_)
  );
  DFF_X1 \ex_reg_inst[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00436_),
    .Q(ex_reg_inst[12]),
    .QN(_10036_)
  );
  DFF_X1 \ex_reg_inst[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00437_),
    .Q(ex_reg_inst[13]),
    .QN(_10035_)
  );
  DFF_X1 \ex_reg_inst[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00438_),
    .Q(ex_reg_inst[14]),
    .QN(io_dmem_req_bits_signed)
  );
  DFF_X1 \ex_reg_inst[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00439_),
    .Q(ex_reg_inst[15]),
    .QN(_10034_)
  );
  DFF_X1 \ex_reg_inst[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00440_),
    .Q(ex_reg_inst[16]),
    .QN(_10033_)
  );
  DFF_X1 \ex_reg_inst[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00441_),
    .Q(ex_reg_inst[17]),
    .QN(_10032_)
  );
  DFF_X1 \ex_reg_inst[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00442_),
    .Q(ex_reg_inst[18]),
    .QN(_10031_)
  );
  DFF_X1 \ex_reg_inst[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00443_),
    .Q(ex_reg_inst[19]),
    .QN(_10030_)
  );
  DFF_X1 \ex_reg_inst[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00444_),
    .Q(ex_reg_inst[20]),
    .QN(_10029_)
  );
  DFF_X1 \ex_reg_inst[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00445_),
    .Q(ex_reg_inst[21]),
    .QN(_10028_)
  );
  DFF_X1 \ex_reg_inst[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00446_),
    .Q(ex_reg_inst[22]),
    .QN(_10027_)
  );
  DFF_X1 \ex_reg_inst[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00447_),
    .Q(ex_reg_inst[23]),
    .QN(_10026_)
  );
  DFF_X1 \ex_reg_inst[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00448_),
    .Q(ex_reg_inst[24]),
    .QN(_10025_)
  );
  DFF_X1 \ex_reg_inst[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00449_),
    .Q(ex_reg_inst[25]),
    .QN(_10024_)
  );
  DFF_X1 \ex_reg_inst[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00450_),
    .Q(ex_reg_inst[26]),
    .QN(_10023_)
  );
  DFF_X1 \ex_reg_inst[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00451_),
    .Q(ex_reg_inst[27]),
    .QN(_10022_)
  );
  DFF_X1 \ex_reg_inst[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00452_),
    .Q(ex_reg_inst[28]),
    .QN(_10021_)
  );
  DFF_X1 \ex_reg_inst[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00453_),
    .Q(ex_reg_inst[29]),
    .QN(_10020_)
  );
  DFF_X1 \ex_reg_inst[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00454_),
    .Q(ex_reg_inst[30]),
    .QN(_10019_)
  );
  DFF_X1 \ex_reg_inst[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00455_),
    .Q(ex_reg_inst[31]),
    .QN(_10018_)
  );
  DFF_X1 \ex_reg_inst[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00431_),
    .Q(ex_reg_inst[7]),
    .QN(_10041_)
  );
  DFF_X1 \ex_reg_inst[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00432_),
    .Q(ex_reg_inst[8]),
    .QN(_10040_)
  );
  DFF_X1 \ex_reg_inst[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00433_),
    .Q(ex_reg_inst[9]),
    .QN(_10039_)
  );
  DFF_X1 \ex_reg_load_use$_DFFE_PN_  (
    .CK(clock),
    .D(_00517_),
    .Q(ex_reg_load_use),
    .QN(_10438_)
  );
  DFF_X1 \ex_reg_mem_size[0]$_DFFE_PN_  (
    .CK(clock),
    .D(_00456_),
    .Q(ex_reg_mem_size[0]),
    .QN(_10441_[0])
  );
  DFF_X1 \ex_reg_mem_size[1]$_DFFE_PN_  (
    .CK(clock),
    .D(_00457_),
    .Q(ex_reg_mem_size[1]),
    .QN(_10442_[1])
  );
  DFF_X1 \ex_reg_pc[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00485_),
    .Q(ex_reg_pc[0]),
    .QN(_09989_)
  );
  DFF_X1 \ex_reg_pc[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00495_),
    .Q(ex_reg_pc[10]),
    .QN(_09979_)
  );
  DFF_X1 \ex_reg_pc[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00496_),
    .Q(ex_reg_pc[11]),
    .QN(_09978_)
  );
  DFF_X1 \ex_reg_pc[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00497_),
    .Q(ex_reg_pc[12]),
    .QN(_09977_)
  );
  DFF_X1 \ex_reg_pc[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00498_),
    .Q(ex_reg_pc[13]),
    .QN(_09976_)
  );
  DFF_X1 \ex_reg_pc[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00499_),
    .Q(ex_reg_pc[14]),
    .QN(_09975_)
  );
  DFF_X1 \ex_reg_pc[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00500_),
    .Q(ex_reg_pc[15]),
    .QN(_09974_)
  );
  DFF_X1 \ex_reg_pc[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00501_),
    .Q(ex_reg_pc[16]),
    .QN(_09973_)
  );
  DFF_X1 \ex_reg_pc[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00502_),
    .Q(ex_reg_pc[17]),
    .QN(_09972_)
  );
  DFF_X1 \ex_reg_pc[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00503_),
    .Q(ex_reg_pc[18]),
    .QN(_09971_)
  );
  DFF_X1 \ex_reg_pc[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00504_),
    .Q(ex_reg_pc[19]),
    .QN(_09970_)
  );
  DFF_X1 \ex_reg_pc[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00486_),
    .Q(ex_reg_pc[1]),
    .QN(_09988_)
  );
  DFF_X1 \ex_reg_pc[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00505_),
    .Q(ex_reg_pc[20]),
    .QN(_09969_)
  );
  DFF_X1 \ex_reg_pc[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00506_),
    .Q(ex_reg_pc[21]),
    .QN(_09968_)
  );
  DFF_X1 \ex_reg_pc[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00507_),
    .Q(ex_reg_pc[22]),
    .QN(_09967_)
  );
  DFF_X1 \ex_reg_pc[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00508_),
    .Q(ex_reg_pc[23]),
    .QN(_09966_)
  );
  DFF_X1 \ex_reg_pc[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00509_),
    .Q(ex_reg_pc[24]),
    .QN(_09965_)
  );
  DFF_X1 \ex_reg_pc[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00510_),
    .Q(ex_reg_pc[25]),
    .QN(_09964_)
  );
  DFF_X1 \ex_reg_pc[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00511_),
    .Q(ex_reg_pc[26]),
    .QN(_09963_)
  );
  DFF_X1 \ex_reg_pc[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00512_),
    .Q(ex_reg_pc[27]),
    .QN(_09962_)
  );
  DFF_X1 \ex_reg_pc[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00513_),
    .Q(ex_reg_pc[28]),
    .QN(_09961_)
  );
  DFF_X1 \ex_reg_pc[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00514_),
    .Q(ex_reg_pc[29]),
    .QN(_09960_)
  );
  DFF_X1 \ex_reg_pc[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00487_),
    .Q(ex_reg_pc[2]),
    .QN(_09987_)
  );
  DFF_X1 \ex_reg_pc[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00515_),
    .Q(ex_reg_pc[30]),
    .QN(_09959_)
  );
  DFF_X1 \ex_reg_pc[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00516_),
    .Q(ex_reg_pc[31]),
    .QN(_09958_)
  );
  DFF_X1 \ex_reg_pc[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00488_),
    .Q(ex_reg_pc[3]),
    .QN(_09986_)
  );
  DFF_X1 \ex_reg_pc[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00489_),
    .Q(ex_reg_pc[4]),
    .QN(_09985_)
  );
  DFF_X1 \ex_reg_pc[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00490_),
    .Q(ex_reg_pc[5]),
    .QN(_09984_)
  );
  DFF_X1 \ex_reg_pc[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00491_),
    .Q(ex_reg_pc[6]),
    .QN(_09983_)
  );
  DFF_X1 \ex_reg_pc[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00492_),
    .Q(ex_reg_pc[7]),
    .QN(_09982_)
  );
  DFF_X1 \ex_reg_pc[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00493_),
    .Q(ex_reg_pc[8]),
    .QN(_09981_)
  );
  DFF_X1 \ex_reg_pc[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00494_),
    .Q(ex_reg_pc[9]),
    .QN(_09980_)
  );
  DFF_X1 \ex_reg_raw_inst[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00415_),
    .Q(ex_reg_raw_inst[0]),
    .QN(_10057_)
  );
  DFF_X1 \ex_reg_raw_inst[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00425_),
    .Q(ex_reg_raw_inst[10]),
    .QN(_10047_)
  );
  DFF_X1 \ex_reg_raw_inst[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00426_),
    .Q(ex_reg_raw_inst[11]),
    .QN(_10046_)
  );
  DFF_X1 \ex_reg_raw_inst[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00427_),
    .Q(ex_reg_raw_inst[12]),
    .QN(_10045_)
  );
  DFF_X1 \ex_reg_raw_inst[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00428_),
    .Q(ex_reg_raw_inst[13]),
    .QN(_10044_)
  );
  DFF_X1 \ex_reg_raw_inst[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00429_),
    .Q(ex_reg_raw_inst[14]),
    .QN(_10043_)
  );
  DFF_X1 \ex_reg_raw_inst[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00430_),
    .Q(ex_reg_raw_inst[15]),
    .QN(_10042_)
  );
  DFF_X1 \ex_reg_raw_inst[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00416_),
    .Q(ex_reg_raw_inst[1]),
    .QN(_10056_)
  );
  DFF_X1 \ex_reg_raw_inst[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00417_),
    .Q(ex_reg_raw_inst[2]),
    .QN(_10055_)
  );
  DFF_X1 \ex_reg_raw_inst[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00418_),
    .Q(ex_reg_raw_inst[3]),
    .QN(_10054_)
  );
  DFF_X1 \ex_reg_raw_inst[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00419_),
    .Q(ex_reg_raw_inst[4]),
    .QN(_10053_)
  );
  DFF_X1 \ex_reg_raw_inst[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00420_),
    .Q(ex_reg_raw_inst[5]),
    .QN(_10052_)
  );
  DFF_X1 \ex_reg_raw_inst[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00421_),
    .Q(ex_reg_raw_inst[6]),
    .QN(_10051_)
  );
  DFF_X1 \ex_reg_raw_inst[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00422_),
    .Q(ex_reg_raw_inst[7]),
    .QN(_10050_)
  );
  DFF_X1 \ex_reg_raw_inst[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00423_),
    .Q(ex_reg_raw_inst[8]),
    .QN(_10049_)
  );
  DFF_X1 \ex_reg_raw_inst[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00424_),
    .Q(ex_reg_raw_inst[9]),
    .QN(_10048_)
  );
  DFF_X1 \ex_reg_replay$_DFF_P_  (
    .CK(clock),
    .D(_00002_),
    .Q(ex_reg_replay),
    .QN(_10017_)
  );
  DFF_X1 \ex_reg_rs_bypass_0$_SDFFCE_PP0N_  (
    .CK(clock),
    .D(_00100_),
    .Q(ex_reg_rs_bypass_0),
    .QN(_10368_)
  );
  DFF_X1 \ex_reg_rs_bypass_1$_DFFE_PN_  (
    .CK(clock),
    .D(_00099_),
    .Q(ex_reg_rs_bypass_1),
    .QN(_10369_)
  );
  DFF_X1 \ex_reg_rs_lsb_0[0]$_DFFE_PN_  (
    .CK(clock),
    .D(_00097_),
    .Q(ex_reg_rs_lsb_0[0]),
    .QN(_00032_)
  );
  DFF_X1 \ex_reg_rs_lsb_0[1]$_DFFE_PN_  (
    .CK(clock),
    .D(_00098_),
    .Q(ex_reg_rs_lsb_0[1]),
    .QN(_00031_)
  );
  DFF_X1 \ex_reg_rs_lsb_1[0]$_DFFE_PN_  (
    .CK(clock),
    .D(_00580_),
    .Q(ex_reg_rs_lsb_1[0]),
    .QN(_00017_)
  );
  DFF_X1 \ex_reg_rs_lsb_1[1]$_DFFE_PN_  (
    .CK(clock),
    .D(_00581_),
    .Q(ex_reg_rs_lsb_1[1]),
    .QN(_00035_)
  );
  DFF_X1 \ex_reg_rs_msb_0[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00067_),
    .Q(ex_reg_rs_msb_0[0]),
    .QN(_10399_)
  );
  DFF_X1 \ex_reg_rs_msb_0[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00077_),
    .Q(ex_reg_rs_msb_0[10]),
    .QN(_10389_)
  );
  DFF_X1 \ex_reg_rs_msb_0[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00078_),
    .Q(ex_reg_rs_msb_0[11]),
    .QN(_10388_)
  );
  DFF_X1 \ex_reg_rs_msb_0[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00079_),
    .Q(ex_reg_rs_msb_0[12]),
    .QN(_10387_)
  );
  DFF_X1 \ex_reg_rs_msb_0[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00080_),
    .Q(ex_reg_rs_msb_0[13]),
    .QN(_10386_)
  );
  DFF_X1 \ex_reg_rs_msb_0[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00081_),
    .Q(ex_reg_rs_msb_0[14]),
    .QN(_10385_)
  );
  DFF_X1 \ex_reg_rs_msb_0[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00082_),
    .Q(ex_reg_rs_msb_0[15]),
    .QN(_10384_)
  );
  DFF_X1 \ex_reg_rs_msb_0[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00083_),
    .Q(ex_reg_rs_msb_0[16]),
    .QN(_10383_)
  );
  DFF_X1 \ex_reg_rs_msb_0[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00084_),
    .Q(ex_reg_rs_msb_0[17]),
    .QN(_10382_)
  );
  DFF_X1 \ex_reg_rs_msb_0[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00085_),
    .Q(ex_reg_rs_msb_0[18]),
    .QN(_10381_)
  );
  DFF_X1 \ex_reg_rs_msb_0[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00086_),
    .Q(ex_reg_rs_msb_0[19]),
    .QN(_10380_)
  );
  DFF_X1 \ex_reg_rs_msb_0[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00068_),
    .Q(ex_reg_rs_msb_0[1]),
    .QN(_10398_)
  );
  DFF_X1 \ex_reg_rs_msb_0[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00087_),
    .Q(ex_reg_rs_msb_0[20]),
    .QN(_10379_)
  );
  DFF_X1 \ex_reg_rs_msb_0[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00088_),
    .Q(ex_reg_rs_msb_0[21]),
    .QN(_10378_)
  );
  DFF_X1 \ex_reg_rs_msb_0[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00089_),
    .Q(ex_reg_rs_msb_0[22]),
    .QN(_10377_)
  );
  DFF_X1 \ex_reg_rs_msb_0[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00090_),
    .Q(ex_reg_rs_msb_0[23]),
    .QN(_10376_)
  );
  DFF_X1 \ex_reg_rs_msb_0[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00091_),
    .Q(ex_reg_rs_msb_0[24]),
    .QN(_10375_)
  );
  DFF_X1 \ex_reg_rs_msb_0[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00092_),
    .Q(ex_reg_rs_msb_0[25]),
    .QN(_10374_)
  );
  DFF_X1 \ex_reg_rs_msb_0[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00093_),
    .Q(ex_reg_rs_msb_0[26]),
    .QN(_10373_)
  );
  DFF_X1 \ex_reg_rs_msb_0[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00094_),
    .Q(ex_reg_rs_msb_0[27]),
    .QN(_10372_)
  );
  DFF_X1 \ex_reg_rs_msb_0[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00095_),
    .Q(ex_reg_rs_msb_0[28]),
    .QN(_10371_)
  );
  DFF_X1 \ex_reg_rs_msb_0[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00096_),
    .Q(ex_reg_rs_msb_0[29]),
    .QN(_10370_)
  );
  DFF_X1 \ex_reg_rs_msb_0[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00069_),
    .Q(ex_reg_rs_msb_0[2]),
    .QN(_10397_)
  );
  DFF_X1 \ex_reg_rs_msb_0[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00070_),
    .Q(ex_reg_rs_msb_0[3]),
    .QN(_10396_)
  );
  DFF_X1 \ex_reg_rs_msb_0[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00071_),
    .Q(ex_reg_rs_msb_0[4]),
    .QN(_10395_)
  );
  DFF_X1 \ex_reg_rs_msb_0[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00072_),
    .Q(ex_reg_rs_msb_0[5]),
    .QN(_10394_)
  );
  DFF_X1 \ex_reg_rs_msb_0[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00073_),
    .Q(ex_reg_rs_msb_0[6]),
    .QN(_10393_)
  );
  DFF_X1 \ex_reg_rs_msb_0[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00074_),
    .Q(ex_reg_rs_msb_0[7]),
    .QN(_10392_)
  );
  DFF_X1 \ex_reg_rs_msb_0[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00075_),
    .Q(ex_reg_rs_msb_0[8]),
    .QN(_10391_)
  );
  DFF_X1 \ex_reg_rs_msb_0[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00076_),
    .Q(ex_reg_rs_msb_0[9]),
    .QN(_10390_)
  );
  DFF_X1 \ex_reg_rs_msb_1[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00149_),
    .Q(ex_reg_rs_msb_1[0]),
    .QN(_10319_)
  );
  DFF_X1 \ex_reg_rs_msb_1[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00159_),
    .Q(ex_reg_rs_msb_1[10]),
    .QN(_10309_)
  );
  DFF_X1 \ex_reg_rs_msb_1[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00160_),
    .Q(ex_reg_rs_msb_1[11]),
    .QN(_10308_)
  );
  DFF_X1 \ex_reg_rs_msb_1[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00161_),
    .Q(ex_reg_rs_msb_1[12]),
    .QN(_10307_)
  );
  DFF_X1 \ex_reg_rs_msb_1[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00162_),
    .Q(ex_reg_rs_msb_1[13]),
    .QN(_10306_)
  );
  DFF_X1 \ex_reg_rs_msb_1[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00163_),
    .Q(ex_reg_rs_msb_1[14]),
    .QN(_10305_)
  );
  DFF_X1 \ex_reg_rs_msb_1[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00164_),
    .Q(ex_reg_rs_msb_1[15]),
    .QN(_10304_)
  );
  DFF_X1 \ex_reg_rs_msb_1[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00165_),
    .Q(ex_reg_rs_msb_1[16]),
    .QN(_10303_)
  );
  DFF_X1 \ex_reg_rs_msb_1[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00166_),
    .Q(ex_reg_rs_msb_1[17]),
    .QN(_10302_)
  );
  DFF_X1 \ex_reg_rs_msb_1[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00167_),
    .Q(ex_reg_rs_msb_1[18]),
    .QN(_10301_)
  );
  DFF_X1 \ex_reg_rs_msb_1[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00168_),
    .Q(ex_reg_rs_msb_1[19]),
    .QN(_10300_)
  );
  DFF_X1 \ex_reg_rs_msb_1[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00150_),
    .Q(ex_reg_rs_msb_1[1]),
    .QN(_10318_)
  );
  DFF_X1 \ex_reg_rs_msb_1[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00169_),
    .Q(ex_reg_rs_msb_1[20]),
    .QN(_10299_)
  );
  DFF_X1 \ex_reg_rs_msb_1[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00170_),
    .Q(ex_reg_rs_msb_1[21]),
    .QN(_10298_)
  );
  DFF_X1 \ex_reg_rs_msb_1[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00171_),
    .Q(ex_reg_rs_msb_1[22]),
    .QN(_10297_)
  );
  DFF_X1 \ex_reg_rs_msb_1[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00172_),
    .Q(ex_reg_rs_msb_1[23]),
    .QN(_10296_)
  );
  DFF_X1 \ex_reg_rs_msb_1[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00173_),
    .Q(ex_reg_rs_msb_1[24]),
    .QN(_10295_)
  );
  DFF_X1 \ex_reg_rs_msb_1[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00174_),
    .Q(ex_reg_rs_msb_1[25]),
    .QN(_10294_)
  );
  DFF_X1 \ex_reg_rs_msb_1[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00175_),
    .Q(ex_reg_rs_msb_1[26]),
    .QN(_10293_)
  );
  DFF_X1 \ex_reg_rs_msb_1[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00176_),
    .Q(ex_reg_rs_msb_1[27]),
    .QN(_10292_)
  );
  DFF_X1 \ex_reg_rs_msb_1[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00177_),
    .Q(ex_reg_rs_msb_1[28]),
    .QN(_10291_)
  );
  DFF_X1 \ex_reg_rs_msb_1[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00178_),
    .Q(ex_reg_rs_msb_1[29]),
    .QN(_10290_)
  );
  DFF_X1 \ex_reg_rs_msb_1[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00151_),
    .Q(ex_reg_rs_msb_1[2]),
    .QN(_10317_)
  );
  DFF_X1 \ex_reg_rs_msb_1[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00152_),
    .Q(ex_reg_rs_msb_1[3]),
    .QN(_10316_)
  );
  DFF_X1 \ex_reg_rs_msb_1[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00153_),
    .Q(ex_reg_rs_msb_1[4]),
    .QN(_10315_)
  );
  DFF_X1 \ex_reg_rs_msb_1[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00154_),
    .Q(ex_reg_rs_msb_1[5]),
    .QN(_10314_)
  );
  DFF_X1 \ex_reg_rs_msb_1[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00155_),
    .Q(ex_reg_rs_msb_1[6]),
    .QN(_10313_)
  );
  DFF_X1 \ex_reg_rs_msb_1[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00156_),
    .Q(ex_reg_rs_msb_1[7]),
    .QN(_10312_)
  );
  DFF_X1 \ex_reg_rs_msb_1[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00157_),
    .Q(ex_reg_rs_msb_1[8]),
    .QN(_10311_)
  );
  DFF_X1 \ex_reg_rs_msb_1[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00158_),
    .Q(ex_reg_rs_msb_1[9]),
    .QN(_10310_)
  );
  DFF_X1 \ex_reg_rvc$_DFFE_PN_  (
    .CK(clock),
    .D(_00179_),
    .Q(ex_reg_rvc),
    .QN(_ex_op2_T_1[2])
  );
  DFF_X1 \ex_reg_valid$_DFF_P_  (
    .CK(clock),
    .D(_ex_reg_valid_T),
    .Q(ex_reg_valid),
    .QN(_00034_)
  );
  DFF_X1 \ex_reg_xcpt$_DFF_P_  (
    .CK(clock),
    .D(_00003_),
    .Q(ex_reg_xcpt),
    .QN(_09957_)
  );
  DFF_X1 \ex_reg_xcpt_interrupt$_DFF_P_  (
    .CK(clock),
    .D(_00004_),
    .Q(ex_reg_xcpt_interrupt),
    .QN(_09956_)
  );
  IBuf ibuf (
    .clock(clock),
    .io_imem_bits_data(io_imem_resp_bits_data),
    .io_imem_bits_pc(io_imem_resp_bits_pc),
    .io_imem_bits_replay(io_imem_resp_bits_replay),
    .io_imem_bits_xcpt_ae_inst(io_imem_resp_bits_xcpt_ae_inst),
    .io_imem_ready(ibuf_io_imem_ready),
    .io_imem_valid(io_imem_resp_valid),
    .io_inst_0_bits_inst_bits(csr_io_decode_0_inst),
    .io_inst_0_bits_inst_rd(ibuf_io_inst_0_bits_inst_rd),
    .io_inst_0_bits_inst_rs1(ibuf_io_inst_0_bits_inst_rs1),
    .io_inst_0_bits_inst_rs2(ibuf_io_inst_0_bits_inst_rs2),
    .io_inst_0_bits_raw(ibuf_io_inst_0_bits_raw),
    .io_inst_0_bits_replay(ibuf_io_inst_0_bits_replay),
    .io_inst_0_bits_rvc(ibuf_io_inst_0_bits_rvc),
    .io_inst_0_bits_xcpt0_ae_inst(ibuf_io_inst_0_bits_xcpt0_ae_inst),
    .io_inst_0_bits_xcpt1_ae_inst(ibuf_io_inst_0_bits_xcpt1_ae_inst),
    .io_inst_0_bits_xcpt1_gf_inst(ibuf_io_inst_0_bits_xcpt1_gf_inst),
    .io_inst_0_bits_xcpt1_pf_inst(ibuf_io_inst_0_bits_xcpt1_pf_inst),
    .io_inst_0_ready(ibuf_io_inst_0_ready),
    .io_inst_0_valid(ibuf_io_inst_0_valid),
    .io_kill(ibuf_io_kill),
    .io_pc(bpu_io_pc),
    .reset(reset)
  );
  DFF_X1 \id_reg_fence$_SDFF_PP0_  (
    .CK(clock),
    .D(_00583_),
    .Q(id_reg_fence),
    .QN(_09904_)
  );
  DFF_X1 \id_reg_pause$_SDFFE_PP0N_  (
    .CK(clock),
    .D(_00582_),
    .Q(id_reg_pause),
    .QN(_09905_)
  );
  DFF_X1 \imem_might_request_reg$_DFF_P_  (
    .CK(clock),
    .D(_00005_),
    .Q(imem_might_request_reg),
    .QN(_09906_)
  );
  DFF_X1 \mem_br_taken$_DFFE_PP_  (
    .CK(clock),
    .D(_00240_),
    .Q(mem_br_taken),
    .QN(_10230_)
  );
  DFF_X1 \mem_ctrl_branch$_DFFE_PP_  (
    .CK(clock),
    .D(_00556_),
    .Q(mem_ctrl_branch),
    .QN(_09920_)
  );
  DFF_X1 \mem_ctrl_csr[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00548_),
    .Q(mem_ctrl_csr[0]),
    .QN(_09927_)
  );
  DFF_X1 \mem_ctrl_csr[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00549_),
    .Q(mem_ctrl_csr[1]),
    .QN(_09926_)
  );
  DFF_X1 \mem_ctrl_csr[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00550_),
    .Q(mem_ctrl_csr[2]),
    .QN(_09925_)
  );
  DFF_X1 \mem_ctrl_div$_DFFE_PP_  (
    .CK(clock),
    .D(_00552_),
    .Q(mem_ctrl_div),
    .QN(_09923_)
  );
  DFF_X1 \mem_ctrl_fence_i$_DFFE_PP_  (
    .CK(clock),
    .D(_00547_),
    .Q(mem_ctrl_fence_i),
    .QN(_09928_)
  );
  DFF_X1 \mem_ctrl_jal$_DFFE_PP_  (
    .CK(clock),
    .D(_00555_),
    .Q(mem_ctrl_jal),
    .QN(_09921_)
  );
  DFF_X1 \mem_ctrl_jalr$_DFFE_PP_  (
    .CK(clock),
    .D(_00554_),
    .Q(mem_ctrl_jalr),
    .QN(_09922_)
  );
  DFF_X1 \mem_ctrl_mem$_DFFE_PP_  (
    .CK(clock),
    .D(_00553_),
    .Q(mem_ctrl_mem),
    .QN(_00028_)
  );
  DFF_X1 \mem_ctrl_wxd$_DFFE_PP_  (
    .CK(clock),
    .D(_00551_),
    .Q(mem_ctrl_wxd),
    .QN(_09924_)
  );
  DFF_X1 \mem_reg_cause[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00381_),
    .Q(mem_reg_cause[0]),
    .QN(_10089_)
  );
  DFF_X1 \mem_reg_cause[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00391_),
    .Q(mem_reg_cause[10]),
    .QN(_10079_)
  );
  DFF_X1 \mem_reg_cause[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00392_),
    .Q(mem_reg_cause[11]),
    .QN(_10078_)
  );
  DFF_X1 \mem_reg_cause[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00393_),
    .Q(mem_reg_cause[12]),
    .QN(_10077_)
  );
  DFF_X1 \mem_reg_cause[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00394_),
    .Q(mem_reg_cause[13]),
    .QN(_10076_)
  );
  DFF_X1 \mem_reg_cause[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00395_),
    .Q(mem_reg_cause[14]),
    .QN(_10075_)
  );
  DFF_X1 \mem_reg_cause[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00396_),
    .Q(mem_reg_cause[15]),
    .QN(_10074_)
  );
  DFF_X1 \mem_reg_cause[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00397_),
    .Q(mem_reg_cause[16]),
    .QN(_10073_)
  );
  DFF_X1 \mem_reg_cause[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00398_),
    .Q(mem_reg_cause[17]),
    .QN(_10072_)
  );
  DFF_X1 \mem_reg_cause[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00399_),
    .Q(mem_reg_cause[18]),
    .QN(_10071_)
  );
  DFF_X1 \mem_reg_cause[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00400_),
    .Q(mem_reg_cause[19]),
    .QN(_10070_)
  );
  DFF_X1 \mem_reg_cause[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00382_),
    .Q(mem_reg_cause[1]),
    .QN(_10088_)
  );
  DFF_X1 \mem_reg_cause[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00401_),
    .Q(mem_reg_cause[20]),
    .QN(_10069_)
  );
  DFF_X1 \mem_reg_cause[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00402_),
    .Q(mem_reg_cause[21]),
    .QN(_10068_)
  );
  DFF_X1 \mem_reg_cause[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00403_),
    .Q(mem_reg_cause[22]),
    .QN(_10067_)
  );
  DFF_X1 \mem_reg_cause[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00404_),
    .Q(mem_reg_cause[23]),
    .QN(_10066_)
  );
  DFF_X1 \mem_reg_cause[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00405_),
    .Q(mem_reg_cause[24]),
    .QN(_10065_)
  );
  DFF_X1 \mem_reg_cause[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00406_),
    .Q(mem_reg_cause[25]),
    .QN(_10064_)
  );
  DFF_X1 \mem_reg_cause[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00407_),
    .Q(mem_reg_cause[26]),
    .QN(_10063_)
  );
  DFF_X1 \mem_reg_cause[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00408_),
    .Q(mem_reg_cause[27]),
    .QN(_10062_)
  );
  DFF_X1 \mem_reg_cause[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00409_),
    .Q(mem_reg_cause[28]),
    .QN(_10061_)
  );
  DFF_X1 \mem_reg_cause[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00410_),
    .Q(mem_reg_cause[29]),
    .QN(_10060_)
  );
  DFF_X1 \mem_reg_cause[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00383_),
    .Q(mem_reg_cause[2]),
    .QN(_10087_)
  );
  DFF_X1 \mem_reg_cause[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00411_),
    .Q(mem_reg_cause[30]),
    .QN(_10059_)
  );
  DFF_X1 \mem_reg_cause[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00412_),
    .Q(mem_reg_cause[31]),
    .QN(_10435_)
  );
  DFF_X1 \mem_reg_cause[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00384_),
    .Q(mem_reg_cause[3]),
    .QN(_10086_)
  );
  DFF_X1 \mem_reg_cause[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00385_),
    .Q(mem_reg_cause[4]),
    .QN(_10085_)
  );
  DFF_X1 \mem_reg_cause[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00386_),
    .Q(mem_reg_cause[5]),
    .QN(_10084_)
  );
  DFF_X1 \mem_reg_cause[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00387_),
    .Q(mem_reg_cause[6]),
    .QN(_10083_)
  );
  DFF_X1 \mem_reg_cause[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00388_),
    .Q(mem_reg_cause[7]),
    .QN(_10082_)
  );
  DFF_X1 \mem_reg_cause[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00389_),
    .Q(mem_reg_cause[8]),
    .QN(_10081_)
  );
  DFF_X1 \mem_reg_cause[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00390_),
    .Q(mem_reg_cause[9]),
    .QN(_10080_)
  );
  DFF_X1 \mem_reg_flush_pipe$_DFFE_PP_  (
    .CK(clock),
    .D(_00413_),
    .Q(mem_reg_flush_pipe),
    .QN(_10437_)
  );
  DFF_X1 \mem_reg_inst[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00324_),
    .Q(mem_reg_inst[10]),
    .QN(_10146_)
  );
  DFF_X1 \mem_reg_inst[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00325_),
    .Q(mem_reg_inst[11]),
    .QN(_10145_)
  );
  DFF_X1 \mem_reg_inst[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00326_),
    .Q(mem_reg_inst[12]),
    .QN(_10144_)
  );
  DFF_X1 \mem_reg_inst[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00327_),
    .Q(mem_reg_inst[13]),
    .QN(_10143_)
  );
  DFF_X1 \mem_reg_inst[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00328_),
    .Q(mem_reg_inst[14]),
    .QN(_10142_)
  );
  DFF_X1 \mem_reg_inst[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00329_),
    .Q(mem_reg_inst[15]),
    .QN(_10141_)
  );
  DFF_X1 \mem_reg_inst[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00330_),
    .Q(mem_reg_inst[16]),
    .QN(_10140_)
  );
  DFF_X1 \mem_reg_inst[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00331_),
    .Q(mem_reg_inst[17]),
    .QN(_10139_)
  );
  DFF_X1 \mem_reg_inst[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00332_),
    .Q(mem_reg_inst[18]),
    .QN(_10138_)
  );
  DFF_X1 \mem_reg_inst[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00333_),
    .Q(mem_reg_inst[19]),
    .QN(_10137_)
  );
  DFF_X1 \mem_reg_inst[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00334_),
    .Q(mem_reg_inst[20]),
    .QN(_10136_)
  );
  DFF_X1 \mem_reg_inst[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00335_),
    .Q(mem_reg_inst[21]),
    .QN(_10135_)
  );
  DFF_X1 \mem_reg_inst[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00336_),
    .Q(mem_reg_inst[22]),
    .QN(_10134_)
  );
  DFF_X1 \mem_reg_inst[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00337_),
    .Q(mem_reg_inst[23]),
    .QN(_10133_)
  );
  DFF_X1 \mem_reg_inst[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00338_),
    .Q(mem_reg_inst[24]),
    .QN(_10132_)
  );
  DFF_X1 \mem_reg_inst[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00339_),
    .Q(mem_reg_inst[25]),
    .QN(_10131_)
  );
  DFF_X1 \mem_reg_inst[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00340_),
    .Q(mem_reg_inst[26]),
    .QN(_10130_)
  );
  DFF_X1 \mem_reg_inst[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00341_),
    .Q(mem_reg_inst[27]),
    .QN(_10129_)
  );
  DFF_X1 \mem_reg_inst[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00342_),
    .Q(mem_reg_inst[28]),
    .QN(_10128_)
  );
  DFF_X1 \mem_reg_inst[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00343_),
    .Q(mem_reg_inst[29]),
    .QN(_10127_)
  );
  DFF_X1 \mem_reg_inst[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00344_),
    .Q(mem_reg_inst[30]),
    .QN(_10126_)
  );
  DFF_X1 \mem_reg_inst[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00345_),
    .Q(mem_reg_inst[31]),
    .QN(_10125_)
  );
  DFF_X1 \mem_reg_inst[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00321_),
    .Q(mem_reg_inst[7]),
    .QN(_10149_)
  );
  DFF_X1 \mem_reg_inst[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00322_),
    .Q(mem_reg_inst[8]),
    .QN(_10148_)
  );
  DFF_X1 \mem_reg_inst[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00323_),
    .Q(mem_reg_inst[9]),
    .QN(_10147_)
  );
  DFF_X1 \mem_reg_load$_DFFE_PP_  (
    .CK(clock),
    .D(_00379_),
    .Q(mem_reg_load),
    .QN(_10091_)
  );
  DFF_X1 \mem_reg_pc[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00346_),
    .Q(mem_reg_pc[0]),
    .QN(_10124_)
  );
  DFF_X1 \mem_reg_pc[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00356_),
    .Q(mem_reg_pc[10]),
    .QN(_10114_)
  );
  DFF_X1 \mem_reg_pc[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00357_),
    .Q(mem_reg_pc[11]),
    .QN(_10113_)
  );
  DFF_X1 \mem_reg_pc[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00358_),
    .Q(mem_reg_pc[12]),
    .QN(_10112_)
  );
  DFF_X1 \mem_reg_pc[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00359_),
    .Q(mem_reg_pc[13]),
    .QN(_10111_)
  );
  DFF_X1 \mem_reg_pc[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00360_),
    .Q(mem_reg_pc[14]),
    .QN(_10110_)
  );
  DFF_X1 \mem_reg_pc[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00361_),
    .Q(mem_reg_pc[15]),
    .QN(_10109_)
  );
  DFF_X1 \mem_reg_pc[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00362_),
    .Q(mem_reg_pc[16]),
    .QN(_10108_)
  );
  DFF_X1 \mem_reg_pc[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00363_),
    .Q(mem_reg_pc[17]),
    .QN(_10107_)
  );
  DFF_X1 \mem_reg_pc[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00364_),
    .Q(mem_reg_pc[18]),
    .QN(_10106_)
  );
  DFF_X1 \mem_reg_pc[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00365_),
    .Q(mem_reg_pc[19]),
    .QN(_10105_)
  );
  DFF_X1 \mem_reg_pc[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00347_),
    .Q(mem_reg_pc[1]),
    .QN(_10123_)
  );
  DFF_X1 \mem_reg_pc[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00366_),
    .Q(mem_reg_pc[20]),
    .QN(_10104_)
  );
  DFF_X1 \mem_reg_pc[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00367_),
    .Q(mem_reg_pc[21]),
    .QN(_10103_)
  );
  DFF_X1 \mem_reg_pc[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00368_),
    .Q(mem_reg_pc[22]),
    .QN(_10102_)
  );
  DFF_X1 \mem_reg_pc[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00369_),
    .Q(mem_reg_pc[23]),
    .QN(_10101_)
  );
  DFF_X1 \mem_reg_pc[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00370_),
    .Q(mem_reg_pc[24]),
    .QN(_10100_)
  );
  DFF_X1 \mem_reg_pc[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00371_),
    .Q(mem_reg_pc[25]),
    .QN(_10099_)
  );
  DFF_X1 \mem_reg_pc[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00372_),
    .Q(mem_reg_pc[26]),
    .QN(_10098_)
  );
  DFF_X1 \mem_reg_pc[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00373_),
    .Q(mem_reg_pc[27]),
    .QN(_10097_)
  );
  DFF_X1 \mem_reg_pc[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00374_),
    .Q(mem_reg_pc[28]),
    .QN(_10096_)
  );
  DFF_X1 \mem_reg_pc[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00375_),
    .Q(mem_reg_pc[29]),
    .QN(_10095_)
  );
  DFF_X1 \mem_reg_pc[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00348_),
    .Q(mem_reg_pc[2]),
    .QN(_10122_)
  );
  DFF_X1 \mem_reg_pc[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00376_),
    .Q(mem_reg_pc[30]),
    .QN(_10094_)
  );
  DFF_X1 \mem_reg_pc[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00377_),
    .Q(mem_reg_pc[31]),
    .QN(_10093_)
  );
  DFF_X1 \mem_reg_pc[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00349_),
    .Q(mem_reg_pc[3]),
    .QN(_10121_)
  );
  DFF_X1 \mem_reg_pc[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00350_),
    .Q(mem_reg_pc[4]),
    .QN(_10120_)
  );
  DFF_X1 \mem_reg_pc[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00351_),
    .Q(mem_reg_pc[5]),
    .QN(_10119_)
  );
  DFF_X1 \mem_reg_pc[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00352_),
    .Q(mem_reg_pc[6]),
    .QN(_10118_)
  );
  DFF_X1 \mem_reg_pc[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00353_),
    .Q(mem_reg_pc[7]),
    .QN(_10117_)
  );
  DFF_X1 \mem_reg_pc[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00354_),
    .Q(mem_reg_pc[8]),
    .QN(_10116_)
  );
  DFF_X1 \mem_reg_pc[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00355_),
    .Q(mem_reg_pc[9]),
    .QN(_10115_)
  );
  DFF_X1 \mem_reg_raw_inst[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00305_),
    .Q(mem_reg_raw_inst[0]),
    .QN(_10165_)
  );
  DFF_X1 \mem_reg_raw_inst[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00315_),
    .Q(mem_reg_raw_inst[10]),
    .QN(_10155_)
  );
  DFF_X1 \mem_reg_raw_inst[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00316_),
    .Q(mem_reg_raw_inst[11]),
    .QN(_10154_)
  );
  DFF_X1 \mem_reg_raw_inst[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00317_),
    .Q(mem_reg_raw_inst[12]),
    .QN(_10153_)
  );
  DFF_X1 \mem_reg_raw_inst[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00318_),
    .Q(mem_reg_raw_inst[13]),
    .QN(_10152_)
  );
  DFF_X1 \mem_reg_raw_inst[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00319_),
    .Q(mem_reg_raw_inst[14]),
    .QN(_10151_)
  );
  DFF_X1 \mem_reg_raw_inst[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00320_),
    .Q(mem_reg_raw_inst[15]),
    .QN(_10150_)
  );
  DFF_X1 \mem_reg_raw_inst[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00306_),
    .Q(mem_reg_raw_inst[1]),
    .QN(_10164_)
  );
  DFF_X1 \mem_reg_raw_inst[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00307_),
    .Q(mem_reg_raw_inst[2]),
    .QN(_10163_)
  );
  DFF_X1 \mem_reg_raw_inst[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00308_),
    .Q(mem_reg_raw_inst[3]),
    .QN(_10162_)
  );
  DFF_X1 \mem_reg_raw_inst[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00309_),
    .Q(mem_reg_raw_inst[4]),
    .QN(_10161_)
  );
  DFF_X1 \mem_reg_raw_inst[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00310_),
    .Q(mem_reg_raw_inst[5]),
    .QN(_10160_)
  );
  DFF_X1 \mem_reg_raw_inst[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00311_),
    .Q(mem_reg_raw_inst[6]),
    .QN(_10159_)
  );
  DFF_X1 \mem_reg_raw_inst[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00312_),
    .Q(mem_reg_raw_inst[7]),
    .QN(_10158_)
  );
  DFF_X1 \mem_reg_raw_inst[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00313_),
    .Q(mem_reg_raw_inst[8]),
    .QN(_10157_)
  );
  DFF_X1 \mem_reg_raw_inst[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00314_),
    .Q(mem_reg_raw_inst[9]),
    .QN(_10156_)
  );
  DFF_X1 \mem_reg_replay$_DFF_P_  (
    .CK(clock),
    .D(_00006_),
    .Q(mem_reg_replay),
    .QN(_10436_)
  );
  DFF_X1 \mem_reg_rs2[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00241_),
    .Q(mem_reg_rs2[0]),
    .QN(_10229_)
  );
  DFF_X1 \mem_reg_rs2[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00251_),
    .Q(mem_reg_rs2[10]),
    .QN(_10219_)
  );
  DFF_X1 \mem_reg_rs2[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00252_),
    .Q(mem_reg_rs2[11]),
    .QN(_10218_)
  );
  DFF_X1 \mem_reg_rs2[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00253_),
    .Q(mem_reg_rs2[12]),
    .QN(_10217_)
  );
  DFF_X1 \mem_reg_rs2[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00254_),
    .Q(mem_reg_rs2[13]),
    .QN(_10216_)
  );
  DFF_X1 \mem_reg_rs2[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00255_),
    .Q(mem_reg_rs2[14]),
    .QN(_10215_)
  );
  DFF_X1 \mem_reg_rs2[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00256_),
    .Q(mem_reg_rs2[15]),
    .QN(_10214_)
  );
  DFF_X1 \mem_reg_rs2[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00257_),
    .Q(mem_reg_rs2[16]),
    .QN(_10213_)
  );
  DFF_X1 \mem_reg_rs2[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00258_),
    .Q(mem_reg_rs2[17]),
    .QN(_10212_)
  );
  DFF_X1 \mem_reg_rs2[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00259_),
    .Q(mem_reg_rs2[18]),
    .QN(_10211_)
  );
  DFF_X1 \mem_reg_rs2[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00260_),
    .Q(mem_reg_rs2[19]),
    .QN(_10210_)
  );
  DFF_X1 \mem_reg_rs2[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00242_),
    .Q(mem_reg_rs2[1]),
    .QN(_10228_)
  );
  DFF_X1 \mem_reg_rs2[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00261_),
    .Q(mem_reg_rs2[20]),
    .QN(_10209_)
  );
  DFF_X1 \mem_reg_rs2[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00262_),
    .Q(mem_reg_rs2[21]),
    .QN(_10208_)
  );
  DFF_X1 \mem_reg_rs2[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00263_),
    .Q(mem_reg_rs2[22]),
    .QN(_10207_)
  );
  DFF_X1 \mem_reg_rs2[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00264_),
    .Q(mem_reg_rs2[23]),
    .QN(_10206_)
  );
  DFF_X1 \mem_reg_rs2[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00265_),
    .Q(mem_reg_rs2[24]),
    .QN(_10205_)
  );
  DFF_X1 \mem_reg_rs2[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00266_),
    .Q(mem_reg_rs2[25]),
    .QN(_10204_)
  );
  DFF_X1 \mem_reg_rs2[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00267_),
    .Q(mem_reg_rs2[26]),
    .QN(_10203_)
  );
  DFF_X1 \mem_reg_rs2[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00268_),
    .Q(mem_reg_rs2[27]),
    .QN(_10202_)
  );
  DFF_X1 \mem_reg_rs2[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00269_),
    .Q(mem_reg_rs2[28]),
    .QN(_10201_)
  );
  DFF_X1 \mem_reg_rs2[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00270_),
    .Q(mem_reg_rs2[29]),
    .QN(_10200_)
  );
  DFF_X1 \mem_reg_rs2[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00243_),
    .Q(mem_reg_rs2[2]),
    .QN(_10227_)
  );
  DFF_X1 \mem_reg_rs2[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00271_),
    .Q(mem_reg_rs2[30]),
    .QN(_10199_)
  );
  DFF_X1 \mem_reg_rs2[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00272_),
    .Q(mem_reg_rs2[31]),
    .QN(_10198_)
  );
  DFF_X1 \mem_reg_rs2[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00244_),
    .Q(mem_reg_rs2[3]),
    .QN(_10226_)
  );
  DFF_X1 \mem_reg_rs2[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00245_),
    .Q(mem_reg_rs2[4]),
    .QN(_10225_)
  );
  DFF_X1 \mem_reg_rs2[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00246_),
    .Q(mem_reg_rs2[5]),
    .QN(_10224_)
  );
  DFF_X1 \mem_reg_rs2[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00247_),
    .Q(mem_reg_rs2[6]),
    .QN(_10223_)
  );
  DFF_X1 \mem_reg_rs2[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00248_),
    .Q(mem_reg_rs2[7]),
    .QN(_10222_)
  );
  DFF_X1 \mem_reg_rs2[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00249_),
    .Q(mem_reg_rs2[8]),
    .QN(_10221_)
  );
  DFF_X1 \mem_reg_rs2[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00250_),
    .Q(mem_reg_rs2[9]),
    .QN(_10220_)
  );
  DFF_X1 \mem_reg_rvc$_DFFE_PP_  (
    .CK(clock),
    .D(_00414_),
    .Q(mem_reg_rvc),
    .QN(_mem_br_target_T_6[2])
  );
  DFF_X1 \mem_reg_slow_bypass$_DFFE_PP_  (
    .CK(clock),
    .D(_00380_),
    .Q(mem_reg_slow_bypass),
    .QN(_10090_)
  );
  DFF_X1 \mem_reg_store$_DFFE_PP_  (
    .CK(clock),
    .D(_00378_),
    .Q(mem_reg_store),
    .QN(_10092_)
  );
  DFF_X1 \mem_reg_valid$_DFF_P_  (
    .CK(clock),
    .D(_mem_reg_valid_T),
    .Q(mem_reg_valid),
    .QN(_00033_)
  );
  DFF_X1 \mem_reg_wdata[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00273_),
    .Q(mem_reg_wdata[0]),
    .QN(_10197_)
  );
  DFF_X1 \mem_reg_wdata[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00283_),
    .Q(mem_reg_wdata[10]),
    .QN(_10187_)
  );
  DFF_X1 \mem_reg_wdata[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00284_),
    .Q(mem_reg_wdata[11]),
    .QN(_10186_)
  );
  DFF_X1 \mem_reg_wdata[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00285_),
    .Q(mem_reg_wdata[12]),
    .QN(_10185_)
  );
  DFF_X1 \mem_reg_wdata[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00286_),
    .Q(mem_reg_wdata[13]),
    .QN(_10184_)
  );
  DFF_X1 \mem_reg_wdata[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00287_),
    .Q(mem_reg_wdata[14]),
    .QN(_10183_)
  );
  DFF_X1 \mem_reg_wdata[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00288_),
    .Q(mem_reg_wdata[15]),
    .QN(_10182_)
  );
  DFF_X1 \mem_reg_wdata[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00289_),
    .Q(mem_reg_wdata[16]),
    .QN(_10181_)
  );
  DFF_X1 \mem_reg_wdata[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00290_),
    .Q(mem_reg_wdata[17]),
    .QN(_10180_)
  );
  DFF_X1 \mem_reg_wdata[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00291_),
    .Q(mem_reg_wdata[18]),
    .QN(_10179_)
  );
  DFF_X1 \mem_reg_wdata[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00292_),
    .Q(mem_reg_wdata[19]),
    .QN(_10178_)
  );
  DFF_X1 \mem_reg_wdata[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00274_),
    .Q(mem_reg_wdata[1]),
    .QN(_10196_)
  );
  DFF_X1 \mem_reg_wdata[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00293_),
    .Q(mem_reg_wdata[20]),
    .QN(_10177_)
  );
  DFF_X1 \mem_reg_wdata[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00294_),
    .Q(mem_reg_wdata[21]),
    .QN(_10176_)
  );
  DFF_X1 \mem_reg_wdata[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00295_),
    .Q(mem_reg_wdata[22]),
    .QN(_10175_)
  );
  DFF_X1 \mem_reg_wdata[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00296_),
    .Q(mem_reg_wdata[23]),
    .QN(_10174_)
  );
  DFF_X1 \mem_reg_wdata[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00297_),
    .Q(mem_reg_wdata[24]),
    .QN(_10173_)
  );
  DFF_X1 \mem_reg_wdata[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00298_),
    .Q(mem_reg_wdata[25]),
    .QN(_10172_)
  );
  DFF_X1 \mem_reg_wdata[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00299_),
    .Q(mem_reg_wdata[26]),
    .QN(_10171_)
  );
  DFF_X1 \mem_reg_wdata[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00300_),
    .Q(mem_reg_wdata[27]),
    .QN(_10170_)
  );
  DFF_X1 \mem_reg_wdata[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00301_),
    .Q(mem_reg_wdata[28]),
    .QN(_10169_)
  );
  DFF_X1 \mem_reg_wdata[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00302_),
    .Q(mem_reg_wdata[29]),
    .QN(_10168_)
  );
  DFF_X1 \mem_reg_wdata[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00275_),
    .Q(mem_reg_wdata[2]),
    .QN(_10195_)
  );
  DFF_X1 \mem_reg_wdata[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00303_),
    .Q(mem_reg_wdata[30]),
    .QN(_10167_)
  );
  DFF_X1 \mem_reg_wdata[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00304_),
    .Q(mem_reg_wdata[31]),
    .QN(_10166_)
  );
  DFF_X1 \mem_reg_wdata[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00276_),
    .Q(mem_reg_wdata[3]),
    .QN(_10194_)
  );
  DFF_X1 \mem_reg_wdata[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00277_),
    .Q(mem_reg_wdata[4]),
    .QN(_10193_)
  );
  DFF_X1 \mem_reg_wdata[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00278_),
    .Q(mem_reg_wdata[5]),
    .QN(_10192_)
  );
  DFF_X1 \mem_reg_wdata[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00279_),
    .Q(mem_reg_wdata[6]),
    .QN(_10191_)
  );
  DFF_X1 \mem_reg_wdata[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00280_),
    .Q(mem_reg_wdata[7]),
    .QN(_10190_)
  );
  DFF_X1 \mem_reg_wdata[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00281_),
    .Q(mem_reg_wdata[8]),
    .QN(_10189_)
  );
  DFF_X1 \mem_reg_wdata[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00282_),
    .Q(mem_reg_wdata[9]),
    .QN(_10188_)
  );
  DFF_X1 \mem_reg_xcpt$_DFF_P_  (
    .CK(clock),
    .D(_00007_),
    .Q(mem_reg_xcpt),
    .QN(_take_pc_mem_T)
  );
  DFF_X1 \mem_reg_xcpt_interrupt$_DFF_P_  (
    .CK(clock),
    .D(_00008_),
    .Q(mem_reg_xcpt_interrupt),
    .QN(_10058_)
  );
  DFF_X1 \rf[0][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00751_),
    .Q(\rf[0] [0]),
    .QN(_09741_)
  );
  DFF_X1 \rf[0][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00761_),
    .Q(\rf[0] [10]),
    .QN(_09731_)
  );
  DFF_X1 \rf[0][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00762_),
    .Q(\rf[0] [11]),
    .QN(_09730_)
  );
  DFF_X1 \rf[0][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00763_),
    .Q(\rf[0] [12]),
    .QN(_09729_)
  );
  DFF_X1 \rf[0][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00764_),
    .Q(\rf[0] [13]),
    .QN(_09728_)
  );
  DFF_X1 \rf[0][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00765_),
    .Q(\rf[0] [14]),
    .QN(_09727_)
  );
  DFF_X1 \rf[0][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00766_),
    .Q(\rf[0] [15]),
    .QN(_09726_)
  );
  DFF_X1 \rf[0][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00767_),
    .Q(\rf[0] [16]),
    .QN(_09725_)
  );
  DFF_X1 \rf[0][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00768_),
    .Q(\rf[0] [17]),
    .QN(_09724_)
  );
  DFF_X1 \rf[0][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00769_),
    .Q(\rf[0] [18]),
    .QN(_09723_)
  );
  DFF_X1 \rf[0][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00770_),
    .Q(\rf[0] [19]),
    .QN(_09722_)
  );
  DFF_X1 \rf[0][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00752_),
    .Q(\rf[0] [1]),
    .QN(_09740_)
  );
  DFF_X1 \rf[0][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00771_),
    .Q(\rf[0] [20]),
    .QN(_09721_)
  );
  DFF_X1 \rf[0][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00772_),
    .Q(\rf[0] [21]),
    .QN(_09720_)
  );
  DFF_X1 \rf[0][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00773_),
    .Q(\rf[0] [22]),
    .QN(_09719_)
  );
  DFF_X1 \rf[0][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00774_),
    .Q(\rf[0] [23]),
    .QN(_09718_)
  );
  DFF_X1 \rf[0][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00775_),
    .Q(\rf[0] [24]),
    .QN(_09717_)
  );
  DFF_X1 \rf[0][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00776_),
    .Q(\rf[0] [25]),
    .QN(_09716_)
  );
  DFF_X1 \rf[0][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00777_),
    .Q(\rf[0] [26]),
    .QN(_09715_)
  );
  DFF_X1 \rf[0][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00778_),
    .Q(\rf[0] [27]),
    .QN(_09714_)
  );
  DFF_X1 \rf[0][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00779_),
    .Q(\rf[0] [28]),
    .QN(_09713_)
  );
  DFF_X1 \rf[0][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00780_),
    .Q(\rf[0] [29]),
    .QN(_09712_)
  );
  DFF_X1 \rf[0][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00753_),
    .Q(\rf[0] [2]),
    .QN(_09739_)
  );
  DFF_X1 \rf[0][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00781_),
    .Q(\rf[0] [30]),
    .QN(_09711_)
  );
  DFF_X1 \rf[0][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00625_),
    .Q(\rf[0] [31]),
    .QN(_09866_)
  );
  DFF_X1 \rf[0][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00754_),
    .Q(\rf[0] [3]),
    .QN(_09738_)
  );
  DFF_X1 \rf[0][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00755_),
    .Q(\rf[0] [4]),
    .QN(_09737_)
  );
  DFF_X1 \rf[0][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00756_),
    .Q(\rf[0] [5]),
    .QN(_09736_)
  );
  DFF_X1 \rf[0][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00757_),
    .Q(\rf[0] [6]),
    .QN(_09735_)
  );
  DFF_X1 \rf[0][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00758_),
    .Q(\rf[0] [7]),
    .QN(_09734_)
  );
  DFF_X1 \rf[0][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00759_),
    .Q(\rf[0] [8]),
    .QN(_09733_)
  );
  DFF_X1 \rf[0][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00760_),
    .Q(\rf[0] [9]),
    .QN(_09732_)
  );
  DFF_X1 \rf[10][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00906_),
    .Q(\rf[10] [0]),
    .QN(_09586_)
  );
  DFF_X1 \rf[10][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00916_),
    .Q(\rf[10] [10]),
    .QN(_09576_)
  );
  DFF_X1 \rf[10][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00917_),
    .Q(\rf[10] [11]),
    .QN(_09575_)
  );
  DFF_X1 \rf[10][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00918_),
    .Q(\rf[10] [12]),
    .QN(_09574_)
  );
  DFF_X1 \rf[10][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00919_),
    .Q(\rf[10] [13]),
    .QN(_09573_)
  );
  DFF_X1 \rf[10][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00920_),
    .Q(\rf[10] [14]),
    .QN(_09572_)
  );
  DFF_X1 \rf[10][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00921_),
    .Q(\rf[10] [15]),
    .QN(_09571_)
  );
  DFF_X1 \rf[10][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00922_),
    .Q(\rf[10] [16]),
    .QN(_09570_)
  );
  DFF_X1 \rf[10][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00923_),
    .Q(\rf[10] [17]),
    .QN(_09569_)
  );
  DFF_X1 \rf[10][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00924_),
    .Q(\rf[10] [18]),
    .QN(_09568_)
  );
  DFF_X1 \rf[10][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00925_),
    .Q(\rf[10] [19]),
    .QN(_09567_)
  );
  DFF_X1 \rf[10][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00907_),
    .Q(\rf[10] [1]),
    .QN(_09585_)
  );
  DFF_X1 \rf[10][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00926_),
    .Q(\rf[10] [20]),
    .QN(_09566_)
  );
  DFF_X1 \rf[10][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00927_),
    .Q(\rf[10] [21]),
    .QN(_09565_)
  );
  DFF_X1 \rf[10][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00928_),
    .Q(\rf[10] [22]),
    .QN(_09564_)
  );
  DFF_X1 \rf[10][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00929_),
    .Q(\rf[10] [23]),
    .QN(_09563_)
  );
  DFF_X1 \rf[10][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00930_),
    .Q(\rf[10] [24]),
    .QN(_09562_)
  );
  DFF_X1 \rf[10][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00931_),
    .Q(\rf[10] [25]),
    .QN(_09561_)
  );
  DFF_X1 \rf[10][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00932_),
    .Q(\rf[10] [26]),
    .QN(_09560_)
  );
  DFF_X1 \rf[10][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00933_),
    .Q(\rf[10] [27]),
    .QN(_09559_)
  );
  DFF_X1 \rf[10][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00934_),
    .Q(\rf[10] [28]),
    .QN(_09558_)
  );
  DFF_X1 \rf[10][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00935_),
    .Q(\rf[10] [29]),
    .QN(_09557_)
  );
  DFF_X1 \rf[10][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00908_),
    .Q(\rf[10] [2]),
    .QN(_09584_)
  );
  DFF_X1 \rf[10][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00936_),
    .Q(\rf[10] [30]),
    .QN(_09556_)
  );
  DFF_X1 \rf[10][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00624_),
    .Q(\rf[10] [31]),
    .QN(_09867_)
  );
  DFF_X1 \rf[10][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00909_),
    .Q(\rf[10] [3]),
    .QN(_09583_)
  );
  DFF_X1 \rf[10][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00910_),
    .Q(\rf[10] [4]),
    .QN(_09582_)
  );
  DFF_X1 \rf[10][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00911_),
    .Q(\rf[10] [5]),
    .QN(_09581_)
  );
  DFF_X1 \rf[10][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00912_),
    .Q(\rf[10] [6]),
    .QN(_09580_)
  );
  DFF_X1 \rf[10][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00913_),
    .Q(\rf[10] [7]),
    .QN(_09579_)
  );
  DFF_X1 \rf[10][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00914_),
    .Q(\rf[10] [8]),
    .QN(_09578_)
  );
  DFF_X1 \rf[10][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00915_),
    .Q(\rf[10] [9]),
    .QN(_09577_)
  );
  DFF_X1 \rf[11][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00968_),
    .Q(\rf[11] [0]),
    .QN(_09524_)
  );
  DFF_X1 \rf[11][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00978_),
    .Q(\rf[11] [10]),
    .QN(_09514_)
  );
  DFF_X1 \rf[11][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00979_),
    .Q(\rf[11] [11]),
    .QN(_09513_)
  );
  DFF_X1 \rf[11][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00980_),
    .Q(\rf[11] [12]),
    .QN(_09512_)
  );
  DFF_X1 \rf[11][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00981_),
    .Q(\rf[11] [13]),
    .QN(_09511_)
  );
  DFF_X1 \rf[11][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00982_),
    .Q(\rf[11] [14]),
    .QN(_09510_)
  );
  DFF_X1 \rf[11][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00983_),
    .Q(\rf[11] [15]),
    .QN(_09509_)
  );
  DFF_X1 \rf[11][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00984_),
    .Q(\rf[11] [16]),
    .QN(_09508_)
  );
  DFF_X1 \rf[11][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00985_),
    .Q(\rf[11] [17]),
    .QN(_09507_)
  );
  DFF_X1 \rf[11][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00986_),
    .Q(\rf[11] [18]),
    .QN(_09506_)
  );
  DFF_X1 \rf[11][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00987_),
    .Q(\rf[11] [19]),
    .QN(_09505_)
  );
  DFF_X1 \rf[11][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00969_),
    .Q(\rf[11] [1]),
    .QN(_09523_)
  );
  DFF_X1 \rf[11][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00988_),
    .Q(\rf[11] [20]),
    .QN(_09504_)
  );
  DFF_X1 \rf[11][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00989_),
    .Q(\rf[11] [21]),
    .QN(_09503_)
  );
  DFF_X1 \rf[11][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00990_),
    .Q(\rf[11] [22]),
    .QN(_09502_)
  );
  DFF_X1 \rf[11][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00991_),
    .Q(\rf[11] [23]),
    .QN(_09501_)
  );
  DFF_X1 \rf[11][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00992_),
    .Q(\rf[11] [24]),
    .QN(_09500_)
  );
  DFF_X1 \rf[11][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00993_),
    .Q(\rf[11] [25]),
    .QN(_09499_)
  );
  DFF_X1 \rf[11][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00994_),
    .Q(\rf[11] [26]),
    .QN(_09498_)
  );
  DFF_X1 \rf[11][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00995_),
    .Q(\rf[11] [27]),
    .QN(_09497_)
  );
  DFF_X1 \rf[11][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00996_),
    .Q(\rf[11] [28]),
    .QN(_09496_)
  );
  DFF_X1 \rf[11][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00997_),
    .Q(\rf[11] [29]),
    .QN(_09495_)
  );
  DFF_X1 \rf[11][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00970_),
    .Q(\rf[11] [2]),
    .QN(_09522_)
  );
  DFF_X1 \rf[11][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00998_),
    .Q(\rf[11] [30]),
    .QN(_09494_)
  );
  DFF_X1 \rf[11][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00623_),
    .Q(\rf[11] [31]),
    .QN(_09868_)
  );
  DFF_X1 \rf[11][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00971_),
    .Q(\rf[11] [3]),
    .QN(_09521_)
  );
  DFF_X1 \rf[11][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00972_),
    .Q(\rf[11] [4]),
    .QN(_09520_)
  );
  DFF_X1 \rf[11][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00973_),
    .Q(\rf[11] [5]),
    .QN(_09519_)
  );
  DFF_X1 \rf[11][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00974_),
    .Q(\rf[11] [6]),
    .QN(_09518_)
  );
  DFF_X1 \rf[11][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00975_),
    .Q(\rf[11] [7]),
    .QN(_09517_)
  );
  DFF_X1 \rf[11][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00976_),
    .Q(\rf[11] [8]),
    .QN(_09516_)
  );
  DFF_X1 \rf[11][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00977_),
    .Q(\rf[11] [9]),
    .QN(_09515_)
  );
  DFF_X1 \rf[12][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01030_),
    .Q(\rf[12] [0]),
    .QN(_09462_)
  );
  DFF_X1 \rf[12][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01040_),
    .Q(\rf[12] [10]),
    .QN(_09452_)
  );
  DFF_X1 \rf[12][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01041_),
    .Q(\rf[12] [11]),
    .QN(_09451_)
  );
  DFF_X1 \rf[12][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01042_),
    .Q(\rf[12] [12]),
    .QN(_09450_)
  );
  DFF_X1 \rf[12][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01043_),
    .Q(\rf[12] [13]),
    .QN(_09449_)
  );
  DFF_X1 \rf[12][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01044_),
    .Q(\rf[12] [14]),
    .QN(_09448_)
  );
  DFF_X1 \rf[12][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01045_),
    .Q(\rf[12] [15]),
    .QN(_09447_)
  );
  DFF_X1 \rf[12][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01046_),
    .Q(\rf[12] [16]),
    .QN(_09446_)
  );
  DFF_X1 \rf[12][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01047_),
    .Q(\rf[12] [17]),
    .QN(_09445_)
  );
  DFF_X1 \rf[12][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01048_),
    .Q(\rf[12] [18]),
    .QN(_09444_)
  );
  DFF_X1 \rf[12][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01049_),
    .Q(\rf[12] [19]),
    .QN(_09443_)
  );
  DFF_X1 \rf[12][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01031_),
    .Q(\rf[12] [1]),
    .QN(_09461_)
  );
  DFF_X1 \rf[12][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01050_),
    .Q(\rf[12] [20]),
    .QN(_09442_)
  );
  DFF_X1 \rf[12][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01051_),
    .Q(\rf[12] [21]),
    .QN(_09441_)
  );
  DFF_X1 \rf[12][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01052_),
    .Q(\rf[12] [22]),
    .QN(_09440_)
  );
  DFF_X1 \rf[12][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01053_),
    .Q(\rf[12] [23]),
    .QN(_09439_)
  );
  DFF_X1 \rf[12][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01054_),
    .Q(\rf[12] [24]),
    .QN(_09438_)
  );
  DFF_X1 \rf[12][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01055_),
    .Q(\rf[12] [25]),
    .QN(_09437_)
  );
  DFF_X1 \rf[12][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01056_),
    .Q(\rf[12] [26]),
    .QN(_09436_)
  );
  DFF_X1 \rf[12][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01057_),
    .Q(\rf[12] [27]),
    .QN(_09435_)
  );
  DFF_X1 \rf[12][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01058_),
    .Q(\rf[12] [28]),
    .QN(_09434_)
  );
  DFF_X1 \rf[12][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01059_),
    .Q(\rf[12] [29]),
    .QN(_09433_)
  );
  DFF_X1 \rf[12][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01032_),
    .Q(\rf[12] [2]),
    .QN(_09460_)
  );
  DFF_X1 \rf[12][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01060_),
    .Q(\rf[12] [30]),
    .QN(_09432_)
  );
  DFF_X1 \rf[12][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00622_),
    .Q(\rf[12] [31]),
    .QN(_09869_)
  );
  DFF_X1 \rf[12][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01033_),
    .Q(\rf[12] [3]),
    .QN(_09459_)
  );
  DFF_X1 \rf[12][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01034_),
    .Q(\rf[12] [4]),
    .QN(_09458_)
  );
  DFF_X1 \rf[12][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01035_),
    .Q(\rf[12] [5]),
    .QN(_09457_)
  );
  DFF_X1 \rf[12][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01036_),
    .Q(\rf[12] [6]),
    .QN(_09456_)
  );
  DFF_X1 \rf[12][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01037_),
    .Q(\rf[12] [7]),
    .QN(_09455_)
  );
  DFF_X1 \rf[12][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01038_),
    .Q(\rf[12] [8]),
    .QN(_09454_)
  );
  DFF_X1 \rf[12][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01039_),
    .Q(\rf[12] [9]),
    .QN(_09453_)
  );
  DFF_X1 \rf[13][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01154_),
    .Q(\rf[13] [0]),
    .QN(_09338_)
  );
  DFF_X1 \rf[13][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01164_),
    .Q(\rf[13] [10]),
    .QN(_09328_)
  );
  DFF_X1 \rf[13][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01165_),
    .Q(\rf[13] [11]),
    .QN(_09327_)
  );
  DFF_X1 \rf[13][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01166_),
    .Q(\rf[13] [12]),
    .QN(_09326_)
  );
  DFF_X1 \rf[13][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01167_),
    .Q(\rf[13] [13]),
    .QN(_09325_)
  );
  DFF_X1 \rf[13][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01168_),
    .Q(\rf[13] [14]),
    .QN(_09324_)
  );
  DFF_X1 \rf[13][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01169_),
    .Q(\rf[13] [15]),
    .QN(_09323_)
  );
  DFF_X1 \rf[13][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01170_),
    .Q(\rf[13] [16]),
    .QN(_09322_)
  );
  DFF_X1 \rf[13][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01171_),
    .Q(\rf[13] [17]),
    .QN(_09321_)
  );
  DFF_X1 \rf[13][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01172_),
    .Q(\rf[13] [18]),
    .QN(_09320_)
  );
  DFF_X1 \rf[13][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01173_),
    .Q(\rf[13] [19]),
    .QN(_09319_)
  );
  DFF_X1 \rf[13][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01155_),
    .Q(\rf[13] [1]),
    .QN(_09337_)
  );
  DFF_X1 \rf[13][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01174_),
    .Q(\rf[13] [20]),
    .QN(_09318_)
  );
  DFF_X1 \rf[13][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01175_),
    .Q(\rf[13] [21]),
    .QN(_09317_)
  );
  DFF_X1 \rf[13][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01176_),
    .Q(\rf[13] [22]),
    .QN(_09316_)
  );
  DFF_X1 \rf[13][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01177_),
    .Q(\rf[13] [23]),
    .QN(_09315_)
  );
  DFF_X1 \rf[13][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01178_),
    .Q(\rf[13] [24]),
    .QN(_09314_)
  );
  DFF_X1 \rf[13][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01179_),
    .Q(\rf[13] [25]),
    .QN(_09313_)
  );
  DFF_X1 \rf[13][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01180_),
    .Q(\rf[13] [26]),
    .QN(_09312_)
  );
  DFF_X1 \rf[13][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01181_),
    .Q(\rf[13] [27]),
    .QN(_09311_)
  );
  DFF_X1 \rf[13][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01182_),
    .Q(\rf[13] [28]),
    .QN(_09310_)
  );
  DFF_X1 \rf[13][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01183_),
    .Q(\rf[13] [29]),
    .QN(_09309_)
  );
  DFF_X1 \rf[13][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01156_),
    .Q(\rf[13] [2]),
    .QN(_09336_)
  );
  DFF_X1 \rf[13][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01184_),
    .Q(\rf[13] [30]),
    .QN(_09308_)
  );
  DFF_X1 \rf[13][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00621_),
    .Q(\rf[13] [31]),
    .QN(_09870_)
  );
  DFF_X1 \rf[13][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01157_),
    .Q(\rf[13] [3]),
    .QN(_09335_)
  );
  DFF_X1 \rf[13][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01158_),
    .Q(\rf[13] [4]),
    .QN(_09334_)
  );
  DFF_X1 \rf[13][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01159_),
    .Q(\rf[13] [5]),
    .QN(_09333_)
  );
  DFF_X1 \rf[13][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01160_),
    .Q(\rf[13] [6]),
    .QN(_09332_)
  );
  DFF_X1 \rf[13][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01161_),
    .Q(\rf[13] [7]),
    .QN(_09331_)
  );
  DFF_X1 \rf[13][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01162_),
    .Q(\rf[13] [8]),
    .QN(_09330_)
  );
  DFF_X1 \rf[13][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01163_),
    .Q(\rf[13] [9]),
    .QN(_09329_)
  );
  DFF_X1 \rf[14][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01278_),
    .Q(\rf[14] [0]),
    .QN(_09214_)
  );
  DFF_X1 \rf[14][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01288_),
    .Q(\rf[14] [10]),
    .QN(_09204_)
  );
  DFF_X1 \rf[14][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01289_),
    .Q(\rf[14] [11]),
    .QN(_09203_)
  );
  DFF_X1 \rf[14][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01290_),
    .Q(\rf[14] [12]),
    .QN(_09202_)
  );
  DFF_X1 \rf[14][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01291_),
    .Q(\rf[14] [13]),
    .QN(_09201_)
  );
  DFF_X1 \rf[14][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01292_),
    .Q(\rf[14] [14]),
    .QN(_09200_)
  );
  DFF_X1 \rf[14][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01293_),
    .Q(\rf[14] [15]),
    .QN(_09199_)
  );
  DFF_X1 \rf[14][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01294_),
    .Q(\rf[14] [16]),
    .QN(_09198_)
  );
  DFF_X1 \rf[14][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01295_),
    .Q(\rf[14] [17]),
    .QN(_09197_)
  );
  DFF_X1 \rf[14][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01296_),
    .Q(\rf[14] [18]),
    .QN(_09196_)
  );
  DFF_X1 \rf[14][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01297_),
    .Q(\rf[14] [19]),
    .QN(_09195_)
  );
  DFF_X1 \rf[14][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01279_),
    .Q(\rf[14] [1]),
    .QN(_09213_)
  );
  DFF_X1 \rf[14][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01298_),
    .Q(\rf[14] [20]),
    .QN(_09194_)
  );
  DFF_X1 \rf[14][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01299_),
    .Q(\rf[14] [21]),
    .QN(_09193_)
  );
  DFF_X1 \rf[14][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01300_),
    .Q(\rf[14] [22]),
    .QN(_09192_)
  );
  DFF_X1 \rf[14][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01301_),
    .Q(\rf[14] [23]),
    .QN(_09191_)
  );
  DFF_X1 \rf[14][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01302_),
    .Q(\rf[14] [24]),
    .QN(_09190_)
  );
  DFF_X1 \rf[14][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01303_),
    .Q(\rf[14] [25]),
    .QN(_09189_)
  );
  DFF_X1 \rf[14][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01304_),
    .Q(\rf[14] [26]),
    .QN(_09188_)
  );
  DFF_X1 \rf[14][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01305_),
    .Q(\rf[14] [27]),
    .QN(_09187_)
  );
  DFF_X1 \rf[14][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01306_),
    .Q(\rf[14] [28]),
    .QN(_09186_)
  );
  DFF_X1 \rf[14][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01307_),
    .Q(\rf[14] [29]),
    .QN(_09185_)
  );
  DFF_X1 \rf[14][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01280_),
    .Q(\rf[14] [2]),
    .QN(_09212_)
  );
  DFF_X1 \rf[14][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01308_),
    .Q(\rf[14] [30]),
    .QN(_09184_)
  );
  DFF_X1 \rf[14][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00620_),
    .Q(\rf[14] [31]),
    .QN(_09871_)
  );
  DFF_X1 \rf[14][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01281_),
    .Q(\rf[14] [3]),
    .QN(_09211_)
  );
  DFF_X1 \rf[14][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01282_),
    .Q(\rf[14] [4]),
    .QN(_09210_)
  );
  DFF_X1 \rf[14][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01283_),
    .Q(\rf[14] [5]),
    .QN(_09209_)
  );
  DFF_X1 \rf[14][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01284_),
    .Q(\rf[14] [6]),
    .QN(_09208_)
  );
  DFF_X1 \rf[14][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01285_),
    .Q(\rf[14] [7]),
    .QN(_09207_)
  );
  DFF_X1 \rf[14][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01286_),
    .Q(\rf[14] [8]),
    .QN(_09206_)
  );
  DFF_X1 \rf[14][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01287_),
    .Q(\rf[14] [9]),
    .QN(_09205_)
  );
  DFF_X1 \rf[15][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00782_),
    .Q(\rf[15] [0]),
    .QN(_09710_)
  );
  DFF_X1 \rf[15][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00792_),
    .Q(\rf[15] [10]),
    .QN(_09700_)
  );
  DFF_X1 \rf[15][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00793_),
    .Q(\rf[15] [11]),
    .QN(_09699_)
  );
  DFF_X1 \rf[15][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00794_),
    .Q(\rf[15] [12]),
    .QN(_09698_)
  );
  DFF_X1 \rf[15][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00795_),
    .Q(\rf[15] [13]),
    .QN(_09697_)
  );
  DFF_X1 \rf[15][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00796_),
    .Q(\rf[15] [14]),
    .QN(_09696_)
  );
  DFF_X1 \rf[15][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00797_),
    .Q(\rf[15] [15]),
    .QN(_09695_)
  );
  DFF_X1 \rf[15][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00798_),
    .Q(\rf[15] [16]),
    .QN(_09694_)
  );
  DFF_X1 \rf[15][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00799_),
    .Q(\rf[15] [17]),
    .QN(_09693_)
  );
  DFF_X1 \rf[15][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00800_),
    .Q(\rf[15] [18]),
    .QN(_09692_)
  );
  DFF_X1 \rf[15][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00801_),
    .Q(\rf[15] [19]),
    .QN(_09691_)
  );
  DFF_X1 \rf[15][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00783_),
    .Q(\rf[15] [1]),
    .QN(_09709_)
  );
  DFF_X1 \rf[15][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00802_),
    .Q(\rf[15] [20]),
    .QN(_09690_)
  );
  DFF_X1 \rf[15][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00803_),
    .Q(\rf[15] [21]),
    .QN(_09689_)
  );
  DFF_X1 \rf[15][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00804_),
    .Q(\rf[15] [22]),
    .QN(_09688_)
  );
  DFF_X1 \rf[15][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00805_),
    .Q(\rf[15] [23]),
    .QN(_09687_)
  );
  DFF_X1 \rf[15][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00806_),
    .Q(\rf[15] [24]),
    .QN(_09686_)
  );
  DFF_X1 \rf[15][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00807_),
    .Q(\rf[15] [25]),
    .QN(_09685_)
  );
  DFF_X1 \rf[15][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00808_),
    .Q(\rf[15] [26]),
    .QN(_09684_)
  );
  DFF_X1 \rf[15][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00809_),
    .Q(\rf[15] [27]),
    .QN(_09683_)
  );
  DFF_X1 \rf[15][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00810_),
    .Q(\rf[15] [28]),
    .QN(_09682_)
  );
  DFF_X1 \rf[15][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00811_),
    .Q(\rf[15] [29]),
    .QN(_09681_)
  );
  DFF_X1 \rf[15][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00784_),
    .Q(\rf[15] [2]),
    .QN(_09708_)
  );
  DFF_X1 \rf[15][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00812_),
    .Q(\rf[15] [30]),
    .QN(_09680_)
  );
  DFF_X1 \rf[15][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00619_),
    .Q(\rf[15] [31]),
    .QN(_09872_)
  );
  DFF_X1 \rf[15][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00785_),
    .Q(\rf[15] [3]),
    .QN(_09707_)
  );
  DFF_X1 \rf[15][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00786_),
    .Q(\rf[15] [4]),
    .QN(_09706_)
  );
  DFF_X1 \rf[15][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00787_),
    .Q(\rf[15] [5]),
    .QN(_09705_)
  );
  DFF_X1 \rf[15][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00788_),
    .Q(\rf[15] [6]),
    .QN(_09704_)
  );
  DFF_X1 \rf[15][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00789_),
    .Q(\rf[15] [7]),
    .QN(_09703_)
  );
  DFF_X1 \rf[15][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00790_),
    .Q(\rf[15] [8]),
    .QN(_09702_)
  );
  DFF_X1 \rf[15][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00791_),
    .Q(\rf[15] [9]),
    .QN(_09701_)
  );
  DFF_X1 \rf[16][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00844_),
    .Q(\rf[16] [0]),
    .QN(_09648_)
  );
  DFF_X1 \rf[16][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00854_),
    .Q(\rf[16] [10]),
    .QN(_09638_)
  );
  DFF_X1 \rf[16][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00855_),
    .Q(\rf[16] [11]),
    .QN(_09637_)
  );
  DFF_X1 \rf[16][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00856_),
    .Q(\rf[16] [12]),
    .QN(_09636_)
  );
  DFF_X1 \rf[16][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00857_),
    .Q(\rf[16] [13]),
    .QN(_09635_)
  );
  DFF_X1 \rf[16][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00858_),
    .Q(\rf[16] [14]),
    .QN(_09634_)
  );
  DFF_X1 \rf[16][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00859_),
    .Q(\rf[16] [15]),
    .QN(_09633_)
  );
  DFF_X1 \rf[16][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00860_),
    .Q(\rf[16] [16]),
    .QN(_09632_)
  );
  DFF_X1 \rf[16][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00861_),
    .Q(\rf[16] [17]),
    .QN(_09631_)
  );
  DFF_X1 \rf[16][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00862_),
    .Q(\rf[16] [18]),
    .QN(_09630_)
  );
  DFF_X1 \rf[16][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00863_),
    .Q(\rf[16] [19]),
    .QN(_09629_)
  );
  DFF_X1 \rf[16][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00845_),
    .Q(\rf[16] [1]),
    .QN(_09647_)
  );
  DFF_X1 \rf[16][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00864_),
    .Q(\rf[16] [20]),
    .QN(_09628_)
  );
  DFF_X1 \rf[16][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00865_),
    .Q(\rf[16] [21]),
    .QN(_09627_)
  );
  DFF_X1 \rf[16][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00866_),
    .Q(\rf[16] [22]),
    .QN(_09626_)
  );
  DFF_X1 \rf[16][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00867_),
    .Q(\rf[16] [23]),
    .QN(_09625_)
  );
  DFF_X1 \rf[16][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00868_),
    .Q(\rf[16] [24]),
    .QN(_09624_)
  );
  DFF_X1 \rf[16][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00869_),
    .Q(\rf[16] [25]),
    .QN(_09623_)
  );
  DFF_X1 \rf[16][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00870_),
    .Q(\rf[16] [26]),
    .QN(_09622_)
  );
  DFF_X1 \rf[16][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00871_),
    .Q(\rf[16] [27]),
    .QN(_09621_)
  );
  DFF_X1 \rf[16][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00872_),
    .Q(\rf[16] [28]),
    .QN(_09620_)
  );
  DFF_X1 \rf[16][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00873_),
    .Q(\rf[16] [29]),
    .QN(_09619_)
  );
  DFF_X1 \rf[16][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00846_),
    .Q(\rf[16] [2]),
    .QN(_09646_)
  );
  DFF_X1 \rf[16][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00874_),
    .Q(\rf[16] [30]),
    .QN(_09618_)
  );
  DFF_X1 \rf[16][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00618_),
    .Q(\rf[16] [31]),
    .QN(_09873_)
  );
  DFF_X1 \rf[16][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00847_),
    .Q(\rf[16] [3]),
    .QN(_09645_)
  );
  DFF_X1 \rf[16][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00848_),
    .Q(\rf[16] [4]),
    .QN(_09644_)
  );
  DFF_X1 \rf[16][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00849_),
    .Q(\rf[16] [5]),
    .QN(_09643_)
  );
  DFF_X1 \rf[16][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00850_),
    .Q(\rf[16] [6]),
    .QN(_09642_)
  );
  DFF_X1 \rf[16][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00851_),
    .Q(\rf[16] [7]),
    .QN(_09641_)
  );
  DFF_X1 \rf[16][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00852_),
    .Q(\rf[16] [8]),
    .QN(_09640_)
  );
  DFF_X1 \rf[16][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00853_),
    .Q(\rf[16] [9]),
    .QN(_09639_)
  );
  DFF_X1 \rf[17][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00875_),
    .Q(\rf[17] [0]),
    .QN(_09617_)
  );
  DFF_X1 \rf[17][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00885_),
    .Q(\rf[17] [10]),
    .QN(_09607_)
  );
  DFF_X1 \rf[17][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00886_),
    .Q(\rf[17] [11]),
    .QN(_09606_)
  );
  DFF_X1 \rf[17][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00887_),
    .Q(\rf[17] [12]),
    .QN(_09605_)
  );
  DFF_X1 \rf[17][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00888_),
    .Q(\rf[17] [13]),
    .QN(_09604_)
  );
  DFF_X1 \rf[17][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00889_),
    .Q(\rf[17] [14]),
    .QN(_09603_)
  );
  DFF_X1 \rf[17][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00890_),
    .Q(\rf[17] [15]),
    .QN(_09602_)
  );
  DFF_X1 \rf[17][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00891_),
    .Q(\rf[17] [16]),
    .QN(_09601_)
  );
  DFF_X1 \rf[17][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00892_),
    .Q(\rf[17] [17]),
    .QN(_09600_)
  );
  DFF_X1 \rf[17][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00893_),
    .Q(\rf[17] [18]),
    .QN(_09599_)
  );
  DFF_X1 \rf[17][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00894_),
    .Q(\rf[17] [19]),
    .QN(_09598_)
  );
  DFF_X1 \rf[17][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00876_),
    .Q(\rf[17] [1]),
    .QN(_09616_)
  );
  DFF_X1 \rf[17][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00895_),
    .Q(\rf[17] [20]),
    .QN(_09597_)
  );
  DFF_X1 \rf[17][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00896_),
    .Q(\rf[17] [21]),
    .QN(_09596_)
  );
  DFF_X1 \rf[17][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00897_),
    .Q(\rf[17] [22]),
    .QN(_09595_)
  );
  DFF_X1 \rf[17][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00898_),
    .Q(\rf[17] [23]),
    .QN(_09594_)
  );
  DFF_X1 \rf[17][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00899_),
    .Q(\rf[17] [24]),
    .QN(_09593_)
  );
  DFF_X1 \rf[17][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00900_),
    .Q(\rf[17] [25]),
    .QN(_09592_)
  );
  DFF_X1 \rf[17][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00901_),
    .Q(\rf[17] [26]),
    .QN(_09591_)
  );
  DFF_X1 \rf[17][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00902_),
    .Q(\rf[17] [27]),
    .QN(_09590_)
  );
  DFF_X1 \rf[17][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00903_),
    .Q(\rf[17] [28]),
    .QN(_09589_)
  );
  DFF_X1 \rf[17][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00904_),
    .Q(\rf[17] [29]),
    .QN(_09588_)
  );
  DFF_X1 \rf[17][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00877_),
    .Q(\rf[17] [2]),
    .QN(_09615_)
  );
  DFF_X1 \rf[17][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00905_),
    .Q(\rf[17] [30]),
    .QN(_09587_)
  );
  DFF_X1 \rf[17][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00617_),
    .Q(\rf[17] [31]),
    .QN(_09874_)
  );
  DFF_X1 \rf[17][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00878_),
    .Q(\rf[17] [3]),
    .QN(_09614_)
  );
  DFF_X1 \rf[17][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00879_),
    .Q(\rf[17] [4]),
    .QN(_09613_)
  );
  DFF_X1 \rf[17][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00880_),
    .Q(\rf[17] [5]),
    .QN(_09612_)
  );
  DFF_X1 \rf[17][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00881_),
    .Q(\rf[17] [6]),
    .QN(_09611_)
  );
  DFF_X1 \rf[17][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00882_),
    .Q(\rf[17] [7]),
    .QN(_09610_)
  );
  DFF_X1 \rf[17][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00883_),
    .Q(\rf[17] [8]),
    .QN(_09609_)
  );
  DFF_X1 \rf[17][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00884_),
    .Q(\rf[17] [9]),
    .QN(_09608_)
  );
  DFF_X1 \rf[18][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00937_),
    .Q(\rf[18] [0]),
    .QN(_09555_)
  );
  DFF_X1 \rf[18][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00947_),
    .Q(\rf[18] [10]),
    .QN(_09545_)
  );
  DFF_X1 \rf[18][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00948_),
    .Q(\rf[18] [11]),
    .QN(_09544_)
  );
  DFF_X1 \rf[18][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00949_),
    .Q(\rf[18] [12]),
    .QN(_09543_)
  );
  DFF_X1 \rf[18][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00950_),
    .Q(\rf[18] [13]),
    .QN(_09542_)
  );
  DFF_X1 \rf[18][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00951_),
    .Q(\rf[18] [14]),
    .QN(_09541_)
  );
  DFF_X1 \rf[18][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00952_),
    .Q(\rf[18] [15]),
    .QN(_09540_)
  );
  DFF_X1 \rf[18][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00953_),
    .Q(\rf[18] [16]),
    .QN(_09539_)
  );
  DFF_X1 \rf[18][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00954_),
    .Q(\rf[18] [17]),
    .QN(_09538_)
  );
  DFF_X1 \rf[18][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00955_),
    .Q(\rf[18] [18]),
    .QN(_09537_)
  );
  DFF_X1 \rf[18][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00956_),
    .Q(\rf[18] [19]),
    .QN(_09536_)
  );
  DFF_X1 \rf[18][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00938_),
    .Q(\rf[18] [1]),
    .QN(_09554_)
  );
  DFF_X1 \rf[18][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00957_),
    .Q(\rf[18] [20]),
    .QN(_09535_)
  );
  DFF_X1 \rf[18][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00958_),
    .Q(\rf[18] [21]),
    .QN(_09534_)
  );
  DFF_X1 \rf[18][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00959_),
    .Q(\rf[18] [22]),
    .QN(_09533_)
  );
  DFF_X1 \rf[18][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00960_),
    .Q(\rf[18] [23]),
    .QN(_09532_)
  );
  DFF_X1 \rf[18][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00961_),
    .Q(\rf[18] [24]),
    .QN(_09531_)
  );
  DFF_X1 \rf[18][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00962_),
    .Q(\rf[18] [25]),
    .QN(_09530_)
  );
  DFF_X1 \rf[18][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00963_),
    .Q(\rf[18] [26]),
    .QN(_09529_)
  );
  DFF_X1 \rf[18][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00964_),
    .Q(\rf[18] [27]),
    .QN(_09528_)
  );
  DFF_X1 \rf[18][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00965_),
    .Q(\rf[18] [28]),
    .QN(_09527_)
  );
  DFF_X1 \rf[18][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00966_),
    .Q(\rf[18] [29]),
    .QN(_09526_)
  );
  DFF_X1 \rf[18][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00939_),
    .Q(\rf[18] [2]),
    .QN(_09553_)
  );
  DFF_X1 \rf[18][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00967_),
    .Q(\rf[18] [30]),
    .QN(_09525_)
  );
  DFF_X1 \rf[18][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00616_),
    .Q(\rf[18] [31]),
    .QN(_09875_)
  );
  DFF_X1 \rf[18][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00940_),
    .Q(\rf[18] [3]),
    .QN(_09552_)
  );
  DFF_X1 \rf[18][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00941_),
    .Q(\rf[18] [4]),
    .QN(_09551_)
  );
  DFF_X1 \rf[18][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00942_),
    .Q(\rf[18] [5]),
    .QN(_09550_)
  );
  DFF_X1 \rf[18][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00943_),
    .Q(\rf[18] [6]),
    .QN(_09549_)
  );
  DFF_X1 \rf[18][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00944_),
    .Q(\rf[18] [7]),
    .QN(_09548_)
  );
  DFF_X1 \rf[18][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00945_),
    .Q(\rf[18] [8]),
    .QN(_09547_)
  );
  DFF_X1 \rf[18][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00946_),
    .Q(\rf[18] [9]),
    .QN(_09546_)
  );
  DFF_X1 \rf[19][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00999_),
    .Q(\rf[19] [0]),
    .QN(_09493_)
  );
  DFF_X1 \rf[19][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01009_),
    .Q(\rf[19] [10]),
    .QN(_09483_)
  );
  DFF_X1 \rf[19][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01010_),
    .Q(\rf[19] [11]),
    .QN(_09482_)
  );
  DFF_X1 \rf[19][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01011_),
    .Q(\rf[19] [12]),
    .QN(_09481_)
  );
  DFF_X1 \rf[19][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01012_),
    .Q(\rf[19] [13]),
    .QN(_09480_)
  );
  DFF_X1 \rf[19][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01013_),
    .Q(\rf[19] [14]),
    .QN(_09479_)
  );
  DFF_X1 \rf[19][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01014_),
    .Q(\rf[19] [15]),
    .QN(_09478_)
  );
  DFF_X1 \rf[19][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01015_),
    .Q(\rf[19] [16]),
    .QN(_09477_)
  );
  DFF_X1 \rf[19][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01016_),
    .Q(\rf[19] [17]),
    .QN(_09476_)
  );
  DFF_X1 \rf[19][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01017_),
    .Q(\rf[19] [18]),
    .QN(_09475_)
  );
  DFF_X1 \rf[19][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01018_),
    .Q(\rf[19] [19]),
    .QN(_09474_)
  );
  DFF_X1 \rf[19][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01000_),
    .Q(\rf[19] [1]),
    .QN(_09492_)
  );
  DFF_X1 \rf[19][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01019_),
    .Q(\rf[19] [20]),
    .QN(_09473_)
  );
  DFF_X1 \rf[19][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01020_),
    .Q(\rf[19] [21]),
    .QN(_09472_)
  );
  DFF_X1 \rf[19][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01021_),
    .Q(\rf[19] [22]),
    .QN(_09471_)
  );
  DFF_X1 \rf[19][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01022_),
    .Q(\rf[19] [23]),
    .QN(_09470_)
  );
  DFF_X1 \rf[19][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01023_),
    .Q(\rf[19] [24]),
    .QN(_09469_)
  );
  DFF_X1 \rf[19][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01024_),
    .Q(\rf[19] [25]),
    .QN(_09468_)
  );
  DFF_X1 \rf[19][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01025_),
    .Q(\rf[19] [26]),
    .QN(_09467_)
  );
  DFF_X1 \rf[19][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01026_),
    .Q(\rf[19] [27]),
    .QN(_09466_)
  );
  DFF_X1 \rf[19][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01027_),
    .Q(\rf[19] [28]),
    .QN(_09465_)
  );
  DFF_X1 \rf[19][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01028_),
    .Q(\rf[19] [29]),
    .QN(_09464_)
  );
  DFF_X1 \rf[19][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01001_),
    .Q(\rf[19] [2]),
    .QN(_09491_)
  );
  DFF_X1 \rf[19][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01029_),
    .Q(\rf[19] [30]),
    .QN(_09463_)
  );
  DFF_X1 \rf[19][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00615_),
    .Q(\rf[19] [31]),
    .QN(_09876_)
  );
  DFF_X1 \rf[19][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01002_),
    .Q(\rf[19] [3]),
    .QN(_09490_)
  );
  DFF_X1 \rf[19][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01003_),
    .Q(\rf[19] [4]),
    .QN(_09489_)
  );
  DFF_X1 \rf[19][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01004_),
    .Q(\rf[19] [5]),
    .QN(_09488_)
  );
  DFF_X1 \rf[19][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01005_),
    .Q(\rf[19] [6]),
    .QN(_09487_)
  );
  DFF_X1 \rf[19][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01006_),
    .Q(\rf[19] [7]),
    .QN(_09486_)
  );
  DFF_X1 \rf[19][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01007_),
    .Q(\rf[19] [8]),
    .QN(_09485_)
  );
  DFF_X1 \rf[19][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01008_),
    .Q(\rf[19] [9]),
    .QN(_09484_)
  );
  DFF_X1 \rf[1][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01557_),
    .Q(\rf[1] [0]),
    .QN(_08935_)
  );
  DFF_X1 \rf[1][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01567_),
    .Q(\rf[1] [10]),
    .QN(_08925_)
  );
  DFF_X1 \rf[1][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01568_),
    .Q(\rf[1] [11]),
    .QN(_08924_)
  );
  DFF_X1 \rf[1][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01569_),
    .Q(\rf[1] [12]),
    .QN(_08923_)
  );
  DFF_X1 \rf[1][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01570_),
    .Q(\rf[1] [13]),
    .QN(_08922_)
  );
  DFF_X1 \rf[1][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01571_),
    .Q(\rf[1] [14]),
    .QN(_08921_)
  );
  DFF_X1 \rf[1][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01572_),
    .Q(\rf[1] [15]),
    .QN(_08920_)
  );
  DFF_X1 \rf[1][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01573_),
    .Q(\rf[1] [16]),
    .QN(_08919_)
  );
  DFF_X1 \rf[1][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01574_),
    .Q(\rf[1] [17]),
    .QN(_08918_)
  );
  DFF_X1 \rf[1][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01575_),
    .Q(\rf[1] [18]),
    .QN(_08917_)
  );
  DFF_X1 \rf[1][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01576_),
    .Q(\rf[1] [19]),
    .QN(_08916_)
  );
  DFF_X1 \rf[1][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01558_),
    .Q(\rf[1] [1]),
    .QN(_08934_)
  );
  DFF_X1 \rf[1][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01577_),
    .Q(\rf[1] [20]),
    .QN(_08915_)
  );
  DFF_X1 \rf[1][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01578_),
    .Q(\rf[1] [21]),
    .QN(_08914_)
  );
  DFF_X1 \rf[1][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01579_),
    .Q(\rf[1] [22]),
    .QN(_08913_)
  );
  DFF_X1 \rf[1][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01580_),
    .Q(\rf[1] [23]),
    .QN(_08912_)
  );
  DFF_X1 \rf[1][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01581_),
    .Q(\rf[1] [24]),
    .QN(_08911_)
  );
  DFF_X1 \rf[1][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01582_),
    .Q(\rf[1] [25]),
    .QN(_08910_)
  );
  DFF_X1 \rf[1][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01583_),
    .Q(\rf[1] [26]),
    .QN(_08909_)
  );
  DFF_X1 \rf[1][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01584_),
    .Q(\rf[1] [27]),
    .QN(_08908_)
  );
  DFF_X1 \rf[1][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01585_),
    .Q(\rf[1] [28]),
    .QN(_08907_)
  );
  DFF_X1 \rf[1][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01586_),
    .Q(\rf[1] [29]),
    .QN(_08906_)
  );
  DFF_X1 \rf[1][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01559_),
    .Q(\rf[1] [2]),
    .QN(_08933_)
  );
  DFF_X1 \rf[1][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01587_),
    .Q(\rf[1] [30]),
    .QN(_10440_)
  );
  DFF_X1 \rf[1][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00614_),
    .Q(\rf[1] [31]),
    .QN(_09877_)
  );
  DFF_X1 \rf[1][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01560_),
    .Q(\rf[1] [3]),
    .QN(_08932_)
  );
  DFF_X1 \rf[1][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01561_),
    .Q(\rf[1] [4]),
    .QN(_08931_)
  );
  DFF_X1 \rf[1][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01562_),
    .Q(\rf[1] [5]),
    .QN(_08930_)
  );
  DFF_X1 \rf[1][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01563_),
    .Q(\rf[1] [6]),
    .QN(_08929_)
  );
  DFF_X1 \rf[1][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01564_),
    .Q(\rf[1] [7]),
    .QN(_08928_)
  );
  DFF_X1 \rf[1][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01565_),
    .Q(\rf[1] [8]),
    .QN(_08927_)
  );
  DFF_X1 \rf[1][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01566_),
    .Q(\rf[1] [9]),
    .QN(_08926_)
  );
  DFF_X1 \rf[20][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01061_),
    .Q(\rf[20] [0]),
    .QN(_09431_)
  );
  DFF_X1 \rf[20][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01071_),
    .Q(\rf[20] [10]),
    .QN(_09421_)
  );
  DFF_X1 \rf[20][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01072_),
    .Q(\rf[20] [11]),
    .QN(_09420_)
  );
  DFF_X1 \rf[20][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01073_),
    .Q(\rf[20] [12]),
    .QN(_09419_)
  );
  DFF_X1 \rf[20][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01074_),
    .Q(\rf[20] [13]),
    .QN(_09418_)
  );
  DFF_X1 \rf[20][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01075_),
    .Q(\rf[20] [14]),
    .QN(_09417_)
  );
  DFF_X1 \rf[20][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01076_),
    .Q(\rf[20] [15]),
    .QN(_09416_)
  );
  DFF_X1 \rf[20][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01077_),
    .Q(\rf[20] [16]),
    .QN(_09415_)
  );
  DFF_X1 \rf[20][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01078_),
    .Q(\rf[20] [17]),
    .QN(_09414_)
  );
  DFF_X1 \rf[20][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01079_),
    .Q(\rf[20] [18]),
    .QN(_09413_)
  );
  DFF_X1 \rf[20][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01080_),
    .Q(\rf[20] [19]),
    .QN(_09412_)
  );
  DFF_X1 \rf[20][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01062_),
    .Q(\rf[20] [1]),
    .QN(_09430_)
  );
  DFF_X1 \rf[20][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01081_),
    .Q(\rf[20] [20]),
    .QN(_09411_)
  );
  DFF_X1 \rf[20][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01082_),
    .Q(\rf[20] [21]),
    .QN(_09410_)
  );
  DFF_X1 \rf[20][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01083_),
    .Q(\rf[20] [22]),
    .QN(_09409_)
  );
  DFF_X1 \rf[20][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01084_),
    .Q(\rf[20] [23]),
    .QN(_09408_)
  );
  DFF_X1 \rf[20][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01085_),
    .Q(\rf[20] [24]),
    .QN(_09407_)
  );
  DFF_X1 \rf[20][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01086_),
    .Q(\rf[20] [25]),
    .QN(_09406_)
  );
  DFF_X1 \rf[20][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01087_),
    .Q(\rf[20] [26]),
    .QN(_09405_)
  );
  DFF_X1 \rf[20][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01088_),
    .Q(\rf[20] [27]),
    .QN(_09404_)
  );
  DFF_X1 \rf[20][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01089_),
    .Q(\rf[20] [28]),
    .QN(_09403_)
  );
  DFF_X1 \rf[20][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01090_),
    .Q(\rf[20] [29]),
    .QN(_09402_)
  );
  DFF_X1 \rf[20][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01063_),
    .Q(\rf[20] [2]),
    .QN(_09429_)
  );
  DFF_X1 \rf[20][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01091_),
    .Q(\rf[20] [30]),
    .QN(_09401_)
  );
  DFF_X1 \rf[20][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00613_),
    .Q(\rf[20] [31]),
    .QN(_09878_)
  );
  DFF_X1 \rf[20][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01064_),
    .Q(\rf[20] [3]),
    .QN(_09428_)
  );
  DFF_X1 \rf[20][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01065_),
    .Q(\rf[20] [4]),
    .QN(_09427_)
  );
  DFF_X1 \rf[20][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01066_),
    .Q(\rf[20] [5]),
    .QN(_09426_)
  );
  DFF_X1 \rf[20][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01067_),
    .Q(\rf[20] [6]),
    .QN(_09425_)
  );
  DFF_X1 \rf[20][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01068_),
    .Q(\rf[20] [7]),
    .QN(_09424_)
  );
  DFF_X1 \rf[20][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01069_),
    .Q(\rf[20] [8]),
    .QN(_09423_)
  );
  DFF_X1 \rf[20][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01070_),
    .Q(\rf[20] [9]),
    .QN(_09422_)
  );
  DFF_X1 \rf[21][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01123_),
    .Q(\rf[21] [0]),
    .QN(_09369_)
  );
  DFF_X1 \rf[21][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01133_),
    .Q(\rf[21] [10]),
    .QN(_09359_)
  );
  DFF_X1 \rf[21][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01134_),
    .Q(\rf[21] [11]),
    .QN(_09358_)
  );
  DFF_X1 \rf[21][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01135_),
    .Q(\rf[21] [12]),
    .QN(_09357_)
  );
  DFF_X1 \rf[21][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01136_),
    .Q(\rf[21] [13]),
    .QN(_09356_)
  );
  DFF_X1 \rf[21][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01137_),
    .Q(\rf[21] [14]),
    .QN(_09355_)
  );
  DFF_X1 \rf[21][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01138_),
    .Q(\rf[21] [15]),
    .QN(_09354_)
  );
  DFF_X1 \rf[21][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01139_),
    .Q(\rf[21] [16]),
    .QN(_09353_)
  );
  DFF_X1 \rf[21][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01140_),
    .Q(\rf[21] [17]),
    .QN(_09352_)
  );
  DFF_X1 \rf[21][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01141_),
    .Q(\rf[21] [18]),
    .QN(_09351_)
  );
  DFF_X1 \rf[21][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01142_),
    .Q(\rf[21] [19]),
    .QN(_09350_)
  );
  DFF_X1 \rf[21][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01124_),
    .Q(\rf[21] [1]),
    .QN(_09368_)
  );
  DFF_X1 \rf[21][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01143_),
    .Q(\rf[21] [20]),
    .QN(_09349_)
  );
  DFF_X1 \rf[21][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01144_),
    .Q(\rf[21] [21]),
    .QN(_09348_)
  );
  DFF_X1 \rf[21][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01145_),
    .Q(\rf[21] [22]),
    .QN(_09347_)
  );
  DFF_X1 \rf[21][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01146_),
    .Q(\rf[21] [23]),
    .QN(_09346_)
  );
  DFF_X1 \rf[21][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01147_),
    .Q(\rf[21] [24]),
    .QN(_09345_)
  );
  DFF_X1 \rf[21][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01148_),
    .Q(\rf[21] [25]),
    .QN(_09344_)
  );
  DFF_X1 \rf[21][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01149_),
    .Q(\rf[21] [26]),
    .QN(_09343_)
  );
  DFF_X1 \rf[21][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01150_),
    .Q(\rf[21] [27]),
    .QN(_09342_)
  );
  DFF_X1 \rf[21][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01151_),
    .Q(\rf[21] [28]),
    .QN(_09341_)
  );
  DFF_X1 \rf[21][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01152_),
    .Q(\rf[21] [29]),
    .QN(_09340_)
  );
  DFF_X1 \rf[21][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01125_),
    .Q(\rf[21] [2]),
    .QN(_09367_)
  );
  DFF_X1 \rf[21][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01153_),
    .Q(\rf[21] [30]),
    .QN(_09339_)
  );
  DFF_X1 \rf[21][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00612_),
    .Q(\rf[21] [31]),
    .QN(_09879_)
  );
  DFF_X1 \rf[21][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01126_),
    .Q(\rf[21] [3]),
    .QN(_09366_)
  );
  DFF_X1 \rf[21][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01127_),
    .Q(\rf[21] [4]),
    .QN(_09365_)
  );
  DFF_X1 \rf[21][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01128_),
    .Q(\rf[21] [5]),
    .QN(_09364_)
  );
  DFF_X1 \rf[21][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01129_),
    .Q(\rf[21] [6]),
    .QN(_09363_)
  );
  DFF_X1 \rf[21][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01130_),
    .Q(\rf[21] [7]),
    .QN(_09362_)
  );
  DFF_X1 \rf[21][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01131_),
    .Q(\rf[21] [8]),
    .QN(_09361_)
  );
  DFF_X1 \rf[21][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01132_),
    .Q(\rf[21] [9]),
    .QN(_09360_)
  );
  DFF_X1 \rf[22][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01309_),
    .Q(\rf[22] [0]),
    .QN(_09183_)
  );
  DFF_X1 \rf[22][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01319_),
    .Q(\rf[22] [10]),
    .QN(_09173_)
  );
  DFF_X1 \rf[22][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01320_),
    .Q(\rf[22] [11]),
    .QN(_09172_)
  );
  DFF_X1 \rf[22][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01321_),
    .Q(\rf[22] [12]),
    .QN(_09171_)
  );
  DFF_X1 \rf[22][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01322_),
    .Q(\rf[22] [13]),
    .QN(_09170_)
  );
  DFF_X1 \rf[22][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01323_),
    .Q(\rf[22] [14]),
    .QN(_09169_)
  );
  DFF_X1 \rf[22][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01324_),
    .Q(\rf[22] [15]),
    .QN(_09168_)
  );
  DFF_X1 \rf[22][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01325_),
    .Q(\rf[22] [16]),
    .QN(_09167_)
  );
  DFF_X1 \rf[22][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01326_),
    .Q(\rf[22] [17]),
    .QN(_09166_)
  );
  DFF_X1 \rf[22][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01327_),
    .Q(\rf[22] [18]),
    .QN(_09165_)
  );
  DFF_X1 \rf[22][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01328_),
    .Q(\rf[22] [19]),
    .QN(_09164_)
  );
  DFF_X1 \rf[22][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01310_),
    .Q(\rf[22] [1]),
    .QN(_09182_)
  );
  DFF_X1 \rf[22][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01329_),
    .Q(\rf[22] [20]),
    .QN(_09163_)
  );
  DFF_X1 \rf[22][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01330_),
    .Q(\rf[22] [21]),
    .QN(_09162_)
  );
  DFF_X1 \rf[22][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01331_),
    .Q(\rf[22] [22]),
    .QN(_09161_)
  );
  DFF_X1 \rf[22][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01332_),
    .Q(\rf[22] [23]),
    .QN(_09160_)
  );
  DFF_X1 \rf[22][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01333_),
    .Q(\rf[22] [24]),
    .QN(_09159_)
  );
  DFF_X1 \rf[22][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01334_),
    .Q(\rf[22] [25]),
    .QN(_09158_)
  );
  DFF_X1 \rf[22][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01335_),
    .Q(\rf[22] [26]),
    .QN(_09157_)
  );
  DFF_X1 \rf[22][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01336_),
    .Q(\rf[22] [27]),
    .QN(_09156_)
  );
  DFF_X1 \rf[22][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01337_),
    .Q(\rf[22] [28]),
    .QN(_09155_)
  );
  DFF_X1 \rf[22][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01338_),
    .Q(\rf[22] [29]),
    .QN(_09154_)
  );
  DFF_X1 \rf[22][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01311_),
    .Q(\rf[22] [2]),
    .QN(_09181_)
  );
  DFF_X1 \rf[22][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01339_),
    .Q(\rf[22] [30]),
    .QN(_09153_)
  );
  DFF_X1 \rf[22][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00611_),
    .Q(\rf[22] [31]),
    .QN(_09880_)
  );
  DFF_X1 \rf[22][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01312_),
    .Q(\rf[22] [3]),
    .QN(_09180_)
  );
  DFF_X1 \rf[22][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01313_),
    .Q(\rf[22] [4]),
    .QN(_09179_)
  );
  DFF_X1 \rf[22][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01314_),
    .Q(\rf[22] [5]),
    .QN(_09178_)
  );
  DFF_X1 \rf[22][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01315_),
    .Q(\rf[22] [6]),
    .QN(_09177_)
  );
  DFF_X1 \rf[22][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01316_),
    .Q(\rf[22] [7]),
    .QN(_09176_)
  );
  DFF_X1 \rf[22][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01317_),
    .Q(\rf[22] [8]),
    .QN(_09175_)
  );
  DFF_X1 \rf[22][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01318_),
    .Q(\rf[22] [9]),
    .QN(_09174_)
  );
  DFF_X1 \rf[23][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00657_),
    .Q(\rf[23] [0]),
    .QN(_09834_)
  );
  DFF_X1 \rf[23][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00667_),
    .Q(\rf[23] [10]),
    .QN(_09824_)
  );
  DFF_X1 \rf[23][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00668_),
    .Q(\rf[23] [11]),
    .QN(_09823_)
  );
  DFF_X1 \rf[23][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00669_),
    .Q(\rf[23] [12]),
    .QN(_09822_)
  );
  DFF_X1 \rf[23][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00670_),
    .Q(\rf[23] [13]),
    .QN(_09821_)
  );
  DFF_X1 \rf[23][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00671_),
    .Q(\rf[23] [14]),
    .QN(_09820_)
  );
  DFF_X1 \rf[23][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00672_),
    .Q(\rf[23] [15]),
    .QN(_09819_)
  );
  DFF_X1 \rf[23][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00673_),
    .Q(\rf[23] [16]),
    .QN(_09818_)
  );
  DFF_X1 \rf[23][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00674_),
    .Q(\rf[23] [17]),
    .QN(_09817_)
  );
  DFF_X1 \rf[23][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00675_),
    .Q(\rf[23] [18]),
    .QN(_09816_)
  );
  DFF_X1 \rf[23][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00676_),
    .Q(\rf[23] [19]),
    .QN(_09815_)
  );
  DFF_X1 \rf[23][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00658_),
    .Q(\rf[23] [1]),
    .QN(_09833_)
  );
  DFF_X1 \rf[23][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00677_),
    .Q(\rf[23] [20]),
    .QN(_09814_)
  );
  DFF_X1 \rf[23][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00678_),
    .Q(\rf[23] [21]),
    .QN(_09813_)
  );
  DFF_X1 \rf[23][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00679_),
    .Q(\rf[23] [22]),
    .QN(_09812_)
  );
  DFF_X1 \rf[23][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00680_),
    .Q(\rf[23] [23]),
    .QN(_09811_)
  );
  DFF_X1 \rf[23][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00681_),
    .Q(\rf[23] [24]),
    .QN(_09810_)
  );
  DFF_X1 \rf[23][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00682_),
    .Q(\rf[23] [25]),
    .QN(_09809_)
  );
  DFF_X1 \rf[23][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00683_),
    .Q(\rf[23] [26]),
    .QN(_09808_)
  );
  DFF_X1 \rf[23][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00684_),
    .Q(\rf[23] [27]),
    .QN(_09807_)
  );
  DFF_X1 \rf[23][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00685_),
    .Q(\rf[23] [28]),
    .QN(_09806_)
  );
  DFF_X1 \rf[23][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00686_),
    .Q(\rf[23] [29]),
    .QN(_09805_)
  );
  DFF_X1 \rf[23][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00659_),
    .Q(\rf[23] [2]),
    .QN(_09832_)
  );
  DFF_X1 \rf[23][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00687_),
    .Q(\rf[23] [30]),
    .QN(_09804_)
  );
  DFF_X1 \rf[23][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00610_),
    .Q(\rf[23] [31]),
    .QN(_09881_)
  );
  DFF_X1 \rf[23][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00660_),
    .Q(\rf[23] [3]),
    .QN(_09831_)
  );
  DFF_X1 \rf[23][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00661_),
    .Q(\rf[23] [4]),
    .QN(_09830_)
  );
  DFF_X1 \rf[23][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00662_),
    .Q(\rf[23] [5]),
    .QN(_09829_)
  );
  DFF_X1 \rf[23][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00663_),
    .Q(\rf[23] [6]),
    .QN(_09828_)
  );
  DFF_X1 \rf[23][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00664_),
    .Q(\rf[23] [7]),
    .QN(_09827_)
  );
  DFF_X1 \rf[23][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00665_),
    .Q(\rf[23] [8]),
    .QN(_09826_)
  );
  DFF_X1 \rf[23][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00666_),
    .Q(\rf[23] [9]),
    .QN(_09825_)
  );
  DFF_X1 \rf[24][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01433_),
    .Q(\rf[24] [0]),
    .QN(_09059_)
  );
  DFF_X1 \rf[24][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01443_),
    .Q(\rf[24] [10]),
    .QN(_09049_)
  );
  DFF_X1 \rf[24][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01444_),
    .Q(\rf[24] [11]),
    .QN(_09048_)
  );
  DFF_X1 \rf[24][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01445_),
    .Q(\rf[24] [12]),
    .QN(_09047_)
  );
  DFF_X1 \rf[24][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01446_),
    .Q(\rf[24] [13]),
    .QN(_09046_)
  );
  DFF_X1 \rf[24][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01447_),
    .Q(\rf[24] [14]),
    .QN(_09045_)
  );
  DFF_X1 \rf[24][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01448_),
    .Q(\rf[24] [15]),
    .QN(_09044_)
  );
  DFF_X1 \rf[24][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01449_),
    .Q(\rf[24] [16]),
    .QN(_09043_)
  );
  DFF_X1 \rf[24][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01450_),
    .Q(\rf[24] [17]),
    .QN(_09042_)
  );
  DFF_X1 \rf[24][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01451_),
    .Q(\rf[24] [18]),
    .QN(_09041_)
  );
  DFF_X1 \rf[24][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01452_),
    .Q(\rf[24] [19]),
    .QN(_09040_)
  );
  DFF_X1 \rf[24][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01434_),
    .Q(\rf[24] [1]),
    .QN(_09058_)
  );
  DFF_X1 \rf[24][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01453_),
    .Q(\rf[24] [20]),
    .QN(_09039_)
  );
  DFF_X1 \rf[24][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01454_),
    .Q(\rf[24] [21]),
    .QN(_09038_)
  );
  DFF_X1 \rf[24][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01455_),
    .Q(\rf[24] [22]),
    .QN(_09037_)
  );
  DFF_X1 \rf[24][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01456_),
    .Q(\rf[24] [23]),
    .QN(_09036_)
  );
  DFF_X1 \rf[24][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01457_),
    .Q(\rf[24] [24]),
    .QN(_09035_)
  );
  DFF_X1 \rf[24][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01458_),
    .Q(\rf[24] [25]),
    .QN(_09034_)
  );
  DFF_X1 \rf[24][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01459_),
    .Q(\rf[24] [26]),
    .QN(_09033_)
  );
  DFF_X1 \rf[24][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01460_),
    .Q(\rf[24] [27]),
    .QN(_09032_)
  );
  DFF_X1 \rf[24][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01461_),
    .Q(\rf[24] [28]),
    .QN(_09031_)
  );
  DFF_X1 \rf[24][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01462_),
    .Q(\rf[24] [29]),
    .QN(_09030_)
  );
  DFF_X1 \rf[24][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01435_),
    .Q(\rf[24] [2]),
    .QN(_09057_)
  );
  DFF_X1 \rf[24][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01463_),
    .Q(\rf[24] [30]),
    .QN(_09029_)
  );
  DFF_X1 \rf[24][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00609_),
    .Q(\rf[24] [31]),
    .QN(_09882_)
  );
  DFF_X1 \rf[24][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01436_),
    .Q(\rf[24] [3]),
    .QN(_09056_)
  );
  DFF_X1 \rf[24][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01437_),
    .Q(\rf[24] [4]),
    .QN(_09055_)
  );
  DFF_X1 \rf[24][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01438_),
    .Q(\rf[24] [5]),
    .QN(_09054_)
  );
  DFF_X1 \rf[24][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01439_),
    .Q(\rf[24] [6]),
    .QN(_09053_)
  );
  DFF_X1 \rf[24][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01440_),
    .Q(\rf[24] [7]),
    .QN(_09052_)
  );
  DFF_X1 \rf[24][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01441_),
    .Q(\rf[24] [8]),
    .QN(_09051_)
  );
  DFF_X1 \rf[24][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01442_),
    .Q(\rf[24] [9]),
    .QN(_09050_)
  );
  DFF_X1 \rf[25][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00626_),
    .Q(\rf[25] [0]),
    .QN(_09865_)
  );
  DFF_X1 \rf[25][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00636_),
    .Q(\rf[25] [10]),
    .QN(_09855_)
  );
  DFF_X1 \rf[25][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00637_),
    .Q(\rf[25] [11]),
    .QN(_09854_)
  );
  DFF_X1 \rf[25][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00638_),
    .Q(\rf[25] [12]),
    .QN(_09853_)
  );
  DFF_X1 \rf[25][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00639_),
    .Q(\rf[25] [13]),
    .QN(_09852_)
  );
  DFF_X1 \rf[25][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00640_),
    .Q(\rf[25] [14]),
    .QN(_09851_)
  );
  DFF_X1 \rf[25][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00641_),
    .Q(\rf[25] [15]),
    .QN(_09850_)
  );
  DFF_X1 \rf[25][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00642_),
    .Q(\rf[25] [16]),
    .QN(_09849_)
  );
  DFF_X1 \rf[25][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00643_),
    .Q(\rf[25] [17]),
    .QN(_09848_)
  );
  DFF_X1 \rf[25][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00644_),
    .Q(\rf[25] [18]),
    .QN(_09847_)
  );
  DFF_X1 \rf[25][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00645_),
    .Q(\rf[25] [19]),
    .QN(_09846_)
  );
  DFF_X1 \rf[25][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00627_),
    .Q(\rf[25] [1]),
    .QN(_09864_)
  );
  DFF_X1 \rf[25][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00646_),
    .Q(\rf[25] [20]),
    .QN(_09845_)
  );
  DFF_X1 \rf[25][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00647_),
    .Q(\rf[25] [21]),
    .QN(_09844_)
  );
  DFF_X1 \rf[25][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00648_),
    .Q(\rf[25] [22]),
    .QN(_09843_)
  );
  DFF_X1 \rf[25][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00649_),
    .Q(\rf[25] [23]),
    .QN(_09842_)
  );
  DFF_X1 \rf[25][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00650_),
    .Q(\rf[25] [24]),
    .QN(_09841_)
  );
  DFF_X1 \rf[25][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00651_),
    .Q(\rf[25] [25]),
    .QN(_09840_)
  );
  DFF_X1 \rf[25][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00652_),
    .Q(\rf[25] [26]),
    .QN(_09839_)
  );
  DFF_X1 \rf[25][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00653_),
    .Q(\rf[25] [27]),
    .QN(_09838_)
  );
  DFF_X1 \rf[25][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00654_),
    .Q(\rf[25] [28]),
    .QN(_09837_)
  );
  DFF_X1 \rf[25][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00655_),
    .Q(\rf[25] [29]),
    .QN(_09836_)
  );
  DFF_X1 \rf[25][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00628_),
    .Q(\rf[25] [2]),
    .QN(_09863_)
  );
  DFF_X1 \rf[25][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00656_),
    .Q(\rf[25] [30]),
    .QN(_09835_)
  );
  DFF_X1 \rf[25][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00608_),
    .Q(\rf[25] [31]),
    .QN(_09883_)
  );
  DFF_X1 \rf[25][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00629_),
    .Q(\rf[25] [3]),
    .QN(_09862_)
  );
  DFF_X1 \rf[25][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00630_),
    .Q(\rf[25] [4]),
    .QN(_09861_)
  );
  DFF_X1 \rf[25][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00631_),
    .Q(\rf[25] [5]),
    .QN(_09860_)
  );
  DFF_X1 \rf[25][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00632_),
    .Q(\rf[25] [6]),
    .QN(_09859_)
  );
  DFF_X1 \rf[25][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00633_),
    .Q(\rf[25] [7]),
    .QN(_09858_)
  );
  DFF_X1 \rf[25][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00634_),
    .Q(\rf[25] [8]),
    .QN(_09857_)
  );
  DFF_X1 \rf[25][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00635_),
    .Q(\rf[25] [9]),
    .QN(_09856_)
  );
  DFF_X1 \rf[26][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01340_),
    .Q(\rf[26] [0]),
    .QN(_09152_)
  );
  DFF_X1 \rf[26][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01350_),
    .Q(\rf[26] [10]),
    .QN(_09142_)
  );
  DFF_X1 \rf[26][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01351_),
    .Q(\rf[26] [11]),
    .QN(_09141_)
  );
  DFF_X1 \rf[26][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01352_),
    .Q(\rf[26] [12]),
    .QN(_09140_)
  );
  DFF_X1 \rf[26][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01353_),
    .Q(\rf[26] [13]),
    .QN(_09139_)
  );
  DFF_X1 \rf[26][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01354_),
    .Q(\rf[26] [14]),
    .QN(_09138_)
  );
  DFF_X1 \rf[26][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01355_),
    .Q(\rf[26] [15]),
    .QN(_09137_)
  );
  DFF_X1 \rf[26][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01356_),
    .Q(\rf[26] [16]),
    .QN(_09136_)
  );
  DFF_X1 \rf[26][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01357_),
    .Q(\rf[26] [17]),
    .QN(_09135_)
  );
  DFF_X1 \rf[26][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01358_),
    .Q(\rf[26] [18]),
    .QN(_09134_)
  );
  DFF_X1 \rf[26][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01359_),
    .Q(\rf[26] [19]),
    .QN(_09133_)
  );
  DFF_X1 \rf[26][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01341_),
    .Q(\rf[26] [1]),
    .QN(_09151_)
  );
  DFF_X1 \rf[26][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01360_),
    .Q(\rf[26] [20]),
    .QN(_09132_)
  );
  DFF_X1 \rf[26][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01361_),
    .Q(\rf[26] [21]),
    .QN(_09131_)
  );
  DFF_X1 \rf[26][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01362_),
    .Q(\rf[26] [22]),
    .QN(_09130_)
  );
  DFF_X1 \rf[26][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01363_),
    .Q(\rf[26] [23]),
    .QN(_09129_)
  );
  DFF_X1 \rf[26][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01364_),
    .Q(\rf[26] [24]),
    .QN(_09128_)
  );
  DFF_X1 \rf[26][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01365_),
    .Q(\rf[26] [25]),
    .QN(_09127_)
  );
  DFF_X1 \rf[26][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01366_),
    .Q(\rf[26] [26]),
    .QN(_09126_)
  );
  DFF_X1 \rf[26][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01367_),
    .Q(\rf[26] [27]),
    .QN(_09125_)
  );
  DFF_X1 \rf[26][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01368_),
    .Q(\rf[26] [28]),
    .QN(_09124_)
  );
  DFF_X1 \rf[26][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01369_),
    .Q(\rf[26] [29]),
    .QN(_09123_)
  );
  DFF_X1 \rf[26][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01342_),
    .Q(\rf[26] [2]),
    .QN(_09150_)
  );
  DFF_X1 \rf[26][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01370_),
    .Q(\rf[26] [30]),
    .QN(_09122_)
  );
  DFF_X1 \rf[26][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00607_),
    .Q(\rf[26] [31]),
    .QN(_09884_)
  );
  DFF_X1 \rf[26][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01343_),
    .Q(\rf[26] [3]),
    .QN(_09149_)
  );
  DFF_X1 \rf[26][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01344_),
    .Q(\rf[26] [4]),
    .QN(_09148_)
  );
  DFF_X1 \rf[26][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01345_),
    .Q(\rf[26] [5]),
    .QN(_09147_)
  );
  DFF_X1 \rf[26][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01346_),
    .Q(\rf[26] [6]),
    .QN(_09146_)
  );
  DFF_X1 \rf[26][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01347_),
    .Q(\rf[26] [7]),
    .QN(_09145_)
  );
  DFF_X1 \rf[26][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01348_),
    .Q(\rf[26] [8]),
    .QN(_09144_)
  );
  DFF_X1 \rf[26][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01349_),
    .Q(\rf[26] [9]),
    .QN(_09143_)
  );
  DFF_X1 \rf[27][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01402_),
    .Q(\rf[27] [0]),
    .QN(_09090_)
  );
  DFF_X1 \rf[27][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01412_),
    .Q(\rf[27] [10]),
    .QN(_09080_)
  );
  DFF_X1 \rf[27][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01413_),
    .Q(\rf[27] [11]),
    .QN(_09079_)
  );
  DFF_X1 \rf[27][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01414_),
    .Q(\rf[27] [12]),
    .QN(_09078_)
  );
  DFF_X1 \rf[27][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01415_),
    .Q(\rf[27] [13]),
    .QN(_09077_)
  );
  DFF_X1 \rf[27][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01416_),
    .Q(\rf[27] [14]),
    .QN(_09076_)
  );
  DFF_X1 \rf[27][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01417_),
    .Q(\rf[27] [15]),
    .QN(_09075_)
  );
  DFF_X1 \rf[27][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01418_),
    .Q(\rf[27] [16]),
    .QN(_09074_)
  );
  DFF_X1 \rf[27][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01419_),
    .Q(\rf[27] [17]),
    .QN(_09073_)
  );
  DFF_X1 \rf[27][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01420_),
    .Q(\rf[27] [18]),
    .QN(_09072_)
  );
  DFF_X1 \rf[27][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01421_),
    .Q(\rf[27] [19]),
    .QN(_09071_)
  );
  DFF_X1 \rf[27][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01403_),
    .Q(\rf[27] [1]),
    .QN(_09089_)
  );
  DFF_X1 \rf[27][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01422_),
    .Q(\rf[27] [20]),
    .QN(_09070_)
  );
  DFF_X1 \rf[27][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01423_),
    .Q(\rf[27] [21]),
    .QN(_09069_)
  );
  DFF_X1 \rf[27][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01424_),
    .Q(\rf[27] [22]),
    .QN(_09068_)
  );
  DFF_X1 \rf[27][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01425_),
    .Q(\rf[27] [23]),
    .QN(_09067_)
  );
  DFF_X1 \rf[27][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01426_),
    .Q(\rf[27] [24]),
    .QN(_09066_)
  );
  DFF_X1 \rf[27][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01427_),
    .Q(\rf[27] [25]),
    .QN(_09065_)
  );
  DFF_X1 \rf[27][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01428_),
    .Q(\rf[27] [26]),
    .QN(_09064_)
  );
  DFF_X1 \rf[27][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01429_),
    .Q(\rf[27] [27]),
    .QN(_09063_)
  );
  DFF_X1 \rf[27][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01430_),
    .Q(\rf[27] [28]),
    .QN(_09062_)
  );
  DFF_X1 \rf[27][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01431_),
    .Q(\rf[27] [29]),
    .QN(_09061_)
  );
  DFF_X1 \rf[27][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01404_),
    .Q(\rf[27] [2]),
    .QN(_09088_)
  );
  DFF_X1 \rf[27][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01432_),
    .Q(\rf[27] [30]),
    .QN(_09060_)
  );
  DFF_X1 \rf[27][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00606_),
    .Q(\rf[27] [31]),
    .QN(_09885_)
  );
  DFF_X1 \rf[27][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01405_),
    .Q(\rf[27] [3]),
    .QN(_09087_)
  );
  DFF_X1 \rf[27][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01406_),
    .Q(\rf[27] [4]),
    .QN(_09086_)
  );
  DFF_X1 \rf[27][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01407_),
    .Q(\rf[27] [5]),
    .QN(_09085_)
  );
  DFF_X1 \rf[27][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01408_),
    .Q(\rf[27] [6]),
    .QN(_09084_)
  );
  DFF_X1 \rf[27][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01409_),
    .Q(\rf[27] [7]),
    .QN(_09083_)
  );
  DFF_X1 \rf[27][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01410_),
    .Q(\rf[27] [8]),
    .QN(_09082_)
  );
  DFF_X1 \rf[27][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01411_),
    .Q(\rf[27] [9]),
    .QN(_09081_)
  );
  DFF_X1 \rf[28][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01185_),
    .Q(\rf[28] [0]),
    .QN(_09307_)
  );
  DFF_X1 \rf[28][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01195_),
    .Q(\rf[28] [10]),
    .QN(_09297_)
  );
  DFF_X1 \rf[28][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01196_),
    .Q(\rf[28] [11]),
    .QN(_09296_)
  );
  DFF_X1 \rf[28][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01197_),
    .Q(\rf[28] [12]),
    .QN(_09295_)
  );
  DFF_X1 \rf[28][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01198_),
    .Q(\rf[28] [13]),
    .QN(_09294_)
  );
  DFF_X1 \rf[28][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01199_),
    .Q(\rf[28] [14]),
    .QN(_09293_)
  );
  DFF_X1 \rf[28][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01200_),
    .Q(\rf[28] [15]),
    .QN(_09292_)
  );
  DFF_X1 \rf[28][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01201_),
    .Q(\rf[28] [16]),
    .QN(_09291_)
  );
  DFF_X1 \rf[28][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01202_),
    .Q(\rf[28] [17]),
    .QN(_09290_)
  );
  DFF_X1 \rf[28][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01203_),
    .Q(\rf[28] [18]),
    .QN(_09289_)
  );
  DFF_X1 \rf[28][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01204_),
    .Q(\rf[28] [19]),
    .QN(_09288_)
  );
  DFF_X1 \rf[28][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01186_),
    .Q(\rf[28] [1]),
    .QN(_09306_)
  );
  DFF_X1 \rf[28][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01205_),
    .Q(\rf[28] [20]),
    .QN(_09287_)
  );
  DFF_X1 \rf[28][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01206_),
    .Q(\rf[28] [21]),
    .QN(_09286_)
  );
  DFF_X1 \rf[28][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01207_),
    .Q(\rf[28] [22]),
    .QN(_09285_)
  );
  DFF_X1 \rf[28][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01208_),
    .Q(\rf[28] [23]),
    .QN(_09284_)
  );
  DFF_X1 \rf[28][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01209_),
    .Q(\rf[28] [24]),
    .QN(_09283_)
  );
  DFF_X1 \rf[28][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01210_),
    .Q(\rf[28] [25]),
    .QN(_09282_)
  );
  DFF_X1 \rf[28][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01211_),
    .Q(\rf[28] [26]),
    .QN(_09281_)
  );
  DFF_X1 \rf[28][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01212_),
    .Q(\rf[28] [27]),
    .QN(_09280_)
  );
  DFF_X1 \rf[28][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01213_),
    .Q(\rf[28] [28]),
    .QN(_09279_)
  );
  DFF_X1 \rf[28][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01214_),
    .Q(\rf[28] [29]),
    .QN(_09278_)
  );
  DFF_X1 \rf[28][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01187_),
    .Q(\rf[28] [2]),
    .QN(_09305_)
  );
  DFF_X1 \rf[28][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01215_),
    .Q(\rf[28] [30]),
    .QN(_09277_)
  );
  DFF_X1 \rf[28][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00605_),
    .Q(\rf[28] [31]),
    .QN(_09886_)
  );
  DFF_X1 \rf[28][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01188_),
    .Q(\rf[28] [3]),
    .QN(_09304_)
  );
  DFF_X1 \rf[28][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01189_),
    .Q(\rf[28] [4]),
    .QN(_09303_)
  );
  DFF_X1 \rf[28][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01190_),
    .Q(\rf[28] [5]),
    .QN(_09302_)
  );
  DFF_X1 \rf[28][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01191_),
    .Q(\rf[28] [6]),
    .QN(_09301_)
  );
  DFF_X1 \rf[28][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01192_),
    .Q(\rf[28] [7]),
    .QN(_09300_)
  );
  DFF_X1 \rf[28][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01193_),
    .Q(\rf[28] [8]),
    .QN(_09299_)
  );
  DFF_X1 \rf[28][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01194_),
    .Q(\rf[28] [9]),
    .QN(_09298_)
  );
  DFF_X1 \rf[29][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01216_),
    .Q(\rf[29] [0]),
    .QN(_09276_)
  );
  DFF_X1 \rf[29][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01226_),
    .Q(\rf[29] [10]),
    .QN(_09266_)
  );
  DFF_X1 \rf[29][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01227_),
    .Q(\rf[29] [11]),
    .QN(_09265_)
  );
  DFF_X1 \rf[29][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01228_),
    .Q(\rf[29] [12]),
    .QN(_09264_)
  );
  DFF_X1 \rf[29][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01229_),
    .Q(\rf[29] [13]),
    .QN(_09263_)
  );
  DFF_X1 \rf[29][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01230_),
    .Q(\rf[29] [14]),
    .QN(_09262_)
  );
  DFF_X1 \rf[29][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01231_),
    .Q(\rf[29] [15]),
    .QN(_09261_)
  );
  DFF_X1 \rf[29][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01232_),
    .Q(\rf[29] [16]),
    .QN(_09260_)
  );
  DFF_X1 \rf[29][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01233_),
    .Q(\rf[29] [17]),
    .QN(_09259_)
  );
  DFF_X1 \rf[29][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01234_),
    .Q(\rf[29] [18]),
    .QN(_09258_)
  );
  DFF_X1 \rf[29][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01235_),
    .Q(\rf[29] [19]),
    .QN(_09257_)
  );
  DFF_X1 \rf[29][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01217_),
    .Q(\rf[29] [1]),
    .QN(_09275_)
  );
  DFF_X1 \rf[29][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01236_),
    .Q(\rf[29] [20]),
    .QN(_09256_)
  );
  DFF_X1 \rf[29][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01237_),
    .Q(\rf[29] [21]),
    .QN(_09255_)
  );
  DFF_X1 \rf[29][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01238_),
    .Q(\rf[29] [22]),
    .QN(_09254_)
  );
  DFF_X1 \rf[29][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01239_),
    .Q(\rf[29] [23]),
    .QN(_09253_)
  );
  DFF_X1 \rf[29][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01240_),
    .Q(\rf[29] [24]),
    .QN(_09252_)
  );
  DFF_X1 \rf[29][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01241_),
    .Q(\rf[29] [25]),
    .QN(_09251_)
  );
  DFF_X1 \rf[29][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01242_),
    .Q(\rf[29] [26]),
    .QN(_09250_)
  );
  DFF_X1 \rf[29][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01243_),
    .Q(\rf[29] [27]),
    .QN(_09249_)
  );
  DFF_X1 \rf[29][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01244_),
    .Q(\rf[29] [28]),
    .QN(_09248_)
  );
  DFF_X1 \rf[29][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01245_),
    .Q(\rf[29] [29]),
    .QN(_09247_)
  );
  DFF_X1 \rf[29][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01218_),
    .Q(\rf[29] [2]),
    .QN(_09274_)
  );
  DFF_X1 \rf[29][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01246_),
    .Q(\rf[29] [30]),
    .QN(_09246_)
  );
  DFF_X1 \rf[29][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00604_),
    .Q(\rf[29] [31]),
    .QN(_09887_)
  );
  DFF_X1 \rf[29][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01219_),
    .Q(\rf[29] [3]),
    .QN(_09273_)
  );
  DFF_X1 \rf[29][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01220_),
    .Q(\rf[29] [4]),
    .QN(_09272_)
  );
  DFF_X1 \rf[29][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01221_),
    .Q(\rf[29] [5]),
    .QN(_09271_)
  );
  DFF_X1 \rf[29][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01222_),
    .Q(\rf[29] [6]),
    .QN(_09270_)
  );
  DFF_X1 \rf[29][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01223_),
    .Q(\rf[29] [7]),
    .QN(_09269_)
  );
  DFF_X1 \rf[29][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01224_),
    .Q(\rf[29] [8]),
    .QN(_09268_)
  );
  DFF_X1 \rf[29][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01225_),
    .Q(\rf[29] [9]),
    .QN(_09267_)
  );
  DFF_X1 \rf[2][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01371_),
    .Q(\rf[2] [0]),
    .QN(_09121_)
  );
  DFF_X1 \rf[2][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01381_),
    .Q(\rf[2] [10]),
    .QN(_09111_)
  );
  DFF_X1 \rf[2][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01382_),
    .Q(\rf[2] [11]),
    .QN(_09110_)
  );
  DFF_X1 \rf[2][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01383_),
    .Q(\rf[2] [12]),
    .QN(_09109_)
  );
  DFF_X1 \rf[2][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01384_),
    .Q(\rf[2] [13]),
    .QN(_09108_)
  );
  DFF_X1 \rf[2][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01385_),
    .Q(\rf[2] [14]),
    .QN(_09107_)
  );
  DFF_X1 \rf[2][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01386_),
    .Q(\rf[2] [15]),
    .QN(_09106_)
  );
  DFF_X1 \rf[2][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01387_),
    .Q(\rf[2] [16]),
    .QN(_09105_)
  );
  DFF_X1 \rf[2][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01388_),
    .Q(\rf[2] [17]),
    .QN(_09104_)
  );
  DFF_X1 \rf[2][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01389_),
    .Q(\rf[2] [18]),
    .QN(_09103_)
  );
  DFF_X1 \rf[2][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01390_),
    .Q(\rf[2] [19]),
    .QN(_09102_)
  );
  DFF_X1 \rf[2][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01372_),
    .Q(\rf[2] [1]),
    .QN(_09120_)
  );
  DFF_X1 \rf[2][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01391_),
    .Q(\rf[2] [20]),
    .QN(_09101_)
  );
  DFF_X1 \rf[2][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01392_),
    .Q(\rf[2] [21]),
    .QN(_09100_)
  );
  DFF_X1 \rf[2][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01393_),
    .Q(\rf[2] [22]),
    .QN(_09099_)
  );
  DFF_X1 \rf[2][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01394_),
    .Q(\rf[2] [23]),
    .QN(_09098_)
  );
  DFF_X1 \rf[2][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01395_),
    .Q(\rf[2] [24]),
    .QN(_09097_)
  );
  DFF_X1 \rf[2][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01396_),
    .Q(\rf[2] [25]),
    .QN(_09096_)
  );
  DFF_X1 \rf[2][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01397_),
    .Q(\rf[2] [26]),
    .QN(_09095_)
  );
  DFF_X1 \rf[2][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01398_),
    .Q(\rf[2] [27]),
    .QN(_09094_)
  );
  DFF_X1 \rf[2][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01399_),
    .Q(\rf[2] [28]),
    .QN(_09093_)
  );
  DFF_X1 \rf[2][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01400_),
    .Q(\rf[2] [29]),
    .QN(_09092_)
  );
  DFF_X1 \rf[2][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01373_),
    .Q(\rf[2] [2]),
    .QN(_09119_)
  );
  DFF_X1 \rf[2][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01401_),
    .Q(\rf[2] [30]),
    .QN(_09091_)
  );
  DFF_X1 \rf[2][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00603_),
    .Q(\rf[2] [31]),
    .QN(_09888_)
  );
  DFF_X1 \rf[2][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01374_),
    .Q(\rf[2] [3]),
    .QN(_09118_)
  );
  DFF_X1 \rf[2][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01375_),
    .Q(\rf[2] [4]),
    .QN(_09117_)
  );
  DFF_X1 \rf[2][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01376_),
    .Q(\rf[2] [5]),
    .QN(_09116_)
  );
  DFF_X1 \rf[2][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01377_),
    .Q(\rf[2] [6]),
    .QN(_09115_)
  );
  DFF_X1 \rf[2][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01378_),
    .Q(\rf[2] [7]),
    .QN(_09114_)
  );
  DFF_X1 \rf[2][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01379_),
    .Q(\rf[2] [8]),
    .QN(_09113_)
  );
  DFF_X1 \rf[2][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01380_),
    .Q(\rf[2] [9]),
    .QN(_09112_)
  );
  DFF_X1 \rf[30][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01247_),
    .Q(\rf[30] [0]),
    .QN(_09245_)
  );
  DFF_X1 \rf[30][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01257_),
    .Q(\rf[30] [10]),
    .QN(_09235_)
  );
  DFF_X1 \rf[30][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01258_),
    .Q(\rf[30] [11]),
    .QN(_09234_)
  );
  DFF_X1 \rf[30][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01259_),
    .Q(\rf[30] [12]),
    .QN(_09233_)
  );
  DFF_X1 \rf[30][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01260_),
    .Q(\rf[30] [13]),
    .QN(_09232_)
  );
  DFF_X1 \rf[30][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01261_),
    .Q(\rf[30] [14]),
    .QN(_09231_)
  );
  DFF_X1 \rf[30][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01262_),
    .Q(\rf[30] [15]),
    .QN(_09230_)
  );
  DFF_X1 \rf[30][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01263_),
    .Q(\rf[30] [16]),
    .QN(_09229_)
  );
  DFF_X1 \rf[30][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01264_),
    .Q(\rf[30] [17]),
    .QN(_09228_)
  );
  DFF_X1 \rf[30][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01265_),
    .Q(\rf[30] [18]),
    .QN(_09227_)
  );
  DFF_X1 \rf[30][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01266_),
    .Q(\rf[30] [19]),
    .QN(_09226_)
  );
  DFF_X1 \rf[30][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01248_),
    .Q(\rf[30] [1]),
    .QN(_09244_)
  );
  DFF_X1 \rf[30][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01267_),
    .Q(\rf[30] [20]),
    .QN(_09225_)
  );
  DFF_X1 \rf[30][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01268_),
    .Q(\rf[30] [21]),
    .QN(_09224_)
  );
  DFF_X1 \rf[30][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01269_),
    .Q(\rf[30] [22]),
    .QN(_09223_)
  );
  DFF_X1 \rf[30][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01270_),
    .Q(\rf[30] [23]),
    .QN(_09222_)
  );
  DFF_X1 \rf[30][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01271_),
    .Q(\rf[30] [24]),
    .QN(_09221_)
  );
  DFF_X1 \rf[30][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01272_),
    .Q(\rf[30] [25]),
    .QN(_09220_)
  );
  DFF_X1 \rf[30][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01273_),
    .Q(\rf[30] [26]),
    .QN(_09219_)
  );
  DFF_X1 \rf[30][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01274_),
    .Q(\rf[30] [27]),
    .QN(_09218_)
  );
  DFF_X1 \rf[30][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01275_),
    .Q(\rf[30] [28]),
    .QN(_09217_)
  );
  DFF_X1 \rf[30][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01276_),
    .Q(\rf[30] [29]),
    .QN(_09216_)
  );
  DFF_X1 \rf[30][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01249_),
    .Q(\rf[30] [2]),
    .QN(_09243_)
  );
  DFF_X1 \rf[30][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01277_),
    .Q(\rf[30] [30]),
    .QN(_09215_)
  );
  DFF_X1 \rf[30][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00602_),
    .Q(\rf[30] [31]),
    .QN(_09889_)
  );
  DFF_X1 \rf[30][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01250_),
    .Q(\rf[30] [3]),
    .QN(_09242_)
  );
  DFF_X1 \rf[30][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01251_),
    .Q(\rf[30] [4]),
    .QN(_09241_)
  );
  DFF_X1 \rf[30][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01252_),
    .Q(\rf[30] [5]),
    .QN(_09240_)
  );
  DFF_X1 \rf[30][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01253_),
    .Q(\rf[30] [6]),
    .QN(_09239_)
  );
  DFF_X1 \rf[30][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01254_),
    .Q(\rf[30] [7]),
    .QN(_09238_)
  );
  DFF_X1 \rf[30][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01255_),
    .Q(\rf[30] [8]),
    .QN(_09237_)
  );
  DFF_X1 \rf[30][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01256_),
    .Q(\rf[30] [9]),
    .QN(_09236_)
  );
  DFF_X1 \rf[3][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01526_),
    .Q(\rf[3] [0]),
    .QN(_08966_)
  );
  DFF_X1 \rf[3][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01536_),
    .Q(\rf[3] [10]),
    .QN(_08956_)
  );
  DFF_X1 \rf[3][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01537_),
    .Q(\rf[3] [11]),
    .QN(_08955_)
  );
  DFF_X1 \rf[3][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01538_),
    .Q(\rf[3] [12]),
    .QN(_08954_)
  );
  DFF_X1 \rf[3][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01539_),
    .Q(\rf[3] [13]),
    .QN(_08953_)
  );
  DFF_X1 \rf[3][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01540_),
    .Q(\rf[3] [14]),
    .QN(_08952_)
  );
  DFF_X1 \rf[3][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01541_),
    .Q(\rf[3] [15]),
    .QN(_08951_)
  );
  DFF_X1 \rf[3][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01542_),
    .Q(\rf[3] [16]),
    .QN(_08950_)
  );
  DFF_X1 \rf[3][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01543_),
    .Q(\rf[3] [17]),
    .QN(_08949_)
  );
  DFF_X1 \rf[3][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01544_),
    .Q(\rf[3] [18]),
    .QN(_08948_)
  );
  DFF_X1 \rf[3][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01545_),
    .Q(\rf[3] [19]),
    .QN(_08947_)
  );
  DFF_X1 \rf[3][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01527_),
    .Q(\rf[3] [1]),
    .QN(_08965_)
  );
  DFF_X1 \rf[3][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01546_),
    .Q(\rf[3] [20]),
    .QN(_08946_)
  );
  DFF_X1 \rf[3][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01547_),
    .Q(\rf[3] [21]),
    .QN(_08945_)
  );
  DFF_X1 \rf[3][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01548_),
    .Q(\rf[3] [22]),
    .QN(_08944_)
  );
  DFF_X1 \rf[3][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01549_),
    .Q(\rf[3] [23]),
    .QN(_08943_)
  );
  DFF_X1 \rf[3][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01550_),
    .Q(\rf[3] [24]),
    .QN(_08942_)
  );
  DFF_X1 \rf[3][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01551_),
    .Q(\rf[3] [25]),
    .QN(_08941_)
  );
  DFF_X1 \rf[3][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01552_),
    .Q(\rf[3] [26]),
    .QN(_08940_)
  );
  DFF_X1 \rf[3][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01553_),
    .Q(\rf[3] [27]),
    .QN(_08939_)
  );
  DFF_X1 \rf[3][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01554_),
    .Q(\rf[3] [28]),
    .QN(_08938_)
  );
  DFF_X1 \rf[3][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01555_),
    .Q(\rf[3] [29]),
    .QN(_08937_)
  );
  DFF_X1 \rf[3][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01528_),
    .Q(\rf[3] [2]),
    .QN(_08964_)
  );
  DFF_X1 \rf[3][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01556_),
    .Q(\rf[3] [30]),
    .QN(_08936_)
  );
  DFF_X1 \rf[3][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00601_),
    .Q(\rf[3] [31]),
    .QN(_09890_)
  );
  DFF_X1 \rf[3][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01529_),
    .Q(\rf[3] [3]),
    .QN(_08963_)
  );
  DFF_X1 \rf[3][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01530_),
    .Q(\rf[3] [4]),
    .QN(_08962_)
  );
  DFF_X1 \rf[3][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01531_),
    .Q(\rf[3] [5]),
    .QN(_08961_)
  );
  DFF_X1 \rf[3][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01532_),
    .Q(\rf[3] [6]),
    .QN(_08960_)
  );
  DFF_X1 \rf[3][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01533_),
    .Q(\rf[3] [7]),
    .QN(_08959_)
  );
  DFF_X1 \rf[3][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01534_),
    .Q(\rf[3] [8]),
    .QN(_08958_)
  );
  DFF_X1 \rf[3][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01535_),
    .Q(\rf[3] [9]),
    .QN(_08957_)
  );
  DFF_X1 \rf[4][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00722_),
    .Q(\rf[4] [0]),
    .QN(_09769_)
  );
  DFF_X1 \rf[4][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00732_),
    .Q(\rf[4] [10]),
    .QN(_09759_)
  );
  DFF_X1 \rf[4][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00733_),
    .Q(\rf[4] [11]),
    .QN(_09758_)
  );
  DFF_X1 \rf[4][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00734_),
    .Q(\rf[4] [12]),
    .QN(_09757_)
  );
  DFF_X1 \rf[4][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00735_),
    .Q(\rf[4] [13]),
    .QN(_09756_)
  );
  DFF_X1 \rf[4][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00736_),
    .Q(\rf[4] [14]),
    .QN(_09755_)
  );
  DFF_X1 \rf[4][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00737_),
    .Q(\rf[4] [15]),
    .QN(_09754_)
  );
  DFF_X1 \rf[4][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00738_),
    .Q(\rf[4] [16]),
    .QN(_09753_)
  );
  DFF_X1 \rf[4][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00739_),
    .Q(\rf[4] [17]),
    .QN(_09752_)
  );
  DFF_X1 \rf[4][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00740_),
    .Q(\rf[4] [18]),
    .QN(_09751_)
  );
  DFF_X1 \rf[4][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00741_),
    .Q(\rf[4] [19]),
    .QN(_09750_)
  );
  DFF_X1 \rf[4][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00723_),
    .Q(\rf[4] [1]),
    .QN(_09768_)
  );
  DFF_X1 \rf[4][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00742_),
    .Q(\rf[4] [20]),
    .QN(_09749_)
  );
  DFF_X1 \rf[4][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00743_),
    .Q(\rf[4] [21]),
    .QN(_09748_)
  );
  DFF_X1 \rf[4][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00746_),
    .Q(\rf[4] [22]),
    .QN(_09745_)
  );
  DFF_X1 \rf[4][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00744_),
    .Q(\rf[4] [23]),
    .QN(_09747_)
  );
  DFF_X1 \rf[4][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00745_),
    .Q(\rf[4] [24]),
    .QN(_09746_)
  );
  DFF_X1 \rf[4][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00748_),
    .Q(\rf[4] [25]),
    .QN(_09744_)
  );
  DFF_X1 \rf[4][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00688_),
    .Q(\rf[4] [26]),
    .QN(_09803_)
  );
  DFF_X1 \rf[4][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00749_),
    .Q(\rf[4] [27]),
    .QN(_09743_)
  );
  DFF_X1 \rf[4][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00689_),
    .Q(\rf[4] [28]),
    .QN(_09802_)
  );
  DFF_X1 \rf[4][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00750_),
    .Q(\rf[4] [29]),
    .QN(_09742_)
  );
  DFF_X1 \rf[4][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00724_),
    .Q(\rf[4] [2]),
    .QN(_09767_)
  );
  DFF_X1 \rf[4][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00690_),
    .Q(\rf[4] [30]),
    .QN(_09801_)
  );
  DFF_X1 \rf[4][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00600_),
    .Q(\rf[4] [31]),
    .QN(_09891_)
  );
  DFF_X1 \rf[4][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00725_),
    .Q(\rf[4] [3]),
    .QN(_09766_)
  );
  DFF_X1 \rf[4][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00726_),
    .Q(\rf[4] [4]),
    .QN(_09765_)
  );
  DFF_X1 \rf[4][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00727_),
    .Q(\rf[4] [5]),
    .QN(_09764_)
  );
  DFF_X1 \rf[4][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00728_),
    .Q(\rf[4] [6]),
    .QN(_09763_)
  );
  DFF_X1 \rf[4][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00729_),
    .Q(\rf[4] [7]),
    .QN(_09762_)
  );
  DFF_X1 \rf[4][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00730_),
    .Q(\rf[4] [8]),
    .QN(_09761_)
  );
  DFF_X1 \rf[4][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00731_),
    .Q(\rf[4] [9]),
    .QN(_09760_)
  );
  DFF_X1 \rf[5][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01464_),
    .Q(\rf[5] [0]),
    .QN(_09028_)
  );
  DFF_X1 \rf[5][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01474_),
    .Q(\rf[5] [10]),
    .QN(_09018_)
  );
  DFF_X1 \rf[5][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01475_),
    .Q(\rf[5] [11]),
    .QN(_09017_)
  );
  DFF_X1 \rf[5][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01476_),
    .Q(\rf[5] [12]),
    .QN(_09016_)
  );
  DFF_X1 \rf[5][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01477_),
    .Q(\rf[5] [13]),
    .QN(_09015_)
  );
  DFF_X1 \rf[5][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01478_),
    .Q(\rf[5] [14]),
    .QN(_09014_)
  );
  DFF_X1 \rf[5][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01479_),
    .Q(\rf[5] [15]),
    .QN(_09013_)
  );
  DFF_X1 \rf[5][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01480_),
    .Q(\rf[5] [16]),
    .QN(_09012_)
  );
  DFF_X1 \rf[5][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01481_),
    .Q(\rf[5] [17]),
    .QN(_09011_)
  );
  DFF_X1 \rf[5][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01482_),
    .Q(\rf[5] [18]),
    .QN(_09010_)
  );
  DFF_X1 \rf[5][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01483_),
    .Q(\rf[5] [19]),
    .QN(_09009_)
  );
  DFF_X1 \rf[5][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01465_),
    .Q(\rf[5] [1]),
    .QN(_09027_)
  );
  DFF_X1 \rf[5][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01484_),
    .Q(\rf[5] [20]),
    .QN(_09008_)
  );
  DFF_X1 \rf[5][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01485_),
    .Q(\rf[5] [21]),
    .QN(_09007_)
  );
  DFF_X1 \rf[5][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01486_),
    .Q(\rf[5] [22]),
    .QN(_09006_)
  );
  DFF_X1 \rf[5][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01487_),
    .Q(\rf[5] [23]),
    .QN(_09005_)
  );
  DFF_X1 \rf[5][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01488_),
    .Q(\rf[5] [24]),
    .QN(_09004_)
  );
  DFF_X1 \rf[5][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01489_),
    .Q(\rf[5] [25]),
    .QN(_09003_)
  );
  DFF_X1 \rf[5][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01490_),
    .Q(\rf[5] [26]),
    .QN(_09002_)
  );
  DFF_X1 \rf[5][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01491_),
    .Q(\rf[5] [27]),
    .QN(_09001_)
  );
  DFF_X1 \rf[5][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01492_),
    .Q(\rf[5] [28]),
    .QN(_09000_)
  );
  DFF_X1 \rf[5][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01493_),
    .Q(\rf[5] [29]),
    .QN(_08999_)
  );
  DFF_X1 \rf[5][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01466_),
    .Q(\rf[5] [2]),
    .QN(_09026_)
  );
  DFF_X1 \rf[5][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01494_),
    .Q(\rf[5] [30]),
    .QN(_08998_)
  );
  DFF_X1 \rf[5][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00599_),
    .Q(\rf[5] [31]),
    .QN(_09892_)
  );
  DFF_X1 \rf[5][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01467_),
    .Q(\rf[5] [3]),
    .QN(_09025_)
  );
  DFF_X1 \rf[5][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01468_),
    .Q(\rf[5] [4]),
    .QN(_09024_)
  );
  DFF_X1 \rf[5][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01469_),
    .Q(\rf[5] [5]),
    .QN(_09023_)
  );
  DFF_X1 \rf[5][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01470_),
    .Q(\rf[5] [6]),
    .QN(_09022_)
  );
  DFF_X1 \rf[5][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01471_),
    .Q(\rf[5] [7]),
    .QN(_09021_)
  );
  DFF_X1 \rf[5][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01472_),
    .Q(\rf[5] [8]),
    .QN(_09020_)
  );
  DFF_X1 \rf[5][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01473_),
    .Q(\rf[5] [9]),
    .QN(_09019_)
  );
  DFF_X1 \rf[6][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00691_),
    .Q(\rf[6] [0]),
    .QN(_09800_)
  );
  DFF_X1 \rf[6][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00701_),
    .Q(\rf[6] [10]),
    .QN(_09790_)
  );
  DFF_X1 \rf[6][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00702_),
    .Q(\rf[6] [11]),
    .QN(_09789_)
  );
  DFF_X1 \rf[6][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00703_),
    .Q(\rf[6] [12]),
    .QN(_09788_)
  );
  DFF_X1 \rf[6][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00704_),
    .Q(\rf[6] [13]),
    .QN(_09787_)
  );
  DFF_X1 \rf[6][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00705_),
    .Q(\rf[6] [14]),
    .QN(_09786_)
  );
  DFF_X1 \rf[6][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00706_),
    .Q(\rf[6] [15]),
    .QN(_09785_)
  );
  DFF_X1 \rf[6][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00707_),
    .Q(\rf[6] [16]),
    .QN(_09784_)
  );
  DFF_X1 \rf[6][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00708_),
    .Q(\rf[6] [17]),
    .QN(_09783_)
  );
  DFF_X1 \rf[6][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00709_),
    .Q(\rf[6] [18]),
    .QN(_09782_)
  );
  DFF_X1 \rf[6][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00710_),
    .Q(\rf[6] [19]),
    .QN(_09781_)
  );
  DFF_X1 \rf[6][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00692_),
    .Q(\rf[6] [1]),
    .QN(_09799_)
  );
  DFF_X1 \rf[6][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00711_),
    .Q(\rf[6] [20]),
    .QN(_09780_)
  );
  DFF_X1 \rf[6][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00712_),
    .Q(\rf[6] [21]),
    .QN(_09779_)
  );
  DFF_X1 \rf[6][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00713_),
    .Q(\rf[6] [22]),
    .QN(_09778_)
  );
  DFF_X1 \rf[6][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00714_),
    .Q(\rf[6] [23]),
    .QN(_09777_)
  );
  DFF_X1 \rf[6][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00715_),
    .Q(\rf[6] [24]),
    .QN(_09776_)
  );
  DFF_X1 \rf[6][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00716_),
    .Q(\rf[6] [25]),
    .QN(_09775_)
  );
  DFF_X1 \rf[6][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00717_),
    .Q(\rf[6] [26]),
    .QN(_09774_)
  );
  DFF_X1 \rf[6][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00718_),
    .Q(\rf[6] [27]),
    .QN(_09773_)
  );
  DFF_X1 \rf[6][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00719_),
    .Q(\rf[6] [28]),
    .QN(_09772_)
  );
  DFF_X1 \rf[6][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00720_),
    .Q(\rf[6] [29]),
    .QN(_09771_)
  );
  DFF_X1 \rf[6][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00693_),
    .Q(\rf[6] [2]),
    .QN(_09798_)
  );
  DFF_X1 \rf[6][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00721_),
    .Q(\rf[6] [30]),
    .QN(_09770_)
  );
  DFF_X1 \rf[6][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00598_),
    .Q(\rf[6] [31]),
    .QN(_09893_)
  );
  DFF_X1 \rf[6][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00694_),
    .Q(\rf[6] [3]),
    .QN(_09797_)
  );
  DFF_X1 \rf[6][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00695_),
    .Q(\rf[6] [4]),
    .QN(_09796_)
  );
  DFF_X1 \rf[6][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00696_),
    .Q(\rf[6] [5]),
    .QN(_09795_)
  );
  DFF_X1 \rf[6][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00697_),
    .Q(\rf[6] [6]),
    .QN(_09794_)
  );
  DFF_X1 \rf[6][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00698_),
    .Q(\rf[6] [7]),
    .QN(_09793_)
  );
  DFF_X1 \rf[6][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00699_),
    .Q(\rf[6] [8]),
    .QN(_09792_)
  );
  DFF_X1 \rf[6][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00700_),
    .Q(\rf[6] [9]),
    .QN(_09791_)
  );
  DFF_X1 \rf[7][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01495_),
    .Q(\rf[7] [0]),
    .QN(_08997_)
  );
  DFF_X1 \rf[7][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01505_),
    .Q(\rf[7] [10]),
    .QN(_08987_)
  );
  DFF_X1 \rf[7][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01506_),
    .Q(\rf[7] [11]),
    .QN(_08986_)
  );
  DFF_X1 \rf[7][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01507_),
    .Q(\rf[7] [12]),
    .QN(_08985_)
  );
  DFF_X1 \rf[7][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01508_),
    .Q(\rf[7] [13]),
    .QN(_08984_)
  );
  DFF_X1 \rf[7][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01509_),
    .Q(\rf[7] [14]),
    .QN(_08983_)
  );
  DFF_X1 \rf[7][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01510_),
    .Q(\rf[7] [15]),
    .QN(_08982_)
  );
  DFF_X1 \rf[7][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01511_),
    .Q(\rf[7] [16]),
    .QN(_08981_)
  );
  DFF_X1 \rf[7][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01512_),
    .Q(\rf[7] [17]),
    .QN(_08980_)
  );
  DFF_X1 \rf[7][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01513_),
    .Q(\rf[7] [18]),
    .QN(_08979_)
  );
  DFF_X1 \rf[7][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01514_),
    .Q(\rf[7] [19]),
    .QN(_08978_)
  );
  DFF_X1 \rf[7][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01496_),
    .Q(\rf[7] [1]),
    .QN(_08996_)
  );
  DFF_X1 \rf[7][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01515_),
    .Q(\rf[7] [20]),
    .QN(_08977_)
  );
  DFF_X1 \rf[7][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01516_),
    .Q(\rf[7] [21]),
    .QN(_08976_)
  );
  DFF_X1 \rf[7][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01517_),
    .Q(\rf[7] [22]),
    .QN(_08975_)
  );
  DFF_X1 \rf[7][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01518_),
    .Q(\rf[7] [23]),
    .QN(_08974_)
  );
  DFF_X1 \rf[7][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01519_),
    .Q(\rf[7] [24]),
    .QN(_08973_)
  );
  DFF_X1 \rf[7][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01520_),
    .Q(\rf[7] [25]),
    .QN(_08972_)
  );
  DFF_X1 \rf[7][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01521_),
    .Q(\rf[7] [26]),
    .QN(_08971_)
  );
  DFF_X1 \rf[7][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01522_),
    .Q(\rf[7] [27]),
    .QN(_08970_)
  );
  DFF_X1 \rf[7][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01523_),
    .Q(\rf[7] [28]),
    .QN(_08969_)
  );
  DFF_X1 \rf[7][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01524_),
    .Q(\rf[7] [29]),
    .QN(_08968_)
  );
  DFF_X1 \rf[7][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01497_),
    .Q(\rf[7] [2]),
    .QN(_08995_)
  );
  DFF_X1 \rf[7][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01525_),
    .Q(\rf[7] [30]),
    .QN(_08967_)
  );
  DFF_X1 \rf[7][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00597_),
    .Q(\rf[7] [31]),
    .QN(_09894_)
  );
  DFF_X1 \rf[7][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01498_),
    .Q(\rf[7] [3]),
    .QN(_08994_)
  );
  DFF_X1 \rf[7][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01499_),
    .Q(\rf[7] [4]),
    .QN(_08993_)
  );
  DFF_X1 \rf[7][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01500_),
    .Q(\rf[7] [5]),
    .QN(_08992_)
  );
  DFF_X1 \rf[7][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01501_),
    .Q(\rf[7] [6]),
    .QN(_08991_)
  );
  DFF_X1 \rf[7][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01502_),
    .Q(\rf[7] [7]),
    .QN(_08990_)
  );
  DFF_X1 \rf[7][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01503_),
    .Q(\rf[7] [8]),
    .QN(_08989_)
  );
  DFF_X1 \rf[7][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01504_),
    .Q(\rf[7] [9]),
    .QN(_08988_)
  );
  DFF_X1 \rf[8][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00813_),
    .Q(\rf[8] [0]),
    .QN(_09679_)
  );
  DFF_X1 \rf[8][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00823_),
    .Q(\rf[8] [10]),
    .QN(_09669_)
  );
  DFF_X1 \rf[8][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00824_),
    .Q(\rf[8] [11]),
    .QN(_09668_)
  );
  DFF_X1 \rf[8][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00825_),
    .Q(\rf[8] [12]),
    .QN(_09667_)
  );
  DFF_X1 \rf[8][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00826_),
    .Q(\rf[8] [13]),
    .QN(_09666_)
  );
  DFF_X1 \rf[8][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00827_),
    .Q(\rf[8] [14]),
    .QN(_09665_)
  );
  DFF_X1 \rf[8][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00828_),
    .Q(\rf[8] [15]),
    .QN(_09664_)
  );
  DFF_X1 \rf[8][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00829_),
    .Q(\rf[8] [16]),
    .QN(_09663_)
  );
  DFF_X1 \rf[8][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00830_),
    .Q(\rf[8] [17]),
    .QN(_09662_)
  );
  DFF_X1 \rf[8][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00831_),
    .Q(\rf[8] [18]),
    .QN(_09661_)
  );
  DFF_X1 \rf[8][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00832_),
    .Q(\rf[8] [19]),
    .QN(_09660_)
  );
  DFF_X1 \rf[8][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00814_),
    .Q(\rf[8] [1]),
    .QN(_09678_)
  );
  DFF_X1 \rf[8][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00833_),
    .Q(\rf[8] [20]),
    .QN(_09659_)
  );
  DFF_X1 \rf[8][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00834_),
    .Q(\rf[8] [21]),
    .QN(_09658_)
  );
  DFF_X1 \rf[8][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00835_),
    .Q(\rf[8] [22]),
    .QN(_09657_)
  );
  DFF_X1 \rf[8][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00836_),
    .Q(\rf[8] [23]),
    .QN(_09656_)
  );
  DFF_X1 \rf[8][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00837_),
    .Q(\rf[8] [24]),
    .QN(_09655_)
  );
  DFF_X1 \rf[8][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00838_),
    .Q(\rf[8] [25]),
    .QN(_09654_)
  );
  DFF_X1 \rf[8][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00839_),
    .Q(\rf[8] [26]),
    .QN(_09653_)
  );
  DFF_X1 \rf[8][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00840_),
    .Q(\rf[8] [27]),
    .QN(_09652_)
  );
  DFF_X1 \rf[8][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00841_),
    .Q(\rf[8] [28]),
    .QN(_09651_)
  );
  DFF_X1 \rf[8][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00842_),
    .Q(\rf[8] [29]),
    .QN(_09650_)
  );
  DFF_X1 \rf[8][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00815_),
    .Q(\rf[8] [2]),
    .QN(_09677_)
  );
  DFF_X1 \rf[8][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00843_),
    .Q(\rf[8] [30]),
    .QN(_09649_)
  );
  DFF_X1 \rf[8][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00596_),
    .Q(\rf[8] [31]),
    .QN(_09895_)
  );
  DFF_X1 \rf[8][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00816_),
    .Q(\rf[8] [3]),
    .QN(_09676_)
  );
  DFF_X1 \rf[8][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00817_),
    .Q(\rf[8] [4]),
    .QN(_09675_)
  );
  DFF_X1 \rf[8][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00818_),
    .Q(\rf[8] [5]),
    .QN(_09674_)
  );
  DFF_X1 \rf[8][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00819_),
    .Q(\rf[8] [6]),
    .QN(_09673_)
  );
  DFF_X1 \rf[8][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00820_),
    .Q(\rf[8] [7]),
    .QN(_09672_)
  );
  DFF_X1 \rf[8][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00821_),
    .Q(\rf[8] [8]),
    .QN(_09671_)
  );
  DFF_X1 \rf[8][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00822_),
    .Q(\rf[8] [9]),
    .QN(_09670_)
  );
  DFF_X1 \rf[9][0]$_DFFE_PP_  (
    .CK(clock),
    .D(_01092_),
    .Q(\rf[9] [0]),
    .QN(_09400_)
  );
  DFF_X1 \rf[9][10]$_DFFE_PP_  (
    .CK(clock),
    .D(_01102_),
    .Q(\rf[9] [10]),
    .QN(_09390_)
  );
  DFF_X1 \rf[9][11]$_DFFE_PP_  (
    .CK(clock),
    .D(_01103_),
    .Q(\rf[9] [11]),
    .QN(_09389_)
  );
  DFF_X1 \rf[9][12]$_DFFE_PP_  (
    .CK(clock),
    .D(_01104_),
    .Q(\rf[9] [12]),
    .QN(_09388_)
  );
  DFF_X1 \rf[9][13]$_DFFE_PP_  (
    .CK(clock),
    .D(_01105_),
    .Q(\rf[9] [13]),
    .QN(_09387_)
  );
  DFF_X1 \rf[9][14]$_DFFE_PP_  (
    .CK(clock),
    .D(_01106_),
    .Q(\rf[9] [14]),
    .QN(_09386_)
  );
  DFF_X1 \rf[9][15]$_DFFE_PP_  (
    .CK(clock),
    .D(_01107_),
    .Q(\rf[9] [15]),
    .QN(_09385_)
  );
  DFF_X1 \rf[9][16]$_DFFE_PP_  (
    .CK(clock),
    .D(_01108_),
    .Q(\rf[9] [16]),
    .QN(_09384_)
  );
  DFF_X1 \rf[9][17]$_DFFE_PP_  (
    .CK(clock),
    .D(_01109_),
    .Q(\rf[9] [17]),
    .QN(_09383_)
  );
  DFF_X1 \rf[9][18]$_DFFE_PP_  (
    .CK(clock),
    .D(_01110_),
    .Q(\rf[9] [18]),
    .QN(_09382_)
  );
  DFF_X1 \rf[9][19]$_DFFE_PP_  (
    .CK(clock),
    .D(_01111_),
    .Q(\rf[9] [19]),
    .QN(_09381_)
  );
  DFF_X1 \rf[9][1]$_DFFE_PP_  (
    .CK(clock),
    .D(_01093_),
    .Q(\rf[9] [1]),
    .QN(_09399_)
  );
  DFF_X1 \rf[9][20]$_DFFE_PP_  (
    .CK(clock),
    .D(_01112_),
    .Q(\rf[9] [20]),
    .QN(_09380_)
  );
  DFF_X1 \rf[9][21]$_DFFE_PP_  (
    .CK(clock),
    .D(_01113_),
    .Q(\rf[9] [21]),
    .QN(_09379_)
  );
  DFF_X1 \rf[9][22]$_DFFE_PP_  (
    .CK(clock),
    .D(_01114_),
    .Q(\rf[9] [22]),
    .QN(_09378_)
  );
  DFF_X1 \rf[9][23]$_DFFE_PP_  (
    .CK(clock),
    .D(_01115_),
    .Q(\rf[9] [23]),
    .QN(_09377_)
  );
  DFF_X1 \rf[9][24]$_DFFE_PP_  (
    .CK(clock),
    .D(_01116_),
    .Q(\rf[9] [24]),
    .QN(_09376_)
  );
  DFF_X1 \rf[9][25]$_DFFE_PP_  (
    .CK(clock),
    .D(_01117_),
    .Q(\rf[9] [25]),
    .QN(_09375_)
  );
  DFF_X1 \rf[9][26]$_DFFE_PP_  (
    .CK(clock),
    .D(_01118_),
    .Q(\rf[9] [26]),
    .QN(_09374_)
  );
  DFF_X1 \rf[9][27]$_DFFE_PP_  (
    .CK(clock),
    .D(_01119_),
    .Q(\rf[9] [27]),
    .QN(_09373_)
  );
  DFF_X1 \rf[9][28]$_DFFE_PP_  (
    .CK(clock),
    .D(_01120_),
    .Q(\rf[9] [28]),
    .QN(_09372_)
  );
  DFF_X1 \rf[9][29]$_DFFE_PP_  (
    .CK(clock),
    .D(_01121_),
    .Q(\rf[9] [29]),
    .QN(_09371_)
  );
  DFF_X1 \rf[9][2]$_DFFE_PP_  (
    .CK(clock),
    .D(_01094_),
    .Q(\rf[9] [2]),
    .QN(_09398_)
  );
  DFF_X1 \rf[9][30]$_DFFE_PP_  (
    .CK(clock),
    .D(_01122_),
    .Q(\rf[9] [30]),
    .QN(_09370_)
  );
  DFF_X1 \rf[9][31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00595_),
    .Q(\rf[9] [31]),
    .QN(_09896_)
  );
  DFF_X1 \rf[9][3]$_DFFE_PP_  (
    .CK(clock),
    .D(_01095_),
    .Q(\rf[9] [3]),
    .QN(_09397_)
  );
  DFF_X1 \rf[9][4]$_DFFE_PP_  (
    .CK(clock),
    .D(_01096_),
    .Q(\rf[9] [4]),
    .QN(_09396_)
  );
  DFF_X1 \rf[9][5]$_DFFE_PP_  (
    .CK(clock),
    .D(_01097_),
    .Q(\rf[9] [5]),
    .QN(_09395_)
  );
  DFF_X1 \rf[9][6]$_DFFE_PP_  (
    .CK(clock),
    .D(_01098_),
    .Q(\rf[9] [6]),
    .QN(_09394_)
  );
  DFF_X1 \rf[9][7]$_DFFE_PP_  (
    .CK(clock),
    .D(_01099_),
    .Q(\rf[9] [7]),
    .QN(_09393_)
  );
  DFF_X1 \rf[9][8]$_DFFE_PP_  (
    .CK(clock),
    .D(_01100_),
    .Q(\rf[9] [8]),
    .QN(_09392_)
  );
  DFF_X1 \rf[9][9]$_DFFE_PP_  (
    .CK(clock),
    .D(_01101_),
    .Q(\rf[9] [9]),
    .QN(_09391_)
  );
  DFF_X1 \wb_ctrl_csr[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00520_),
    .Q(wb_ctrl_csr[0]),
    .QN(_09954_)
  );
  DFF_X1 \wb_ctrl_csr[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00521_),
    .Q(wb_ctrl_csr[1]),
    .QN(_09953_)
  );
  DFF_X1 \wb_ctrl_csr[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00522_),
    .Q(wb_ctrl_csr[2]),
    .QN(_09952_)
  );
  DFF_X1 \wb_ctrl_div$_DFFE_PP_  (
    .CK(clock),
    .D(_00524_),
    .Q(wb_ctrl_div),
    .QN(_09950_)
  );
  DFF_X1 \wb_ctrl_fence_i$_DFFE_PP_  (
    .CK(clock),
    .D(_00519_),
    .Q(wb_ctrl_fence_i),
    .QN(_09955_)
  );
  DFF_X1 \wb_ctrl_mem$_DFFE_PP_  (
    .CK(clock),
    .D(_00525_),
    .Q(wb_ctrl_mem),
    .QN(_09949_)
  );
  DFF_X1 \wb_ctrl_wxd$_DFFE_PP_  (
    .CK(clock),
    .D(_00523_),
    .Q(wb_ctrl_wxd),
    .QN(_09951_)
  );
  DFF_X1 \wb_reg_cause[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00591_),
    .Q(wb_reg_cause[0]),
    .QN(_00016_)
  );
  DFF_X1 \wb_reg_cause[10]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00186_),
    .Q(wb_reg_cause[10]),
    .QN(_10284_)
  );
  DFF_X1 \wb_reg_cause[11]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00187_),
    .Q(wb_reg_cause[11]),
    .QN(_10283_)
  );
  DFF_X1 \wb_reg_cause[12]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00188_),
    .Q(wb_reg_cause[12]),
    .QN(_10282_)
  );
  DFF_X1 \wb_reg_cause[13]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00189_),
    .Q(wb_reg_cause[13]),
    .QN(_10281_)
  );
  DFF_X1 \wb_reg_cause[14]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00190_),
    .Q(wb_reg_cause[14]),
    .QN(_10280_)
  );
  DFF_X1 \wb_reg_cause[15]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00191_),
    .Q(wb_reg_cause[15]),
    .QN(_10279_)
  );
  DFF_X1 \wb_reg_cause[16]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00192_),
    .Q(wb_reg_cause[16]),
    .QN(_10278_)
  );
  DFF_X1 \wb_reg_cause[17]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00193_),
    .Q(wb_reg_cause[17]),
    .QN(_10277_)
  );
  DFF_X1 \wb_reg_cause[18]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00194_),
    .Q(wb_reg_cause[18]),
    .QN(_10276_)
  );
  DFF_X1 \wb_reg_cause[19]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00195_),
    .Q(wb_reg_cause[19]),
    .QN(_10275_)
  );
  DFF_X1 \wb_reg_cause[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00592_),
    .Q(wb_reg_cause[1]),
    .QN(_00015_)
  );
  DFF_X1 \wb_reg_cause[20]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00196_),
    .Q(wb_reg_cause[20]),
    .QN(_10274_)
  );
  DFF_X1 \wb_reg_cause[21]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00197_),
    .Q(wb_reg_cause[21]),
    .QN(_10273_)
  );
  DFF_X1 \wb_reg_cause[22]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00198_),
    .Q(wb_reg_cause[22]),
    .QN(_10272_)
  );
  DFF_X1 \wb_reg_cause[23]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00199_),
    .Q(wb_reg_cause[23]),
    .QN(_10271_)
  );
  DFF_X1 \wb_reg_cause[24]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00200_),
    .Q(wb_reg_cause[24]),
    .QN(_10270_)
  );
  DFF_X1 \wb_reg_cause[25]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00201_),
    .Q(wb_reg_cause[25]),
    .QN(_10269_)
  );
  DFF_X1 \wb_reg_cause[26]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00202_),
    .Q(wb_reg_cause[26]),
    .QN(_10268_)
  );
  DFF_X1 \wb_reg_cause[27]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00203_),
    .Q(wb_reg_cause[27]),
    .QN(_10267_)
  );
  DFF_X1 \wb_reg_cause[28]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00204_),
    .Q(wb_reg_cause[28]),
    .QN(_10266_)
  );
  DFF_X1 \wb_reg_cause[29]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00205_),
    .Q(wb_reg_cause[29]),
    .QN(_10265_)
  );
  DFF_X1 \wb_reg_cause[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00593_),
    .Q(wb_reg_cause[2]),
    .QN(_00014_)
  );
  DFF_X1 \wb_reg_cause[30]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00206_),
    .Q(wb_reg_cause[30]),
    .QN(_10264_)
  );
  DFF_X1 \wb_reg_cause[31]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00207_),
    .Q(wb_reg_cause[31]),
    .QN(_10432_)
  );
  DFF_X1 \wb_reg_cause[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00594_),
    .Q(wb_reg_cause[3]),
    .QN(_00013_)
  );
  DFF_X1 \wb_reg_cause[4]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00180_),
    .Q(wb_reg_cause[4]),
    .QN(_00030_)
  );
  DFF_X1 \wb_reg_cause[5]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00181_),
    .Q(wb_reg_cause[5]),
    .QN(_10289_)
  );
  DFF_X1 \wb_reg_cause[6]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00182_),
    .Q(wb_reg_cause[6]),
    .QN(_10288_)
  );
  DFF_X1 \wb_reg_cause[7]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00183_),
    .Q(wb_reg_cause[7]),
    .QN(_10287_)
  );
  DFF_X1 \wb_reg_cause[8]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00184_),
    .Q(wb_reg_cause[8]),
    .QN(_10286_)
  );
  DFF_X1 \wb_reg_cause[9]$_SDFFCE_PN0P_  (
    .CK(clock),
    .D(_00185_),
    .Q(wb_reg_cause[9]),
    .QN(_10285_)
  );
  DFF_X1 \wb_reg_flush_pipe$_DFF_P_  (
    .CK(clock),
    .D(_00009_),
    .Q(wb_reg_flush_pipe),
    .QN(_10433_)
  );
  DFF_X1 \wb_reg_inst[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00529_),
    .Q(wb_reg_inst[10]),
    .QN(_09946_)
  );
  DFF_X1 \wb_reg_inst[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00530_),
    .Q(wb_reg_inst[11]),
    .QN(_09945_)
  );
  DFF_X1 \wb_reg_inst[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00531_),
    .Q(wb_reg_inst[16]),
    .QN(_09944_)
  );
  DFF_X1 \wb_reg_inst[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00532_),
    .Q(wb_reg_inst[17]),
    .QN(_09943_)
  );
  DFF_X1 \wb_reg_inst[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00533_),
    .Q(wb_reg_inst[18]),
    .QN(_09942_)
  );
  DFF_X1 \wb_reg_inst[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00534_),
    .Q(wb_reg_inst[19]),
    .QN(_09941_)
  );
  DFF_X1 \wb_reg_inst[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00535_),
    .Q(wb_reg_inst[20]),
    .QN(_09940_)
  );
  DFF_X1 \wb_reg_inst[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00536_),
    .Q(wb_reg_inst[21]),
    .QN(_09939_)
  );
  DFF_X1 \wb_reg_inst[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00537_),
    .Q(wb_reg_inst[22]),
    .QN(_09938_)
  );
  DFF_X1 \wb_reg_inst[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00538_),
    .Q(wb_reg_inst[23]),
    .QN(_09937_)
  );
  DFF_X1 \wb_reg_inst[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00539_),
    .Q(wb_reg_inst[24]),
    .QN(_09936_)
  );
  DFF_X1 \wb_reg_inst[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00540_),
    .Q(wb_reg_inst[25]),
    .QN(_09935_)
  );
  DFF_X1 \wb_reg_inst[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00541_),
    .Q(wb_reg_inst[26]),
    .QN(_09934_)
  );
  DFF_X1 \wb_reg_inst[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00542_),
    .Q(wb_reg_inst[27]),
    .QN(_09933_)
  );
  DFF_X1 \wb_reg_inst[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00543_),
    .Q(wb_reg_inst[28]),
    .QN(_09932_)
  );
  DFF_X1 \wb_reg_inst[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00544_),
    .Q(wb_reg_inst[29]),
    .QN(_09931_)
  );
  DFF_X1 \wb_reg_inst[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00545_),
    .Q(wb_reg_inst[30]),
    .QN(_09930_)
  );
  DFF_X1 \wb_reg_inst[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00546_),
    .Q(wb_reg_inst[31]),
    .QN(_09929_)
  );
  DFF_X1 \wb_reg_inst[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00526_),
    .Q(wb_reg_inst[7]),
    .QN(_00029_)
  );
  DFF_X1 \wb_reg_inst[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00527_),
    .Q(wb_reg_inst[8]),
    .QN(_09948_)
  );
  DFF_X1 \wb_reg_inst[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00528_),
    .Q(wb_reg_inst[9]),
    .QN(_09947_)
  );
  DFF_X1 \wb_reg_pc[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00208_),
    .Q(wb_reg_pc[0]),
    .QN(_10262_)
  );
  DFF_X1 \wb_reg_pc[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00218_),
    .Q(wb_reg_pc[10]),
    .QN(_10252_)
  );
  DFF_X1 \wb_reg_pc[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00219_),
    .Q(wb_reg_pc[11]),
    .QN(_10251_)
  );
  DFF_X1 \wb_reg_pc[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00220_),
    .Q(wb_reg_pc[12]),
    .QN(_10250_)
  );
  DFF_X1 \wb_reg_pc[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00221_),
    .Q(wb_reg_pc[13]),
    .QN(_10249_)
  );
  DFF_X1 \wb_reg_pc[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00222_),
    .Q(wb_reg_pc[14]),
    .QN(_10248_)
  );
  DFF_X1 \wb_reg_pc[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00223_),
    .Q(wb_reg_pc[15]),
    .QN(_10247_)
  );
  DFF_X1 \wb_reg_pc[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00224_),
    .Q(wb_reg_pc[16]),
    .QN(_10246_)
  );
  DFF_X1 \wb_reg_pc[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00225_),
    .Q(wb_reg_pc[17]),
    .QN(_10245_)
  );
  DFF_X1 \wb_reg_pc[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00226_),
    .Q(wb_reg_pc[18]),
    .QN(_10244_)
  );
  DFF_X1 \wb_reg_pc[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00227_),
    .Q(wb_reg_pc[19]),
    .QN(_10243_)
  );
  DFF_X1 \wb_reg_pc[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00209_),
    .Q(wb_reg_pc[1]),
    .QN(_10261_)
  );
  DFF_X1 \wb_reg_pc[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00228_),
    .Q(wb_reg_pc[20]),
    .QN(_10242_)
  );
  DFF_X1 \wb_reg_pc[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00229_),
    .Q(wb_reg_pc[21]),
    .QN(_10241_)
  );
  DFF_X1 \wb_reg_pc[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00230_),
    .Q(wb_reg_pc[22]),
    .QN(_10240_)
  );
  DFF_X1 \wb_reg_pc[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00231_),
    .Q(wb_reg_pc[23]),
    .QN(_10239_)
  );
  DFF_X1 \wb_reg_pc[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00232_),
    .Q(wb_reg_pc[24]),
    .QN(_10238_)
  );
  DFF_X1 \wb_reg_pc[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00233_),
    .Q(wb_reg_pc[25]),
    .QN(_10237_)
  );
  DFF_X1 \wb_reg_pc[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00234_),
    .Q(wb_reg_pc[26]),
    .QN(_10236_)
  );
  DFF_X1 \wb_reg_pc[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00235_),
    .Q(wb_reg_pc[27]),
    .QN(_10235_)
  );
  DFF_X1 \wb_reg_pc[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00236_),
    .Q(wb_reg_pc[28]),
    .QN(_10234_)
  );
  DFF_X1 \wb_reg_pc[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00237_),
    .Q(wb_reg_pc[29]),
    .QN(_10233_)
  );
  DFF_X1 \wb_reg_pc[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00210_),
    .Q(wb_reg_pc[2]),
    .QN(_10260_)
  );
  DFF_X1 \wb_reg_pc[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00238_),
    .Q(wb_reg_pc[30]),
    .QN(_10232_)
  );
  DFF_X1 \wb_reg_pc[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00239_),
    .Q(wb_reg_pc[31]),
    .QN(_10231_)
  );
  DFF_X1 \wb_reg_pc[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00211_),
    .Q(wb_reg_pc[3]),
    .QN(_10259_)
  );
  DFF_X1 \wb_reg_pc[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00212_),
    .Q(wb_reg_pc[4]),
    .QN(_10258_)
  );
  DFF_X1 \wb_reg_pc[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00213_),
    .Q(wb_reg_pc[5]),
    .QN(_10257_)
  );
  DFF_X1 \wb_reg_pc[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00214_),
    .Q(wb_reg_pc[6]),
    .QN(_10256_)
  );
  DFF_X1 \wb_reg_pc[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00215_),
    .Q(wb_reg_pc[7]),
    .QN(_10255_)
  );
  DFF_X1 \wb_reg_pc[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00216_),
    .Q(wb_reg_pc[8]),
    .QN(_10254_)
  );
  DFF_X1 \wb_reg_pc[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00217_),
    .Q(wb_reg_pc[9]),
    .QN(_10253_)
  );
  DFF_X1 \wb_reg_raw_inst[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00101_),
    .Q(wb_reg_raw_inst[0]),
    .QN(_10367_)
  );
  DFF_X1 \wb_reg_raw_inst[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00111_),
    .Q(wb_reg_raw_inst[10]),
    .QN(_10357_)
  );
  DFF_X1 \wb_reg_raw_inst[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00112_),
    .Q(wb_reg_raw_inst[11]),
    .QN(_10356_)
  );
  DFF_X1 \wb_reg_raw_inst[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00113_),
    .Q(wb_reg_raw_inst[12]),
    .QN(_10355_)
  );
  DFF_X1 \wb_reg_raw_inst[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00114_),
    .Q(wb_reg_raw_inst[13]),
    .QN(_10354_)
  );
  DFF_X1 \wb_reg_raw_inst[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00115_),
    .Q(wb_reg_raw_inst[14]),
    .QN(_10353_)
  );
  DFF_X1 \wb_reg_raw_inst[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00116_),
    .Q(wb_reg_raw_inst[15]),
    .QN(_10352_)
  );
  DFF_X1 \wb_reg_raw_inst[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00102_),
    .Q(wb_reg_raw_inst[1]),
    .QN(_10366_)
  );
  DFF_X1 \wb_reg_raw_inst[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00103_),
    .Q(wb_reg_raw_inst[2]),
    .QN(_10365_)
  );
  DFF_X1 \wb_reg_raw_inst[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00104_),
    .Q(wb_reg_raw_inst[3]),
    .QN(_10364_)
  );
  DFF_X1 \wb_reg_raw_inst[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00105_),
    .Q(wb_reg_raw_inst[4]),
    .QN(_10363_)
  );
  DFF_X1 \wb_reg_raw_inst[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00106_),
    .Q(wb_reg_raw_inst[5]),
    .QN(_10362_)
  );
  DFF_X1 \wb_reg_raw_inst[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00107_),
    .Q(wb_reg_raw_inst[6]),
    .QN(_10361_)
  );
  DFF_X1 \wb_reg_raw_inst[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00108_),
    .Q(wb_reg_raw_inst[7]),
    .QN(_10360_)
  );
  DFF_X1 \wb_reg_raw_inst[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00109_),
    .Q(wb_reg_raw_inst[8]),
    .QN(_10359_)
  );
  DFF_X1 \wb_reg_raw_inst[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00110_),
    .Q(wb_reg_raw_inst[9]),
    .QN(_10358_)
  );
  DFF_X1 \wb_reg_replay$_DFF_P_  (
    .CK(clock),
    .D(_00010_),
    .Q(wb_reg_replay),
    .QN(_10434_)
  );
  DFF_X1 \wb_reg_valid$_DFF_P_  (
    .CK(clock),
    .D(_wb_reg_valid_T),
    .Q(wb_reg_valid),
    .QN(_10263_)
  );
  DFF_X1 \wb_reg_wdata[0]$_DFFE_PP_  (
    .CK(clock),
    .D(_00117_),
    .Q(wb_reg_wdata[0]),
    .QN(_10351_)
  );
  DFF_X1 \wb_reg_wdata[10]$_DFFE_PP_  (
    .CK(clock),
    .D(_00127_),
    .Q(wb_reg_wdata[10]),
    .QN(_10341_)
  );
  DFF_X1 \wb_reg_wdata[11]$_DFFE_PP_  (
    .CK(clock),
    .D(_00128_),
    .Q(wb_reg_wdata[11]),
    .QN(_10340_)
  );
  DFF_X1 \wb_reg_wdata[12]$_DFFE_PP_  (
    .CK(clock),
    .D(_00129_),
    .Q(wb_reg_wdata[12]),
    .QN(_10339_)
  );
  DFF_X1 \wb_reg_wdata[13]$_DFFE_PP_  (
    .CK(clock),
    .D(_00130_),
    .Q(wb_reg_wdata[13]),
    .QN(_10338_)
  );
  DFF_X1 \wb_reg_wdata[14]$_DFFE_PP_  (
    .CK(clock),
    .D(_00131_),
    .Q(wb_reg_wdata[14]),
    .QN(_10337_)
  );
  DFF_X1 \wb_reg_wdata[15]$_DFFE_PP_  (
    .CK(clock),
    .D(_00132_),
    .Q(wb_reg_wdata[15]),
    .QN(_10336_)
  );
  DFF_X1 \wb_reg_wdata[16]$_DFFE_PP_  (
    .CK(clock),
    .D(_00133_),
    .Q(wb_reg_wdata[16]),
    .QN(_10335_)
  );
  DFF_X1 \wb_reg_wdata[17]$_DFFE_PP_  (
    .CK(clock),
    .D(_00134_),
    .Q(wb_reg_wdata[17]),
    .QN(_10334_)
  );
  DFF_X1 \wb_reg_wdata[18]$_DFFE_PP_  (
    .CK(clock),
    .D(_00135_),
    .Q(wb_reg_wdata[18]),
    .QN(_10333_)
  );
  DFF_X1 \wb_reg_wdata[19]$_DFFE_PP_  (
    .CK(clock),
    .D(_00136_),
    .Q(wb_reg_wdata[19]),
    .QN(_10332_)
  );
  DFF_X1 \wb_reg_wdata[1]$_DFFE_PP_  (
    .CK(clock),
    .D(_00118_),
    .Q(wb_reg_wdata[1]),
    .QN(_10350_)
  );
  DFF_X1 \wb_reg_wdata[20]$_DFFE_PP_  (
    .CK(clock),
    .D(_00137_),
    .Q(wb_reg_wdata[20]),
    .QN(_10331_)
  );
  DFF_X1 \wb_reg_wdata[21]$_DFFE_PP_  (
    .CK(clock),
    .D(_00138_),
    .Q(wb_reg_wdata[21]),
    .QN(_10330_)
  );
  DFF_X1 \wb_reg_wdata[22]$_DFFE_PP_  (
    .CK(clock),
    .D(_00139_),
    .Q(wb_reg_wdata[22]),
    .QN(_10329_)
  );
  DFF_X1 \wb_reg_wdata[23]$_DFFE_PP_  (
    .CK(clock),
    .D(_00140_),
    .Q(wb_reg_wdata[23]),
    .QN(_10328_)
  );
  DFF_X1 \wb_reg_wdata[24]$_DFFE_PP_  (
    .CK(clock),
    .D(_00141_),
    .Q(wb_reg_wdata[24]),
    .QN(_10327_)
  );
  DFF_X1 \wb_reg_wdata[25]$_DFFE_PP_  (
    .CK(clock),
    .D(_00142_),
    .Q(wb_reg_wdata[25]),
    .QN(_10326_)
  );
  DFF_X1 \wb_reg_wdata[26]$_DFFE_PP_  (
    .CK(clock),
    .D(_00143_),
    .Q(wb_reg_wdata[26]),
    .QN(_10325_)
  );
  DFF_X1 \wb_reg_wdata[27]$_DFFE_PP_  (
    .CK(clock),
    .D(_00144_),
    .Q(wb_reg_wdata[27]),
    .QN(_10324_)
  );
  DFF_X1 \wb_reg_wdata[28]$_DFFE_PP_  (
    .CK(clock),
    .D(_00145_),
    .Q(wb_reg_wdata[28]),
    .QN(_10323_)
  );
  DFF_X1 \wb_reg_wdata[29]$_DFFE_PP_  (
    .CK(clock),
    .D(_00146_),
    .Q(wb_reg_wdata[29]),
    .QN(_10322_)
  );
  DFF_X1 \wb_reg_wdata[2]$_DFFE_PP_  (
    .CK(clock),
    .D(_00119_),
    .Q(wb_reg_wdata[2]),
    .QN(_10349_)
  );
  DFF_X1 \wb_reg_wdata[30]$_DFFE_PP_  (
    .CK(clock),
    .D(_00147_),
    .Q(wb_reg_wdata[30]),
    .QN(_10321_)
  );
  DFF_X1 \wb_reg_wdata[31]$_DFFE_PP_  (
    .CK(clock),
    .D(_00148_),
    .Q(wb_reg_wdata[31]),
    .QN(_10320_)
  );
  DFF_X1 \wb_reg_wdata[3]$_DFFE_PP_  (
    .CK(clock),
    .D(_00120_),
    .Q(wb_reg_wdata[3]),
    .QN(_10348_)
  );
  DFF_X1 \wb_reg_wdata[4]$_DFFE_PP_  (
    .CK(clock),
    .D(_00121_),
    .Q(wb_reg_wdata[4]),
    .QN(_10347_)
  );
  DFF_X1 \wb_reg_wdata[5]$_DFFE_PP_  (
    .CK(clock),
    .D(_00122_),
    .Q(wb_reg_wdata[5]),
    .QN(_10346_)
  );
  DFF_X1 \wb_reg_wdata[6]$_DFFE_PP_  (
    .CK(clock),
    .D(_00123_),
    .Q(wb_reg_wdata[6]),
    .QN(_10345_)
  );
  DFF_X1 \wb_reg_wdata[7]$_DFFE_PP_  (
    .CK(clock),
    .D(_00124_),
    .Q(wb_reg_wdata[7]),
    .QN(_10344_)
  );
  DFF_X1 \wb_reg_wdata[8]$_DFFE_PP_  (
    .CK(clock),
    .D(_00125_),
    .Q(wb_reg_wdata[8]),
    .QN(_10343_)
  );
  DFF_X1 \wb_reg_wdata[9]$_DFFE_PP_  (
    .CK(clock),
    .D(_00126_),
    .Q(wb_reg_wdata[9]),
    .QN(_10342_)
  );
  DFF_X1 \wb_reg_xcpt$_DFF_P_  (
    .CK(clock),
    .D(_00011_),
    .Q(wb_reg_xcpt),
    .QN(tval_dmem_addr)
  );
  assign _10441_[1] = ex_reg_mem_size[1];
  assign _10442_[0] = ex_reg_mem_size[0];
  assign PlusArgTimeout_clock = clock;
  assign PlusArgTimeout_io_count = csr_io_time;
  assign PlusArgTimeout_reset = reset;
  assign { _T_11[4:2], _T_11[0] } = { 3'h0, ibuf_io_inst_0_bits_xcpt1_ae_inst };
  assign { _T_113[2], _T_113[0] } = 2'h2;
  assign _T_114[2] = 1'h1;
  assign _T_115[2] = 1'h1;
  assign _T_116 = { 3'h1, _T_115[1:0] };
  assign { _T_118[4], _T_118[2] } = 2'h1;
  assign { _T_119[4], _T_119[2] } = 2'h1;
  assign _T_12[4:2] = { ibuf_io_inst_0_bits_xcpt1_gf_inst, 1'h0, ibuf_io_inst_0_bits_xcpt1_gf_inst };
  assign _T_13[3] = ibuf_io_inst_0_bits_xcpt1_pf_inst;
  assign _T_143[0] = 1'h0;
  assign _T_35 = { ibuf_io_inst_0_bits_xcpt1_pf_inst, ibuf_io_inst_0_bits_xcpt1_gf_inst, ibuf_io_inst_0_bits_xcpt1_ae_inst };
  assign _T_37 = { 2'h0, ibuf_io_inst_0_bits_xcpt0_ae_inst };
  assign _T_40 = 1'h0;
  assign _T_41 = 1'h0;
  assign _T_42 = 1'h0;
  assign _T_74[2] = _T_74[3];
  assign _T_93 = _T_118[3];
  assign _bypass_src_T[1] = 1'h1;
  assign _bypass_src_T_2[1] = 1'h1;
  assign _csr_io_rw_cmd_T[1:0] = 2'h0;
  assign _csr_io_rw_cmd_T_1 = { wb_reg_valid, 2'h3 };
  assign _ctrl_stalld_T_15 = 1'h0;
  assign _ex_imm_b11_T_5 = ex_reg_inst[20];
  assign _ex_imm_b11_T_8 = ex_reg_inst[7];
  assign _ex_imm_b19_12_T_4 = ex_reg_inst[19:12];
  assign _ex_imm_b30_20_T_2 = ex_reg_inst[30:20];
  assign _ex_imm_sign_T_2 = ex_reg_inst[31];
  assign { _ex_op2_T_1[3], _ex_op2_T_1[1:0] } = { 1'h0, ex_reg_rvc, 1'h0 };
  assign _ex_rs_T_13 = { ex_reg_rs_msb_1, ex_reg_rs_lsb_1 };
  assign _ex_rs_T_6 = { ex_reg_rs_msb_0, ex_reg_rs_lsb_0 };
  assign _id_ctrl_decoder_decoded_T[7:6] = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1] };
  assign _id_ctrl_decoder_decoded_T_10[8:1] = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], csr_io_decode_0_inst[3], _id_ctrl_decoder_decoded_T[3:0] };
  assign _id_ctrl_decoder_decoded_T_100 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:3], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], csr_io_decode_0_inst[13], csr_io_decode_0_inst[14] };
  assign _id_ctrl_decoder_decoded_T_102 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], csr_io_decode_0_inst[13], csr_io_decode_0_inst[14] };
  assign _id_ctrl_decoder_decoded_T_104 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], _id_ctrl_decoder_decoded_T[2:1], csr_io_decode_0_inst[12], csr_io_decode_0_inst[13], csr_io_decode_0_inst[14] };
  assign _id_ctrl_decoder_decoded_T_106[13:6] = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[25] };
  assign _id_ctrl_decoder_decoded_T_108 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[12], csr_io_decode_0_inst[25], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign _id_ctrl_decoder_decoded_T_110 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[13], csr_io_decode_0_inst[25], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign { _id_ctrl_decoder_decoded_T_112[13:7], _id_ctrl_decoder_decoded_T_112[5:0] } = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], csr_io_decode_0_inst[3], _id_ctrl_decoder_decoded_T[3], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0], csr_io_decode_0_inst[27], _id_ctrl_decoder_decoded_T_106[2:0] };
  assign { _id_ctrl_decoder_decoded_T_114[16:10], _id_ctrl_decoder_decoded_T_114[4:0] } = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], csr_io_decode_0_inst[3], _id_ctrl_decoder_decoded_T[3], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T_106[4], csr_io_decode_0_inst[28], _id_ctrl_decoder_decoded_T_106[2:0] };
  assign _id_ctrl_decoder_decoded_T_116 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], csr_io_decode_0_inst[3], _id_ctrl_decoder_decoded_T[3], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T_112[6], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_114[9:5], _id_ctrl_decoder_decoded_T_106[4], csr_io_decode_0_inst[28], _id_ctrl_decoder_decoded_T_106[2:0] };
  assign { _id_ctrl_decoder_decoded_T_118[27:24], _id_ctrl_decoder_decoded_T_118[18:16], _id_ctrl_decoder_decoded_T_118[10:6], _id_ctrl_decoder_decoded_T_118[4:0] } = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0], csr_io_decode_0_inst[20], _id_ctrl_decoder_decoded_T_114[8], csr_io_decode_0_inst[22], _id_ctrl_decoder_decoded_T_114[6:5], _id_ctrl_decoder_decoded_T_106[5:4], csr_io_decode_0_inst[28], _id_ctrl_decoder_decoded_T_106[1:0] };
  assign _id_ctrl_decoder_decoded_T_12 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], _id_ctrl_decoder_decoded_T[4], csr_io_decode_0_inst[4], _id_ctrl_decoder_decoded_T[1] };
  assign _id_ctrl_decoder_decoded_T_120 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], _id_ctrl_decoder_decoded_T_118[23:19], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[15:11], csr_io_decode_0_inst[20], _id_ctrl_decoder_decoded_T_114[8], csr_io_decode_0_inst[22], _id_ctrl_decoder_decoded_T_114[6:5], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:4], csr_io_decode_0_inst[28], _id_ctrl_decoder_decoded_T_106[1:0] };
  assign _id_ctrl_decoder_decoded_T_122 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], csr_io_decode_0_inst[3], _id_ctrl_decoder_decoded_T[3], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T_112[6], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0], csr_io_decode_0_inst[27], csr_io_decode_0_inst[28], _id_ctrl_decoder_decoded_T_106[2:0] };
  assign _id_ctrl_decoder_decoded_T_124 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], csr_io_decode_0_inst[3], _id_ctrl_decoder_decoded_T[3], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T_112[6], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_106[4:3], csr_io_decode_0_inst[29] };
  assign _id_ctrl_decoder_decoded_T_126 = { csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], _id_ctrl_decoder_decoded_T_118[23:19], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[15:11], _id_ctrl_decoder_decoded_T_114[9], csr_io_decode_0_inst[21], _id_ctrl_decoder_decoded_T_114[7:5], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:4], csr_io_decode_0_inst[28], csr_io_decode_0_inst[29], _id_ctrl_decoder_decoded_T_106[1:0] };
  assign _id_ctrl_decoder_decoded_T_128 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], _id_ctrl_decoder_decoded_T_118[23:19], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[15:11], _id_ctrl_decoder_decoded_T_114[9], csr_io_decode_0_inst[21], _id_ctrl_decoder_decoded_T_114[7:5], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:4], csr_io_decode_0_inst[28], csr_io_decode_0_inst[29], _id_ctrl_decoder_decoded_T_106[1:0] };
  assign _id_ctrl_decoder_decoded_T_130 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:2], csr_io_decode_0_inst[30], _id_ctrl_decoder_decoded_T_106[0] };
  assign _id_ctrl_decoder_decoded_T_132 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], csr_io_decode_0_inst[3], _id_ctrl_decoder_decoded_T[3], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T_112[6], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_106[4:3], csr_io_decode_0_inst[30] };
  assign _id_ctrl_decoder_decoded_T_134 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[12], _id_ctrl_decoder_decoded_T[0], csr_io_decode_0_inst[14], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:2], csr_io_decode_0_inst[30], _id_ctrl_decoder_decoded_T_106[0] };
  assign _id_ctrl_decoder_decoded_T_136 = { csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], _id_ctrl_decoder_decoded_T_118[23:19], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[15:11], _id_ctrl_decoder_decoded_T_114[9], csr_io_decode_0_inst[21], _id_ctrl_decoder_decoded_T_114[7:6], csr_io_decode_0_inst[24], csr_io_decode_0_inst[25], _id_ctrl_decoder_decoded_T_106[5], csr_io_decode_0_inst[27], csr_io_decode_0_inst[28], csr_io_decode_0_inst[29], csr_io_decode_0_inst[30], _id_ctrl_decoder_decoded_T_106[0] };
  assign _id_ctrl_decoder_decoded_T_138 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], _id_ctrl_decoder_decoded_T_118[23:19], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[15:11], _id_ctrl_decoder_decoded_T_114[9], csr_io_decode_0_inst[21], _id_ctrl_decoder_decoded_T_114[7:6], csr_io_decode_0_inst[24], csr_io_decode_0_inst[25], _id_ctrl_decoder_decoded_T_106[5], csr_io_decode_0_inst[27], csr_io_decode_0_inst[28], csr_io_decode_0_inst[29], csr_io_decode_0_inst[30], _id_ctrl_decoder_decoded_T_106[0] };
  assign _id_ctrl_decoder_decoded_T_14 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], _id_ctrl_decoder_decoded_T[4], csr_io_decode_0_inst[4], _id_ctrl_decoder_decoded_T[2:1] };
  assign _id_ctrl_decoder_decoded_T_140 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], csr_io_decode_0_inst[3], _id_ctrl_decoder_decoded_T[3], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T_112[6], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_106[4:3], csr_io_decode_0_inst[31] };
  assign _id_ctrl_decoder_decoded_T_16 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:3], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T_10[0] };
  assign _id_ctrl_decoder_decoded_T_18 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:3], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0] };
  assign _id_ctrl_decoder_decoded_T_2 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], _id_ctrl_decoder_decoded_T[2:1], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0] };
  assign _id_ctrl_decoder_decoded_T_20 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:3], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1:0], _id_ctrl_decoder_decoded_T_10[0] };
  assign _id_ctrl_decoder_decoded_T_22 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:2], _id_ctrl_decoder_decoded_T_106[0] };
  assign _id_ctrl_decoder_decoded_T_24 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign _id_ctrl_decoder_decoded_T_26 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:3], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], _id_ctrl_decoder_decoded_T[0] };
  assign _id_ctrl_decoder_decoded_T_28 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:3], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0] };
  assign _id_ctrl_decoder_decoded_T_30 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[4:3], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0] };
  assign _id_ctrl_decoder_decoded_T_32 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], _id_ctrl_decoder_decoded_T[4:3], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0] };
  assign _id_ctrl_decoder_decoded_T_34 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], csr_io_decode_0_inst[3], _id_ctrl_decoder_decoded_T[3], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6] };
  assign _id_ctrl_decoder_decoded_T_36 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], _id_ctrl_decoder_decoded_T_118[23:19], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[15:11], _id_ctrl_decoder_decoded_T_114[8:5], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign _id_ctrl_decoder_decoded_T_38 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], _id_ctrl_decoder_decoded_T_118[23:19], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[15:11], _id_ctrl_decoder_decoded_T_114[8:5], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign _id_ctrl_decoder_decoded_T_4 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:3], _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T_10[0] };
  assign _id_ctrl_decoder_decoded_T_40 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], csr_io_decode_0_inst[3], _id_ctrl_decoder_decoded_T[3:1], csr_io_decode_0_inst[12], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0] };
  assign _id_ctrl_decoder_decoded_T_42 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[12], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign _id_ctrl_decoder_decoded_T_44 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], _id_ctrl_decoder_decoded_T[2:1], csr_io_decode_0_inst[12], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign _id_ctrl_decoder_decoded_T_46 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], csr_io_decode_0_inst[12], _id_ctrl_decoder_decoded_T[0] };
  assign _id_ctrl_decoder_decoded_T_48 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:3], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], csr_io_decode_0_inst[12], _id_ctrl_decoder_decoded_T[0] };
  assign _id_ctrl_decoder_decoded_T_50 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], csr_io_decode_0_inst[12], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0] };
  assign _id_ctrl_decoder_decoded_T_52 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], csr_io_decode_0_inst[12] };
  assign _id_ctrl_decoder_decoded_T_54 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], _id_ctrl_decoder_decoded_T[2:1], csr_io_decode_0_inst[13] };
  assign _id_ctrl_decoder_decoded_T_56 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], _id_ctrl_decoder_decoded_T[2:1], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0] };
  assign _id_ctrl_decoder_decoded_T_58 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], csr_io_decode_0_inst[3], _id_ctrl_decoder_decoded_T[3], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T_112[6], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_106[4:3] };
  assign _id_ctrl_decoder_decoded_T_6 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], _id_ctrl_decoder_decoded_T[2:1], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T_10[0] };
  assign _id_ctrl_decoder_decoded_T_60 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign _id_ctrl_decoder_decoded_T_62 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign _id_ctrl_decoder_decoded_T_64 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], csr_io_decode_0_inst[13] };
  assign _id_ctrl_decoder_decoded_T_66 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0] };
  assign _id_ctrl_decoder_decoded_T_68 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], _id_ctrl_decoder_decoded_T[2:1], csr_io_decode_0_inst[12], csr_io_decode_0_inst[13] };
  assign _id_ctrl_decoder_decoded_T_70 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[12], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign _id_ctrl_decoder_decoded_T_72 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], _id_ctrl_decoder_decoded_T[2:1], _id_ctrl_decoder_decoded_T_112[6], csr_io_decode_0_inst[14] };
  assign _id_ctrl_decoder_decoded_T_74 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[14], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign _id_ctrl_decoder_decoded_T_76 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:3], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], csr_io_decode_0_inst[14] };
  assign _id_ctrl_decoder_decoded_T_78 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[12], _id_ctrl_decoder_decoded_T[0], csr_io_decode_0_inst[14], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:2], _id_ctrl_decoder_decoded_T_106[0] };
  assign _id_ctrl_decoder_decoded_T_8 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:3], _id_ctrl_decoder_decoded_T[1:0], _id_ctrl_decoder_decoded_T_10[0] };
  assign _id_ctrl_decoder_decoded_T_80 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], _id_ctrl_decoder_decoded_T[2:1], csr_io_decode_0_inst[12], _id_ctrl_decoder_decoded_T[0], csr_io_decode_0_inst[14], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:2], _id_ctrl_decoder_decoded_T_106[0] };
  assign _id_ctrl_decoder_decoded_T_82 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[12], _id_ctrl_decoder_decoded_T[0], csr_io_decode_0_inst[14], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign _id_ctrl_decoder_decoded_T_84 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[12], _id_ctrl_decoder_decoded_T[0], csr_io_decode_0_inst[14], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:2], _id_ctrl_decoder_decoded_T_106[0] };
  assign _id_ctrl_decoder_decoded_T_86 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[12], csr_io_decode_0_inst[14], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign _id_ctrl_decoder_decoded_T_88 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], csr_io_decode_0_inst[12], csr_io_decode_0_inst[14] };
  assign _id_ctrl_decoder_decoded_T_90 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:3], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], csr_io_decode_0_inst[12], csr_io_decode_0_inst[14] };
  assign _id_ctrl_decoder_decoded_T_92 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], csr_io_decode_0_inst[12], csr_io_decode_0_inst[14] };
  assign _id_ctrl_decoder_decoded_T_94 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], _id_ctrl_decoder_decoded_T[2:1], csr_io_decode_0_inst[13], csr_io_decode_0_inst[14] };
  assign _id_ctrl_decoder_decoded_T_96 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[4], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], csr_io_decode_0_inst[13], csr_io_decode_0_inst[14], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign _id_ctrl_decoder_decoded_T_98 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], _id_ctrl_decoder_decoded_T[5:4], csr_io_decode_0_inst[5], csr_io_decode_0_inst[6], csr_io_decode_0_inst[13], csr_io_decode_0_inst[14] };
  assign _id_illegal_insn_T_11 = 1'h0;
  assign _id_illegal_insn_T_15 = 1'h0;
  assign _id_illegal_insn_T_33 = 1'h0;
  assign _io_fpu_time_T = csr_io_time;
  assign _mem_br_target_T_3 = { mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[7], mem_reg_inst[30:25], mem_reg_inst[11:8], 1'h0 };
  assign _mem_br_target_T_5 = { mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[19:12], mem_reg_inst[20], mem_reg_inst[30:21], 1'h0 };
  assign { _mem_br_target_T_6[3], _mem_br_target_T_6[1:0] } = { 1'h0, mem_reg_rvc, 1'h0 };
  assign { _mem_br_target_T_7[30:20], _mem_br_target_T_7[0] } = { _mem_br_target_T_7[31], _mem_br_target_T_7[31], _mem_br_target_T_7[31], _mem_br_target_T_7[31], _mem_br_target_T_7[31], _mem_br_target_T_7[31], _mem_br_target_T_7[31], _mem_br_target_T_7[31], _mem_br_target_T_7[31], _mem_br_target_T_7[31], _mem_br_target_T_7[31], 1'h0 };
  assign { _mem_br_target_T_8[30:20], _mem_br_target_T_8[0] } = { _mem_br_target_T_8[31], _mem_br_target_T_8[31], _mem_br_target_T_8[31], _mem_br_target_T_8[31], _mem_br_target_T_8[31], _mem_br_target_T_8[31], _mem_br_target_T_8[31], _mem_br_target_T_8[31], _mem_br_target_T_8[31], _mem_br_target_T_8[31], _mem_br_target_T_8[31], 1'h0 };
  assign _mem_reg_load_T_1 = 1'h0;
  assign _mem_reg_rs2_T_3 = { _ex_op2_T[7:0], _ex_op2_T[7:0], _ex_op2_T[7:0], _ex_op2_T[7:0] };
  assign _mem_reg_rs2_T_6 = { _ex_op2_T[15:0], _ex_op2_T[15:0] };
  assign _mem_reg_rs2_T_7[15:0] = _ex_op2_T[15:0];
  assign _mem_reg_wdata_T = alu_io_out;
  assign _wb_reg_replay_T = io_imem_req_bits_speculative;
  assign alu_io_fn = ex_ctrl_alu_fn;
  assign bpu_io_ea = mem_reg_wdata;
  assign coreMonitorBundle_inst = csr_io_trace_0_insn;
  assign coreMonitorBundle_pc = csr_io_trace_0_iaddr;
  assign csr_clock = clock;
  assign csr_io_bp_0_address = bpu_io_bp_0_address;
  assign csr_io_bp_0_control_action = bpu_io_bp_0_control_action;
  assign csr_io_bp_0_control_r = bpu_io_bp_0_control_r;
  assign csr_io_bp_0_control_tmatch = bpu_io_bp_0_control_tmatch;
  assign csr_io_bp_0_control_w = bpu_io_bp_0_control_w;
  assign csr_io_bp_0_control_x = bpu_io_bp_0_control_x;
  assign csr_io_customCSRs_0_value[1] = io_ptw_customCSRs_csrs_0_value[1];
  assign csr_io_gva = 1'h0;
  assign csr_io_hartid = io_hartid;
  assign csr_io_inst_0 = { _csr_io_inst_0_T_3, wb_reg_raw_inst[15:0] };
  assign csr_io_interrupts_debug = io_interrupts_debug;
  assign csr_io_interrupts_meip = io_interrupts_meip;
  assign csr_io_interrupts_msip = io_interrupts_msip;
  assign csr_io_interrupts_mtip = io_interrupts_mtip;
  assign csr_io_pc = wb_reg_pc;
  assign csr_io_rw_addr = wb_reg_inst[31:20];
  assign csr_io_rw_cmd[1:0] = wb_ctrl_csr[1:0];
  assign csr_io_rw_wdata = wb_reg_wdata;
  assign csr_io_status_debug = bpu_io_status_debug;
  assign csr_io_ungated_clock = clock;
  assign csr_reset = reset;
  assign div_clock = clock;
  assign div_io_req_bits_fn = ex_ctrl_alu_fn;
  assign div_io_req_bits_in1 = _ex_op1_T;
  assign div_io_req_bits_in2 = _ex_op2_T;
  assign div_io_req_bits_tag = ex_reg_inst[11:7];
  assign div_reset = reset;
  assign dmem_resp_waddr = io_dmem_resp_bits_tag[5:1];
  assign ex_ctrl_fp = 1'h0;
  assign ex_ctrl_mem_cmd[4] = 1'h0;
  assign ex_ctrl_mul = 1'h0;
  assign ex_ctrl_rfs1 = 1'h0;
  assign ex_ctrl_rfs2 = 1'h0;
  assign ex_ctrl_rocc = 1'h0;
  assign ex_ctrl_wfd = 1'h0;
  assign ex_dcache_tag = { ex_reg_inst[11:7], 1'h0 };
  assign ex_rs_1 = _ex_op2_T;
  assign ex_waddr = ex_reg_inst[11:7];
  assign ibuf_clock = clock;
  assign ibuf_io_imem_bits_data = io_imem_resp_bits_data;
  assign ibuf_io_imem_bits_pc = io_imem_resp_bits_pc;
  assign ibuf_io_imem_bits_replay = io_imem_resp_bits_replay;
  assign ibuf_io_imem_bits_xcpt_ae_inst = io_imem_resp_bits_xcpt_ae_inst;
  assign ibuf_io_imem_valid = io_imem_resp_valid;
  assign ibuf_io_inst_0_bits_inst_bits = csr_io_decode_0_inst;
  assign ibuf_io_pc = bpu_io_pc;
  assign ibuf_reset = reset;
  assign id_amo_aq = csr_io_decode_0_inst[26];
  assign id_amo_rl = csr_io_decode_0_inst[25];
  assign id_ctrl_decoder_1 = 1'h0;
  assign id_ctrl_decoder_15[4] = 1'h0;
  assign id_ctrl_decoder_16 = 1'h0;
  assign id_ctrl_decoder_17 = 1'h0;
  assign id_ctrl_decoder_19 = 1'h0;
  assign id_ctrl_decoder_2 = 1'h0;
  assign id_ctrl_decoder_20 = 1'h0;
  assign id_ctrl_decoder_27 = 1'h0;
  assign id_ctrl_decoder_8 = 1'h0;
  assign id_ctrl_decoder_decoded_andMatrixInput_0 = csr_io_decode_0_inst[0];
  assign id_ctrl_decoder_decoded_andMatrixInput_1 = csr_io_decode_0_inst[1];
  assign id_ctrl_decoder_decoded_andMatrixInput_10 = _id_ctrl_decoder_decoded_T_118[5];
  assign id_ctrl_decoder_decoded_andMatrixInput_10_20 = csr_io_decode_0_inst[27];
  assign id_ctrl_decoder_decoded_andMatrixInput_11 = _id_ctrl_decoder_decoded_T_106[5];
  assign id_ctrl_decoder_decoded_andMatrixInput_11_1 = _id_ctrl_decoder_decoded_T_106[1];
  assign id_ctrl_decoder_decoded_andMatrixInput_12 = _id_ctrl_decoder_decoded_T_106[4];
  assign id_ctrl_decoder_decoded_andMatrixInput_12_2 = _id_ctrl_decoder_decoded_T_118[15];
  assign id_ctrl_decoder_decoded_andMatrixInput_12_25 = csr_io_decode_0_inst[29];
  assign id_ctrl_decoder_decoded_andMatrixInput_12_33 = csr_io_decode_0_inst[31];
  assign id_ctrl_decoder_decoded_andMatrixInput_13 = _id_ctrl_decoder_decoded_T_106[3];
  assign id_ctrl_decoder_decoded_andMatrixInput_13_1 = _id_ctrl_decoder_decoded_T_118[14];
  assign id_ctrl_decoder_decoded_andMatrixInput_13_19 = csr_io_decode_0_inst[28];
  assign id_ctrl_decoder_decoded_andMatrixInput_14 = _id_ctrl_decoder_decoded_T_106[2];
  assign id_ctrl_decoder_decoded_andMatrixInput_14_1 = _id_ctrl_decoder_decoded_T_118[13];
  assign id_ctrl_decoder_decoded_andMatrixInput_15 = _id_ctrl_decoder_decoded_T_106[0];
  assign id_ctrl_decoder_decoded_andMatrixInput_15_1 = _id_ctrl_decoder_decoded_T_118[12];
  assign id_ctrl_decoder_decoded_andMatrixInput_15_14 = csr_io_decode_0_inst[30];
  assign id_ctrl_decoder_decoded_andMatrixInput_16 = _id_ctrl_decoder_decoded_T_118[11];
  assign id_ctrl_decoder_decoded_andMatrixInput_17 = _id_ctrl_decoder_decoded_T_114[8];
  assign id_ctrl_decoder_decoded_andMatrixInput_17_3 = csr_io_decode_0_inst[20];
  assign id_ctrl_decoder_decoded_andMatrixInput_17_5 = csr_io_decode_0_inst[21];
  assign id_ctrl_decoder_decoded_andMatrixInput_18 = _id_ctrl_decoder_decoded_T_114[7];
  assign id_ctrl_decoder_decoded_andMatrixInput_19 = _id_ctrl_decoder_decoded_T_114[6];
  assign id_ctrl_decoder_decoded_andMatrixInput_19_3 = csr_io_decode_0_inst[22];
  assign id_ctrl_decoder_decoded_andMatrixInput_2 = _id_ctrl_decoder_decoded_T[5];
  assign id_ctrl_decoder_decoded_andMatrixInput_20 = _id_ctrl_decoder_decoded_T_114[5];
  assign id_ctrl_decoder_decoded_andMatrixInput_20_6 = csr_io_decode_0_inst[24];
  assign id_ctrl_decoder_decoded_andMatrixInput_2_5 = csr_io_decode_0_inst[2];
  assign id_ctrl_decoder_decoded_andMatrixInput_3 = _id_ctrl_decoder_decoded_T[4];
  assign id_ctrl_decoder_decoded_andMatrixInput_3_5 = csr_io_decode_0_inst[3];
  assign id_ctrl_decoder_decoded_andMatrixInput_4 = _id_ctrl_decoder_decoded_T[3];
  assign id_ctrl_decoder_decoded_andMatrixInput_4_18 = _id_ctrl_decoder_decoded_T_118[23];
  assign id_ctrl_decoder_decoded_andMatrixInput_4_6 = csr_io_decode_0_inst[4];
  assign id_ctrl_decoder_decoded_andMatrixInput_5 = _id_ctrl_decoder_decoded_T[2];
  assign id_ctrl_decoder_decoded_andMatrixInput_5_18 = _id_ctrl_decoder_decoded_T_118[22];
  assign id_ctrl_decoder_decoded_andMatrixInput_5_8 = csr_io_decode_0_inst[5];
  assign id_ctrl_decoder_decoded_andMatrixInput_6 = _id_ctrl_decoder_decoded_T[1];
  assign id_ctrl_decoder_decoded_andMatrixInput_6_1 = _id_ctrl_decoder_decoded_T_112[6];
  assign id_ctrl_decoder_decoded_andMatrixInput_6_12 = csr_io_decode_0_inst[6];
  assign id_ctrl_decoder_decoded_andMatrixInput_6_17 = _id_ctrl_decoder_decoded_T_118[21];
  assign id_ctrl_decoder_decoded_andMatrixInput_7 = _id_ctrl_decoder_decoded_T[0];
  assign id_ctrl_decoder_decoded_andMatrixInput_7_15 = _id_ctrl_decoder_decoded_T_118[20];
  assign id_ctrl_decoder_decoded_andMatrixInput_7_17 = csr_io_decode_0_inst[12];
  assign id_ctrl_decoder_decoded_andMatrixInput_7_2 = _id_ctrl_decoder_decoded_T_10[0];
  assign id_ctrl_decoder_decoded_andMatrixInput_7_24 = csr_io_decode_0_inst[13];
  assign id_ctrl_decoder_decoded_andMatrixInput_7_50 = csr_io_decode_0_inst[25];
  assign id_ctrl_decoder_decoded_andMatrixInput_7_54 = _id_ctrl_decoder_decoded_T_114[9];
  assign id_ctrl_decoder_decoded_andMatrixInput_8_22 = csr_io_decode_0_inst[14];
  assign id_ctrl_decoder_decoded_andMatrixInput_8_8 = _id_ctrl_decoder_decoded_T_118[19];
  assign id_ctrl_decoder_decoded_hi_58 = { csr_io_decode_0_inst[0], csr_io_decode_0_inst[1], csr_io_decode_0_inst[2], csr_io_decode_0_inst[3], _id_ctrl_decoder_decoded_T[3], csr_io_decode_0_inst[5], _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T_112[6], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0] };
  assign id_ctrl_decoder_decoded_hi_lo_17 = { _id_ctrl_decoder_decoded_T_118[20:19], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[15:14] };
  assign id_ctrl_decoder_decoded_hi_lo_18 = { _id_ctrl_decoder_decoded_T_118[22:19], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[15] };
  assign id_ctrl_decoder_decoded_hi_lo_62 = { _id_ctrl_decoder_decoded_T_118[19], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[15:13] };
  assign id_ctrl_decoder_decoded_invInputs[31:2] = { _id_ctrl_decoder_decoded_T_106[0], _id_ctrl_decoder_decoded_T_106[1], _id_ctrl_decoder_decoded_T_106[2], _id_ctrl_decoder_decoded_T_106[3], _id_ctrl_decoder_decoded_T_106[4], _id_ctrl_decoder_decoded_T_106[5], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_114[5], _id_ctrl_decoder_decoded_T_114[6], _id_ctrl_decoder_decoded_T_114[7], _id_ctrl_decoder_decoded_T_114[8], _id_ctrl_decoder_decoded_T_114[9], _id_ctrl_decoder_decoded_T_118[11], _id_ctrl_decoder_decoded_T_118[12], _id_ctrl_decoder_decoded_T_118[13], _id_ctrl_decoder_decoded_T_118[14], _id_ctrl_decoder_decoded_T_118[15], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_112[6], _id_ctrl_decoder_decoded_T_118[19], _id_ctrl_decoder_decoded_T_118[20], _id_ctrl_decoder_decoded_T_118[21], _id_ctrl_decoder_decoded_T_118[22], _id_ctrl_decoder_decoded_T_118[23], _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T[2], _id_ctrl_decoder_decoded_T[3], _id_ctrl_decoder_decoded_T[4], _id_ctrl_decoder_decoded_T[5] };
  assign { id_ctrl_decoder_decoded_invMatrixOutputs[39:38], id_ctrl_decoder_decoded_invMatrixOutputs[32], id_ctrl_decoder_decoded_invMatrixOutputs[18], id_ctrl_decoder_decoded_invMatrixOutputs[13:9], id_ctrl_decoder_decoded_invMatrixOutputs[0] } = 10'h000;
  assign id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_lo[2] = 1'h0;
  assign { id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi[8], id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi[3:0] } = 5'h00;
  assign { id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo[9], id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo[0] } = 2'h0;
  assign id_ctrl_decoder_decoded_lo_11 = { _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:2], _id_ctrl_decoder_decoded_T_106[0] };
  assign id_ctrl_decoder_decoded_lo_12 = _id_ctrl_decoder_decoded_T_106[5:0];
  assign id_ctrl_decoder_decoded_lo_18 = { _id_ctrl_decoder_decoded_T_118[13:11], _id_ctrl_decoder_decoded_T_114[8:5], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign id_ctrl_decoder_decoded_lo_19 = { _id_ctrl_decoder_decoded_T_118[14:11], _id_ctrl_decoder_decoded_T_114[8:5], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign id_ctrl_decoder_decoded_lo_22 = { _id_ctrl_decoder_decoded_T[0], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign id_ctrl_decoder_decoded_lo_29 = { _id_ctrl_decoder_decoded_T[1], _id_ctrl_decoder_decoded_T_112[6], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_106[4:3] };
  assign id_ctrl_decoder_decoded_lo_31 = { _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign id_ctrl_decoder_decoded_lo_35 = { csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign id_ctrl_decoder_decoded_lo_37 = { csr_io_decode_0_inst[14], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign id_ctrl_decoder_decoded_lo_39 = { csr_io_decode_0_inst[14], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:2], _id_ctrl_decoder_decoded_T_106[0] };
  assign id_ctrl_decoder_decoded_lo_40 = { _id_ctrl_decoder_decoded_T[0], csr_io_decode_0_inst[14], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:2], _id_ctrl_decoder_decoded_T_106[0] };
  assign id_ctrl_decoder_decoded_lo_41 = { csr_io_decode_0_inst[14], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign id_ctrl_decoder_decoded_lo_53 = { csr_io_decode_0_inst[25], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign id_ctrl_decoder_decoded_lo_56 = { _id_ctrl_decoder_decoded_T_112[6], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0], csr_io_decode_0_inst[27], _id_ctrl_decoder_decoded_T_106[2:0] };
  assign id_ctrl_decoder_decoded_lo_57 = { _id_ctrl_decoder_decoded_T_114[7:5], _id_ctrl_decoder_decoded_T_106[4], csr_io_decode_0_inst[28], _id_ctrl_decoder_decoded_T_106[2:0] };
  assign id_ctrl_decoder_decoded_lo_58 = { _id_ctrl_decoder_decoded_T_114[9:5], _id_ctrl_decoder_decoded_T_106[4], csr_io_decode_0_inst[28], _id_ctrl_decoder_decoded_T_106[2:0] };
  assign id_ctrl_decoder_decoded_lo_59 = { _id_ctrl_decoder_decoded_T_118[13:11], csr_io_decode_0_inst[20], _id_ctrl_decoder_decoded_T_114[8], csr_io_decode_0_inst[22], _id_ctrl_decoder_decoded_T_114[6:5], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:4], csr_io_decode_0_inst[28], _id_ctrl_decoder_decoded_T_106[1:0] };
  assign id_ctrl_decoder_decoded_lo_60 = { _id_ctrl_decoder_decoded_T_118[14:11], csr_io_decode_0_inst[20], _id_ctrl_decoder_decoded_T_114[8], csr_io_decode_0_inst[22], _id_ctrl_decoder_decoded_T_114[6:5], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:4], csr_io_decode_0_inst[28], _id_ctrl_decoder_decoded_T_106[1:0] };
  assign id_ctrl_decoder_decoded_lo_61 = { csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0], csr_io_decode_0_inst[27], csr_io_decode_0_inst[28], _id_ctrl_decoder_decoded_T_106[2:0] };
  assign id_ctrl_decoder_decoded_lo_62 = { _id_ctrl_decoder_decoded_T_112[6], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_106[4:3], csr_io_decode_0_inst[29] };
  assign id_ctrl_decoder_decoded_lo_63 = { _id_ctrl_decoder_decoded_T_118[12:11], _id_ctrl_decoder_decoded_T_114[9], csr_io_decode_0_inst[21], _id_ctrl_decoder_decoded_T_114[7:5], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:4], csr_io_decode_0_inst[28], csr_io_decode_0_inst[29], _id_ctrl_decoder_decoded_T_106[1:0] };
  assign id_ctrl_decoder_decoded_lo_64 = { _id_ctrl_decoder_decoded_T_118[14:11], _id_ctrl_decoder_decoded_T_114[9], csr_io_decode_0_inst[21], _id_ctrl_decoder_decoded_T_114[7:5], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:4], csr_io_decode_0_inst[28], csr_io_decode_0_inst[29], _id_ctrl_decoder_decoded_T_106[1:0] };
  assign id_ctrl_decoder_decoded_lo_65 = { _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:2], csr_io_decode_0_inst[30], _id_ctrl_decoder_decoded_T_106[0] };
  assign id_ctrl_decoder_decoded_lo_66 = { _id_ctrl_decoder_decoded_T_112[6], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_106[4:3], csr_io_decode_0_inst[30] };
  assign id_ctrl_decoder_decoded_lo_67 = { csr_io_decode_0_inst[14], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:2], csr_io_decode_0_inst[30], _id_ctrl_decoder_decoded_T_106[0] };
  assign id_ctrl_decoder_decoded_lo_68 = { _id_ctrl_decoder_decoded_T_118[12:11], _id_ctrl_decoder_decoded_T_114[9], csr_io_decode_0_inst[21], _id_ctrl_decoder_decoded_T_114[7:6], csr_io_decode_0_inst[24], csr_io_decode_0_inst[25], _id_ctrl_decoder_decoded_T_106[5], csr_io_decode_0_inst[27], csr_io_decode_0_inst[28], csr_io_decode_0_inst[29], csr_io_decode_0_inst[30], _id_ctrl_decoder_decoded_T_106[0] };
  assign id_ctrl_decoder_decoded_lo_69 = { _id_ctrl_decoder_decoded_T_118[14:11], _id_ctrl_decoder_decoded_T_114[9], csr_io_decode_0_inst[21], _id_ctrl_decoder_decoded_T_114[7:6], csr_io_decode_0_inst[24], csr_io_decode_0_inst[25], _id_ctrl_decoder_decoded_T_106[5], csr_io_decode_0_inst[27], csr_io_decode_0_inst[28], csr_io_decode_0_inst[29], csr_io_decode_0_inst[30], _id_ctrl_decoder_decoded_T_106[0] };
  assign id_ctrl_decoder_decoded_lo_70 = { _id_ctrl_decoder_decoded_T_112[6], csr_io_decode_0_inst[13], _id_ctrl_decoder_decoded_T_10[0], _id_ctrl_decoder_decoded_T_106[4:3], csr_io_decode_0_inst[31] };
  assign id_ctrl_decoder_decoded_lo_lo_15 = { _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:0] };
  assign id_ctrl_decoder_decoded_lo_lo_56 = { _id_ctrl_decoder_decoded_T_114[5], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:4], csr_io_decode_0_inst[28], _id_ctrl_decoder_decoded_T_106[1:0] };
  assign id_ctrl_decoder_decoded_lo_lo_60 = { _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:4], csr_io_decode_0_inst[28], csr_io_decode_0_inst[29], _id_ctrl_decoder_decoded_T_106[1:0] };
  assign id_ctrl_decoder_decoded_lo_lo_61 = { _id_ctrl_decoder_decoded_T_114[5], _id_ctrl_decoder_decoded_T_118[5], _id_ctrl_decoder_decoded_T_106[5:4], csr_io_decode_0_inst[28], csr_io_decode_0_inst[29], _id_ctrl_decoder_decoded_T_106[1:0] };
  assign id_ctrl_decoder_decoded_lo_lo_65 = { csr_io_decode_0_inst[25], _id_ctrl_decoder_decoded_T_106[5], csr_io_decode_0_inst[27], csr_io_decode_0_inst[28], csr_io_decode_0_inst[29], csr_io_decode_0_inst[30], _id_ctrl_decoder_decoded_T_106[0] };
  assign id_ctrl_decoder_decoded_lo_lo_66 = { csr_io_decode_0_inst[24], csr_io_decode_0_inst[25], _id_ctrl_decoder_decoded_T_106[5], csr_io_decode_0_inst[27], csr_io_decode_0_inst[28], csr_io_decode_0_inst[29], csr_io_decode_0_inst[30], _id_ctrl_decoder_decoded_T_106[0] };
  assign { id_ctrl_decoder_decoded_orMatrixOutputs[39:38], id_ctrl_decoder_decoded_orMatrixOutputs[32], id_ctrl_decoder_decoded_orMatrixOutputs[18], id_ctrl_decoder_decoded_orMatrixOutputs[13:9], id_ctrl_decoder_decoded_orMatrixOutputs[0] } = 10'h000;
  assign id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_6[2] = 1'h0;
  assign { id_ctrl_decoder_decoded_orMatrixOutputs_lo_17[18], id_ctrl_decoder_decoded_orMatrixOutputs_lo_17[13:9], id_ctrl_decoder_decoded_orMatrixOutputs_lo_17[0] } = 7'h00;
  assign { id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_10[9], id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_10[0] } = 2'h0;
  assign id_ctrl_decoder_decoded_plaInput = csr_io_decode_0_inst;
  assign id_fence_succ = csr_io_decode_0_inst[23:20];
  assign id_raddr1 = ibuf_io_inst_0_bits_inst_rs1;
  assign id_raddr2 = ibuf_io_inst_0_bits_inst_rs2;
  assign id_waddr = ibuf_io_inst_0_bits_inst_rd;
  assign inst[15:0] = ibuf_io_inst_0_bits_raw[15:0];
  assign io_dmem_req_bits_addr = alu_io_adder_out;
  assign io_dmem_req_bits_cmd = { 1'h0, ex_ctrl_mem_cmd[3:0] };
  assign io_dmem_req_bits_dv = 1'h0;
  assign io_dmem_req_bits_size = ex_reg_mem_size;
  assign io_dmem_req_bits_tag = { 1'h0, ex_reg_inst[11:7], 1'h0 };
  assign io_dmem_s1_data_data = mem_reg_rs2;
  assign io_imem_might_request = imem_might_request_reg;
  assign io_imem_req_valid = ibuf_io_kill;
  assign io_imem_resp_ready = ibuf_io_imem_ready;
  assign { io_ptw_customCSRs_csrs_0_value[31:2], io_ptw_customCSRs_csrs_0_value[0] } = { csr_io_customCSRs_0_value[31:2], csr_io_customCSRs_0_value[0] };
  assign io_ptw_pmp_0_addr = csr_io_pmp_0_addr;
  assign io_ptw_pmp_0_cfg_a = csr_io_pmp_0_cfg_a;
  assign io_ptw_pmp_0_cfg_l = csr_io_pmp_0_cfg_l;
  assign io_ptw_pmp_0_cfg_r = csr_io_pmp_0_cfg_r;
  assign io_ptw_pmp_0_cfg_w = csr_io_pmp_0_cfg_w;
  assign io_ptw_pmp_0_cfg_x = csr_io_pmp_0_cfg_x;
  assign io_ptw_pmp_0_mask = csr_io_pmp_0_mask;
  assign io_ptw_pmp_1_addr = csr_io_pmp_1_addr;
  assign io_ptw_pmp_1_cfg_a = csr_io_pmp_1_cfg_a;
  assign io_ptw_pmp_1_cfg_l = csr_io_pmp_1_cfg_l;
  assign io_ptw_pmp_1_cfg_r = csr_io_pmp_1_cfg_r;
  assign io_ptw_pmp_1_cfg_w = csr_io_pmp_1_cfg_w;
  assign io_ptw_pmp_1_cfg_x = csr_io_pmp_1_cfg_x;
  assign io_ptw_pmp_1_mask = csr_io_pmp_1_mask;
  assign io_ptw_pmp_2_addr = csr_io_pmp_2_addr;
  assign io_ptw_pmp_2_cfg_a = csr_io_pmp_2_cfg_a;
  assign io_ptw_pmp_2_cfg_l = csr_io_pmp_2_cfg_l;
  assign io_ptw_pmp_2_cfg_r = csr_io_pmp_2_cfg_r;
  assign io_ptw_pmp_2_cfg_w = csr_io_pmp_2_cfg_w;
  assign io_ptw_pmp_2_cfg_x = csr_io_pmp_2_cfg_x;
  assign io_ptw_pmp_2_mask = csr_io_pmp_2_mask;
  assign io_ptw_pmp_3_addr = csr_io_pmp_3_addr;
  assign io_ptw_pmp_3_cfg_a = csr_io_pmp_3_cfg_a;
  assign io_ptw_pmp_3_cfg_l = csr_io_pmp_3_cfg_l;
  assign io_ptw_pmp_3_cfg_r = csr_io_pmp_3_cfg_r;
  assign io_ptw_pmp_3_cfg_w = csr_io_pmp_3_cfg_w;
  assign io_ptw_pmp_3_cfg_x = csr_io_pmp_3_cfg_x;
  assign io_ptw_pmp_3_mask = csr_io_pmp_3_mask;
  assign io_ptw_pmp_4_addr = csr_io_pmp_4_addr;
  assign io_ptw_pmp_4_cfg_a = csr_io_pmp_4_cfg_a;
  assign io_ptw_pmp_4_cfg_l = csr_io_pmp_4_cfg_l;
  assign io_ptw_pmp_4_cfg_r = csr_io_pmp_4_cfg_r;
  assign io_ptw_pmp_4_cfg_w = csr_io_pmp_4_cfg_w;
  assign io_ptw_pmp_4_cfg_x = csr_io_pmp_4_cfg_x;
  assign io_ptw_pmp_4_mask = csr_io_pmp_4_mask;
  assign io_ptw_pmp_5_addr = csr_io_pmp_5_addr;
  assign io_ptw_pmp_5_cfg_a = csr_io_pmp_5_cfg_a;
  assign io_ptw_pmp_5_cfg_l = csr_io_pmp_5_cfg_l;
  assign io_ptw_pmp_5_cfg_r = csr_io_pmp_5_cfg_r;
  assign io_ptw_pmp_5_cfg_w = csr_io_pmp_5_cfg_w;
  assign io_ptw_pmp_5_cfg_x = csr_io_pmp_5_cfg_x;
  assign io_ptw_pmp_5_mask = csr_io_pmp_5_mask;
  assign io_ptw_pmp_6_addr = csr_io_pmp_6_addr;
  assign io_ptw_pmp_6_cfg_a = csr_io_pmp_6_cfg_a;
  assign io_ptw_pmp_6_cfg_l = csr_io_pmp_6_cfg_l;
  assign io_ptw_pmp_6_cfg_r = csr_io_pmp_6_cfg_r;
  assign io_ptw_pmp_6_cfg_w = csr_io_pmp_6_cfg_w;
  assign io_ptw_pmp_6_cfg_x = csr_io_pmp_6_cfg_x;
  assign io_ptw_pmp_6_mask = csr_io_pmp_6_mask;
  assign io_ptw_pmp_7_addr = csr_io_pmp_7_addr;
  assign io_ptw_pmp_7_cfg_a = csr_io_pmp_7_cfg_a;
  assign io_ptw_pmp_7_cfg_l = csr_io_pmp_7_cfg_l;
  assign io_ptw_pmp_7_cfg_r = csr_io_pmp_7_cfg_r;
  assign io_ptw_pmp_7_cfg_w = csr_io_pmp_7_cfg_w;
  assign io_ptw_pmp_7_cfg_x = csr_io_pmp_7_cfg_x;
  assign io_ptw_pmp_7_mask = csr_io_pmp_7_mask;
  assign io_ptw_status_debug = bpu_io_status_debug;
  assign io_rocc_cmd_valid = 1'h0;
  assign io_wfi = csr_io_status_wfi;
  assign ll_wdata = div_io_resp_bits_data;
  assign mem_br_target[0] = mem_reg_pc[0];
  assign mem_br_target_b10_5 = mem_reg_inst[30:25];
  assign mem_br_target_b4_1 = mem_reg_inst[11:8];
  assign mem_br_target_hi_hi_hi = mem_reg_inst[31];
  assign mem_br_target_hi_hi_lo = { mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31] };
  assign mem_br_target_hi_lo_hi = { mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31], mem_reg_inst[31] };
  assign mem_br_target_hi_lo_hi_1 = mem_reg_inst[19:12];
  assign mem_br_target_hi_lo_lo = mem_reg_inst[7];
  assign mem_br_target_hi_lo_lo_1 = mem_reg_inst[20];
  assign mem_br_target_sign = mem_reg_inst[31];
  assign mem_ctrl_fp = 1'h0;
  assign mem_ctrl_mul = 1'h0;
  assign mem_ctrl_rocc = 1'h0;
  assign mem_ldst_cause[1] = 1'h1;
  assign mem_npc[0] = 1'h0;
  assign mem_reg_hls_or_dv = 1'h0;
  assign mem_waddr = mem_reg_inst[11:7];
  assign r = { _r[31:1], 1'h0 };
  assign replay_wb_rocc = 1'h0;
  assign rf_MPORT_mask = 1'h1;
  assign rf_id_rs_MPORT_1_en = 1'h1;
  assign rf_id_rs_MPORT_en = 1'h1;
  assign size = ex_reg_mem_size;
  assign take_pc_mem_wb = ibuf_io_kill;
  assign wb_ctrl_rocc = 1'h0;
  assign wb_reg_hls_or_dv = 1'h0;
  assign wb_valid = csr_io_retire;
  assign wb_waddr = wb_reg_inst[11:7];
  assign wb_xcpt = csr_io_exception;
endmodule
